-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Zezlmd/LTABzDx7rT0lAZJBFfElFathgwD9/6SrI4b6VIxEg+dM16SixnCqALGl7
9VTD8EscOfBrM2l6uYKocunolFmjY2RIxCbVqF8YJSOGwlvZ3KsvHONvrFkKWOi2
KM3RJkS3Y0m2h/UFCy75Kgh1KhHKkNBzw28oqedBo5mjLTDAcgEUnQ==
--pragma protect end_key_block
--pragma protect digest_block
zUXW8wMDDFfqT2g5/dT6yF+fHdQ=
--pragma protect end_digest_block
--pragma protect data_block
HuBCtV1crkAUF0wJOacUUKHpFLyCcPS0ReHQJdqGUU23gaZ6Y7Jh9LvPlC5hAbtZ
uPWtM/mtgF7NYJBBnfxAnlrEEtI9Pj5zNxV+ESoVJD8IfskmTaYMfpOLETwwjp4o
Pmou4HeBrPBMZsRwsb3+MBFUxYrtkr1o7phDRP/SxzxSij1Odyd5ObyFhL5ZS8fn
8OGoBUYUFEo1ocwF+PGAdiu/r143yPbUb0Adtk4VDSUeSHbpUYOepcLRNSf+8zea
Vaa6uGPio9hfTa1g1VBWzZj1H1co4gzhg9IaTKi+44gSUvSSLFWWYByjDdzZYwux
3CfL+A4J3e7o63OBS7UbBt7JyhDG5k1nzMGsC/t8G9IcboKvUNJ6yNZV+qHQYtto
yxLU6l4LPl7OuZSc+dsblHhSrnGZ6wAV2PKFTgpKBZmmelQTZegrZ+EQcAv7Xpwo
4Hqqz8hyWTDm6m7jxlx+sVFnICFbsqSWrSITx4xFGsInAf/OumtW11VETzIhkR34
dsPlqF5z5P3ppnNVxoQviLYKXKQfK8XBEp11a+LJKjVxCInMGezbR2xSff6VDRrW
ZY/DmQXEVyAGlbmyTp5etuouwh6YSgATsQNLLlxdSCXxjX0o+w2d1EdBfxUcdIxd
r1JWL4mHy7XzA0J2L9Y3eQBR7H/KLACRYPzPZm+Kpi9lMsDoXxCbTQYXwnkhPJnI
CEiMm7mxQQ5lB4/0RzlAdAfBHfWvfQoOyOOqSoj+ed1jm/bsUV+f4ahaJacvEOK5
UUuossdn5/jsVYtWd8uApw+mFHDaQQVR3N6WVyoNf1fXiX+zhqowEI24vEiuLDxg
NqqZ2WyVwI6FbfFbfuVzo6JMTylM1AXh9P+RYuC0dzcN17PVS6NiTeSsWJjyyhV8
Bh/aKYX3U/2D9oSgoqqvj01O1GzMh+m1lURTACKxoltMzfQB4sRkgmgebonogqCc
+pplDbSItdjngkNnVxDSq7h++dC3arBIWlO8r3kw57gJRLLd/+mu7XY45QqdZ/Wt
3gtvHDIRNMRTImMJiJpcX3e8jttya3XB+GwCmqDmb+zv0dmjy0cSoMFG2Ph1Wydp
VVxWSdI2y92jpYCCSzYbO+z/Foo0u8kTbrxk3WefTUUln5ggA6/7f21fH+SpY/PV
nWl52abMkuH2ste8mMqhP7E4M76/ZkL4Y2heew/Rt9CIBEGFLEQLAK2GE3jwUV6w
USUYMMrPfneDaiuxbN0adrpfYs05H2OXanAeg8lEHuIm0n3zpWq2yUt0cOflkj6Y
tVeDEEEny4i7wGoVyk4qvKG54HhlkvrNkRg4hy5DhOPbRj/UNczW53yTv+1n4DPn
O1kaDY5TpXl6ACF9FBkHuTfU3dUqU8GXCRLs+fka/3Falxa/VHLNOPs1yz/A/3ZB
TTqNgDbq2LXS9MEOh0UCs+Gd05zq/7PNkyqtq6jUsZTXT5u1rZC94O1MXgyVCree
tf3n5RoJUe2ivhqE1iDSJOnizUaqm+WBnPHxn4CPZKek+szi6b4NmSF+HF9LKtjU
VQwfmtGuXT6d2IFr6f9wrJjQqtpMHbUHyVl0sUKpRyHFYlBdDIb06c6yYoyc0EVs
KvnqZYhxxHadbWLVQbtZIROI2JgJSfslfigoliphq12jucE5VaF0hT9UCNFGbuOH
v7hBIbOsggaNYLTfdeUywUxEFk1efQ5hbdZ4V3afOV8EkzF67M/8AzY0q9SUIj6k
BptvoVpnE/6yvqtxw5Hta+VJBaIZCpg6xi6Me2A35ax++M3HN2EWOqdNYXq00FoG
B8rRj4HqYmKUpGJNBk6N9BoU55taRs3eXngpCsjx4V78lm8MDUHOi0waynKcLRxF
bWK6L3QFEuXdYYF/N32JxPFw2OeZ/YZmJHE8D44WRfH8cwFp6Hua5PsP+wY5Q/ov
Mx0M7mZ9/AvwSqYceZ6qDzy5L+Hq29SJibhlKRSOISGNpC/B+n65zY3tB/y5Q5/7
n3pHfVve6zdKDVvrPqsfl1fOYxBw5KK1J+bNmQoETo1ZtWJH6xWB2PgFhQ+PFP4l
UDIekKfc4MqqddE0TpoYDA0vg1DrFwQle44w8SS6dzquwwDAxDLjjCUiPK3Uttlv
b3Cpd2/KvAmEZ8pdA8SbETbFPVlKIEz0qyIBWg9xyoE7BDhly0CBXfOY9rCkscJB
GrMMwPSh3Yg594VcKtX6WC0Xv8/Mb3qdSQbiPAQlkih0/3hzMtiJsKoJNaSPk+iV
/vEd+u3ntlwQ7/CEgDiUlDTei6CLzNhgQw7TacTO1EUzq4q0HRv3bu4QgJx5cNV1
J96qfuG/QjClHM/eciMDoqK1L4ZsmALrubp+QMBEIIdPUfIWUrps4JjQ67T0bZU+
kB+2R+TJdGjrGZsCwclOiovCGL9iPt+6OSQR8DafGZZzUxzQOPncJ9/zWkPMVVBc
NRY9dUanaJb0iRVj0ZDRltoWGbIbs1M3REXjhoqHl24VCLSK0xgYaJBFCW/06OcP
g44xxDldSHUedAoFo4nz0qvBYCKOcNglW1Zegxqqsi6cRJVbYW18YCA7MuchCzpI
sA0VgBYvpcXzUniT0odsxfvaNzLXpbEGyLvXO7egQMosokAl0C/EyfpbuYYVuKkx
T9ifFEYZVlRXeQ3Br6nuARc7M1We1HYHBfvg4TvshBYN0KojQu56A91h+IikCgLi
I9jOfJNssrmuZsuOQ7GOEaKHrwECbm58kFLVf7VxU3nkJ2SZz5Qz2R8dZwgMpzwS
4Rvm0ACEpZvferRssYUPYvKFzH3zlSPobmYDZJV2FXHateNomifkjfLPzqGxRuQF
9h6mMA0/lUtIEB420aV7/sqOKtZg2aLw2e0b5jj64R2Vqv+Hr9EXWTXPH2ns6Sm3
hXu/NlsAtSmT3uDTjztYkP1JEnwfgcv7nkBwprqgyTgSH6L0R61H3xwbO+zox48F
udJn4swkr9dEPWuocioY3CB2zHoQlx6dXA19KW4RKb2zn3+1OpgVTZm8wPQziPll
IXWq2jUlxlSR4+1qvl/DW2tGz2uy7Gkf111ZB3Sd26KFJoI3ZCWsuFGBka22xbzc
KvQt7Fz0X0WrB6EfJ/aDvJnFf0F2+KbnbGqpuvvC4XOAZkZ8/B6Yly8YdWeIdsq9
04XxZK3d3wGArJSK/dn/QjroNI6LE8Ficda8gHC/ZQJkOU6nbp9g+QWlHHL8yIOe
gjMhMaFkw6kLC6a9Vydty9wrn3z53TAI7UNJzaxpAu7zvNg1EihOa10BItLNO9Ja
L0HubhdS/k43NW9orTP17hnXkukkd4i9OCfoRSLcDDD4vGOtAtJ6s2FvShgbZn0+
+TyArRNrMlmIKsWI7lpD/yIGOYiGTAkmNhvS4unTEjAN/L4F4zTHkPvHdtPK9b7g
pcBUn5XFk02Kzm8dNy64uaC4kOY6RFAKm7lpmNU5BWfxibd7dXZgtN8Aao9oP6tP
bJ5iCr8wDDckEI4WJTpnyTXAVQxkDokOxlGMMdQfDZ7c4b56qRWyn4+4LmajHaup
HykLoo6888eYcfirtDrGAtVRAgOQxIeG2/xQDDRbDGwAS/xw7OKG66TsFa8vUJGr
HglTm6ks61JH8E+G8HM34tzFVYYdwI+AU9GwurX/ikld5+WpETf8Uv4EW784spzh
uLcTLVi4HUrXranHeaVelRymy6hWJ0KLVkmd9USD9w6/Yk66Fs9ntRejIOfCHb5t
BdygErFqrH6R6LAWqubDDcs/W30RvgDjcLUJ65hHCj/ZKGF9LuEf5cMeTrLNLD6D
/UdHo8ED2q55F05FDEXf5EAtWE73TG65HzrF8lhPYdKiuv97BjEFs73/5RmqambW
uxGSOvb7Kn848zKPc+czAy+xgvc7VeZ99IxQc5LtTw8LI+UnVI719dnjQHQang3R
3oWACwNdhSYEuczF6xFGuQrJ6s+Uu0odDybQp/YlxbF84K4kv3bADG1A1Egae3Yz
kRBeVeg3d6ev5sufTVaYSMlwfsYBUftdTh44Qs4VNwb8BHm0XR9ZjgW6jFZMDcP5
VNm6w0wF34OxZRrsL/K/zpegEY4CQYOAceJoeC3qvC1NLXYaZUeOMbbfAJ67cVsS
jgPqsVlIsKkcpWcZwGDTScv93hycCPTtd8jjxpD9e1J5iUsxxSsZfQNoz6rtOuyc
p+09eXQIN/cbnF3i/9THtZTNeD/LnrRV43VJc/IXB5RgIq+ex1bwOOZmTYyjTR08
WpjU1n3IQpj6D0Ik3ZKtMs8SVirJ6Sx5i71ach4Od56VR8380v2s5yxp2uec0O2B
jXYcqBR2RTVEAHRJAVPR46tLWWiWimdFNDwiIYuXNbVHYN5kGgQivETH79k/2UIW
zKfhLVGJU4inSd+8D4Q80WUWdmE67MB3Yg5lVoJuVnTc93wdHSLB/rvyQSutNDHX
o2dtTtzcSYBRCEBBcyOa12z/WVSEzoTrE94r9IQR0CSZYJw7xQ+e3cI0/uZk160L
T7LCCW6zrH5vjI126DB0d14pc+f3O95swI83uic877/RkLLKz4YDpLIZFoz/iWNs
YorNsQ5S3RRc+2ZH6OsiVngCgxEjs66mI8I9aB9yWaMU+GzwcbyR17wnS2DhAuFd
OS7DcBWokRwy02NaSuODajxsDeWskVQ6/4exIUY07WIWi8dR74UFwOBdN7wSwv0W
+wrXtC4XFbLCtTQdt0KV4DaWLnlAiqv4jD35DlfHEctV2gEZVG8OFFWVs4uP5XOZ
NNDnpGrYlN2fJC+AdpROjb84AbiXPX6UXYySS7ZF1+WWddxiuESV/n5BjfjIwHYJ
xPJfqZRvP5lgVLHww8pQRGmsZkRmsCGTqWGOwkXkFDcrYBBXarW/onyg2roHXYk8
UtcrEEf0lPNnI/FNZuTgOygK7xWcFhGzcO/Jyec5NJ7jizjDIOt4P/JIopt1WOqH
uNPbmTAPO/jV/Mg4SWbeVHCi0dGrf7g0svADHcesLPnxpKT//K0v5oMDYXRbvT4+
JpN0zNg1WimqCK89XkVG7JD+GGTotlP60yPoTpBYaLqvTiFc6qVwK/wO6jlT3yoY
CltCXlCGxk8VtIcIjn+GQreLA8xvbkm0lEcU9rhOExn3DyyXagmvkoNqjMnpGyxi
oEzUmLFCjdsX2KdYkcSvuuwTTz3E4Ay3NSWZPBhIsd0vxsn8zXtuVXlJZnCaBGEs
cnDHmFJWvmhYtBIuZgstevwHQ6LuYgGk3jvRRv1N6de278jpEOXI6MxexnJo/Z3I
vvzJE0PryNFD6FozdVkP95dUQPUtLRDPlDbDuxEOkovNRqFv66lrmEMZQ/mx/gqP
sLuVqbRuUfNlgoCesWJIhNjjVPKFstrpBajZn0hX7ZCD+BihHZWyhH5jl90KABrK
sM6DqIiw5jOZ5libivk6rpDY0t7yb7facXThUnB1H0PqgdhCqCroeZDJnibVmpkR
vnWmzuONqLwepTOs9uVfDw67PxGRtp1HtF0sW71fApohDGeOuk+pYdfHutfDbolw
Q7IThi3uvWw0QXh4lzObZxWE2TXE40SLJdiE4+wKJDjKVjVfFbfGn4JzKQapkIVE
pOd4bUEh65OG36Nz8IdAKD6roepN7wjrgoGKmSiv5FRLdkRHFA8gepyJjmvgiYFz
uiDiN8aV4kuPLhnq3aAL0V0q5PEySA0/D2GdzfepzAaKj6svjFBpXS6Ry2opaKR4
bUf/K+pZT7XouTw5kv9JuNlBMuZTEL3+BC2vQSMXMahcdkjLJKRuKM/69eXb/TeQ
rxQB+3UXJ3ajJZ8HRgF8KaCaUI7xKPkp9BTXYu3EfoBYFgYc5CbsS+SbIKGCXE9R
D2tG4bFt9Nxg2UdjSNll+9bee+Fd18K2YQAQH875hhmBK/dj11ZohasXnJ/zNcvT
z+/ZPECG8Xt9ZsukG4Px/vT350JCcDVsdRIAu2NGnufnIV4gzNGieNfitV5a9GBG
7iIenKY4OIHTWNaHEF+aa5u3qxQ0B2cSITYP7ItsFJywvQl2MiD/GOdRfDRZwPqE
NnUzQaoFVkyXNN3WVl/aJWOGKaF5+Yt6dYnsqkoNw5YxJPmF+uN7hrsqWA8Qbypk
8N3+GVYfoW7b66OasVQOJrbLe5zR/b4BcJ1jcXBaaQFNi4c0lgLKDd3fxDXqoiIK
oVrJmDtYVK04pt8knDdp+ogCTWMsw6AI52gHmIEABVPMzI3jBrp6RFivEVME4cpR
nPb96uuE3MD8K3E561Rl7GQEP6+wO+arYSZmbpL7INdZlTPQ716v2EsdI313f+V2
jAexIBbS6+proS/qOMh9rsUrn65NGFB+sJs11eb5XQ+86jR4j8F7y2OZHkCldTuT
TDD4v/fwR+DNOAYIFQbeiCsqjL+rWnsqQy4Hdk9DuNpRPTO7q+ber6V67bl7T4TE
T/t8NYmLEjp46W9i4YQcgfe4ufkz+lvNCFkzVgpTfjXunX/Vot54SD/8xIU/iHMf
75piI5GKPLOs7EgcEfRz0xpVTcUn5OSKszKUhxCKY4APDNTatCwhjskA/yroAYpn
lwxrA8NrJPLd9a/zcq6kqMqcOoEuddEYPcrCPim+cbXtBePwzoWLjrgmMrCry5TM
kr5DhaZ3IRSZm6DPPTWNAT5ti2scqtkaXsmWGdfBtgueOP1tTptnxKBZhsg4Z5tM
Hd5A4dMcvATNE/+o4Fm5RwXxOUpdgnkBZD94jvwIKs+0S5u2ljKNVWwAzkfI1IN4
e/wm7Z+z8eKmvAa9VTbl6NzfD9bOdr4WxLYuzFhBCNqwC0IppzPMnvGKqf6OB8CF
11sp9h4lCJTXhpWeBkONBjTnTFgj4zbB6t+ci95nhrJceSrxEDrGyVA5Mu3mJJq4
zUy9nzMSL5JSaeXc7PGt3IDKYmVypzDEAFQ8O6yWJjO2JuGQb/7zpbFca4ph6dHy
MUBpwNlbaWkt8/dccr0EkSbRlYWSqlRCPOMfru9AY+Bs/bG1Cd1hsSz1Mlwg5BJ0
Z4yEU4OJ9r0rq92btKIl/SesFqnh2JXCIL23yroj4I5j7nr9zck57FBgvj1V3335
3IeB+7Ky19NTMy4wUSYbBh25VvAP1XEWlfWwdIY7aw/92S/NiDSSPHTwX61RJd1S
n+wFHzJfmvQ+wfxAq9EOVZPP04C4U6vUpkfi1g/DKMxyudK+P8TqSxDJMObvvrCn
rT3KeydWzVGP5o4+btHLXqpyrjNBEGdJpFkxrVnaWGlaBoSkkF2vuLqhDUqPfcGV
HDoiBXJGeY6z370ZjLdBollInqOJN9j57BQoxuaoNW8vZmsGy2LTkzpjt43GQxBK
wt95nlTJvAzQOBuPnYPfUYLJUVY+96G0OPgQxIb6ShCoP9Aj835CCXRZwgYvzYfZ
vU+4MHr1LTS5cOUXrXDFryzpCEVe1D6bvfDdMTIAGiWezRqlYP1iG6VXutnuFEls
J/Nt/ymAfdsdiKt93NQO7qlRC7C7gChxPycr79fmQGE61lAMQtQVANvUKraCzfnX
Cm7lzNZs2yJShjrJdNT4wnCQzvgGPrhB1efp6GMKaU9ozwYqXz1bkEevQBObrJKA
7GirX8BcmIlhn59bWKMRAfLwycBUXNVUCNWY570ShkZK3OAVxqwOrGz4nhdtMq88
IcaAmm9EtC1urolUMHkMdTh5jin1WTH8yOWul3TVu75D1X8+BSYwimrdh7isuJfA
SCTOO2SHxKEpKBisviNlS+0MjHY0UX1SFV1szSE8KHBS7zngTK9YH2y1eXcAh1tU
wYKpLzwaHCxaE6zZR8s+eolZkGpgkw8zD2wCv5qduajJj+CCNf/8o1RfKcXFPDcL
GZq+bQXw9aFh05PWYorxRcsrLLTxJQk+jSK7XHqeJOnEVLCZrHyrHJQA9BitMcUl
+1oUiXyRBaJYm41urNaH3hKopih0m+2eRnW/Uob44IcX7n0ixUrAmnSE/lD+mpHU
Xg+DjtOoqYaf+Ppjv6fCoA5e6wMk4E9+Mbnl6z7TEqO+HQZoY9seYUJvIyvp6O1r
eo0meZdgWjCAuxnyO6EZqb5GH6N/wqovYosX/QCbL3R3j3TB1WAYbWBmmsJeIH9t
+OVKjoJLiPGHAn93vNcc4mua/BTvUyHeHl8jR9yLdZUHhTkheKlai8l9vOE6P0kM
3UnvKhQjPv1p1jAeA5aBatnZI5ovo5FRixb+sV8wllr5YFsOWXgmrJotEXsL8Mrg
PUsh6lqhZlbL0z9kTHhQ89mufQc5YGLeZh7pAzDcmKajhuq1l84a+nSyTBARBcB6
FWHxfEI6NO4zx3p6AJ0Z4y/Akq1anXvaa86w7G04ZN8RHqCvPIkH6yVMb6t7oZK7
CyPSvPxvVFzYYKbZYGleafOTIZZAePA95ivb9ocWfmB4tDApeKVl3XF8bvyPJt7w
9ClPCxKxGMVlh3iLZ0CLC6kr+pzwoWXMz9C6Rtjjj+ifkYvmeQxly0Znr5ggwzxw
6MWcL51ymQrHSYnBK6esraKu4iHIqjtfK++zaXXZa9ARoFvXqH3oA4o4ALHWonOZ
dnCJuajVKlhFuslYG5qUQy83V7mnI3j511V7vomBDh7oYqO3KMf/aZviql16+Ina
k4Nb7KXbnGAT1Vl3CeFKEY/PHx8cYXD6bSeFbV1s6znczVonYTapcAbRR7IN47XQ
tL8QXQ4gg4tI7Y1VZtGVrqzwQkMj3HK057dnSEv+pQh55v+l1dQE8mF3uyuPwXQh
zbNtfdiHkH6+8yvsM+TZQjLAi49DgGvbK8KY9C4qKmmaq2cNtdxtg+2gI8YCFm6g
Py/5H6InYciaazpd13q0m+SqmdZr3Uv01Y3K+xdI5UvPtrpejp+doJARGClr37iA
ZOJilODe3IyOUFgEO2KkM1a7hOZMhd3MKuci1W68XaJsZrwvAsn7ajpYlyNB/jqx
9YmRfvLnJqYiM60zETJRt6k5NQQqSY4kk4S7o6cY3q64Ld5qqp9d2IyZUOB4QqIa
1mxf6exhYyK3GlZ5LvKL2TOCmLi8tdYApYj4zJZsmcSISTMCs1XnbjNvqAZuolZW
qlSTWHNscKgaZQWeTnUgVcmq/teXyB+0hL7dJrDdcuIww7qk98TdeUsew8iGujoa
RtAvnPptRWC7rHbV4+BDEsk3eTGoNLbahmEvb+NgDOiX6LiEulassA5GHWJI13p6
LxqtK/to3VKeDCEq5m+z1PIx7220x2OAL3Cd6f7Uz1gpziQRNeqOZk+3zgBg+t20
s6fkL/RYGKJ/QPlSbasF0tWUGoUhsAHBKKQuAUsGLXRQPTPNEl2olB/CRAE50yjf
/v9vSE2eS6v1njWpdzv/FN/AJfbVqsZo4NMhX0/AR1za4fXfvIgMiHub+o5+rGNQ
aVPBfqGkxXuru0x4ruIOaWqFQt9E7MDeDqYoIabVbtyT/07Yykled+VpHGwrNuj1
BTC7a/2k4OyvyLGbuSz2dyxlpTIjqiNUHCSbOKpsB73Y7dKBDjyfWi9E1vcllLhi
ufX9Od3WvY1GI4QUfp3+bNrDAZInJGm8/O/wID/VmPznQ9p6tRtA/PHDk7QLIIjp
xIPKhC6KIaqb99aijnqkdeRMEya2PKTF262+52xSj0ITBs4xgePqRzmw3ycqmaIX
Z89BGObCb9bI5pA7/H8EGYjMNn3T8yN/dTmYCEqhnWMRrz28mzNe57Xg9SB9rgRt
VvdXiI7e8Ou9taYe+F8mSEP858AcvYWWZYCPaXmG3EUDxqLPis7bfDy001Uhppdp
2Y37qfNCf9fVEIKhVxbRIqdO61ZO/s6B/DF9JxQjShLvW4LAXEWj/OfnW9VEyD2/
xgRe/IPV5zXvx3LqCHUQcq7tjXYjQMVggQLmLfmduMwYRplpNkN3OHDJSXq8v6AQ
zKGinOseTyEKbVOA6WIrap/nU+PO0FwuAWjklji3WD32rW13SAUqs3LRFTRmj63o
SGARh6B64g4rVrKpq5xkUsd7VRmjj0SVOWtvsRj5pq3sKkAM0PoMP5HBeOvF9fHz
xVXZP3rOQrCMhV6uQ/8EepD93kd8zjAI5EsG2WWrRc4GVu7vyH2y6vNLOIw/1rwg
Vg+olSp5mzIPWJbkMzJtHD6+pUwB4oKo8lgIoeDTXE9pz8VqQhcTr/ibBKGDb5bn
u1sjw4PYQEMOOwNsKKFs+MCJudeNpw9K0o0OAFDl3ed0+TdWrYv7fRskh2Bed3xH
uPASgGO2S74xIKFXjFtNTWdgP/LukSs9BYMqLZu8hMKPpOQ02QfVBLfXDcJOpetv
67QRjfTIg/A7SAqBDompip2g1E4CxunPVYz3IH/HziMChvKQrlDv4TcIroPvbPlJ
FYicGydSYpp3+rQznNnsWtNlHcCLd/N1IvE2y1omqXEnV6RFHroyFSGKWfYmBNzo
G8Qf87pBNK7JprooljycqutAVOKVRKCpflbJUM89kia7Y7RT5/cxQ3sZM6iupSm0
ld98kfQMEDKfwjbB23dhRgo/cXEc/VjOr+tYPKaTGOQmGhQikR8j6pcq7To0dBj6
wdFlbIBU3QOa01YnCchim9AWQb9P5PM6CH9E+f7ZFt0YO5Ijxaovt8fFXGkDL2Ok
JZ4nvomBus66wRbSOHLBD3oakeHcs/KoucwyAUnA+7Gi76da/obGf6oHrC/Ko7iS
+tL9AYDk3TQ9cTW3iv/DzTFGfWxKz2ojewaq3WW0LTvxQodN8UlCMSCadsAWFmSS
yAtvx2FZk3hbqolSxlfwcRrmKv19a4RoQuE526fyv4KaQgO3L/jRCTh0QmC5KJJB
I6/EbqVkSzuxRQ+nxLkpKV7FQ864I0osskKyujfHrGgEMOOUWW243UtuVMLQnzCF
ZsDgEdMFfiME/5yTuEVBAcr0i6ITRhpHHPSy35C6uxl3OMy6VVFi4X8edSbTya/C
an21HQAdempky5dgLdTjLqNzWe2AnSijAkwXYt+LEdaTk67yUGZ001P8ElUtudH4
AMGXfwGZ6p40C8T345drQkraaMLaiuB0jIQ6bcuDpYmwx0PNyI8J+Ji+D2cuMGjr
8vEwauOdREAO0yZSnKLhk4OtRKYmxIPeS0NYSyFBpsHxoFFsJisQNskfULWubTHK
SE3X/9SY2fAViKKzAibbqg1OK3IwLxZbnpqQt5O1Bdi4TvlCSsBqaUVzxY/AFJWx
p3BalMe5d8ZANm1Kc78jPMTOsjTpqGjTOR8Vv+mEr/O+OPeJadI7323IsY5nk+2q
TnJUxZ4GO7MmGyhiFLDYo+QsyaZo6uTrQ5rltZhRohhlXkXK1v1ph/XlPuu3U4GI
oo7PqHKdooNGqAx/nvifzclRYmFzuebkbsbUSkELBbMM7i6efbr/7f/FUivUs7Yi
LJdoepJ96IyTnmJ1BaSttJa4nfhH0X/MwBdjYv1qHFn6D1iP8axta56bG4W8e09e
iU4urrrQPfTMEodVLQfMSuUtIsbcQ/ptXMveP04bjU6HsyAlrWx7PRDZEX+NxsgJ
rdPfGVQaRU/dHSiCJMZjgP2/JhAb6AJSNO/mray1DAt+2ouFjc2ClScAnKQpsaax
4eiTm9qlVydSt0BBDVmdD2G9hSdIltQmyTmGoUkwTeIpJnKl9h9HGzZ/wWzio2Kh
xLU7w6WNlxm6kzsC/VRvc1+FT5tF8nAEwozV96BBFYLsMGosGRbyuRl6ZDu2vdUe
yHu1P0p6nfkpq1SeqRDLcsNomZXSTtPjQ07QEWbZUKiBttWx0VW7oPciMjIc9zSM
XHqtUXeZVt9D+FxM82wi/9EBpxc//FwmZLkOMimNA4/boqBsugdaFfuMahPW/ibU
OuKWF3jeE6x48AFcFTaPD0oF/fOqSgh0241F4DpQ6gZAyBi1W6PXmnLsf6jKrR7S
gXU16G5kOkHiHfHdpQjC8PySoyr0urh7lfgjU1guPEL85MTziwko5tZL0IuEksay
Vpphc9h6j6rARxs6HYz/eoP7D9jWCjRfeGoBvhK1DIo1q6Q91ZKEj1zHWEsh5hWf
GnvO20QCSIlMc88QquUIyUIY2NK8RLRoO/KO5/6sklG2OIZstqqKwNVB7lno//hX
XJLD16YZe7S7d8Ol/AtC+6G74OEaRjz4iwwXlaqLS1pO81AOV1oEqihNUY9hSVXP
0leN25eul65B0Uqfr12gbr5oCYPwr91/rOPRJwcGugHmKpO6pLTHaAHSNMIbZXJM
8ddwhLpBxKjeo5iX7jfDeZShodE0wTARyL8YHEu6r3LWiayEon8Xxhrb4u4mdIGZ
Lez8tVCyYYCkvFGqmkmLySeM4zErPhq083gGwoLBrXxxyyP+76AG2PUM8e4EDGBq
EeYHxCKCQGPexwBbJ90YON0G90RXulIwlv1aC2F3EEK/otXbinJifqWtQ01eOI2N
xiAs2pBzY93DFXw8stw0WsmzrRvAyWhD1ixdzsMvaVKKQVgeR0+zFfN1VX5sVY+X
rDX2FTXLXkBvceyCOpzQJdf3SsuIbnerTW5ORvmN/44TB2rZm9D9HHYKKtfPshL3
zo/vzmQWPLsrg1oOn25vKjbYCxDNB5hltJRT5uE4eqay3p32jHYk0EP9zW7NmSrp
SBis3zbz06xlGBUriAq4+amQec2FocMIGvaqrS9+9dR8wiGI3kB8m+SXTylZ8UpV
OFqYZ7aaJP/ungw0mnxp0nXA7qrImg43jWmwWH/QhO4SWILivNBqlzToPeffBzro
AS5BO/nFrxLKULmV9WqkaB+UGflerLjQsdbiHZPQO6SHvrJg0EER6NE5bimcgxhk
eqD6dt6eZicuVWM7R2Pkoz3NipIyzVNxSuQHm4cp2IUEkOEJFA1Sdp7TYdLcdIkc
q6g5d1Z62luw0W7FvVW//EkCK4sbYpDC3MDTZ7xSilc94SQ+bmTqfdPs2n611hR6
zh7BlCPKJAfujjJgyXuRTSGDC4blP+TufaASX+jJMywQ7tickk+BAsRocPVQst9L
QyZC/Ng//WZ9FJKI268kKRo9rvyA3YjaTwIVaS7cZu2XybysMrqlM0PvyFbGtjc9
MzHTt1jUCFAob6cnSY/i/0tO1RMsfUhE/w+mo48l6VwW/82NDKkdHHu52PHZRGcY
SGg5lVEl+NFP5q+6BrFRp7CJm8PtRU1I5s6gRwhU9E7EDIg8pu6NyMHfyCGa5bd6
abcDcO9JNX0pufDfSVKi89Uhz399aREjJLuNw2d6b5nx7BC6w59Yv9/CqyGn2u+y
H60Es6hRKG6E3E+xvq6OBzCVo03w2R8bZGxq/h79t/JGqRIAAIPOj5FUYnTQVoSc
Vd/aIn/8AKYyMDc0XDa+9Jd71jQBUUqvEsMu9Dnukm6bGxIVIft1oS96RZS4nHbA
xekgUZhw1TaFJ5NrZlQZKbofpEdUqywMID72aUKAeVr+KNKj7yDlaWp8w3wykpb1
cLVWhLhaLMpT7kUowa1mi1M9Jz4TbbZCnZT2T7H2SS6NDNfFvjxMyCWq6GVNS+EW
vvfm4jhr9YOTwgT3taWlcX0iV9dHAjMXka+nr3nv33YXHe8WeVOzLqlPKmBr1uMB
KywRB9+TuVJgOzhB3cNtnCT4O8u6rCGLKsiraexPyWRiwWFlByVMngT6titeNxZ0
vl7OC8pSC1pCgS0gAeZLwQClX9H21psJoeiGsi2icH8aLYPVYQl3XtseD/WZbVwx
aV9ge1rmfcKYodzY/PN2yRm3nwF24q7Ae7kJbDY/0xDtygKydPue8wIxbKZjts14
knbEgbnQiODVTNFz4EsgGEsxGBK3CdUsggb8l3GOEM65tRokk474l7zZBQMUbX+A
uQi8l5RUN/HKJYmcFbndQHj8urQry15cTDmppyUCrqsIQCjBrE1D2L8/wdjMUOiK
n5CHjs25j2JzZW90Hn7IDPaqLQM50tfKfgY9nzKgcBuArlnkQ1Ifh7wAZj7J0pEO
iLfAXt2TdDFHpQhNLeZFAr0llUAoDu8hmi/QCwYbHL4fD/2Coh32j1MSG2p39QVQ
dFXnpqyP4FATPzOob4tlh2owZBNwk4yWQjzCbn1q/0Y89fzMwEC7MB3KKs+5cfUs
igRw3wH1kcS3DZBWzGFibLgMa1rKHoEzXTZt1NRpsCrabI7j4qi6YWY/oz7QS8WR
0UO1BxfvqoO3HRJHXziWbl6w6HvjdGYSZAWfMBsaFsFRvi+ETnZAT1cPDDni9dja
eedf8TMZZJvQje3A+untJgU88FbOF4W7Hk2VyQOKtHndtIJKOTwnI/eMq1qUQEOO
UdoPcjjfS1bqnwADG5Voiy3ttuO8Kkp7zrjTjFtFmW052A1WQB/riI71F/Ie18Lm
81HUCF2RsvvM+z1Ghxkdr2Zo0UWGLy1u8vLLuAstfOClDDC48QwPAyq3e0D8ciii
ZODCf3R8QgvkPro8rzaI/ZQl3ViCRLzSLnr1jLocsXccvs1e24i0LDhUyOieuDZ3
byS5u0nU4xkpvyi3IaLAXQrMbQtUpWvwHMM0WzShpoGluI1SrU7vEN8uZTF1zVOK
M5pjBYstYSC3Pyd86MPJd9zUXnhjDo/D/EO4IlNy4ran6+NWN1fYXyX+oz5EJARR
EPUbE+Yjlv2wAMaF6dU5nx7C1g9/S0fkVTNpA6UaBcZgDfGemvdNgqBSmM3P0BV+
qrM3xVUQ9z+wdyEowe7vBzwIHJ4idYYVdNzZAPco8ViETY9TeyEUfpqCyaHgy09x
FgUIuLeF8+D3fqe6D85qTZceGovANwHPPgQ2lPRHYcFXqUG8IHn3JUVtMSGN+9Pb
7bMVYNxnAnSN3c0Ct3GUxvGBVgmRemyHF2iK1rlqWtAm8p41s4gVaGjWiotOvdvI
0pZRK1iZA4Xy1jEbi5CTizJTKNN0Mwbqd9t25TpoHvnHo5vu0/zglHrLLEvlsAPs
aco2diOn8tdBJYL+g4yQVJnzcuZLFNwR+SBU+hdmXBU6F9UJB86lSdY0Hk6xvCiD
S71e0FxFzXr7GlfvDAKyVEUUMrxWW/kzRrAGZ0IgOq/Ia51OLnlvLMCPwrBVRBW2
0MsOXDNHn7RtLTZHWMzLQ6aKIQLnbrKjoJVqXfj1W+HJT4zUoXWMejtBdyIQLbGn
OcbRjgGBVRjzJF7/87V4Nh+/iW3P/PLCex0KjY3NCIH4lwfvPYE5eAwtkThNnW55
bouVx+G2zXwOXsiZrfrsOx1Zs4Gp6B62an5HkzrVx4skUAeWRH0S+XJH0YUObaxa
DuLMz3m7U5k/78oQi9elwqZCaJFupkgNugAh0Y02MunZpCF53e7VwwhBWZzLE7p4
IrYrP5ZqMpWT5k/3t5rRdpZf6ythtHQVt/+CwmnJhWdcuZWZjhry9PfiR8qfo6qR
ApWmpEYmgS7BVcKgOndPTnfFavvfgnTaFPXKjKnXs+cYk8z6+9qBYWPG/5Q//mRf
T1d/gmpzTb+6isE+40IGhOVQtZtfgCpZgovoojCFaLgkjIRn/3lvgQi1hodECUk9
gfh6fNoBzkYkNoUZ4QiJ/EQM8TOKPLqsodQIgSkclEZS/D8Zz2XWBD9kABCjc+Bv
z14LuI6jJ34F9IjzT0Gos/FB8+Frz5ZWlYYVoznXRa7ykBOF8Oeh9KiYNhU49K3c
GyuabW5jKsQ62Vkh67pkxzDH1abYEmMl8FstKIhoOA4SICw1mG2F3h1VAkit9JKI
On6M9r+LN3FLCidk759UfJmsvw0HgpRlOdGtZXOuwQOIY+KxPQbF3lwvtciXbGrb
r6nlEIPIvlnrPaXYWfrV8hQYunVJRkwk7JMe/e7596fC8b6CIQO9DQ9JwS6uMOlM
JK79jMBcVo1orn+pS7E0X2AukIlHeftGPB8q9iWXazdJVaBun+ylPYE2duU+KKKS
jFZhuGkAubmfuPV4a2p8iqvT2KRim1qE4sJTp4MNuqHnzWZmQkQ9N0khOOHiao6E
TtsB4eT2QHH0dEojGCYxZ4qFl4YNhpTjuB2O5cT8/eq21xqjHABPcFNqPcIKh4+T
+qZyqBtWReFuCsBeV46mZ+Xzz3pB8qg/oQQonqUQr2/SQejwLwq8iL7AR8JxemKg
WT1txvFrYK1xWpIXL+E3pTRXvSftN9RXvm13fWDDBh8/antBfzkjvR7XlB/aqqWz
AnOb06ZfhaQtPefbRgezTq4oLDgVebGuP65+0cTgGMLVK/QjLIlrt6ZERVWuxTjR
FHVcOooU51xcO4wvI/AgoOEWB85+o0PXVR1p1kvFHGCtiKgURhZzxryT/MCAuKXm
Ntq0+O7Ibv9FK5odmx4rjY8e5TfKIjQXdGuLOxMKmSZCasM0/CwzW/U+FbjvX6u9
N/Ia/fEQnTlNoKNL2Lw0h/s/pJKCVgGY4Y6KPAJK25sthkTqR5qgwm5CFCu/5V/L
BI2cbR0uzskYIT9njNqvJDHkhCmR8Yae25M337HwVvhYCcMtGthKZ1yQ3R8iGM3M
TFESsUrekSZMGLhFyLHFLpGgNsinLmm7VF2pqZu0JqxN8Pt10AQRYMsD8FoGIuv0
F0pd2VeCEDQEzveprWpWXsi0ndy632EjAUW2nXyI0LJqaJMXJzavT7kqYxJ58hyR
kw9zsPNVn0sdXDEuQB/XRKVCOboiexsOMOW1yG74yR3oR4zQOjDPBOSZPEx0dSB/
ursOHb8yuvUsWYvNcE6T5kqyb7P14ZeFUOgEmU4nJNIwRkhmmhkiKQPoyllQXkMo
4jgLkF4ZeASvyR8eCj3t5V6p+M+xHlfIZdPiC/c1085K/shhOkbTKc/0F4c9cAqJ
fQFC/z3HeelyxKhJtnfPkbdIyU/elUcsHkkPoApQb+4by4w9Q2ZkrGWlZGOzstZf
95OnriWT+nBybnrdVbZdRBiQWkEn0UzbfvkAqVvRIJMY+JTGhM53qTi94E4eKsRS
BhDlYZU6PsgTJbFkArOhf+xjQp6solJi79GsLkCOo6n5VCOjt8V96DNoPjjaOGrs
RcT4952mMqt4QGsYHbJeqqQgfPKViOdtPN2SANOdA0kGycdsH0LJMBAL70ZfD+ZZ
Xm0xwYyjWFitBymJkdkPckYdPTZ7c1zIx0fnHYShhk8AtoD/+SBJ3CWuNwjEBRv2
KxygaUN2jCYx5qtcpvxehRsIt6I4wx3DJG4tCGcKc8jtWU1siPYAKJzLXkiYmUdB
/c/qQ7QjN1//oEg9u+tiddrm7pMfF1P9yCr2waSyVsMfA7F5yt3XflCxmgcgvhop
loHpni2lVnbP+GLtF+FYw8QTfFy36ENDl69pxNEOG3az4Zsrym0gnOF3W0l+in0g
RhMZtFyL4O7SJck6kejpRjPXPg7hTyBwYn55gTguUDereat2EYWFMn8lubYUc1qL
dYlHrsEn1+N8dcGHw2FKyhvNAdM3pA2WkmU3vlDXnjaAmDCeKjhT1dc3LvYs2fpw
wKwm03VASvayjzvWmYIcXAB0FjgjB8cbAEQlLVh9x/tHg9ofFLzD7b1isehddAdZ
KWkdS6dJjAzEW2FQozprspbiu5TKDgtb2i35P86PrAGbooQcLlwnQTCzl+yEoD20
4nYhcs/N0E5pGnP2lr9kp8hEiUeKh3AYAfcOtrmXAgVhtnoXRJid5gtD+zBfSIOk
j0J4PcWm4CCFRj7HuwGZP0/KbpYUHMwWvY4vKAy9P2o/5bEjjlr5X6WqPI+5aP6k
UM48ZnNSREPAA3qkgpTyHGsxF+VRlDmZ64z+0XXVpGFym3lm4ji/QOTrcOQ9Uwli
be4gNVfY7B8rj31Luz01CLn6/cQahOtTXihhuxfOeLWJ+SG7l0euVM4SUcaZ/IM/
gPXD5W71sStX3P5J+fVbEm4phrjseN/ngriM47cjvA4n3yDEwaRs3ypbUjkRute8
U2xajNjdQOMDU3uKsKQNJKPI4M2YanWmfb6GzvNme35NeeHnZ5quTClU5gUFVO3k
qZBUAH58gw4GyqWgKd+INZviSPTYu9ra42gZWYsKWKWJmAcsFgWY4S/MOa8tCjpS
68tQJfqgrJbB8F5RtvHOEuaeSp1e8K6c2rmUGN7dqJnwkooRu5QmVct1/j9Wym28
aw8kE8QZBKmPaFcLsyBaXpJHOVaEn1J1j286rm+pNd3j4Kpx135AK6GWDFBuDBdR
PYXpsVPktqOrIic8Ls4HrvWfptDGytPYZ6Oful1ex5vfJhuLs5ZPsz2BZ+qiBjm3
8RJRq8uxfvLTCm3xhuDB3+4xbiQhENw7Ew0a+qe7yz7VDPCkle5H+Uc0/X8vRYqP
Yabv7U33q01Im+gnLTi9v1Rp+t5sOiy/lmjS6DuH4rGWxAiU0ZKQpt47ovxQ2GYz
9cYDwJNrsraO99zVvpuiJr20ALS6FTF7bjvDy0HMaKKBmSHk0TPmD+WtwAiodRun
hPGsckmvrp26OmjyEsSZtoGTJLbJt4dJVbjviPtpVG1FO4LThLVRz9XrXT5VUDsL
kzvjAPm1b7QW/w8Pd+nLc6+ACsxT579v+UvWskRhX+ZL5jdDshGhhkmfbq4YHxsy
VJxF9C8PZqlNRslIc/7VfUfkkwpgsPw5kwwoMuTUoTXPiSpUr4KQkj795DK3Dr5D
FPbsEELi5nvEWFK7bbLqKsphPOJKZ18dCDZJgwB0Qpo0zruU0rd2I7QYqsp+Cppd
RzYK1pFqy6J+WDrL+Gadat6JJQXXHv/xTe7RwSL0PHmlYmYqPhV4Sg0MRRIyAV7o
v63+/tKPLino1rFksGfVriZhj/G/Kn+XtKOB1lIhqjbeYQ6NwaNkxBtx51blG9sq
5uBq4leVBctbtwSF6SJS0bq1uYMzub+duuAKlyz4vORQLHfBd0+5Xis5i8k928l/
faV2ShUS/pqFCG7bWPp/Y+jTb2JIPe5cDcRo8Dh2/vICdMX9k+myBDWQRK0OyNZ0
0fUeyV4uOOe+M4sRRY341IdOUB+bI6gQUxzJCI+fIr4XDGTnfnlPcg7scdv7cjXc
c3JzvD8bNPt8YvzZLOVP5rA881tPGjN9OCNIBzjZ6kpt9EfBkS9JvPjmX0c7rQWO
OfYwaP7BJYbj9WMtGGqtxOBZFId3QkFIoFYeHICuInRU8qZXe7fIuwRt6QS9cB8+
F6MABuaKYXbd/Y9LGMNyZXs1Lm+FIVlK+bRuWqOCEJI2JtUeTmg/ysyXNndG3Cqi
PuJG7FaCocBRYGh4K4FDXIzzse1tS7gcDlPP3ImGWamef47dC9KLzya/T22kNXkO
5PNpYj/hjXa8+25JjbEH+Syf92cgS7anBsQ28axhY11DYhHgMmVqd2mMUpuqNfz8
994m2oy0cR0T3OBzvpRxMH6hCt5wf/APmgSVEVmn0umHJkSyyXZrQMTDGa0SSMUs
Fn5XKxf4mTcFX3WeibKO9rS5DMG1S6PKyQcvoaCRz+pMGE2MwHnldcIHSDbTFSem
lahUhaOJ9BJwMMqGiYVDwLngayX87TfPztUqHkzfuwoHcQ3twrKiAYxu3ewlxvzV
93F8jDS8iKaX5sn3/h1H9BUphOctyh9QrkSlpP2EX/wX3YntKjeGXhj5tb2I4TTE
77DkXZgFOQjsiRHtztIzmYepWBCEDZ+QW+ldE2r1Nba8uV/1tTd1ipNhvVzu8muw
EGC7fZ6QlSKDKzlFrXi7VAEfvKuuanac7eqqZMnRp9nngDH7pLP9olMtU2qRXhpk
Gh6byMyoiFi6oteKqGQWMaI+mWWCtRVb50MovUFVR0KnZ8Q9fysjXzTffihauqlD
HVo/6I3pWUXXwywa2CJZLTbmNX0d7VLyB8fDsb8jn08EYhFaAQbh+CzUY9c9G+Ny
xW65LMd87gC8uQXLuHUAu/RWR4XPTYBHEqVEYLAKp33Zcy5b9mGchPyqD7sJGYgx
omucvhqgKdpEzjiVBsHo2X2yadfpz7inxpEFM8mqfTTY+syVMm1O3KTTqDEX8sqg
aI5KXHK2dKH3fVlb2xk8CxkivRLT8apuZ4dnn7NcMPWJJtvrjSyhjUNPyJNXV4J3
aDhZz4zFj0fQjQQfZgee60anhf9l1JCd93StmfXkyS7Bx+j5cQWiJGyLC9VkL+Dr
DrwQ8Ojxhr0NQfSu9OjrBHENwm70yTHz7tqKkTIHfmukB69aYCJTOJ5D6dIorzpd
rQJOSOH3T9jSZtw+waFIj6D0WZSyDu5NMFb45lRJjZj7qVFg4K1KTi1IufEBp175
1nfoazYKqGu6+NVUEcpinUTS9kp1F1lceQIUKNmUsEOTTz8oHx6jrfrnKK1Gc3nK
dgX+NdPd5FuHCLMUyWmPVegU3nUlvYzPkG7QGBEx4ME9FrCzt9ACf7OQEGRrCEQk
q1ECdhF7ZaD8il02956RWaAqjD5hyNf4dxz6RJEzJNQBOz3tg0J+s9LR5ddszo5o
oYoKCzzx0Gn0QdE9/1L5D9cPVAEPcLSFJibhjo8GHM6l1P2LKVccVgqwU3t5i4an
bjm6Zoqy/Kki2O9Hi2FBVIJo/4TtHnUh+lpLDperI8jTumji7XcUdjhPDFEAMAmH
JS73PNmGRAOhwO/+tophCl7iwKTD/FpRqkeKnYMUHE9LyUoOtBnIvg+lLJ5hyhR4
Nr81veCc3LDFdZfJ5eM1+C0IPYRHJR0JZkmPUwAiysJ4Sl8hR/lcS81UeMobQyLg
i7QX3YHZKcY/lcg6thGRmralB5Ep6ac8pn5X6Ldl/4cJ0i2xa13Ul6h7LfakpZ5p
BNAz/Wb66FXafkfsMbNMk/Nd2w78iHyYzjuEhYkGelrRXadiQtD+Cbalo16ROcF2
I7+6n5loOh9PdtYnaydyx6JC5iBIDdoLyfWBzbtZ95AjhaYWKSQqHl8yH1dN9i66
rPnDIZZ6nY4et+zpaFb7NjLCbDtm40RUX6O/oD5SvDSHtOkNoTO+D3CtM+ENtE0x
v/trWi29gIJUkX4W82scmQGqGit+BjrSAUDbaIspKo6Z1l8Jb9UlzBWAkpkwf6Li
B7R97tDTznf0iIyHdbdfEF9yAHSvEIItcNuufzCIKKHMUqhgUuruQmxlxcNvV3C8
GuMF4/282ilZonqQk27p870y8Gqg57oxheJrjekChUkhCtOAwPlquBFhd12//oqP
LQX3p663+729FDcvxzHnnD4f0Umrhlk75S2EfITSxpYUXzS4QBKXEBZVnlMSYANd
vA2uCvO5lwIA9TQo47dWUwmB7v013XozMLmNJp3dGGbmG3IgGhLa0DVPV99WIsDb
eImUljIA9JG4IG7MdbhJdArPIUHIGs41Ja6XMg8ehTsBfKO2JpZeg0joU2005wVl
U18IwukXS7UOKy137FqfYfxUv9qwb210031RMVk5yVNX1c1QKKgP9CCxdfIp5KuK
xK06UKgKXyOEpUdx2s4RMDijb7l5cf3ka7uK4ljONXZpT2/q6ktAR+KmQAOWPbyn
XtORhd1Fyip+/OZ5axgYVoU8PBzGytS7Bs9gsH67PnivwSe3V786TS5T2JvxYtgm
gnmOE6IQaRorXqQ7kg4lioK7ci6AELcbRnIDhCw6ct1qtx7wjsw4VLuSdRuRy+qD
LF7vqO9Tt2Qf5/3NsaxdiH2g7RvjL+GLdKRJb82Ytf1R21KaPTiy8k/5VBAWC31A
cSXhulskHwESBRQs9a7KU9sAIXO4xCP5GOwXD6uGS4U5MUNM4oV8JqwbRlGd3PpZ
0q12KOtYZushhGLLtTu04HCFiTESni4+F7bW10Pp+7Eys8xaoVHG+LtdKr2SGqGQ
7Z5Aa/YDgxYFrzjc/6cw235ZCiqWf8dHQrDZ05xps3VzHX/kfJ0B1uOtS1wR7pkj
EMQdfunKYQHBL0DroNLz84+pAiFZUx/fhJIK5dS4ToRBoV1Q0hD4PDSU97+S/3DP
REzagwuyjrNuixJLTeCIkUfKVLPX1rQRBcFDfFQgQR0kE+S87FcebuUwtadv+q4m
mkin5lpa1+qyS84HKADlrP5idOvzoXforyZIvnFggKknL1mbKQysuYVBP79mAnOD
vAveMSkWiiOHeo/QKb9l3q+9/ITttbdBfvKr+WKsrv3jwEgH5bOAD+GsD4fPqaH7
jxBhnZAGFU77lUJezwJLVxLJIzETsQadt370e9/HFM4hEASekiMVE5gp4dXRHLZS
5vI8phCX0RX+Ev3a3H6oRD+5y1hrZll/5ze7XckWI3Bwh4cWjOi42GaJ0z5XWkQT
juBDmyr9htOpVusMUg1yd5YaxMxg/IIGUnOb/Od01bg1bqfUeBeBbRTyLxjmAH8P
n3O8+lejUV0PKaC4Q5zIMiQy5NAXBqvDqv2ecqz4vpChuEGegzIDeOyZZPmt4MfZ
9aeBAAAOfwCn3dylsC5+QMNR9kF8MqmwhfT9xk4Ivrj4QI+C1dJXDgpypdrlpNPf
4ouKP90DxBcoqmrmcRtho5VA27kfaJA8ddixh7cZOdz0qPh1jpJ91XeBC4Ola7F/
bBqO1hz4ZbvPUy7+n+2XvqqME3HzHCfaIbP9p4VcWENnKrXkFuH7g7QlaB8J4Tzk
DYHF2TiFxZEYncNlRkfwZCNC9c6JY3gr5fmomrNW8F+yaJ0xnZ6n357MzgNzedbj
+Xxk9ttELEkdZgAj6Ha3tHQgzFXddJuE4JbxsCcRepzaMQ4zAlvkvBBORDGcjvPP
aPjxv5dP4cepIWzbDROeI5cbmEYkWwkbLFBC/n0GeAiOa5IcWW1ZQTgGtyvH1FV+
uGuKOjVtRTfxJu2Xa4as7ZALoMcwk+ISQyesifjLrQfvSomSWW1BxyNERwUdI3yH
SgE0OKscEllCO3HOha3wdaLr+hXpEnKxtf30yjyu/ztFrnuhcRJuExnIj/Pu11Mr
oPnfhBYlyDEbxWrpQDh0lITQApU3o8QChwxbXwcUXl4J6DJf1FVeBcD7LHNXnckw
6o19K6CilWhUyUUj6YpJzdDUBhk7WtyIbu7GqQPU69BZg1IVHjDqkt/AxfwMcBOx
p7Ai8loXD5J/j7LwkHC4HuGWghG3qGF1Y2f6eLc2CqzJGGfavbJ3OlIpWcR4lit5
7Bczm60DZy4cQhPo2+pr+3CcnEG5gsWjYEvOCe3YfZ6p0tNS4CfQ+I5fwv1wgxh9
GTqbhjBIx1Bp+q5xuivEGjj0prdnMsHpGiR9RECU9S3baXCwM7y98iirtDjcSBK9
g74BMJAVoK+DQ8oxg2+oTvX+Nc8RHm0UEuBdvs7XDHHDwS037MlKEBjZ4hCv4rKf
FE8q3/R0JyIY8ZUIMiyVL/ztK/47+0izjdZnkzPfIDENCiT8A15CYfW/1lgt8KJw
BY6rE0934BCwAiW4zpcUmDcG9mpWj80wMDLVMkCjZU5vogcucfNvuHlxtM+zxUXe
hvklO4xwZg88gXyzkgBkM9WnPMbM3jN2qdadzpGAAwypKv/x0xjlAsMTzjidWfiX
5/akGPoxmkgwn0+2wqBj2HBBjju8lpcHU0hWdDF+RKwDn92BksbM4ZQwOJ1BK8GD
kkUCW/iPy1bWbcpEToSW3ANzU+fopQ3xdfajiTNYUE3tKChOES7J+osHBSVU/MqO
FkApdS/BumsvI5Tmo0wwOgWWv12T/eGn3puQGIuzzr4SSdloSLZjuBWc3jkhb74m
hFzntWiULOMSOblczd/LMBuVQX9AtPWTaY4z2EcUTt8LGG92wPppAEeF/K+2npT4
Ka9jFBUkXqixNLAdTg6+/xDR35ffOq/bV319uMEPCuEh2MfwdjrlIGk2mJHKUNZS
4MKKl4BOMDrxmHtEmduwJjvgBixb5P9/9Wb3tNP1SvEjHRnLCMWwtRsVGjlhslul
HeMVMY82PfwMvpwBmcZZ0+imKIuxaZqCHvhsQwMMkbvCbGpDyBz7rjVB+6PBys45
FK3NwW4/NleOeB70dXOXx0VnDMnrXxRTBpEZTQ9yZudX5rK3B5Ju+awDE7mwAfEH
Vn2XtsTjIBo4CO+n5DeFqJkJ+loBukkw+Rbb9zRZ+KCD/NRWht0pxITaeC6Dbv08
axEWbTOOAna3qEHC2vxmUp5CymWQXL7nHrJdBb3N7snRznEXnEfMllwUa5ysaEmm
toLXuuyYB4ue/gewzhiBLwgJFNaJjP876/M4P6/mjOLJKkPFiHYcR6jl6pxOMboB
rBccTMnRx6fvRAP9li0XZgSHvkpIg9iEiY6IF+mV4FWey+jpY3X2U4jK+pcqn02W
aEYkfJJobGtYdkGl+57IBju+MMRtj1JHBpC6UHVD6zaD/NGoeqTw+qzZDVdD0suT
yF8LihRjlSDVf+olKLg/zzjTN+tFgwNw/NrDFKOMyvqmkZJGXMKEci6iIHiR8Y1A
DKtUtgfCivciJiJXSin/gDvsP3jHUSlNf+9teQWfobUlqfcZvuqWnofhVbxAwjU8
qUNWEN+etTf6ZMhM0Ut3ehRo/zFXKLH5M/8knF63XstBm9K0RGaKZuHpFcdHCaZ1
umrLE558pZ54vQ63uoAcrOZ8F86ykjUy1yyNDFxutKCRAVWyBqeG+C+9B0mvuZ5y
ePKItU7+zehE+sp+W4M6QEOb8/85yF1y0xv6Oy0ANyyZptRM/bnq66f93CnhREg8
SoMUEXYzWLUKIUb6Mw++UJVTQ6SvSiWLE6FXuQ+4KieykgkvuNKfN5aZN2v6h8TI
S9FYIX1yOQqoqS13woYQ90MD8YzAwfO+ObZEqxlUpbKzvyoQRKbEa7sZwHJgPSfs
2BY+l1l8q7+iMxq8v8nneOxrjlniGS25PNh9ZBAEg+WMzkympDkjX/TmSPvUdndO
oKkhBuAUJVyXkb6D2N1pVFCm2lmbH2StxpB8ASfowI3SwEq027HwiTweO6GJeRWw
56a9VWPP0hgZThsVvgBOPz0vcp57Yfv+pmi71ug5w0ovT8pQeWeN6aoojSmfZF8p
s34sEVVOahrKRRwnuY0I0J0qUWgicJFEKzBeIZNu/UVji4uBxln4kxwFFOw50dmb
MWIzyhwabhJzEuVNppRyhTY8JT/PBL8AA6rzZ8ocAVqf4Lb3qn8wWT7iNh9a3yRz
MENsGepN18QRZqn/VN3C/YMbChWo9W1aG+gm5GoYGfl4o3L8RQKCdeeLqg9zDQiG
+zm4WwNVfZFHEjJQzPODJhXYH4pTp2QMEy/BzIcbyR6ZlmUng7Dw7gUMtdYpX4Rg
HqsPlEIPcITU/sZqUithnb8g/cGGSTksxN+jz/I6DxAbo3rDo9waNo3z6VR7RUgx
hZzuLnQwQ1sJ7EEVLZcHWrZfVs2wKwCnBzhfS0z54xO0KslaG/Dwmyu0JlF8KSRv
RYf3kC5fC2tbe3AJa0olYBTg3kG4O1Em2flzBBMbAkntGKJp0m1651BQaVSxJ86E
Eff4S5NmMVjpGnCNbiYl1o+GP10g/xZuLdnb0J2DBqVR5RXbqbdEI356JgejJa77
iPlzzDMzPbs+IlpHDBvaRbFrfZE1cPNpaqOOjvPAWyEfEsflrePU7ipW96RfILef
PilZkJLWCL76bwmf6WxEK/IbteScc1WW1sxVhZOGUfSRsAaW7xGhpSoobFx3UzMJ
m00YDdvCir6xezbk+m7DX1fR14RGgaM31hT3wEWPE094J26YHNly8ci6aiJlBEr1
k26UoRj9gWb11MMHTJAIu7jDb2v7QyMK0IVOlKWXwNzUbauh9fQQHzCMkpx7gkjU
Naibn/N1trBUilIzGGk2urILgxng5l2SxgmbvpVE15lngfAhJuhF40Sgarji0tzf
YxT9u0nYn3CzROg22sedKojoDN+fajxsh067W1CILB3HvQpdqrsoheijErtHu3Bh
HgW52BWAzeSC7FovhWo5nEd4mIu4S6H5LNNE1IFx5zDbtSsxDvq/u46Wexpkt4Ho
zG1sI8jFg098m9QRq/pFNC56IgolRzfDJHUXCMXDQv51eV1ScrD4WtcUyAcRUrDm
mHOGSaT0V0Ez/xzPRiWZbfwL+YqkLNkur0yzvc0Shu3caexvxK911c7nePAj/Rp6
KIZ5M0ITnSO7aj6tATbJKdAFpGF8uSbnPBUjuL0JgRVgSVZLk00sB47Z6zLYWCd2
m7SDIIJeOjqjhmGXB9siUszYe33vnsERFST43VpX8Mjk+PLaH9wscSIxbPteueWu
gtTGyjTJ7W3jU48xZz/ncSt7scAW8aJkVi8y64tFqjE7GSgUmCDJ3moeHwxscOym
CS3FsHUHMZyKC8UCc5oCG7cq2DRxQndxA8tpLF+EntYQLlOCp978EfbN58KHEQvV
qCop53WdvmEhkQuqy1cNdnWRJ+eFolt2neGMeUGzhSFzOHOHACU5U4WmPOZHvdMA
qULvaI5BVbiOfQnwMuxa3bKpE8DffuZUn2x9DivLZvUS4JmTuW60pYcWl76FaOv/
qShEMNb65EVAJP3DghNVg01l35u1WAvHm9zJPyEKpCcLlrXjopjCeL/j4j90bQ1W
e/hhwi21f0aq/8uIta1itgm5w3RfKtj+c+5c3FgH5HZ329atukPi1wbofiG+pk0+
66RlO/LW/kX1rtZ+Tj+vL98nNZ0raQD+XRl5k1p/c9gtlydFqiBiDNvmrnIm/ub8
E8Feca+p1Avf3g8r4eKl4+S6zLbEQUOoLgWiCHYBWiKR2GZzIet9vNaWvK+4ckd7
x7QEgng1WrvehDOFqYaDuiPflfAkbWC3nO3cQbBn8agRdZAvcYZeiScY7029stSG
vA88fYDPFktQ8J+8gcvoIJJRt0IF8bshC1f8M9Iu7CrMp7SJd5AJDO5V0P/LigET
cj5EbeqlYikNl+n9Zfj1Ygci6EARlCyNy3kdhiCBZp80syLx2hgEeRvUQWjQ8hh4
WujdnmLFymmbU5TWcixzppgU6PBOrKZn4Ef12KnNciBhmd5mVU+3S8pf6YqzCHCp
2m09xVhBMQMHGEwwD9mbZQMPX9mq5W+HqeeAaQnG2zZUprc+SKgF5TdlpTdGi+Xx
wg2V2hL0G+9tS4gI/6IErXrAKg8iOi1catHs0kYPnPoTfjUE51kfD5xCa5B+Zwbj
IurX7cue+C10v2hXAizCx1YWZ1wRiYP65EOS4Cd7Cm55Ws49KHMUnm+2vzOzGouG
RDRH7Yq2Nava88OqveRcKtGPhlrRe4lC68jmnjrUQOOGHyAxloVShB+Zfus4BWBH
KvkM7pefjogwkJ7dfMcBma60eiKyhUonhNq1whvHFhBx9z/zmV1vNv9mum+ZEiPQ
Jr+fuUMx9890AsHKuR1yWwWkFIsGhkmlZavuLN5Ls4J1CMDpwlt8oYmfTIsuRUmb
Hgiksuz+V0XAAZifUZ/kifjDCwn00ic1W+S/KIBfQSvSRHFjqncwBQEg9sLYYriI
QF2CD8s8ynwpxRiWk4yBYTjFVJ9fdMsk3xJgMML4yaruCQefuT2QS+PWK1ySz3ZA
3zL1Libk+68emEJAKGPLMsHQW8UbruThK4ou4Ifh+IvPC313LWV9xekh+a1GMKpL
3GBIqj6pOKqy1XaxFyTe+jd8UHE+Lm0fdC6WOWoB2hodY0P9y8r/9wIm2+HGBfpD
oXE4GR/b0vdV9U++6Uvu4VvT/71ztXxHPzeKNtShsFe4/AXPC4UQYhOGjcfavlhZ
Rrgix8+NsFOlbB2aIYRD9PrJ+MI4AV86Th+hmSXavt1Ud3WCza0u3mQX8X4vc10X
e3eXMhTqVS/8cFJT09+K/W/KxJn3TPfi/Gq45oAFMe2+19Q6OdiBG3gqf6IFMW7z
7NJ6FP2lICdASlcVt7XYK8Tjv0tScVzH/skjiaxiHInDTkyNl0bEEcPkmJKKfRLD
jfxPggdc5jo2LSk41FmLW09oWsogj1dV4DkqwxAEndUuc7F9LQZg5a1wEthOoB+4
q9EBrW5TM7+frITFb7kokP5LJ4Bur1lAMCGvW7iH0uwQOn9ItFgSI9GyMyUBAZJf
yU1AHXgUL67T1aZgHz83cPy+CiJX64C1y3c4GqzlVTa5FU+HWzPOOeapt7HkYbeg
H9YGS9NacR6VkK/Tzczpe3GoHZIC2VYMsLZ555nCBu24aMvTvnLLWw3shoG7/qrb
LzBg9BifPKrRgT55hPKQIvaPtOwfwPJThPwSLjTCRt94/rCAedg5tKtY9HZkCb85
q4YN6zwUx4h5EfMc1NpzJ+I0f2j8owLZS6gOZRI0VT7riColeBn8nzWK9pGK6zUF
2N3ewFoeygj8aTZUhnVb6K8DiPaVgk4YU36oQiQAdlPEY7TMNTAjafAyZbzSurig
0kXENKqFK6VTqllzpeSt0+vq9zccJlcHVKJOr8f02CrjhLGNnhyBaRFlzfDCDVpa
L0DHeGpdrZmQTo98+e+u9HAq5eIKwFRTT1R0sPCckNGlVZ31l13yuNn8AXNtpnJB
76dwYzW6YRmVE7Fa9FvATJ5fEdsspBU9zdw4IMHBAKOFoGjqMPklOa6P8M3Qz7u1
9eJCjACsl1vI1LPwJ/s/flFD0peOqIb11VDhP29Ir4YI5qMyvkvQ/CL2xbtZu49r
vhuQsDzT6AVNVw/ZXofgtycVWLPyUQx93Q8au/obMqxXcJ6sV3B6O8tDK8EVDgbe
4QZu7n6ySFLoqQXIBP5halqBPmgVkP+JmM/Ubz3kowsauSJtt6BJhRpEuVYpAqka
65OCQxwRD3x4iRxxdtposS3AB2iEuutPEET1cClby66rt6SUut4/wVF9emucixK3
D/a8tQx21ZQVrGJPm07pZsx7MIuvXvgevXNu1w9SNa/o+6wSCQP6eEhpSdzAgh1V
Z6XZGXWS1IMY4geYoriVDipN90SIYLzA/jn7KVKFqP8SbtjuEmPStMptnuwxrpwI
QDE93fxTfnYZ/c2Jqarimo2hcl1BeUIIC/6Fuxkm02N/+ZFABznCuZZjOpIVbVus
KgtmA19+afX0ZWNJFKA4raR8MwLURtoyWKVvmoE2hB3X0NQsJCgK0oHJDTvsBHwF
0n9a4wBcGY+HiykmrsjicqdCgDMuaZC/iSz9XTy5uIpHj5LkipFihVrZS/PAvgEp
y4MySL/JsG9a4xO3xjGyEkbgnFwYzQ/C5zQzmkshWty5y4DTkbnSDgvPgJQguy5g
CjwiynOVa0Hnq86TprYX7clzJK79Jmtd88SdDX6ifXVQikdwQj57G3VGp45prd1r
s0V1qxTDH30f18qh76HnorXl4v9SU1iX0pX26WHsHxbM/qPqsYH4QYQOzPLyvk/Y
TOdI+YPZAg6/xv12rRik2N/sL/aHc2tlyF8lr6xFVHiOR0TZ1gLZ2SHzeaSvuU8J
VA49mkVgoininDfGVANJQsFCvocRmR7ISaNqHcivXZ4tmljPJ9W458vwL6+6s8AA
UxdYfXvWSlg/kE4r6x154Eo2Syt9dv298GsKW0oyYsnqDY+tUnaUMafpbFv8UkfG
NRGHO9sEHk4iLkxsGKzILbJf6r0m03srs2ioy3j3IE8Xr7eqDvC+t6mTa1J75umh
NnQFt/s6+GcBFD23ngnbsmzlms1sAXM2WlI1YcozxmRBlNihmwdmGrhVsBDnuBeq
GLwvJCAgimH+XUNu+k/4tj85diFTKBsLOX3aGmSXJrYTXsPwp9hL8QWSBf8Mei/c
phiA5Ezr1fx0BvFtTAji1fRSN7W6wrBuh4KoH8VPflnRTJC4XYJdFdbLHGd5+TYK
RbLfDWJ1X9rhcJGwc/KC0ezgHcONr87tJEyveC8nyKYkow4Kd/qtCaX3+UFtJ0kK
yZzafV9ZHos0tYAiREX++W3kWg/XZuqct4UQxy19xeIxXjpyU39qRYMZqkk200Ro
rRFcS1Ske5pOJB/AawA4u7pQKknh+MhHH11E5Wqg/mPn6gU8B3o/cYAl5R/VAn57
6kcVDrAR0MGv/zgv7/UVo1ROkYOkNbnyl1ppigQvQijD/1cgaOUzR1jZCP1J+sg6
vu5pv42UD7sw3AJasllzjc/i6idBVv2Gh3gr5VV7M0njEV+VBrYZUAyI+ov075VJ
rv0XIiAUlw5KeZgsd+Ei2ybUR+HAJu04Cr0CKacvPcD/PI/vmJZXzAYG/t8vJR7a
atM1G2rtBY0JtE0YAO5tbGxq7/uxCXDnju2kkor67b2L42SYCOF0CGB+3bmNZTln
L5F/w+sKGPAAD7WnnhK6xWn3QmVp3qrlrbasOqZCp2EhoBF0VC7sS3r9sgxSbYcj
W2qpujRvSitVtU2juppYRpYrvUOPfUBl6MNFHR4cHcldP7RAJM7TRLDIDAYyso0B
MhQfR59maXQdAFTRsUVYTj9nFxGQD+9f7/1GHP+Du66utYDEaAJOcKfKAiVgfSC4
Vgkuso9fCf7npnAPEXfsonIazE75CJQjJBYzIxy2rZThvzoPwuvOKQaSnMqw1Xpc
ZpXNmIBx2AZzpJ3N8B272qABQv2oVCjFX8K8Mqjduh4itBoCi2GFQPYDxu5OZFG4
WbGPvlcTLGkz7RSksjg/X3H6lcG6YyCohrR6a7dhiIdKWOZNrWP6uKCGbX9DMcUz
GBO411nWLxNDPW//nY8fxE4kCVHFuhR+Be0af4IJfCeKG0wde0hlV81RU7wumfn9
ZbMRcXCcSpp/hCJ3fiBk8Mokn83ZHomKIAgdvcz8e/pFiQ7+lbQ4jpNVQuEQ+Khw
EZwHbVGZblYGYZMCVc5y3lc6o2lG/E6ovaWes9rL7ITKjrherXATfMMKFmD8EUmE
3IFKYT2sO0IXnQ5NRJGTyS0T1z4e4jnHJgsYejKDxsRLn7027m4B18ck5izbiPhw
ARAJZ2AFLiu6aa6u76gCYk2juAIK7Cx/AnKyo0QigMWoJync9h4rnBKoHKl86OPq
h4FeMLA44hZ+eS0IfdKMmBmfS4H5rah8Jr3D5VGqwlb+BJnb6EO595dYmppJq92J
T0pCn6638D+zkbgBwpUfHHvSQwZs0gw0phaLJM7elo2rWr9J8bmYw07w9tnWXlHd
mLqeJ8N+cc+3GRK/8hQqR/vZ45ETykq9hNArYDsUz+r2dYsMjKAhA+fMNwiJjnl5
WHzTxJj5sUo+7kCRQVE/pg6G41rIp6t78bJInx5Dd1fpkUrjgpJERz2lsoAJA5l1
olYZBJJTNnd+f8o3swKQ0SocgxTjSUJ8mvfqufHQKJ9LpOY9TCbVzykYlFkpsIHc
3sqdpTIhgwPTSr7/gn+17dySbmu5IJVR0gCqrZcmPjR5hpOEUwv7VrFTIXjzVBq0
rw2cuofyu/hP4C55mzIN38JlOKXDMKhy2cNYZ7QUn40G+vCDuKLY7yUP5mWQSP1Y
ZKMarWcWSVQHLsowNBwycOwnM3VISeA+LXv548rK8vWh652MMnQDPqyaOZW/sCzj
LHku13nH7DT429M/rJPw4VXb5Lu0rk/yyP3ZP62vE8i0sQ9j0d1ui6mb8fwKwwEj
H4q7kHFEOQ2EXJge1kh1ab9YvMp2kc4CVpd7cqRuBBPcMiIlgKonlGNNLEQsUNo4
Fg6G6JeeD2ziXn2uuGzO5x+u/RpxUePstrwAZ01bWAZnJZrJXe5ApJYhSPAbHcPT
6Nquqfo6MkCWT8fupqIfKC2OXYAQVmT5U6c0lHpsxY6YHTmeA+qhQxK4QFyuRKeX
KwCk3WeLElcG+alUiUSSyjvdo0z+bkP94FbSNw0mRGFBVf+xS8UzHEUaEXNqtVL+
RPECCm/ijjMRV80io5iMgDWIvjHIMISBJm41VcA5+6ScFSAZNA6kHCLyMCG+nPCz
Dhfp9wrv1l4B6O+kAPNEn5NRKXBiu1S17TBWJW8g0bSkWle+w0OFLSjwFWuslv3n
03m2sz4qGcdg0nN0CTvdEwLsuqlTO9yAm/fIfPgGJuIJFesmKj4PoDWYLlTS07Od
Ha3qNOpde47YMKuvngP7EKIKfr1D+MhRlWTVXq3QJ21AuBaqqGhRi54Ah6xsNebS
IYJGzPrg8OzaBERRkHP/BbQtWetbkkA6JEwxy5oco9U+1IpIkGIjXGu1FcTXvY2K
Rn6LW3VUzefCHDwiMEUKDzbDwflT2Lh3NI7QQ+2t5w1Ggc3pbEFmSdrTk3u7WeMM
oLzHW5+NHMdtP4uf6ChKPJd4HZ7hZtKYpTA+EPSpRupXFVYvq954suSJiaY8Jn6q
DLOIYoEB5SFsm6K2B4XvEv339RIuBwpSKKeozo5PrXLiHiaVZ+QIV2j/suk3MWnN
izgeUkFSTzdoZuFTK+2NKTPmsjAKXl4bIK1DKKgTrKDCru2hrAFr7j/Cc9Hl0Y3D
WeL3gvYFawP3/qYJHYBHQevuMgYy9G8qzrVZo8EwjC4J8rw4/ccT+0CBgLThMCW1
cL2UWhilTRSaHVKGTjtdr5Pv1lwj7REuo/6fTGmG1kFa4sENRx+a/iphnEhhgIyQ
nN4chDvgRCbHB6MIM8B0c5V+t6a5MLV0lcXNVL+KC9zBFpwpq/kWI/cl2vMvvhHJ
LrZUkZXfnLYTSMuZT9t7bxKQNiFbd1w8NPN0Sq1V8RnyobnYDpZT5fIIbgH76vSK
KABsVuc4kxEcmyukoHHju3okheuEIoWTCDKzwarsyRNnbv+Fwggb7paZnDRQhSrc
2JCcfomGJJ2Pd28myWsEuR2JFkU/knB/u6yz06vwxl/hUzrQAg8yNJ3taEOdd0iz
NNyTFPhU326ypCvBOI0Avojgs2w+yC4CNN7iaBTz24Dx5ZREjFpYMd1O5W5spQS0
sCJd6TRBW4fhJGwpGldEavO4FpXd2hZPAgbJ8p6sCYirCdolwfZ0ApP12/yFgh0x
WG75FRgGEOld3zCu0k5dAmRudxa6V13PBEjr3zK80T0kBVNoeYGIRPLGLTa4Vb17
tRGQGJGQJVA5Qaees46HdKq/UJlxHj0+TonlNO4yGxtPQE6nBY8wGvdJMMF/x9la
ljWXs05wERiqU9jEZuP/0nNGhod8bQtLDX8/Fnt0XFbEo1Lw3dlw82KEuzASM3ap
tMpizEi1BPcnGBHDJorESDbV9fhFnIBRRn0LEX9p9WS4ac8uyDwvBZqbxzPmDyw4
JBHGSc5hCaWEK5NVkI13JnDVMMILUvhT8569OW/f8f/iFN30kjuRBXhSxiF+qY1L
MeaDxtB7kfZ3MgFdyZcLfcEbGrVsZe0h47zPLAKP76KoBK6MH5PE+apxEhALhHfQ
xon9cJ1OCMc3l7UBJo874wdV14hiRyj4gbyECldcJSWQOo2MNtPbj9MYjNkiDoPX
zQKj5JWNu4FNVJrj+fdEKD3NymnGs9RrhkIwpGgt74ce8uRduTivbp4cOjCF+n0I
iiK/IYEoFtUeIfliDo1DP0SHy5nfNXQv9YiGdQzFgyshfKEOR3LF3j2CnSkt5/pf
OnnxkRrJOtsYfyY8lWyEisxb45qV4qN8vASpvGDUs6g1urTApPCNxL7USe9JDuF0
wHME6IWTlrrpyQ3IPO1e4iQxR2LreHgGBlfbgElAa7iOiQO+8WRoEFjxeRjO0Loc
xSMzSzHRSTRZV8bMNxMOOu7CeUhSUmdQVCbv6nRiIj/UlXAlqdp3faVwL7NuACRx
HpdNKcVyyVIU3uhQ8kRqBjQ0tQ7DAEnDcel49J+CGXaSnhqDUIKRndQMzOrfOE0I
FMT1/9RehRRH/kG/dSIfmy7f5MHDV90uWZmjSIMQfnMkjflOidYEnyZ74rO9uP+d
xxOF0TG+ltdKNj54goJuVaNCwGsEpmkGV6kwTjTm/IntmaraLsyDR3WAaIlQ4irX
NpoZ0fJfyQKbjHJHx21HEfZuCIGUfdXMRPQ2+/td0m2Hd+794bVgeYlGSZRuZSbU
ezyIwBZ4WJZ8ekvSZaXFDSgLM6Eq34mlUg8vQdnCMGN4X2lyHB/0qlYGg2Jgpss9
EO62V1kn/52AY5dbWf6DgZ7FQiwC5RvSMD3M/6Gs5l1FkQ1D/smhlCyizDUfpvhI
qxKrsDupf4VfxJ1zZTmse6noeZfJNqXCIwMXXmIqG8xhF3f1U2NpXV043J+noRlW
ahbw8T9wtizh6erBQhsfVgKx8z6d3YZroNDLA8DAbNFMMZCazS4VJBMO+FFmyT5S
vGV7JA8Ny0UVkTeFV/tJCYNo49zOAgz8p1XmXagj6xOwZwjM4/GRMde1sJc7/CfZ
mZEJHWMnGs8uhcDua2vKQM4Ipwz+rP+4tBOnHY9leG0e53QOno/LUaUSgOsQW6io
7d056GIvZILAJBJFK9t/3xNycQIParFZ7J4LV+2yTAnFbvLjXYqVXdP/yUv1cua5
Sua99k8Gpg30dqxiA/IlmXiusLfX/W8QWCPSh4AvNjd46S9g39Dj6OukKcijXVO8
JHee9DwEU7o8tjiPCegPKbKEMEISTKbBjDvETUsle+yqaYxsVJ7Bqb7dUjbRMl8s
mNk+GtjNBTXQc8zMJupMhuobLKsdqldviwQU/o4feIxZ4zDUfZrCpn8eNF35e+EV
gULbTqPmtM8va7kyxzykqqMSz5PKKeDQGguoDUBmZE7g4WyITw6nSZMDAb3T3cfX
g8oWyy+tvG3GnlbttrGPFgpYeemI+52LiQN8XLwRxnCMqGftWRkO8PEr/2NEM1ip
VQ0/QUnNoU3iLnphrvnjp2o9AAU8bbhTatFwT1WM4rqeLH9zWhcqmCYoxfIKgO/O
YcZudtRl364bnb1q2zmEnIAGDKJ9BQ1XhVLXdexeWM7bwmiTRGlqz+bZr3WbstU5
AyHi1PbV6XUGceQZ/KswKx+zw2YX75+RasdXJMHDTnSbtZfusaFjahTtbp7a+Dpa
e/GI7GUWmru00wGm1GsWqQTII/kt/tadDwey5/UCIuG2jtLqOBw3REpgqgaiARm5
0D+ggwTOKJ1pm1ryecznX9V7PML6qkpiIEuXY+1n5/E2pElGJfaFJGci9MroNmqK
0UaT4TSO0knGYV1U2XmeJJNZjtY3xi4yAJWNcchGc1Ci3GVM0SKZcUI0NmhSVDN6
exsA6AfgmFHyIOLqcDy0ItE5c3344l199bhf5FwGTxTq1N9b8MHrgCLojznks2ac
r3pTLf+Vbp9YFCxit0nEtRnFdcFMApeSnTWC01/Pgy1KXFdPHN9rBrkaOmxpBad1
dEnfaymA/OuFE4mHtPh1KHwKiXtIais+/O2u6Rjrtd5kr5JshyVufYINnEOXgRVv
nNpnxmBMHz8V9T9rZxc1O9ZsJcooZFxvmiWpuqGL+p96FkBYhILS29IENxvLx2Cr
nAHn8XNr94ZmT5ZUBezV6+ntRIfUsow+dUCn3SEMGQcILB7VE6y1SErGAL0VeSad
WT+VsYAfaWLj7yWJ/t0SQgPs1QDEYJEoEi6WscolYkvYW8JnnOOZSvlScqXwp3hX
95gqxEhqIC4OlrnzmIjEaOuB+nBkRo+TO1ZM2vDr6ljJ3Z/EvSUxP5ZRdvMh3pkR
LE8zMN8KAO5h14U1LH3ayKevac0kTORcWKdyAmNCS1Xq3BnDAW2nlvKwUTIbrIn5
8uPuguONGaYP5jvidi7hiSX/lIZ608/UpXX0iwQsSpUwJv7vcJuxj74rr/XutzIA
TOLcEUoS4u15VFENu9k/nUvL3sGJTh+/I2bdqUo5bgMK9GiM55Z3yP1OVLS2aqGJ
KRgDgM8yGA7Av0IIR0yVNpaOm/IgyzjV7Yns8p115Ll/DUWHnVUQOo5fzPLqc1W8
8q7DVwMQBO3HWQSXOkVSsss2ouIx1DCaZipRoMmwtYia+IEu/TvFhcsHttluYGMN
qn/dSBzKNaU0Ide25Mf75iB5oIMCKQNi4bCQNECOaYAddXQzqZ3bj6ImHw5MtX6Z
/Q0vLhrELjTkjPjH2U7xmkEYmdmw+AOU9RBkTU0211rSw3Pm4TuR+S+SGELxuav+
z1TMmFgowu6fvpTXgb0Kecgfqb4AclWg3b8fH843/mIL6m0APGnitlvI2u7G18g9
hnq/WH/qb3cPFCQaS8Q2TOQgrzSiZzZoI+sPnq2jBM9WDfLiOEdDVDipwW/RiqlW
mwb6Z3jHHmHd+/mdWvfEGaJFui140AHMZW5omXgMHTAo3tqFVH3uBHof0PZai9qS
Alug752ltf+HHbghuzAnyJc49CVynP2nYxCKXd5Di3NE8WeX/M4fg8KObB4mp1Pt
NeoSS41eq5LjFOzw9+LCYYyamg3OeD6gU78wqnYI9aj99yn/z6YckYTwxqsxN/kc
CRQOKnQfNMKK09b5JHzgu9RJ55ms9YLvvbkBatjcW7Im8HvgUtxfMGDFyLwr6oPh
g+oXInT+nW2Atuj7AqeSfvnSHMDEqYNsrBL2lZELpsXxrg4ZY9W5G0+yjqObZs/5
GxPLBHHhGZOmYdltGf8KXs0hEc1B1qiZdTWehuTdlVdHRbmRnoPaKd6om/gbYsE1
rhjAC95fXxVuThoX7DJfmvtKS1YHf8l7OLDU+RjRiAItMtE4qIbnGMoJJhWyIZQ9
1dSzjkOdERPe4z7pLgdULmb+0SPj4lILzVTMuAnzx9r8/qfZrFmimEoSaeIkY4UT
i6bzjtWvgHh2TAoXKVl+h9xXTpsTH0Y13IYRm+4ffjQHeUKFpAbu48Y5YBpytI/4
ckTkRPXPATPVIJX7LhwOYUZacc3jESox3LIrI3LZpwThf5RTsDlluRJQuaxU1JJv
tbgrpIdiL//XCcZ6ljc/ZevmIacYZAjVhdxd0xp0+wgU2GiDAPRag4epjfniAW+C
jC2SBW8sFBJ026BgGscpRC7TDwFeOv7+4Uuc5u8Ub0YkekeQIHwSEUwyYv2fHXE1
1BDvL2ujRh13qWInj2exuytxHOmf3Onl2jLGZ9DnnHgAQg3o9wbVE/2fpvj9Ng+G
nAp3Q+XTkUKuIyZxdfQVcW8KMcZ5C/ZZpYeKUNcQ3XywMuWAVPA2TDim8jGxI25s
epJUxqccXw5+HXlnQwzQqXY7klYyzlF/fnVXhS0R62Jq+Q18vZjTWZsoVrRiqxdY
t1TeokbK/ia6/9YRjTn3BJE5D25+0chT4EW+pdKkqUC1z3By/5hNx3CaDgR26ON8
Xux8XIDJLP5GRTKrKj6cC+oR9xs3cSydvve0PwGrmplsqWg+7AY9XKr0I8ljlFor
3OwC+yYfLui9xVPU/a6g0xjwIDM6rMqxUKWgWcrROxPwbaDflCKQTnZZ8BOQd4nP
JRG+BoluVHFXYt+v5ttYn6aG2rr4yT7scGafL0whRKsRBv5kxReCdoU5WCqd7kVj
+zzf97OxU29BExHGANVlZZjUmNJnhEEmi13Iwm4Hun4hO/AgIWt0+jBaBFyRREj/
LVZCWK8OHRnDLgkQ0Af0Lb7LbPprwExu5yyoFUjALaoiWfj54COGfvyOIFIr6bvN
xA4vo/BvywdyHztQlAtVDMoSnABxjhRLbPqwX//O4sk8IqhpmSqEuNLnwYw6snGv
RyfHxAlxvrIHpIS2I9+JVwy4ueunJRYFfI2uFgG1o9T/dPqP2Nm5nm5omQpJcuwK
s3n12kDkoB/czOyzqjFB19eIePGhNsh3/OxiGNO7MAAKoL0sul4NT25htNTK4zsq
FM2dp99yIThsAlkeps9BRkK+TxkAv3efbRqV6hbNaqh7uH0p/k1DWoqzNDGpE3va
Q6UppqaI0534Yanb+oK3q64+HVAoF+e/xu7jyqoy2ifJlNMnAD3q4jQLvU5AEOzU
vViremMAg1P4q8EY4X3P7juuSs4Y6x+NsAUU6MqAMXd4gShOE1HWCT5hmop5YKrG
xtOtjyvh5UBQaCymwGa+LYQGsXl58etgcWmBHCfEPdqA5IzETKf8FCb4sAWdj339
CH+7GUBKNq2ZmRren8BhFKoWewVjGJiCG8Nm7t97xsFAEmYg4xNO4RCwr0OKwky+
09s5GJuLjNUD5QMjUqZEhU8U8rBIhze86bfETmG3bKxJwlkf+0k0ekdTsPOHsi3V
zqnORNsj0+rDuLTBV03ES28SCfcf1/kbeFvLhHO+2dRlg7fXLCZ9+YYXOJsTNiXV
JEvWRnrMikqyMUtCV7Yfgo68Me+3d5FdNU+BR8dRpmZi8Oty8yat41arBkFW2MoT
tA0jDPE1s2PyHBRkyt2Qx9QNXMbgkzh4gdlSccWH+DmHbyCEkqpVOoNh6MbUFx96
xQE2KGYZZPo2WrnvTxgJzZOC19phWRimqk4YJrO2TBWEATa4vg7modmauUUIFwo/
yHCKz9nJ3gT5boq23rplO5SdacQIMbRyirAQhnItazDx4MvWNQCL663mmpl406K7
2PKNFGLQZfOCtdsmjOolXUG++G32xplFoZQMk+GV7MBqyEWfUv1Ctk7m51hndUxx
zTHeCW7t5ggjuiY/BwuIfoWnViaxROSLkZhJ7E9RYTGZJf5YWiWD7nmOmA9DSkdh
JR1Rrp7RP7Em+pmFeTcdH6xfeRYVsVdYts+ohDsfAwW/toXBRRnXyS0fmY+2UkJf
HZJxnVNnir9Xpjy29P2Nkgh2azvjs6n35/sdZuO1LnqMYHmEMZyGzTM+5RzW8O6t
deyHhRGN31UYNwX+C5O3EdxtzK2Elxeu4VjxhqjS60suk4CFt4EWSv7M8Sx6S2Ec
IoTpKTUgYAROd5zq+u0ftFu845CFX6GsNzfsFbSVkcYLgmQJQmo73M95J/jcnKdW
LdDQgPwGN2A3KLvLMN3cslhuGAYyLECVw4M5yV/6oDAO2njHsjmogmbg+jHW55Vc
67nwpTzyBXRoFHPruSIEd+D/88bfI41Q0AYZ5SG6YQkwnqaOrFXp0JbNHkNXzrw9
rx+2h33e8yAv1zHdXSf6mijQZFK3s6EAocIMKXUTsQhnjwIS1QcAHzFa7Sy5toRB
XQibunRISvkOBeeXcjvynAgNfZ6wKUwZd91znn1l/90jAg9mrk9DSlZ96JWPUHje
FwLtvE2INHfd6QXNQ/mbqZYUHUeR4ZKkY1FudxUKlJK9q27lpZvBHt6p/o/ruE62
PIHhnyCgnEj4RnOwhqawWROuOU5G6/teVl3B9mHiz4cQGSL22zRqNwNYrnawDOVI
B9EdV4L8OaKbxKvQFDVF9pSFBWKqpTyb2Rqe/ox1AbioAd/J5524Cj/EmLrFRZYE
ExYVsLjqX7y117Mlfe3qO9ulsn+Q5FYE+4l3vQ6cb9PJpSVRApZMqYj7tBJgjwbR
w5N44mjOW5DFTiny2SD5Ax3rdpnO63H4j+l2klCm3k0cq95kwHoAD0kq+t4Wxh0h
nqIJB0KG8KEbN/WmZYPljDYsuOCwg2kVmSotRRp7wxE4n6iQQaxyqEpB4K+8EzkM
NtKmzveyWSJXr/PBAhqG/siGy8OPquW2OJ42L2/Oz7OW8yoAk8akmvNgaBZoHBYY
JL6jK4JmQdFnclpEEgXBFEbD00akukFgqqFexSWipLA6WpSiKC+nOdpDPMXAYLef
Vd0MCet5GNjLS/25Dxn2ngO9/Xn2Htmdb6rs5E6/ys1WXc1hAP5XTbh5hmA3zZk4
Fk/VO0FMtD8IWEJL1oBKAH/uvVqFYMKZvi5Dv2+oEfpz6o/qFnyhg4p0oLyacheF
377oWc2cp5PwW0AnWzXLyNvtDZDnMi9t7yhLKSJJ6VLEXhQEx79QB7ERFPSnnenx
3wG8UQqXk2wKLBFfGIbHGaGAYwazbm8gwsZ3yk7AAfyMipXgUsOMepYLQe0KCA5l
hr3cPDugY3DZvQVsouWlccAXh1jNGfnE/bGui/ywz2ERbwCzhsD02zGeXS346iKr
mqDelByRkHwKli0oyWWymKQW4biGv21NGFoGVhl1V35Eo9qaTwMeEkzzogiUz+Sg
7vuaZNquPRJjjdT9CIvEaNRhYO05A/kxdr+s+CaTKv1oxJDTIFtScdRGkyLK0ZMI
aVNTZiitKm4q5cIaLtvkX9NTl8teJXboUkA4sD9X8ujXFKQPef1pqnUnkBoDlmKV
C+zKeT4h7W2rb/XrNRSEMVmIEdjuKP7GQ1/8YdtMAYEDBjLZkAN+xwIms4XnIZ+G
ToDO9lsVzgvSwSicYEY4LX73cRF7Tw+LTlK4OzoeOkPdsIITDfbW8Tqn++N1y4np
F9T0SfAIj89C9ONWF4lPuca6vkWmxRWC6WPfledetatcdb77xTCqVcep6Q1PCfGp
+W8vHYRJ0AJFVXyY26kbSn8SGpxreiKb14JjsSgv0ukcswchP55C9JNdKOPZnqPf
UskV5QCGopPmKq2WoNXiSj0h4gBCiuhh1cpqUgLGdVqcxtpxhN9YLclqykfBcmIw
SOVSgyFxcGa+bVwaMJS9mliEPD0l2t0bVRnhwUCo3VW2jqgT5s5O6tODEmKjG0Vs
WFzTWs7/TquJVKB4TGdxm/bt9rp9CPiPvmO+l6EfVItnCI7FaZ1BDPFKRHmxFdlG
lGQwmx0bXbnw6f5WXe7HA7Nf6wUV4+iPfHMuyrBbl7aquG6VDpQr1L4oJFbUEChx
oan4S8KmVbyqeNNIaAIW7jilvtOP17xmGaaBSqv6EaRlETgzMzSWQvuvKsBt10rj
ge1ROsowU2I2o73/3XINAhudF3Iw2JDuNvBNAZAzEjzgneY5AR6a9VFQjM1/4kea
sZsEZSQM789Zn9/xXCAuqoFjJ1bC7o/OXSAuEnIqNOvulZcC6iQH94/aasHPRqW2
4yAHw2O66owHmv0jZB01/FugKH+d6d5fjcDtNpCn2ewqGnRYwGCbmMDrCtV32vWp
lENHYJMGrwKBoHjDPUIdq3GIMvPmkwJnH8SWzpUB2W3ytyRWqCxKDbXBIpwBtRDF
fQ8p3wHyNyY2EJQj5+j6oGDfC4J6ZtoKs6Pqi/vM02zopc+U9y6/LGz+0cDrutaK
RHZnLylALJMeZlYsy8PmspIrUvTcAjpodFJm2aK41UOJ/FQ7di5tLOGUhGdGsSf1
BtbOFj8MuMnha8M6M7qIZWcDSuGnZJxhKboirbOmhEUv91Fm0EPoQgr5YQikGdZU
O5Uz0ZsmzlZjxZrM2UQ1A+uG8Ry/s+/HH2+16nzkfrWbAFSVmdoC/OGj4EI0ASqe
/cIbZPs5Uq+tXZ88HmPK+rwfjtZ4dTYfU4VH47SHOG2uZ55AqZUkAJyGmJt3LNzb
dVTNeV2dSSWCeOl9d33Tj0XKTdSmIy5FpSWAFUsgXmiG2GvN1bA6NKgba2ycDHbI
GNCl3oZFAW1zzjrVaZNOwX21EfqsG2b6DtAU45RuKmO7ALhPaHLNS7Cb5QMORJ9Q
XxBp/HbGhDtPVtSxgD34fdRPxSTyY+SWwvwdrjS3U1HBfC3ZOn5da8mt2kstkrxq
sYqN3oPXQAgd0fcyvKx+lL9Ws2wjT6H8Q1q8cEAL8Pzldr4DhzB0b2jZmd1f2JjU
5iTmadAAmsEW8O0Wvx3pI4vViHr7DwOvvMHYY8B7Bx0e3JH7Qrow3S22jw267yPh
ZgG/UNQjUMlX3AuMmvm5VUEcMlOC4jkd1QIHBevDHK/wConCyV3Go8pJX/NBMZvp
HT45642FyI+SMHLa7wO700YU8AZLp8Ng4xWYvL9OhldJbV8fInEqk27AvrBXgGOV
f4o74n3hDPD3kP6GZnvDPtZJ/6Cp//Go1bv4uHFbzZ+TXj7PgZUYiycLGzlrQD09
zim8IQIwW91ZPCHvfH2RVOdI0hX0HtGosBnNkKB8swndXHYjijrQpETHv1xZsZrv
khpJ9QCZ4ZZWkEr2+SDVCpx6HKvRJJKJ3EQ47v1gPDUDisS8wuvux2PC2wJA+hlw
SGtQBHrYErjH2lhJoDFxw4LE7QTfQVKsQjmSiLwOsQuJdpqnzOyaFGGJgw4gi/nv
ZIWSCs0YNQ1j7yLCQR6J9/T+RMwNyftKT8plMWEZ0YbbLO4Fx+lgjF4N/CJdZtzD
RBKiHUAPsxh4DP7R6X74nCHVczi44E6qLV3eiKRe2RuK42cOXxvFCQJMeAAteeYr
qGzeq0xou2DMWKjoHFyH2qUssSF4GAjdvKWgdlj9pTfg4bhSOfdfNolqdJDbIEyh
c/847MD4RQFGhqbW5fCSlGu91wSgjd95zMWOiGE3EqPVE+mvkPmjZxnrkFFQokPj
6cBqJ+nvaYtAKlUEinROO0SpWgqG00C/Sv6QXw+l5VvCi8SodFCnccH2sp1iWQDm
X6X/Kpz9jvlJWbbklJW0tudzlpM2AjpKdBb2W6bzg3baosrIVxfaZDsJWyorEQmk
N2Bfk9sHQNIswTOoFJWV0RrOE4daAwILmxHnprzrdBXhBtROUTt1Fcjc7S1g05qK
xDzAcNrk/LPNu4PRwoQz98wLnVF5kKTa5+6T25bkpyh1gQYDPwAPd8aT4Wr+7EsI
ww8dfseRUdFTbQp03254q4KKqw8X7MYGrr4a2EjtSygLHgIXtFyhPexno19DnPXY
G9L7+DsgioJeGhzz0FKhGVoeeqeviMToxs9Z+NqJhxYtUAnphXYSITaD5Lf+N8XE
SokYZzPRMvea4c1z8Ug19JqSrXvtuuvBb2SRrxDkZMNTkbXMWAJarPDhGDO+1Idd
h+IvhOYcsJR2OjLonLJMNdwNLph4IgUQ5uJyc7/D+6omPRTXDW38GslcSCPnnqG9
K0mk2mPIa1STXPzmLLGf8osf1aBuDLKFg7zi9rLgLQFvtwHatLFDkfrmPUXMx+e6
AMfLONgBsESP6T53HlLDTkePbjqwLgMs11hc8MLAUIek48LHnC8vEwUvKoNEYus8
dLF2WyqjY11MdqNnDeU6TCMscax/VKBTJJ1E+2+DGoU8ueMMpQYioRzikubYUpk+
blOtUd+7fj/6O/scgMs3SO6plKea0WUpRyOWP0NwC77uUijY4jphIK64PBeLZY8i
xbadgZGYTfRF7SqAOQHu5dM0Bl++S8Xs6zAxh1JTDfrcA1OceBPI+tyyJ0ELVpAB
O5ebrcuI6L2i3KtOy2x0vbCpde49hqcSjVRQ9wD79KsNTl5WuFT9Z7V6A9yWKSia
5wsJjKoQ+mrvnn93XyJ/ZQh+I3150VttTwPRHhcNxLxC0em0q0VmpWQq7YUEToGg
jyIw5LuxN1B9DrutlC6rPeGvZPziiQqoUz02FPle3b8rhJlynU/lLZIE/xZlYI7F
FKUUnakAnOhAPB4nRvdwBhUv34zW31sFh5Dv3FYsFFSdDNuL1CNKDKRJZAgYNbXF
C+QCvJNFGI0cTN1SUCodFmOaKSxQNnZ9dv0nKVHeIY49zloB45dx3lNKsi3Xzko2
p/m8iM24HXUJRqL7bEhlLoxv/veRulhtNg7YLJu/yTTv4HORr7FbCs0W0wIVhqCI
5P/e5e7zWRjMbrXa28TvrEGLKl+9mh9JIgR8R1jzJhBjGHjNJVkToiGM3gUj/16P
qRm8wNoDDDUZQMNm/82X4mgbrKDbI5i0gyY6yeyI/Tq0gbX201zehzglwVibhqe3
TtYOIjKLdetYuLdxSZDaDbzD/fidNFmw0z0/x+1VMKVTh5w1US3xCfRRUcgmNJj1
Z6rANN22SNHha6gvL0chzBUr8XuaYB6dsIS+aF4fYtU1lSdQzRlNlZQlbiykoA/Y
nal76rXo2r3E0ZUb77ioXDNrdvWoAhRn4jimiG5ovFMix5QdCT5r2toXmGzmxf7R
wxgt1rbaFLJ2WktakD4sM+U06oAEVHWra2lYNlgTy/1J/pT+rVI3Ivpxs6SOPTsR
2caq0hittaSn8Tg/alaCy/dM7V80D8AntfAZ9VZW8FrzZgyQ30CNO+qMLdrKUKp8
Tgsa++JJB7TCNkyjaw3vv9MQ6+zc5NmAve3lTvrc0lQG/m2BFsrUWGuzVCnK9XlT
hlQ3xS6J8OXHZhfydSeHGmLwd3wFIpyUu1ircDm4sozVn+c8XoDdTog7y8ElB7Vm
RGScDc/13l6kwhA9ANVtD9WlkEKj3OBCcszO0ldcjalX4qqGPuQgtg+qNXh5hUm1
fa5ePTdCFXgrCEg3vIh2yVFzr4HwU+Hq/gZk//yGJdl49qbexht5NbQfwhqLjOdl
YMBbfU5eHBdmjRau2cTiHxubD2hNuKy/zv2GFfEcr16noEedIjaE2PI2R+l0v11w
3BCMTHvtiUjSc6nwV6/EVnEO5hQdXzTELPGuYjm3dh1XaIzFDPo7yAPYTFRZyK7D
8cpKIY+vz8V09RbvBOPxc1QniPUKli0wTlURR7oXMntU/X1zZYXucebb1zgGCahO
dtcqqah+XibMLgaN80PlfKs30tDfk6DSios17zGTLK8jkLHZoEp4Lqh4yNquFaFW
jbuPgissV7I+BxP0xvvOY4xw3d299XAMh35fuuKDodpJDhxVg+H7fiIOfHnQ/aJG
uT3C7vgOrpKJIIyYhvnEdYd6G+rhNmfUbKV1p/11Zkp+y61Asdh0/JsWNOQwQDSB
ytCTBsRBiFJLaszY1Sg+M47JH7kRrlMv8/TMQ+JzVQD+0KepWalaEweifEZriJCc
FKqrnfh8MrKCqW16Jza+dctrXPkuVP3rupO4x3eu+Rjmq3asJkrFf55q/7eLxLo0
5h2wToBHK0soiFg+eYxG5M1kEQ2P7itkDL+GfH1bs8BV6fHuSHEAYbCbrhTpnLyz
Tl764MgPQkBOVhgygiQaFvBzPzW3ecctfsCTDHvudQvLwppJOuiT885YvK5az8VI
Y43MRXhKQ9fsyQU3NJNkPh0ySdgzIHLJy7KkRU0+fzwaxNhoV6M8QvBt/JD83v4g
YefozYwhzY3d858Xtv9P/Al/hOrf0iflu5Ng7gTukGQBXiEoHGXuJuqp1eyPh3Vs
j4QxWXOMBsaekaNHaVtJlG1JxeqXNXaIP7rG9liTbjccVKwtk3qlAoyF8x2gUNSn
x6K635eWEKDBP4SlAgDdaNQpcPswJkQiqlXG0M8vGxCbq23WQrjryTOXzohBDqGl
WN0t6zgq7PySa22Bpt2vIBs0qJGgvaJJIxlp9ZFisxS9M7f4VRDvW96NKphJovZ9
j7m0zJjgjTiGs9+pG2KKBzxteiJAvCL+BsbBILd1fIn36rKX7JgzhZ8+kPNlsOCE
fDAOhxH0OSlb10FLpGSBsXp+NTvqiqqa3wtJC8QVfqYtHn/LLYwXdTSwVKb5EZuL
vjiYcBWz9nBdbO1ZcxsyrCpBebyZFOdhlbLHSWDShqhGrHFJ6bMvrqfkiE8F1I92
A5i9IxObRqm56ZL2448xvlr1SFjPTtgsgouZxKORalvOzQ/C+k9STx0yDCl0Y9wU
R+wjBYDxHWnZhcesQQp/GzPXbNRVR6XsT+TvQV2nhA7zehr5ZEmIeg6yCZWYVrkU
6c4Luwj+XNJiZUV0xBtkNzRGbmGibIwqXq2owDxo88zpXj/pTGPDpZPblA2QWJ63
+6+2CCKuhQ2pw2OsxdPwFYIt8G5h+TD7JG7tH629IvkkLf9839hOhCf3IroSMsia
G0xJyA5TJa38Aobdt6ikIwYfTc1fs8mgsVGRlnOu+4PDdrMgOGGrmEMiq/mRC6Df
2HTPnxWTw/OMgkYjYmDb1pO3Yn409uZ4I47OPwM8tYPk9CDNJNVYaKpLzw0IhJp2
y3HnOhMSVLBWu++IrfFcor7PwASOh1f5N7hum11QjwMkVXUa6rI5PHeamoj0PnbQ
tFkvAjgTHpmIW7mlYY32K1aVoFNrZb34St7r5+mQ7cezSwTPhOBJCizJXC9xMzhS
VasZODtqjmjPQoCsd9MN52ZFM+21UkQ9Ywu9vybFBhfwPJp7oMdOeloNtWo748cp
9dkKU6GOZdYn6m+aOQnLCQ8BtFj1I73J/oRQrmXidYK4QGYUTPQN2C90SdcJj51r
/L9ra7PwyKiQymHaLy9KXrXTA+e0daeTby1aP2WMNFl1iuJj2cjHL23CttSWxTKw
NpIN9w2kanPGlRJEIAbOjHZGHaloDL5u4QJXcvZELnzoL/NfxxToeNWZeHfofg9o
TBIu4mxCpgTKzS7wa4RkqN87e/BiTwI0fPc9754pZFadlxc8vznomKXuSu55IsMk
/c3mwaSNxHzWnN/REGA1JRgISrIJitYKgUxgDQmEjIdG1rMBODXtrSBsbMfDHR2T
eRDKDIuBApIB/4v9H5hJ1HWcAd5ZahHnohl2awbOrXgORXIA1EWRV/8VjBpDs4BX
3w/LR0JOWc0nePrhuWZfUhsiy6L22CCg76SWDKu4v82ldo44Yq68pAlTPvduYEVg
Enc9tckyDfai+/71Tt/tL5R4RlmXwnbv4zmX/UkyE7Cz9TRtszuHh/Yvz9xYMY54
es4Rob8wep8bfLNJwFJs12CrGNlnPwKpYlmWmHK2vJdcR6OslS0KqdvmaEs5LmVl
toRpcgGrXiDKnRfZ5+jSTMTxEpGYA5nEW5TEAyjgMcq6TTCD+xEdRSp6s44yU93v
QPIkagrIdK2NfSOU6xItqW0XYpfZYpjrun+1aAzMlXC1GuTXK447cbHbWxyWaI86
ZJCjnasln03BhPo+q4x5tDIQj/moajKvWTViQ1bGJEa1yz0yXNpApx9KGpeoPxYo
SeDlixbH3A61ph91/fd8EViQhjSonQFclmFjY/WWinUnPBpoCOPh/OJeWBA8Rpg6
qT+yB59jzVRVpMx/gAhLOnG5tutacUkFHvGuFSWIL0cFlonVAq5uMN1u7yXSnbyX
R9EMDx2HDJmnxknpG1ctzKSDtSdWAqVn22mgL3YyI163eKCxjStjwcj8PVDunaxm
0/gVwpyDiUOiSLJugoRHRn+3qyetM/N+GbT/mLGfc0WS313z7TSWk7aRA9V38J99
NmnkTcqMqeBWBMXrGN0e9U3EIb83VygJg7O9uzLCztQXiVartQPWjqkDgzIJyvDa
Sy905iEhck6DAJs3GDbTHZQVtwoQTUW118xDe1P6iYTs/F1VU59RDgTR0BcH2He9
JziNVTh58ap8sTrcuNhJWNHJ5LL1REv17J8HgN0X/Z05HyARsD6kST4buH68WbNi
ci3wty7Am8/9ThF91kiiGdOEZx/ysNrAEOcGCJYt8RyC/ZoESjPvflIDxai9Z4cc
5v5g/6u5dX/VgJlDDBVt9Eym+1eaqaeM0MImL9/6RWcvFQAkZkilp9p1jk7JDHhw
3DNReZXYXod9+yrKg/2kEAzfJbLETzU/51bI4i+NNCC8lhERTxjEOP1s8jYpF2oQ
cRjwCOpvhm9Ojw5UdOsf2uHgLhXin5UiXTNmK4EsfHV+OHn0zxvckdFBNBHFIPbj
UULa4IUf1fN5s4z6XsLJ4rfZYplErx+5/d3ORC7YlPA8nUbbCJNii9qPvM2VqSXt
s19W27uHRLbRHJ1ps9M2JGfcuwcGrpjjLvp874l0Dg+lWCT58RcwdCQbH3cz2Efm
riGgJC4gKJrE4zpn4LP/TpmqfRFwVoxnxuFt7g/kg+QfkeYchqynsbr90Apa52Rt
HlG3d0nDekEgaqQD4WzCYCd8ttFn6hdxLDJ8keA+xHtmPX+dYaTkwGqiyKwyc3/O
kPvZHWYlHdcSQBQTWLFPW/9aE3sStMg/Ix1uNSIxs3+5d+L87iU5Y23Ad1+LGg8/
RjE6q6w3gTkA49PfhnRpl92F2FZ2GmyS/02im7wLuZJLCaI6TOQfPBntinPXh5QW
Yu09OLEDz6jWrV5R8WoZR0vV9bJbEwDX0Z7D7wBzNuWeUk+Sl/PazuH8LTCXzcYA
nHuVGFgeUHHXlnNcayypnr4N8EPIGzQ7Qiml1lEDO29dWfhpw0s/B7k5HjvWqdn8
bIXRria8NZUjzEEe8Guu33UPTftCh++LauDwgfg/ZMB+u4uq91ONAy4U/Ud5wbjT
wrRrLf2DBwQ6FWYsh6ruF41Bjpr8RcIMo+69I14dt2c13OuhNSd0k0cNXr1wnB2N
B/GIkumiA5Bgig120NWhp5Z/lEo7FzUJFx5j7V8wTT1GzCJRxsKxPG+cB4r5YSai
/LHrh6ggFV/EadaaE2Yv2I0xxikOB/TawiksuXjMCtDMh3O1qsLaknK83XZvA82o
/1pHmaOjMpFdb009sDwRwkPhoye31gGei0FcidbP7wklhlz4ahAsY+nzKuUAr/4/
W+WYrVpDHdZFmxOB+PxpMJDmyaIY3NQisbmrZvbNMMrq+7m8OjYmBV/5lNUWSM22
W0wniXJwgtBsjjm6Lys8tJtvjqpAa4GAIkEunh9gcDC2HQFhKZbvRD1APkutZB8S
4uak+N9f0x2B/N13K5JACzMCb40KQx0i2b+YtUGCNDtdg9NjxexHwYBBXO5M+IYy
P7jS5ns/a8Jv5+Dggdl18pqllgs7lsQMfo4BZxn0D0kyyh8ZC0jOXj0JKWFOcjL0
lFwRSCa1vptEy6EAUzY7aadmouVUJM8i1tPF1BO7A1bgrhNwNgEo5s0yum8co4gg
l5S/xXobvRgaIoD9Y67cEx4leVfIC4RYeyHQ8ysQaCA91OvRXZTME/WOFzdJzqK/
jtPTcS9vigSsxmMdrz6v89cNzhtTJUMyTeI3Fnn2PF+9oZixWjWGhp30hilNYCsp
qREwztjrv3MeHjRFNn4yiDBA51bSW7ip0AtGZdjF938yxizdlQUSxdBZpMSGKjvC
WiwNJhLqDsZx8xSl+d5OjkzO4OROkRKdj/OqxEcDhaNpDyN9ysbOds6laglIDtRS
jAwNGM5fDGhpRJmc//Z97vuwgzQ7Xlx9VpRhlWCYMQIPCJoJc1LVXh+mcttJ3HMl
dKql7zu5NH8xybiyaJiHfJTYOSESRI9vlx30FnS85ZN6zuz+bKa9zyQp7bZRwjL3
SJYusDwbnxw5dq2Vir+9EOle0cAzn1tjnHRp3XCJYwR6mnU0Kiru3+ETNbf41q8z
LpU6/ORCZXCKnfKjblAtRniDF0pGGg5WXKH5AOHvCgsB86BpjUwNyeYWge5yKgHX
QEJVArcJ4vsNmMGnidO8c3m6ec63L5Gl8mW1OESdbTyQ/AMey/1BjrN3mniqsbuV
7HUgNZjrnVB84rvVJkH6Rs9OGPT1j9fNVMer4GsnHBoxdxjn3ZjUxJeKR4GzO+23
oxpiEDRF2kctqYSqKUx1aQQoj8rvsFHZDtV3ahdVNfYh0ydcWWVFOB6hskCHhSbg
cnIi/c6Y7YLv9uFN9+76DOKwxK2l94wA3REXtQi2X/0fz+H0o0sydBaonNtImAii
cG9G5nsgCirxN2mEovMgzGBvJXzSLz0eBv5vie0sdbd6UqpYqfyJJERIWogIs3yg
5hkKsXu69CthF5S6g40+kHiV/VhtHnn2/S16Q1a3zE9go/xZkcEFml6n1IuSm5G2
/VSSP5Azw+dUqSOpG2NgHKgODqypOWAKpI0oIoodi1gSlpfgEokJcgfrwFGbugM+
8cxjGdJlEwATXhie2Xg5P+SamzvWYLfvBugxXhprz+s4PwYgpSb/nW92VyRRbGiD
3kVgISXZdexbSqi1opk2xJzdLfqQ7vwkcvc/bDckKmOdUEHGv6SjnPfhzY8Ypk77
qg7ajef6TIYFL2B+X1Z1sReJNaUPhG4xpZHLlD+FWCSN+GACYyLSMmj/asYlbJRh
1tD3AjP2UK2sdWBUcBKVNNNsiG9NsHSNoxdNT68zQhVdIadp6Qb5Tzds5iWD496Y
z7/UWQacR7mRW+JN8qu4pASYppphE5M6Kl2abVjbno0twwQbwgVP3+kgBFAmvliQ
2U2iJXTg6EB74vA11a5YCqqssfR1gkGG0n7BAn5Kp74aIUdGE5bR2JSa9kz9T2sk
Q9kpjwJKuwSlMH7b+t0O1RfRGSS8Nt5bt7cFYkab+TP63R8/CNKESr5xcmixVUen
F8BV9NSJXxtlrvaarpLbCYSKp1tZAGzG3QvUo3Y1AkQa7Yf/HlcZ5ga+vjNSw2Gq
lFwsCapP7N8FsnqFv6jTtgybqGu/+QVQFqX9WHna1389njBgAGz+/I3jrWzM6y2U
CT40HNP5VPEefzp86/C9ydrxBCgE88veTsQPc2JCJh0agOEE5lxxAGnqAid1uMm9
kFeAvB8oOP4m+r9VSx0EByqv1WrEZB2XyppILpNJPv3+5N6UuLjJVhlgwbJD4Oxu
zboqKytUqEdkHDTlWaCm27lzNCNNDUyEvLVZLEIqX4iLDvKb5nsmdtw4jVkJDerV
4Y5+9tlxcZXCZ6AWj0EaoMxAZ2LWs7Kej7kRPNCieiYH97OVyC9om+5eCXKTqsru
W8dfryfvO0/cyp/Tuhu/3xSy9t8rJ4RnaVjtaajkgWRGKkSDV6p7zri6iyKfqeUS
1iBTFD/vBFSluGXD8HrwBtN4onSsz5xhU0Eeqh+9xzobPazLcZPZXVUQXlwySWVy
x2RgxBtjhrQJJO/OpXMbHNyFtFOqu/jVQVIesddpbsiGWmwTZv5+RbfFsFkytJV6
XdgVtAxbbUfaqu4+IlG4ePzfNYZKmJ9GfKA7CQU1OQki2iTPAWvBgKtrrnh0exOf
1snsBdBlFbBlUpfqtwE4o+6m/Dtv8yAgQypQwvOsra2n+VJh+mcu6751FFsOjiny
iv/YYLvRO43CDRjXDBSeGR5Q7VACaNjLQ2SZG93+ogwO1SImGFof0K5g/H0cMD04
P3YWbbWZjDCko2Nnu9zkOqspQUWvoP+LfYLJ278QdASCM7ksfFunhzTE432g/q7B
QCBj5b38J5+DaAvmYFRwxaoTbxTFxFLWcj4Xv7sp8clU7/5lejAtRDF5C5xTD9N8
qBl3TWyfsdFtK7TAQrMW8jLuYOkLauQ+lmPER9Bw02yk2t+Ivoae1F7+gxgUaX6W
St0Vup/1WsmYKNQlqeNq7locuJkbaUzdy6+p7uy4t1wybDzcYkENeNJSVajmyaez
7YTg0NqHgK07jxBITptIiXTS8KR2IUC7FzPO6SKeRqhZA1EC15Nyoz+INaFJ6tEQ
OIcWEhvpZE2O5JXE3gOn9FQc8W15T2J+jOM+AIJmbnI/1F4RSmwKzjpSf9qpVmd3
1FerzRYamO67ktYL1QGpbFAKvWRV6GrphSy9GViAQGqBYVVyZ7yGzjzyBahJnC0a
Ie81cFrmXJNDWPlWPGMyVjsstOwZOuMwsybpMIWlpPsRj8xbUzzexUN8ToKXOGiV
81y2KEDg3BRWddBcCIrZJqSmi3wPxszDVlQiCige0rzCqVPCGuudrU5yZWOqjRvl
iWFGtsqkpFOSnUGMBd1PENXkmkAJUSPhXKVADtCY5pHIPLA525SjmYH3zlhunazV
GzPxtEaTk4XjQUL2ug9Is/WTJ8yVxssuRDx8w3YA8+g1uKZZeXDheNaIrXj9d61P
U9HA47FI4Nm5AQmx3DMTUvhOrMyQmgBgtOd3uinA/CHCk26oKZ9SneRVM/4R+Y3x
94gRZhl6Yt7qeeG1lmTLuJmsa6zf1DqxqTt/j6vNhRyPxLUprmHeEC8rKz1wECwD
diMbXrth/S9ac3RDFxzxSzuB+Ti/BKdz53XO2PyJB1jFDkKRdVsSUD5vb4OvBFuL
U7QipxWOuRUplviG+amGZNMUXqoNFgEzBDtTHHp6xRNkQWLjOOl+yXiBpbRh9X1F
jyk75qbrPuvk7uG20aucCajI1a26qrVjpW7UtZAw5vuAuHL8WJHOMLNkenHt2Pxl
6jGkT150ogbKzdGbunixdFP9mFrpc/tqKgC5rH6K7aaxlvkfv677A7AsCE0ZYYLR
JhfhOijdnSKwYl3oHnIYqj1tmIt0JkzHIwqEsOzj5xdhbnQpj4cge8NR/kKh3Fkz
oRjhW9Hi9hbWcah5kowSyoVVBWPR7PlATuNTm6RvL6JWAN+lu0Fu8Px5h5stDwRA
WGNrdkvK4ixtGi55qCoAgCE2uenZoQOUF6VFjTGX1+YR6I9bFSbyfUg2o4aGNgLt
03+e/41DQxdgheIs59clFdGnEycf3TBXR48fH4IzH0CjpTGfL6uLXjyRwDPl8XuJ
nSHZyAXw+Mf3Y4VaNVwVzUfkefaoUhfFhPcILime1BPjfarickJ7JAaHywl+BU6k
+Zo8VgoQeMk2JM9ROi8vWOedhPd8BuPL7aduhPirR1uP2bKEfOFRL8JXKhrtD4yi
IJDcSNY81Q3vkfkGZocLK8G9aGTey3/Iet+eKhqSFajE8m0+gNRAtQ0ppEaAGl4U
8/w9JFDrnhxH9JnmO9N4JojVoactQp8K72mpZOcrpFdQm/Jvu++Dz2VxrWhYQenP
b7r/a77dF9N30tVMrLwTr89ZhAAXI4a5RkrzTjowz4Tz10SfTPWB/tAciLiSqTfQ
o7SLNuDQr0Wdv2bFdjYM1ELd9EIMxbxN264/ZbYpd69PaFU9j7l7z5hbfHwm71q7
Thg1t7z871kJXcYXelHjpLR01SStSOfW8SlCR0Yc8lorPuysqdLKfHq/r/ioNpG2
NEMr0lNphMZ6UaCFyPS+Dh6mfIu96nFIjvWohl28HS//hXAHOkX9OgsVURw40Iug
at7kfCjyNOqt13a6XHmyQunBfK3cpXQwQHUm66oCDolqwiM6TQhYxSibzfjOSxQL
C+UJ1rZGcmpv1aA8fq7CngPnX1ICdtda/wWShXg/ZMnMJT571e6HRitf6oTLeLmM
MKZQYyrUIXIGK3xhX+yFN+JKQSwQF9DEN0roWdxduFi93BjfUCGMCPgxMnTe28jT
O/pc60ICKLVXButl5f8o7pOaoFEELq505UXLwSkVIndtsi6WcP/86P7sGd+WWkcD
5I55MZYQtFGavB9asQJ7ahCTrud9QSYm/FT1P1ckEOkWOKsqzgkHa5n82RoulMO/
I2iK3Q72QLUe3UWuShDaxtllhQ7iXj8ucX+rhbUm0dlAT13ZeNh1hgmlPhsvmlJP
rPM+Hzl8adNMioixNMmXKuP2p4A8KmRS7CxY6xLErvX8yAi5gOGI/ZpUatyEjtpX
MwLYn6+Xw8PsXTRQZCsWHbVhNhTEemh4FRsDGQ/KqOOxEC/RPdsboI8U68nFZQkc
OtIo6b9UX9tJv7Ptumr/SD6vJCtExlWcc+UMoKfnU7njl0+Nu4ZhCO1XSK2Oj+XX
V8U1jGmhgP3l24LGek0s90SG+Rgdg6ZIIlrVKphgN3wsCMdAKpnX9HTB2pJP2FGn
WnwQh1ZUxMCQmxisHSLFVXBJicuJLMZg4ycV0KAXfkv686Esq/kMdRKR7kGbQem9
w/7413/METETeleGT8wxLCdgbKQ5hK40nX38Ur5uJXBM8GrT6AWzKxMffpYJeydj
V1ZHV0aeH81bjNBT9WfT8wM0tahITNIQoCSKISG8FcOb4ZHMCLrx6BX6ZAOeypk+
JoBf3+cknjF1yp/4jZp03iQEUJ6oKfjUtQprv496Cu0/QOoN9+EfF2b0w0XkonJm
Si8cMHvbTKKg+CLXpQBVfhEEcW3xXfvr603ZUGZpHUcv3PaGkQPYvV9KAF38xF3m
3ZBOGcnxLUlDUf434/7lVvi4AkbQbntcEAyRBrUwK9rtbks53AeNqbjk+Vj4HlUG
sDXoszo3B3r1IvjWsVjLv8k/3cUQ53w6yy59P+Dfh2tWQY3HqbRyo6cvZfM7b88t
+TJbDELb2o3OG0Yn5enJgob0C7dsXf2KOAX4zdoHObvCIR73t9Bzxlo9ueA38G+S
yJR/wIiM4nDx9Vu1ZqZ0uuiSF7eqknA5nopI5iCqbvi5MMLo56YM7JOxiM6Y3t7Y
s6PM20xibb3NniI9bbbXarTkWeMRHsWmXyu/fs5HIstNlXgUZh/7Y/RxQCf/JGgo
IOxtIXiwCmXAOfQ6ZiiLXiXX+bEgVE9alVBL0MEV9okYr0eTkZXsoA8Fwn2UTw9C
1TFCF2b3UPI/yc17AY/8wSS48g1999YPqUJT04xi2Hbewdre1qD1Q61hqdHSYmQX
Q1rXR1Ykqq0AIvT/CN3lD1cWOQLUDBZ+Fgzk94VgJU3yYBZTLdBLVsC6rJeChiIn
DAfw60kT8zmpXIJ5Sk2dvFNny/CxraodqE6WZ+9Mji0jLoOhzKH+xFM2BFgb3dYO
6FCwztJTWY35+U5YZz7Zqa17Iz8uocC3jsxV82D3osud/KNU4okSCE5ITHTNfuHk
kt23tj4BIIs7vtPobDvSkZIZ8+GuzRP5pXEYKFsyKZts+cFXx3ehNwbr1QAhGrOH
MWphTghZsk5eJhDWbFiSktMXdFr3dRpsTWnVFzLXcTdg2qqqy6KC9wDpyrqTC4gG
TW7JzKYIZnU/M7v58ONdbs8C03KQ+EKR/gNxG5WzdSOUou3GdQdkloF3ttckKXZj
3u2R7NVlUooYHAxHP3MUIid5/uR0yRxjTJmZCAOfYNwrmY91AIRYk6Kd5VwnFc7M
lmCVcCeDPCEIddJBDdzmfxKlgplqAAxtMUSa7vXNa1Wdm/FBYjcr6IfQiZr1XXe+
q1ZA1+3gUu30NfCajvkB1/El/Uo+Ufy/eOddKOEvdRS2rcEI1ZLS3E/TGsohYlFD
0MhoiOV5Ler9nFWdR1/hVGKVgaLC+V9L+CAoEdlo34ebMjIZa6dU3DYHAx7Pe8no
yQlRvMia5Zc/WdstOiXvZ2f8ZpE5eWVmX16zPMi5PLhqcZY/MGU556zNbfxcJsWP
TmzQMBxC5Shg4kiljNI5Y+jg2gg0wg0aVNe1jL1F19VKoBWwKpggWu/IuUkgJ/n8
8qIxtBa3wVdYBL8iLst2/RxKH7TIjxp+gR5v05RQnikCbwj5123pFaPk4kyVSvLH
BTGHksME0LgvJq+yTIECGqxEiMaKUkqDKdo5MvwYHPot2zdLkB2U8UfToewQlseC
cp0eM+qE5HmSy0HWznPRqqSMNJKqSb9VP3oivDl2PBb7dasiCrTgoGkxCpZGx03d
JuXMQ9mG65npLTT9tUfpi7I/bCSipvqygnlhPqA/c2r9MHS99b+wuwADmvgHM05V
1gs9fjg5EixRla57k1xXFh3Kx9Dj7wKb96s9Mc6SH1sjW5aT0Kr/j0/+Oy5TdZ0G
IawLLZ6qBXso6qh3to6rLSw/tubIpCKs0RX+VNUYzCyugstWJlYW1gxoxtEcaIxs
Xu42aG5QDgbQRRzjctBgKyGvqfipb1C5vdp3RO3+VgUcheSW6/c5EFKTUGgIHkQG
5Ed3yRTRWD5dDAtM7brxK9ZdBCo4zUWQRf5qvXGPl6hRKBG8U8Y/K5OR4WBvphfG
6yvP8kVizwCnXBSq1ctVCDOKSr0B5a/0apP/gQhhz1zui0CHhh0vNmpl9layPcFQ
n2IUDWo79tu5mR1GUZWCAf2mywSWpt1arHdy8AfTIEwQISg6x/dPJYyGaLHHKxNz
Q17pjSW9i7LOymSyVJk/2v/sSiokYomTDdPSc4qm5Kwtbj/pv2p39FMr60lSVV5A
vHhdMuDAUazZO+R/NIo3vwd2IT+4em0H7AGT+44XqdJ6ubPzH7yYKeNiUb5tCboQ
wdkNlwFSA9CKGFza1QLx01kelH4X/FtgBwe8TvAD5PAo4sVrrxYI0lYEu8J/DfUt
PyqwShDDu4sLlTySUHHtd6BgGjqiMHA2wKHq8R3A+8NQyghTVUlD6dKEnEt6l/9I
bkcg+iOYcgWtuLWDuaYr0QZIXRDtaAxNx7mAst66jvF5BjyBtQlEjQ7tVVhUh2Ni
7GtXRI+FaBXbVRbQ7FiyNN4lC962ypr2p5IarzYez+McPNtIfJHfmOIMvv9T4BMk
CrwEkrEj0fynVpRHvWxtBnkaAUixozeN4X48OcxfFEWAgJ6kpMQ5sVNbNKzFbPBf
d7FZpf0q6JfEcH6IqUlQIkQ7YCNy6NkvJ4iTWM6d7gFHUIWa4Wurxi3o1ZtnI0qi
UzOAbY+bV+hk+Zrf+q4FLc8bXLT4qy0FINif2lwBDub/id8M2VjGrCBdQTCgNrX+
IhsKqpuTEW4pdhleCDf907AIYvFJniBlSFX2c7K+VgoIf3Kc36IKRKDqQGl6SAmV
Puy1WVbOxyRmMivEvttljYMXZjUH8Zt+6qDr/s/pV174eE4TuxPtWAZeCstLN3r5
0oOZHSmJfvpHhZBt0w9zybfvoZr1iQCEZ4jKics2oXGjpZqJ9DTTWl8nHakD2iUT
gvTkGIJWEySlQ0PW5tNh5ltQdy6sbWMV0UaMXVzQhim2Zf4/OQkKaeRVYPAPmayv
jTit9IkG4AFNHRMdblvDXfFhw9sV4Ry/jH9RYoC5Akzwl9UBtrA6o6ZwzLgPbVO0
GfgA05HuGYg8o64EudHKPHdEL+yIkwAYk06y+cOORB6RxeeQexSSoXf+AftqC4pt
5sM+L+NM93LMnJfrtqz5cKsrd8UCGtc/tJEF5tDdFcrSsITixBj+IAfP/1kcZdaP
KVj0aD2eTCCUjTSwobe2tC4favoAgJXCpc2EZ6KLNZ8L/aqYQZfO7VNc2UIHY11o
WFKoKwHLvzRZa3O0Ss4q22Haazr19z2YN+02gdHxyYXCpNm+dUFRWaTOWiJuhp6Q
jTEXzahQ7yz774Uv+dktoCXRw6nOk4DsOlOyC8Ui5HbnjE9XfEnQAkPb9ujXX+bf
GURDPs+LF2nNbg7txMlmjnVI8IgmLbMH6UemjDdJXH6BdjKhuuKMKfs/Ywlk+/yh
ln0N7ado167a9Et8YXCg1k4tEFR7yptaBgy8Cb07DmrmsWkdIie2AWMcVzJzHq41
GmOCFnCaboR1TPZLHJLcbzKfRBkXsyUtGNpg0peG7kAdTCQ1R3BkdBIFEPiadecg
SDKGxsf93JW+zaheRyeLHdHkNiqW0UwS9PgORsY4bumm5X2DNjUOSegqSgmfET2G
fh8Vt+0XFAeNN2sPU8PAX+tbaD+gZRqyAVtt2X5BWDVk5UzIp4XYoi/m+MC1O4od
o1H/NroNFDbmfw/srtOuqxly5bEy2br1bBGpA0rfEDnJ8oFHjqth+H3weCCSGKSG
dzZu0XO+9iLVJxYhJNiwJL6GoQlKR4f8S5NK/zxGhvrtlj6tcaImYBoglWqGFAaY
9R52oZj3k8+ShkJJG6f/cSiFu0i8bZrzoJ28uGZQTjYL9Lr3kxt2Zg1rQqDNHFAH
9LJ609CXmO2LwHd//E3T+RU2RDP+y4PAjLdtHpH0dJtZSmPt9xcnBhlJXCygyPYP
Hh/glDLx3jR8voXc0Glhb4U/RDGPsGDlposUCEsHfkU/uxy0PQbP/9QIutsBkWe+
KibWm7cRmx8wl/qYW9oP3WLxpLoLzZmrQugeZF9F4Yjg7TKnP1TCEx5nfDOQJj/4
2tlkWEQRheUcuxk+F1k4TQSFQg4baAJ/XcQYaH2dv9FWphYTkZUFqn+aQ5GYlLFb
v0vdWfImxzC0BW/5R+hZuM+vU6RsdcGNLXyzD3vQ594QRpVv8lZ0hkvfV3hUa9BG
MvsK5kRDX6l+n0zPDQ0ugKy1MwCglm5ljpIJRW2TJH4X4YFQStLIVojao8Wb2S2l
W0PLsPaNL6UJXboPVJGt2SsBRxy+y2GnUx90Lc/nRvI8Hwh2bL8IySilx1R3OODP
nNqMGxd/0WRnmCYb0SqUZFaERaRRjmtyKkGt96tUeXQq+5VXU1ijm8aDUnCgSwxO
yFRtfJ/X54GqJLS4f+PSYCZwyCV8eFqgEQd4gh6KUfqUtEaI7NPQgFwH/wVz77y7
Ic9AO4URKO2sdsKuu/tBN1TDiTkiiOyde98U98nb5y1GZqqgHEqjnYIlQfUonOgV
MB/o8Gz+rp8LSVTUyAsL/ch0SW2nKtt460nrup5T1khPO04l3j/4DlH2hrnCi1rT
j+CrQzazblTCcaIFZyagAmUGGVyDx5+bnepP3o+HKC96lMXhr/Cj6PiSEyvynO23
1uRsLQD88I2oA09c1r+aYg29/MuWGQzMT/W1hExalNzm0fyu/PBAMqmmtG231HSo
QX+hb9qqaMC2Ha4RxhgsaERmjGoqxad2qUHGOEklEU86S3nOHY4bnDxox+O8Viv9
pTITRvdBeT0sAA6jKHjCVXV+N90b9N5INroem3abbcCfn9S9pRZYeH+dlg/fI330
k2bPiBNX72ELRHTy5tNRH1wH2KKmBT15sQ4fUUBXWRKA77VFZSgR5jHXdX7m5xew
Trro0LYLcKnDnxrEHa9ls6CqdVW57y1k6tntW9UfS7T1phFn8yHG6cSq5rnexZqq
Ase6M29IcQ9Dop5RAfemQoQVmVYdHyg7jszR8GmUsWInNSJdyugkBPbK+Zi1261l
X0ZraGUsyIwCM595LrFoaFdx1jfbddcTTtzxJD2VJt1BpfYIhEkV/PZAUpUcilCC
qBWL5z7S+800IpoSpcX/CsTwkit/IHQL5Wav3Ph4T0sCtfUPQNmNfvFDO6gjrgw8
/re5iWbSQ493c9Iy75tK19Wd+jpEHoZSM5eXJ+lsUX/n7GuUduFIwenGM3bNIxO5
5V7atiVj8J75fuho89YvxkGlvSczhD7yCQiF+jdlrR8iM5gQ4lSRaUKZ9BdaHqgk
lbuLEx8KAWAeurAbqPLUgsMyBh5sRDcg7fZ67SPytE7k5g+A3dKexQRwKf4ppjeJ
VIo0t58/zroRMLvMvzCQyzLOQ6/8IkeltiMHMYF5A5QEMpLop5gz2gww8eTyR3G+
caSyUblCV/wkiI0G6MFmDNLm2s9pkUnd9bw9vrYAgzgIJyZiq3r5Gvq+P+QCR2ve
RQmwQ+EfRlsbE6rnwAarQt9063ECgqoXHHeX4CsLPD0bgHa2BFfKkxmKq/LDIirY
eyrGNoMAVHHzVsaIY1Xlnydakjkr+sflgVY1G77VACGTK5HS9CqTQJ3QuaK4pxwQ
ooObwpRUqjB+HQnXTGbf5bp65LDurmCuJoSonXxah8BjaO1kI08Man3OB9w3xPjm
YRquHDurNG5xMZuF9Tx5UxtJyyVg2E629m4DEgMEXu/+AJDHHxFFf2brSDvwB3zq
EutZj7iA4fOydoxz4E90AftiQ3e6kqwpkymMmXDmWBEgXVqpAylPjm/mqZqMlcHi
LFjMq2VHp8/3qaO5ircOm12LuOnRma06ezTl18JRNj83FzQWZt+onKv3IURpzpPy
CIGhjBq6NM1MrNX9Xh31zmwipSkYCojk/teB91MWR3+D/18koETjxt9rRl18pHE6
gxd60vP1BbUjyATf2SE0vBiXTKeryj4hs2sknkE3dzMoMZEcT4FWAzxV0CA70uGP
h4BMUjx01HX/D4a4T1lry4KnSgs7rlEc09cE7eiBuLh0sqpCg99eUG8OGXHP6zt5
7XmuKrXVEeNHOhZ2B7y76J1ixq6KhduA18NemV5HEJeA9AlZGDpohRM91DAnqDa5
36NJJ33unohMvZkRBsGFQNFlISeDV5J1Fv2WYGSXEKtron3j/srddfnkJ8Us+MpQ
ACs1ZJ8f1/ozTRu9ACvuEExhwS4LcHPt7C2h3nJqTQ6pZhdO+CKOgWdT7z1ohFt1
2DFCJF/Am2iYPsiQZ++O45otjrzDZQS8nHqjNo/H8TQnUmnmp5fxriQaT4bq5Gav
owjqYD4+2FJfG+cs0qWsPdbPPkiEJuf3ZRXDqil96bg08r5hVwlAYsWGkSqy/0Pd
P9RCK1Kr1Bdh02R3JlM1B/JeB3VJKSSBXxfV8HvEdYT3J9wsRtMQgZyouTIbtJfQ
FiSKqMK7KbAV1/Oms1s8XwAttVDxdouVQYMK9qUtft/RFHpeuXXEPjdnCHP7a/Ze
0gEs5g3xx1Y2/Y/P7bcY+k5n7aa1MXgDX4UmnL3sjsyCjxzv9Iy3mpeYYtbzCVbq
2B4fQILsPHNb8ChAox9fzKUQ9iD7Ox7N7MwcwUERFj+/u3jvDiU41FsNg82luqSy
l5ACzgfJOU2iImbkwpJ2uMPF7cPoBBMWvH1VpuOXjt8JtxmDTGq5JNHZ0i+Xabs8
ieIM/YVqxSmE3poAppBQwmYTwndHJiRI+H5KFTMTMg6RGBopO3IaeiaTIs8DLblY
lNBQ7CntxhwPLc6IcJ4rlt6vB/CixiK/pFWwpUrHututmr+o0w45W5OeYkpmdsCq
OK7LQ8wKMB8wVvsHk9uiGeNTTkt7t4i6OkR7UL/Cs1jfUWM/2/Mp7dLMQL+p2Qxk
7fRq+o45suHa85yE1NBNc0PtIMnjfcpmCTaG6Hvv6RQhT533VczK0zpkN0DnwzgL
NhWDHCDlX8ReU9a13M7iUXlNy030UeDUt1NnOwe4WDPpuvGWJNBqxzhevUQ1PmDF
2lsBfPtfLVGx9yRhXgOUfvy1UtbLPukHaUeZ6BPI0rW8uBTM4lj+I3dHgxNyk4hm
whXNoNQ4OMytNxpqk+vV0rMkyWGsbiGaki789FTTHDvgM9NdmLHRWdvYZhX1I7wX
fphlN+s+Yg3hNPxpfi8KK9YARB4pvFtuN9S/M6ILHb50nD/seadwf8K+Zm0XHFDb
CvW5XsYBu+O84Z9fJYJqsR4JZEDVPGBthyqp5IBPQLzDFbq0yKCw48/LTNOhEMaO
slC9Kjs+Fv24GNRDgJewQxrdwV4kUssFcigJm2Xe6dXEXlBb1d65c5sbg9vAW3n2
zfGBvgu38w1K3DqqCD6AoHiBVH4U742nl4ZvyW2FQmrSp9jlAX4Axejmufo2R27i
wy7qxhALw7Dv/rKiISKDqTDAf+qReQRLkehwGV4safZxUcXbXXBkmagwEy2aPkGB
MHtcFjloTRtyDn5eNcbZmK7qae82RUjupomikbtXm/lBShe0QQXPoix0te6Hac65
NSQV9Q6CYZ1DUkWLvsOHFf6vK4JDwh+KRwFsbAm1tUH0fRmkgLlIsyTu+EH6ZJR+
BbtdWjNdec740xFv8hmyiKFLnd2dnCAekIemam++Xs6iRjj9cjUfetmmPFkHq70J
4PflvuGwG7GLEsm0t4l/0ZJ0kkt7p12CzqZL+YIrYVGqXGtNXMBXY7G0YP0uKTzV
qShm2eehKMJ9+BbP/0wO1aibssgtbfFths8w7b0zTsqbvpE/5jJ3W5FnDNDUpS7/
EPasIyCldS4AX38A2XWMrMn/v8fz/hazAGismBnanzFHzTdD77YKyxV0jZHZx7G7
1nbvByAW2BaEZAQjFPUkSHNtXZ62bD8arjJG1A8BAwa5DxjB2uCKxmkUw4rXqAWj
zuuzqT40FguQLcrlbqHbHrR9lEV8KthQ6uEfous6vZzSFKBjlA0ynTSygtbpmruG
2P5qgzyvmo4fPpM3W3pXS03G8fzyLSOdR4feewHWG15AJSTftxcgQfXDt8eXkfd5
IDs3ovZ+ZtwObZWEnUxflYLMCksYBBcgHGO0qWzJuqcaZ2BIaBWZTXoDmQvS3IDV
G9bHqitkahloLZJHm6A/dBQ77QyFohZo3pXphkJWgw799Xk0hjBlPcDEQTJX19Ar
hom86b+8It/XLNE++gdMfeULBCzlIPMAJNQlg/Tf3ebpgygxfzRLGejseECpxcTq
Kioqtmo2gVAmCxE9hxp1aDXaPg9nmb8IGq0IqDoSrKJgFPGSJGVKhFmBVcbAuQ5j
38UKBvKkrG3UetbG0ooLxEGGrpRoTxzlKYeM8uE74h0Mm7SFMoR0B9ikm1e5j9Yo
hSycZNSefb+9HAOAik6yPlCN1MZUKtsGtIqrqCKRy9Du5YxWXklzwiqZGlk5ZYHd
u6bA0+GfWFOsBFhRIyjQG4iNONC9kO/YvHZJEgJQBm2Lj/AcHnOSIzMMH4XLEYiQ
6bL2Rh67G2o1s8IJhD2jTEXkzkY/yMCXYIEaz1BcHxG11cOQnK8NW6vCQAn/J3js
LQcNHK64pEX3Rz7pTRuJVrVDe6BnuyNXZvtS8fqS57sQb7XgjWb0515e4GmJxJaP
fs0OyeE6REzPlsAw3Z228dUDA6upv48WVRMpza2gZfRrC0rA2SA3TdsS0a70zcT3
gQb2IO9YRYr9MlUTDVBIQH1+bItPi+johg5D/gbQ9I1FY29grTmNtzeRk5QvkB+P
d6IAuK02GzRgDxw5qRNGqhhOya9TBywTKjXfUdaVonhObuSIQV3fQHgHGBRZM++T
SazuVb1ufgCFx25LkDBzCvXJbzFhUjOlgJVKINC2srMLhfNsyPuCDLo3+mb03+SZ
SEZLNxa/yU+y7X+ZTNp+MkLkFxaqEOJLMEKoF0RiXr6PGZwQ/vaFqVwodokAVC6J
sSprjQdiqeC1Miegt/T+/SJlMrEfTerGHhZGqXNp3FVXz6LU/Q/KT5YRSXfSYa6R
zCQK/2/+HrJHRQNAnds1ajFDqaRZshiUWnuMtfLoqHqyzKjUs2T42UZsJINF3dB5
bd5Xq2Oix1gwmePN2r/nw5gnwCqJww/mxU/GZ4IpCZWs2b81WZFJNGZAir81etMB
u/S2UZkWiwlX5zPrWL+xtYpb+XgX0GFpeMBJ8BEkGrwH71a6nUvKI8+d9Ew6rjpR
gvOf3iXHQbidknmcRY38qvHZnG9MWc/e6nvrbQUsFxjAh1TOOSQSrKpg4AZR9bkU
N6664PWblFY/gMEYxgO3ygFF62Bzfmx2pNHi2j9zSw/77IP7mSZQ2dBQ9lSxpmpB
CoswYVUoEs7iZq+tKh3dQh2aCB3ZW1Wti5yMG6PW7leqq6aPh61skY5Pcp1RBiXg
gSPNoEQKCT8UY5bvQkIwOILyGGb+TwGva3Tx+MRTO9zN0SpQJE93JE30UfPNOmMj
9NLLx2ZMN8usg5Tms27wJ+sFkr8pZgPN2b24PV4TS6Ua5qoBIly6C2H4Iu4SFji6
Wam+U8UzUT484VjXn5yGpooHAzuhYxarWSRqXzLWuKL5+xL2ZgnakNuTH5egmxg9
2oxXa92DfgnHiwM859IjrxdHEQv/hlY8Bz+kopY/zVMl9nKlGCLdQHVAYqWQ37yJ
L1jP0fVP5TzoadbDSXZwYdVr2To9l/m4xU3TqJ+G/tMdhwp4ort1pl197kYuB1DX
Uy1Vr/hIe4DW9ofDhbu6Tw+Sy17JmMiFdGp/2bfauOg1lPGNjdK+vAvzAt3kXJMc
aYih1P3KDJa34bf/st88mkUTECbJDjnB7Zfbm7nCt4EwrhSCqQF64y9u0Vcd8xYv
yBXEZbefgurkQgyx09zCwoRUrpp9+mUNJWGrzRY6qZeeG4hqHj/6E6SunysSQjvN
Mf1haKWWmLopSem2gCfIq9mzsFRNtJwHBnU2MCqKCHAwrDMPFZ/6+g+4xemR9DA9
4zQJ7juKDtJ9vjpsz0LQojyC5r88CUCcZEdMxgHEBCkShTobbTGFYPTJPTIv4ayf
dq0tPEA6YR/CjjjEL9a2vJjeyvJfQVHgH17o6TFL3UZaadjcuNZrfvhK3GrZswnR
SqCkKeaqkoCzEDSjPC21Kqti8OFqmzz2PhMK/w8g8T9MU1LDCuf0im2f7Fdss0sJ
Rx+pzucDe+au8wH89OwHBjaQgICOw+CCQ7K6ASmvcLekvb958D6xZ4v4XwE3+61e
0LmpaU43pNWUtgfxGq6MBF7l6x05zm+ITNd6+IW/XTPVU+FN2x/I7ONsFkABoO20
K24S7Tsvno52/5L3h+ODJEJtyPIW1jPbKVansYLDxpakQCbyOD9ak43SSkvGxrRI
a2eV9kr+Mi1Qla2YRAdHTgEYlgeEihQ5FnW4xTInmPCuFL8J7sKaCVCJ3Qs1Grh5
Ojb97zU3NJciqNEYYoAce3rOc37YnsJjUrqHHEnny7LYhZU9zAOg03hMxk4FTend
adb0BeoRtI+4ddbcVYQ3CVQSh/oVPhRyqosS9WWH3TmNfqbYlIzOVc0fmP89Ral1
EdEI9FqbCdaeX3V+o62N9Kwv+8OF7Q2It7/s3J8Hi2osd9oe/fSldv/DPTsI6wPg
8Rs32oysBQ1k6GUVtgR5CL7PHRueg7Rg3mud4jyx1QWzMv/YlKkZ/0cA5BvsDn41
wvxua/NnGryQ4zQ0m+DPujArDyd0OdmxQwwOI28Bip+sWBG2CeinxeXgzyh4V5cm
YuBmp9s6GpVG/+OU2qLQPEfNKk/y74SnHW3rUcTeKGKPss7lFCMK5bYN6DzWwgx6
H0o4zG2/wMi6Wgk60GLgcFxLdhHYk1v6QBPUYmOnuWOVFpYkMS3zgD87w0yQASMo
JZry6b+LIEbOUn4ogtq1HH6wOFyUr+1GGZuT1m+YKlUuaREgZZCYA1bQwMyKJKY+
aGWhs6c45+EEChOjegn6JR/R+7xLN1gBj4nMbfck2mEVwHXNgSnlsVf2pkAJSvrO
MOU96jGb3MkRyiHnA2hEW7RYaBd+y8DtuH/w1eIqssh0ACQCeJ0YKHF7tX2H4rzp
GQRRYpQ8/bTjnkvMIr8Vs39NkuC3/2epoSMKn7gb8uR9jp5LhUJE4b4dCFO3RaY9
bcOpP0hD9nmeaXMOEa4ifKgyQqZEZxXpN8REY+Z6H6Wmo7aBG2SsrlALqhN37Ngd
q4FPNEa6bTCy0+e0TIAkIe036qLMjBRebd/cFUsaK7RMmx6LiMkgtzbDXcYQepuX
oHNRtkzQBZDqzSToSFVC+3pOXckHuLDOH76hCE+gswY9Ps3QeAI4lPcajJEzvDrT
0CaneYJwUQuWPeZVtqN4Roz4fex/iQQpFmPewL8VXyl/2Vq0WJ32xPtRedAvDp5O
4ih+oXbsreC0o+khIa/fN6sXEeb8ts6JKZ6nSaWcDm/U1nLh7qhqdvibwcaUQhye
qTb+8YO8EH2mAYYiN23ju2MohPEIZCeZatdsecLJcry0s1IaW84vKb3492FxGNkD
j1Fwv7fIoP3gh8y2ausvcZ/rKq+z4EMTi9DJ2tXO6eoqVIdg70ovDohU7BEGBOrp
nhAxKgPfMnoOY2nFKCgiXZTpWJJWWYITddU6Lkb+Iutn5CJnrFvPDqFQeXAk1vDu
brQvf/ucsdOhcscjMjJfZG+6OW0nvaode6CFcUWEY0lCZ25Re/poQrBAKv13Joa0
OqXVIFg+357ZeIkaWF9z7Ej/6D6yF7b3fH1A/fzQEHbb5ettisTUPJS2HJi4WOBg
2/LcBPdaasEp0oQReJL/o7RvpqxoUN81xs25eGQQYirJUU83J2kw50FnrGnWobzJ
xda3G+DVHvkfptPAJZpaiyFGs4DFl9RAGEhIjkQqGI+nM5ajWS685kSh21VjfK/N
ztTt2cLqa2jGr91t+blCiIgMod9/rUb8c6PecOOD113xgxL6G1zxMQVLf8isNTfu
93g5sFTVCRZph/HzXvm4ANvHaCjzeJ1hz/YY1les4cemPVoXokg1qLCB5ijBC5wL
uCpMvmjH8Qvlbr55lInT750uoV/XyMTVj1e+Pq9EJd6GYo20Zxpar3ySAFovu9tF
wF+/HrCMuEHY3VdJMsns31v4Ash1DA5J1/HOZUWUw+iGMBV8rWlxtOyWWo5IERze
+EkAEFNVsTHl9K6Qcw8yXF7bqvIYgY8EdHVBf//7FOc0S0JYJMIMFDMZoSlyqPHv
A3ejKiwOkUPvQC8nLJO5H5x+f1cMQdhx7R+rtm0gb7a/vIDha513kQMvXhqBn2yv
bYxdgE3kmc/4qoiwOMmVA4FTI45ezJ8p7DYqZbLDwNvFZhfmvE/QFeuAhIFX9/nK
S3xO94QIl4nOgWgQizyx39dpH8RFKaZVpQo7IaQ2kodSRaRCCFAYaA00U33SnyoU
1z3G76q3eHX7xvTW9Maa8sOx88eDjNABv9vRKAc6zF0wdUNjuXYHq751noiKbkA2
yK5mIIPulE94JpgM/4Cy37L7ik5biguP1wopK40Hv849Ij0XdR94EczMDkrzH2wE
09ELbSA+3+ge0kyOYORzAHBHXI13o7ywyOpL9WTgSYwBsTjTHcjwSNM/LGyexL8H
dA34wKsm05ZgaK3XAGHYLP0nwGNbBkGlCLNDyQSATSfggiNiQzfmxBI1kYWiUcoM
Bu413UfnPI13fI6cwPXB0ezbmk8hlyJKZdzZOSzlJh16TG+9o/xQt25GbTud5I4A
KkhKXnnKjLCQzZLDwUJqzAENPtRsKpw1hFphbJPei+Bj5rC7VLOOAEf7qauOHWkf
H+i6Am01iRNhpDrdHAbpYLXAxovI9yilXT2F35Hlag0RKiRW4aC9w2rdQ6xaewjo
sjaEpf3TT3zKP7Q+78GV3suSuCX29rQwOgLo49KKa2WnHJHTKdAi7QVUHM0UUf72
iqnWQAZQEsl4gwTGRaqRia9+trHwHmFgPKpvSnSmUeDD2CPN4TDAHZ5eDN20eyMd
w808jt++mWw9M+niRIiLId5dC1/8j+qwYtwcetgDq9jAByVpIVb1wTM+lGHXhczh
1Y4zIvZVK3PiQ8rtddLwAZeRHjv7CPleHb1QBxQ/ZKYOF8pIXMxrxUaj4pJugNU2
6wIxApT3KVttxSA/KWQNLa6VA1jHydSijJUy88Eabiwa5grs2XFwXDUJLFG/4Os9
1lm3OjNqT9tWlN6KRkRNw6d0WHabh2/NMSB9653seBXnzt1x/lzQcKVs+XgmqIYw
w7GIoXzxvcleyyQ8TtennixoI2h95394489rFMjiQ7G2XxCyx+2SpXwtnM5OOaNh
L3mupaAMUN5nwwfrZKGluHOxo5uCBD0NKOv5iYUf+vYUrdyEUxjl5FFf5+/Ytip6
yOkhjfPoQVaYj8cP+XUtaeOmAAN7H7Q61nOzoAJRHfklhovFGz1R9GjL2vaglo9K
HhE9tentIFWr45gWFwtz2Q2AVzkAz/dJvkoUPtBu5GtKKbbRSZ9Ks1UPfZpJ5lq4
7SLrL27wu4aFn+r5uXpGXNIJVUmT8S9ZooJBOr/bl119McpNNHrMLiwdqfjY11Rj
SgiEteYdsG3GMY76P1+97f5wcj1DVML4GJfEjIs280wXihs3g/8oIlrU+Z9USf8D
ij2Qi4w3vpJAi7XLCmIkTk/DxAKYzAlaRk3hYTRqq8bxLL7DmLro64f35Pi17qbl
JCAZVpvnjij94VucsJ0O0keKMR40/6HPQR1dSATu8RqNT1bVAlrJXL6PpbfF48N9
9+HDWWvfZA3FwUTfU2yzuNY+NODwdhWnvblJCLXhPOYY54VJu6i4RnWieKOjPCid
dnLh3m/n3qBjJsaQSqLLC3nYep86jv4Zo6TXuPcRVatqdqAwbMpY4/uU2h/YatoX
Bdwb26BFLY17pn/MSXg7H5xShdB/YSniQcu4AkI5+3NW3aMFcj/fgW0Pmol2RJJX
V/zXG6BLkGRabMthwIt2rBqQ3/KdSXIsr+xGUnEcQKP2sUNHxyT8Gz/yNIDa52X8
ZvcxqY4+QHD0uHRGszVW7FAkyu22H4E07s+H8Os2v69GL0riHzQ40MU/SasX2aeV
jxFpd4XT/QcGdR/xkxUevQoHpFCYH6Ow31nGDBOLZ5ZBEbWoQEpGFXbyWLjgQpKG
kqFPvpYC8shijgb/5r0Mlq+/uL6c4J5fHbvKmP1cP1YFDUUjyzP6l7XqWxbBzeYL
GZfjPg4hn8KUOYTd9zu3LyloHLp0mh6oti9pTxS5CAbOex5R1GJ8nheQW5SSXnV9
Ei9Vi3BUqn5Y91S1R+m84qEjuKj7aHXL8KvgY6GNkCwZXR6jqY0GadunHPvFMA0a
caZwoM6jHGgdSz5GJ8DDRR06r/MTm3oW/HL6o+ujojtTyd1ICBzmgFSplnB7FyMx
yzd9+kc+QL1HB5KYiF4w/XqASiQ43fw3A5817huXwSLBM2lANVPUgQycq8/GVfqA
2TIREb4iRVrCEvmACUOqe1Sbn89XWDoA3ZDeiq+MXr0Ur1OLpEeLtJAqzQpzqLAE
IgKfW21iodbQEF1zwDBLoFuoofH4f58XA8OBUTQIQovXLeAUt2hv+jT1ScHTncOr
ihABM4XiPZGsoeOZogiZop1vzShNGxfOrycALCnNFpiQWLpVjF6/RfoGflZnzg/g
MI4F2u23P7PneBHAP9UbhAKUEZC+VV/4Wqc/+Pi+gNcF139xosqYMTVFXIQPuBG+
aROI2//lBozzro/afzY6L9zyni4mxN3BpLKD2IFQZutbujytjX3+/9uSBX7Hqp/k
rVnZJWWeTWaCvbSrfhPx11VFSGtMY8/2TQ0Vwi9WI+iMYfe78CwK0K1hZnqZ9d6e
HCnfIFohk8Ic5YFgwyGQapywpRDSIl8EDwB9tVjVx1lv7GKaY8jvaVDgcUuF4/cP
nOmm5S0J3Mzkp4d46EPkFfc6P11gA/4vPBoiCaUt/Qgl+bUmXOD1a2NAQb6N9zM1
Fx+UTOD9HEL/Ogo0fpMUZ36sp9WcooSsLtOKyeIt7or28RTovfaono1AK52pHjUn
qR+ASG1Nhx488K8nPoaop0m30ZY4WsOTJKshV2B2hJM8XcpORx8UyK/NUCOnEJZy
AYv6bWIIkPhiXzX7ufX/9ElLPpb3riAXIk5DWCnWPghrS5b7vjckRhFNB4fCITbV
mkCW0H3IFangDxNf/BbVn0dWNK3TSyWQ4DDya0ZNIxQwCC9RbQrnEndQNu+eMlwH
lMPzTcy+P1rv2ehjVvtuKroYuj1i3AfrI5X+77UfcxIytVmFA6GkJr57X2DDIyfd
2d5JaW5rFvznbkOe47NueFnV+5sQzarXLFBSWm+QuS08kuKgTTBHURVtcOJQOxxv
yrF901Ri2mz2UCdrK2zCKUNNl4qzFz+n6LSktf91/Imo0/RAvDaggzEIYEvO+N/D
UMSXG/+9lgSSiEsLXOd/q/V2k/0hAqvpAtrxv/pPQWyOmBHq1skfU9JInFBlYiKb
KmCjSC0XL5DaOP9xuqDag1FPG+13zcKEbJjJ0a7eKgKuB2h3fTKVbLHnaVtvW46H
QU4XojKbaIMYwYmP/Kzn9YWXuVkAtKXkdsYe6XGVPPyb9ZolKmDbH1BrY+TcQQsv
Kt5SYRnXuuuZqx9oCuLFYfJ6ejs6kkAwbvF1+mnTnAwnEzh+eO3M4JTXlGq2NGRV
Pds3A5ifKM2JhKNTDUsagO+WzzT2mUDCllFel4G+jlB95upn/BMfXryMd47TBKo9
tc6PASncaEDg2Z5HEhWdfFCizfNOHFkcJVnKEmiyH9ojLzz0KMxD+9Erxa6nf2oE
boy+EQBnxiqY5/Vursi8UMgi9SyA7bAVmnrr8r3uRAow2QRUjbrLgMor/IPCi2nZ
IHFRINweOcSV5UrNAubkD/RKWPtpSIa6RXh4xRDQzg59k8LEy6q8NjBqbrOgKAzg
sPwLRYND3GfWjHo7wxGiqGBFs8dt57bZScJBkKi71YmFHaVOYDTDwM8q9lcQSqMi
R4Qv6FBHJf2xTDtRm8dsdgS2l2l+ZpUuWJ35nkRs6iBT1TGn5tRdEQWWeUC98ABd
3dZyjsZGplP/iQ9X0XR/5tAVt//a1sjMu0nlhOBDXlS9KNJWxBVI77VyExc0DUw0
xM7OaBAVFBBAW0miB+F7h8fK7djKi/Tv4s50nAOfwpYQtzY8NEKRWybqyitCFa2f
l1v3ZNmFpZKnjTsExnRUGxgVLb/JdPm4CMCTyMAB3KUcOyaVJrl2Coqey+3f9eTO
8Hiq5rKVQUZLLJZoNgh+F5YTjrwR7tB7l+Li0Y0wifgDuoNSfFan2E7MwzDjQM9S
Cna4UuC9s6F6vQJUv9r9mxYyBSN6xdSL0BoNu+2FLoPzyV2lbSZRTq0NXgmxef6q
0FqQnjZYZnq40yuWPSDDge2EGbWLEP0VfCdIm5CtDfURFTuaAtP//OSOj3m5olOH
odqVYlZehiRftf3PDKy4aHXYzEJP0TJ2VPub3WfZKHXAlpE/klu7XZvY3hMnSSNo
qjYqQh7fdd5cbCWTnze0Sacm/mzcgHgnqIccr1opKHQE7Z83y85rb4tln5cxY+ak
ZwfYB4S3RkGx1jP858wVyW2/D/YDs5ep9znzBhG001Gk1SKAWNV31E+TS/Ku8aP/
aAblvkJvAJK5L+M9C5YkqmK3kwesJoicsqCG95Syc4lM7vgusWVw7hPgLvEljF2S
tCjvfNXTaVAK9o/10nXQAIrzqCF6ERSBaQwlxMgofYtbRiyfkeYXR+F9Vj22mOEs
jVmjurjLalb6X4nl3ChZ0prgf2Zn8IGK++wraRK3SwXjdMIOpwaJs8B0k6LTlHe/
5RuqUXgprSbT3kh6LnOn5mjFwxSC+Ki8Ohb2Mstu3t9RLeOdyR49XeeFmvwbnsd5
E/u9/lfde77D00uJg9HJeDkEpoAIwZUPhLiMDme+SNBB/uk2N0Gg58KhhVBnt0J2
4PiAzHo6l1ddXLQ1xFULQd7JNYZAHLAPHVFQJqy7a7fn4KNG6ymt/uyR1O52gg+k
0Cmx8ls6nLeoAtciAtzNilR4YGcIHQ/UENZ+SSjx+fh3AhVXlbgmDZgnzoQRgoUE
GcxS1eYiBfEjyW3vYBapwNVuKkogvFVcfjicOB6aioLc0qp3xcVLcWB3D4PFcBss
N8XEw8L2g0Zze6DoCptLM3eetNXXbUVR6Fd65uxDkLkzExr7cVe3etipj5wE5oQp
fuOS4ayx4rIHGBaX1J3sxiRCA0KkeR8fxCy5EbCfsy9ms+YPRVrn/srT9C/4S52m
LdLMy8w2VMhrs03TATjsODqCQru35c1itV1q65kG8Y6kltTa9X+PRLDC8ceFnuBE
8ZWRfXnsodO+O0PkzC2yL+k2uRhtCn3VyxzI5AO0HPAvm7vDLNnizfEbETCc6kdT
CH+CSJ8Ek8nslhrxGV5GxuIh4b5I0zNZ/Ik2YtbrMZQ6fQS1au0SVKSPlqM3fvNe
lMsxR8DXoVeU+dYvccRocPzwyTmtpi+HF49m73LMpZgmTKvt/uIcBv07j1v+/bXF
FPzI1UF267bCfemHDpKEi7sOT1ubWleTuKlSwxEIZ0tlO1wcm3ySBYlVL9hrsjj+
ljep8aMZa4AkFraLzk0hPY229iVEZmTL930kgXjLYOJkVBZzn0L06vp0w2nHnbi1
xWcoMPGreJNdHDIyyui81rAbGSlsO8R57NYcSyGKaHiYutgSTUzpq4wxEOcwKFiX
e+GjLNPI/E2fB9+Tt6YV9VELMRIVMujaY1Xi/Bcee3eQf19aGHbSRv2ccVmk0lDs
nZ8g+LFCBft6D7V4wIRPwSUk8nfTFFrJGrSL9lJf5d82/oESmCZ5BFZYJdIpMMh7
RjYEFLHEIxa+arRaGmYumsvRHJopVWhg/dipaGvZyBTt4h6cyL8VgMMwnU4e/oG7
iJvtUVvhtm50Mc8IXEN1qFr+gkLeXAjefoqFTelYmwu/NSJS7vva4nZs4L3iDtLJ
zW4chaS2e3x2Gl7I652IqtyOLcPSRxnIt2/7H7QOG0OlA++qpcSaDw7GNaJTIP0B
uSVmhRbLaBf6hj/6lQNE7FOOMiRZCZ7q/qtGHxuMaOx4pFTEX3LdQT7T9QmCD/w6
bTIkJ90tg/FL9za5CpOh0DjmAwCkHguEltBUzVhOZxh/ToPUAd75bVT6uRNGYxhj
ORgpMgTnZu1gZryAgQ6oSmONf6HIrXpT2/SyumvGkacNRXs4AmnmufQuVbLi2lrO
qoQPyGCSd0IMDwUdB4bS/hz9ozSVCMuh1WYZuJMbRKUKFXkyuJxLCbZTa61ypPAq
bQR+81AGy1SHMVFHPnfKUUPwHFrQufmLGEFEeundF4sC46y4u0dtnP1n/xmWR1m4
NSKZsBhk0OSsgWZNOR1qQoFEW8N5VxUTw/d2yxPKkn3wsqUDisEMV7UeJ+rTsrxH
LAF1oyy3THjMookLTKBPbxpiqqoyxghTH6PDuZ3Tlyg1BD7SWEFu6pAfEQ2g5Ogu
N6uIok8IHxSzOrvHQMuUvFyQ0V/FBPoTDd+BcSqbYXPUMf6qqgC0QGoQ0poPgu3C
06+3eU7uZqm+RfKHxX9mebSz5QKa1x4uAtAncd27jBXrMPsTAONNUWxteUtUHjO6
dVpJaddfbFcdJLAdWefS/xt3VsbWmEKeD/YRpE3/xfCVdvHtZ/tNdnbsw8SfMVCi
44gZ3V39sPExRXutB1hJ7gwrlLXtrPFr8v5HabatsV0y73Bhw4zpJoYy6ptMmSga
zacofjqbzXJAGNTBQpl/QOJ7NGizNk8Z2/Jgsq8RcW3KaD7kTWrafJGuAuDpqTXX
Z1TTGfWzvdd+M3CiG4cnMommur0zlc7fV/MbDS+JhFyRCeeLKW7iuDfpyc2d3eAB
jT5Vl6tFL30PpF+m1Hoe8Jn66Dkz82sG0BnM1tWaejAwCzlqczDbdZ39Cf8VFSem
ovy0BFOeUdiha40FTvtUdrop9NG9YpGrD2grqNj625H78o5U4ziOOhJ5cmUwTkYb
Bn4bwflSXe3rVa7HtoFTVEQtKnt2oebx/glmiTh09NHdthWaTikIRtK5tq1l0DkQ
Uh76rv5NmnUCjIMSEcXdL70KR6eSmzY0xLiBnfWmx8cCdUq6ZCYs0OAr5dS79E8c
OJgDdKRibeyFhuvXs4tP4jRlBOK2VE/7WCaldhaXTuSUScQLrxj2eacuXWlJHTPy
AV4060gdiVGYCJwMfr14qGSo04gSjuVf+E6Oiy7tpEO5RvrxHQy/tVLh61GVcoZ4
RF9hg0W9+zRgoP33zmA/hvpd7ijlR/vdfYVaDeemNcjwbI5MFfs1/1OGXoF6N5Wg
9nOPPYgH8r2xllOV3glhxgc7Gm89EbwWTIURhhmW32Pq36ubVhE2NLX2y2q0LdLS
7AzrSuF5hT4g9WRbRAz8X4v1RfIgfaq6y13ZplJAnvwlAOm/wqYaMYafd2j2UOkp
c0vDkRBmfxdxMsiFZlADjLiLiTXRqstwKZJVbcU2f52NfuRqqghaIISrAIztg5WA
7iWA7eYx1McNqYh3z4uQKLtSl2QMpjWRqUASByvjU4hSR+/0ir+x9OlFIkRjiWnJ
GG2D5V5qTkNFYbyhH2U82i3KA4XWjcw7WcZ2DgkYvq8gpUwao5YyTA9FteJ5X3b5
16bEGdVxuLHS7hQ9UQ4YRs5g+h9pp4VT0Z7bQ6BRGex9v6TX+SISmhyWqWQ9bmJs
UykbPXyF+AcW60T/sfI3WaXqGeZhmoMBLlrfmcDZIqLPCq8+Wgk6Mb3A/27yBQB1
zPRRJX0duVgyetrha/a0R6rf7NtFVZyJPDUQDafdZMu4bR4NvdArg9MiJognOFen
ELCJtcCsDkgSchychRmD/Z078ek7AGHcC33W/lJ7IczmcK1Zq4tyzzUuwTB9JoQ2
QnHC78FmdNARZp8d8yzcxOg+CSFnPyIGverEdwqm9dNYKsCUQVBGFW9UAuMA7yGl
SwgWSjHA4PAYrduFteSDdvhdKupvlkfUigxVd1NpKoQ1XLRQLYaTKP0kbsL4Nt4p
8/FzmJBrcdjKHyGFpgxmS9GcYANOHKAPqldd3whGtzqXg9dm4fQI6hGDP0BqUrrw
bsPePJcpf3wF+hKjd7XDA+0GNr8oW7fQ1rlAC6alxlrphCwmRFNgzSOTtcX9cuyK
57Y1b4y/EUSXaZi9esX3tmJsNyb4b+W1c5gd6J8TM3+SZnufwKxKfweKTM7Rxef8
0J2MI+3i+PrzihUwcNv0w4BejRavA/t9FBCxatlHFHB47rCtp4A/AbjOAffXh+yy
LZRpXKHFN0hSNMq0tzvhQJeMDlmwSsFbgSIX+KYLNckXBfYePm+QaTvNPTAERx/s
eWULrzxHioCW9dZUtTabnQN90jDwZ4KxsZq8oPWE6jJV70/wGXrmofEOUss3k8eb
hGMCWWCu/m5cQ7ha9L8ZFe0jhDVzejrLR2FsdXhtSssutOyulfmI/IMVjKuzgIEv
aXydoVwyD1drrNpoqP+WsYtTn2pHhOXbn9Cn1Raj5yTa8EcT03qupJ/2HaWt427B
Y7esEpe3uXGON+koLu3ykaF10nCkmu6nS+8PwEWewdop/g6ikhAmEETnwFdFE4/l
h/wbZrEgm5qUeiCSYqJFIC0de+Xro7yL4NIFljjLw+38avV/8S4ZV7JpM3LGHDyN
lhS9cW9PqzMlgnf7/y/9Z4OhdZk+pyzaYezx4xC/U82Rq+gBGfJJONUNMK+kQn2+
Cy7lcVyZXqTsAhx5uwpnpVAVgqb6inVVwDc78Zmr6OASk5pXxPzDIQy6A60Hzl8A
NE32BsQvwc9uWnCzfTPqNLGTNCQqK2FVWDJ47IbHzB6pEQBCpX+Tw6I6YPozlNfn
q8/I2GGnFzvPxmg6W9x5UvRHw2hp2kKGy/N9Wui4P/nzHVi1i+KvZq6GNb64Ddzm
gK1DXofic8hVKm+Fsz39ewsRLlVOXgEaAD0IxLNxAB22+PChILPkw7Pgcd80ImkC
P7VGaCtpOAqjjTPtnKV9zyPUKo9hZYtvs3U0juEjxsrvkWS8Ez2RkbUOlweAFdTz
HZDcFRgRX2TzXHpCIMzn2nAJZDMkxmsmtxczfQ23tq3ynlgsa1ksCGPKfKEcpk7h
Gi/cu3mPw9Jfgxc7VnPnhrUGgS0b5LownYWx2zjAw8+p425xlPMMurnCMI4YS3/F
YH8p6cn+2tj0nMLCNDqtjzdNSW/SGn/KrmUUPr235kGkfVhuLjnH2V3F10hjBFBN
Bo7NklTYojgKBPRfVeo34j4HRQyjpw+aYtWnkQlIhaaPCvePnSSEI7wzLksEdJId
Bzfd2dM7KftjavOM18nvdKarUu+QqdDvCTVHdi7yw6GvV7uoVh28kKvxaenM1oXn
RKjm1KTWnpylTg2q95FoE+dhrECMucnl9lbk+w0XX1txtU/+Yj32G12fh1CRl7So
hEuiUngMmQocOX3sC045H1DuJ/fUPLTadukdIiQ/KVWe16pUzAqSvMI5f5w9VthQ
r32l1BzCcy5Xz9Xjz++LQAKw5buHT3T3jxN1KawCA2Plj83bbWZ9decKFI4pLesf
wKukrEW9VvPvu9D/JQJfSGvfVnZNjLJal6dClFbq/rf2w6ZexMfc3pVwunxCY6Gp
lL0fye6EFl8aedZnB+BLtuyK0123SovLlF5A+mOI51TRX4NvLen3za5+bXhfm2Ia
uJ2IUCnoLSdwGRqdBCKuJJNroOpTgIjVKDDTERaI04e7phunQuSSoMe/2XtJpybS
w+wb3O+fPsl1R007AM4jPwsRsYlsSxqMscFPSwr/hlbij3I8jGlrPVCpa6eJqLRy
McYIEXSD1eC3/kJnhCRq5C278uk+cfF6Lcnz+Cq5AaVmdC7kJd1ugzF/KfXY3eM1
MvLsSqxDPNlkhdd69qCGwIVrjyt9T9pVHJ81g5+aC3vvve5ggfvekYTc8LBngDLD
Uon8WZDAXaIZK47iR7i9C+ILECzOpDKS0106GIjnBHUyF+QCoCduPohu/t3QoSCU
gi+7FWEf29hzLyigvvGYRZ7KWz/FD/GYezGMBLiL1miK6Txu4nIKVEKLMbscAfCk
utCK0i26XslISRM6PELyFyhxZoz6itnuYcGfizBkFQ0fcOufY8v0yTcS9gwZTDvW
4PGSECw/sUms70/TR7LhWlsa1rYw0sJ7NvwPNHrtEiOOJhIhQzrQHLHY/EZq+Np6
/1hH3ku0d4eaICTZ2uj3p1M0nSHdtXHxTECmNhagLqJqVRZNlJN4gRPEhhqW5Ekp
p/Oc51pnftXYtE4hQr8NCSSvMTAZF/8P316MdYrnwsiiuOB2I77ruls5pIm11mRI
PwqeVSqDRHopEnT/6ZaZgx5y/oX8rFvjhJTzKvFOI0tLKEH0bqkTbmTrOLwp9cvE
xScGQYszQqHmUKm+TLiDz/oVy2D2iwuPlUq4QiWyzMUErfRlHL142AynpiKajyf1
hLHmjF2rSjEeHQqrUmby86ck0MZ9y3e1/39eIH1LLyoLZ8L1wfPTPPntcXXVHHcp
2sZtgAZR/N0Of5o9m3+BrhTNpST3+0DScB+82IfdUkLD3EcgjOyc0yl8zdBeQgcz
HkwC3CgN130tdmwzGGhpiAhRAnfdbaUWxKGPRGJpPzmOqkOdiooeLx4/FCP97t7l
EEiYufBLuguTIfDSv8ZR7jc5nrZUj1kIrSG44HCL3IHvCPaomB3ttwNQMMQRAeWo
vuCoNp0Jq4pg7CfzU4/86cWTLH+F9QGHd7HN1DFjDJaQpGLgssc0XWohBDixhX3z
LeGRNgv3dCNb4VQrph1eqFnibe5v9jMCYgzTdJTV1qJXS82VN8lCzIUmnQH4n6iB
glYZHLnm+2+u+anVmvGAALX3EOAmfpQo5wRv39dBx0IjiUHhFbJNDqbyikPrItOo
vDO5mLp/3eL44x/IhDygk5hZP2WMgL7ygCLlOsvsR1e5FHzkLFVEvhyYEh9zdy9S
0nbOr9ppJHmX76bwbwhPfEFvxzKGUVpVcaSPQAQgS3Rgt+jMEnAZaPvg9lQPrNao
9+AQJp7uiXVd5ykAHhhibdr1Cc8CkloG4gWJ53k5srWUFrNBNCHaSGRYHKJdHCju
dh7FMu6/QErLtKt2D/jq5U+D3kGfUp2bZyLcc8GGXq0a6Ft6omXyY004RmkU05f1
JtBb7+wSukSNw2D/wW1QSTcWJoWIQ267Y5nvE3+rq3ggL9mST08SWcqmLKFHntMx
OOdE+Zq/uG8iw3gMN+wVSvXv1K0rESrZL7lthRA2CEqhx/kmI4PQ+refcyOGaYKT
5HU9oHav7GLzJurUiVTL25TiVFoUXOIqyDdUNhaNc0Yc5SHQm+18yXFmUN2cPMXr
DyhvsTFXWV8rot+mPWdJ/QRVXEXwi4nQHYko5qKxz4l1ZNk1uL3OK3DoFVyu9sxf
pNXnjsTwIJXBo+aiY0LnSAsWUR/PNZboWfxmGl8U8TYLnLIMZg2NtFVP9NmkOqn0
+SsDm+FBbIHJigBUQwAwyKOJDggVOHzmchxnpgbbBLUNMBAkSwAWFBa0Sa4SXgs9
C+pvEkC7PKj4DFdbtssTM+xMoSghV+C50yI+X/3frgVKPtAEjoJvFNTfFF1t1KLz
F+Bg2zWs+yB9yJGTlT+xisab8ByRCL/Kj7+pEyqd0AUyP01y8aBnoBnFIGaAI6Bl
tXUgR8MfyPZJgc6CTiwNC34AYldS8hxAdEMvFB7uGKwjWsQbfromr1ra8KBPdQSf
SXhkQSlzjoMqGgZgnb0WLWZJfFbv4vTaZk1Oy8QwNwPcjelMzmqCBHRCgIeTfT8A
Mx94pzvOguk4REpYroVZxheslb1/CWBQe3aLgwxsXBUz6WH5jxS9eB0CGe09a4Od
cpEMZpenL9b8SP1oVvLd/sLox1XwVDsGUmgRcD45HRBdyYC3veXIIB3sv5wQoIFj
A1SWQnkwzVngJgrWKXUXEqdxm4IzPkcXBs0Z5STyNhqZqqztEpmVNsCcOU24v04i
LZ3G99mcHDw5p+kxMz6amX22JNcUQg4K7c5hObXxeBhZwCBzH5tnRjkjOdtp5PGA
7mB1PMz46WXxyLUegIvEcm962KZ16/BtC4H4mIr2P9OGsPkC/OPETCl7ve/ViQ0U
/rjMWBECkW35ZhLEfmdsOdpCBC8tYbghAjTEnFuAeaFiUbcvqYHy2v2o4JwwgIlg
il62ShXFTc067/mXu62GE1/7NvRzfm8ivlf+jP7A1GuOIgEy+52cjpWAzk/IvzU8
x9FLpWtO0I23lCR7B4tlokBGcWs83PailAu3FBLMXPapU2Sf0rzy/v8UcOiSRKbs
HqrMnopE9uXp+VMWTbuG4/FrbRgDD7HdLL/vrHzvUMtfGcuFTP1egTuuBHI0p8XM
Zg3WVZyo4RsTfSEVQmzbAP8buND2RJjBpqTH6xj9Gj0SjBELHhzryd32E7sH/J8E
jVGK4zrCbOajhsbNF7LQk0N9RSfGWfTVTz8UU9BGzjQfBZfFhqEB2sD0i/DDYDbK
8zdFtNaKvdJ3aL5LZ1rAJ24iM3zqmd96DldTtEJE2ljolOz6AnYYKjSoOn8rrNGc
k9sVb3rN+ZHPD4x6j+bExvVIzCStl9twlQYbEAuDaSnOHLjZIGmlYU1tkf/nnrDb
t19OAptXfjDLdhqVGYkc11icTTpwc34ILFvtiebpjAu+/KpwUjFu8XYNgQEbgHe4
cCR8VkSULiJxO+B8U85+IvNx9qxvQ4X20c/R371peck9Y9xRASrMZw83VFTJzSrK
fuBeGxR0b+RYJdcn2zcpITiycRRj/8JaOIlQ5LJswoufRh2V/bhju7av6uTd7Zxp
mRruY/xsLTq1Yhgpnca3r9H+lbX9lHxsZkXkU0CBxp5Xegb/EVrWPsi1w5KFHD7/
YXWqW4rVEgUEX73FBgPtkvzJGSsNPGjUQFSQZmxG8fkoxTYjZ6/ezsRdf1ZvKiNc
PLzC2c8zA2uaNi0akwezXCpW737+9wrvL8C6g3PpQYMinuZr2bYDAb0MHSUAvqnZ
OoanblK0d5t0KqnfN/zAciwE2NNArl9T/5gi9/bT7FP2xnEBtWbgN+qyLhCbH+yA
UsqDrhSlrqBzCxP3ov8+706IVy17Kv0LMa0rNW+KP5UEjJwkV/cuWUcEGW2Uc3BL
1MI/Bqjs6CM6VlKemepiW6UJDtj8wS3lmwH2yCtdt9VhBIeQv+0PUy857K5eVtaq
wNvgc0Mt+QSUxGjvNhaVJIPIf0o8WxlzV+Mmknj9qpfl2T6zBmrlKkd2JN0fbww2
GD+X5Et7MPPlLMWt+LpQiePhGjvRIBX/x9eNY4Vu7sU2QyxkiAY+wr91pez3Bh1u
/AZHDrfq7cNH03ExtHsqqr59P/EXiY8xXF8249zlvd2GDXkIukwkrgE22wCF1nYP
iqkQsb29HC7APfw4Rn9I/eD+yT6tTX36LnU07ecAPC38HebwpYSetgjbDmRwe1+8
oKAcunI3cEFS0TQAguild3vulaS1OXBwYcrtZ4CG7MvKhe/fVcoWyj6WctKKmJS3
RVq2sdEMyJTSP/JKa0VMJ0RI0bG27rncBkSO6VuAYlKzTWN2B6wZ/dKSP2Sc+ae6
kuQCbdFnKaMdUInNyPU5Y1T2J+yiU5+V7YsIgQAgCXd/Hgjc4POaWT3dBsT0WEYd
ArVXkwNtxdeABuqofkigO+N8j8FcEWEeL8/5KEL7+s+gpbGvaI5wVY+xpXVnlSUE
ySUhqR2XsxiQVqgR1Fkgojt+fx57GjlN9fRUe9gMLiKDo67U+Gw0nVp5na9eWtmi
3CmDSyR5xLG0Rflpk6K+ePNb5pcI7cZBoNyBIEMxoY6k6irz6vp87aNClXesBOo9
6VIkmX501oCclazo9rYbgfz60lZn1KazgVK8oW2Rsidz1n5/GwUvJkoq5apFQajj
yr6UJ7PKGNn76FcqdfW89s4ic848/MLsgIpZssljvbZm9d7nNSxrvR+fapXn3+KG
51Xg+U6XB8BFCALAOY+iyM9kfO/Pi5BS2az15ipgNQL3W13z++J/E9hKnii0EcOO
R7nDW+uhkORk9fsSXhsk6HsABnl2khS7nFIPUvc6oMLjNfBFYb3L9/RTPHX5gYCV
Whv5muLQF3GG04XLncF5MDyxJTL0OEA5wdujYgfZpd2X2XWOVN7Hc2d+2IIxKklW
k1DMd753swmr5W/PVUAlBlplO06tCmlleK4gzOjmqCDFjoaK1d+nvNIe6YXJ0DWi
I+IrjLz9VenyAXPE9xCererjBMmjttdiRTWT9Dn9eI1NLopZCl33zR4AxlHk5nd+
e48VNKSDBO6JJvnTV2NBgGGRiVVzo3fYsivDMygUHQYtZQqg2ULHxTVe9nT5XbdM
QfHa+cGFMLpVkjo/VFZP7GqKz3WQkQGtna3KqxDWTh8Ap4VXowRJhhL+9M6YclPQ
vB/g6yoeEPnvBAhMW9h/ftWvnbFsBVO64DBdedQkXuCGdLhWM+F7BCLi+trmxQo7
uN/fnSBrZHzAfDHpQIPkjKsXmR83TQgSTx7L3LolLZqQJzf717VWJynkgHWwhAPM
FSthcbBdKvRF9NdhenMzhkX0j4uAueJRetotKEkvHi38Zb8cUjiWm8fRAcykYcIs
ooMZkKXUG5asYEi0Zj8MK25WLHbaRYzE7boAJtyMKswc6NsbJz1dBRlj4BBAmMAK
pemAmj2CNpKlOHbdeQ1+NKVRgSkbNidjkTNuCO2vOTIsnt4KG0spaApUdurLuZ7O
hJInS9NnUGQA/tN1fGN5xjfw/dXIFWPto6fOhh9qJrHSR24RNeKVKg7rZCXzQGfj
8ctvb/6yKUej97DC1OQnFlKHkhJHqoasMF1Kila2kKXqt7oRVkEQVSuBsuo5JI10
IgE+Woj9xShcCJugH7f8t4lqSvxNTgPp8lPQGCAG66gzPJ6Y3+2h8HEyDEDblzap
rFeMNsl4hPMaP5eoo+b5360hdT44/U+AS/kTa7619XJhKrSKNeKb0HQD12cph9hV
glqV+FV7lxXqLHgTHXMXOiOFxSPGxfb9OeaPizUeNcPYyLInuPB3YWhs0xwbPQhJ
09VHyzlH61f0xUJlRgn61FvZ2aH3IhXJZqqQ7Hyv07Tr7EoR7SOD15YSwbSeiTb9
c927A5D3NdPn+bWbruBvXgWDiJfN4MoSNK0F0CIT44y8F+DxHQYgs6/u8f4IO7i1
bXwkDlyqEFEpO3NUp87pHWDYDm0Cq9Aacez6NTDyf92XbTKIAANkvf71e7TiKpNf
TLNTZ76tOwtvgwmzveJqkRAUYZbZd5qNrAzR2QDyTtDjMzWu4RgFXT9U1j0zYDBF
AzdQ/8dQWbXE5baFrU80olR+tUKLOMQgixGBBNGQSrasOg0lRaADaHEBr1X85EMg
ndqjIvZAumQz9hcHpMgmc5JkKwjpwKzLNtGghgsjCpXaOiIgsL4flM27WMsQSZAo
V2fIOqyyV4Uv20tCTTVIPuu3N4e4FlkhyUgcrNAiqUaZFwh06PvHuA/cRGmytBRJ
j9Nq7mRR/o/VyH06Bd/FZFp7VM2RRlfAQwsBJKE9Wsoyp7N6GrUh5Wal3+pvjTn5
nNauTUItStwCkIng89cLrvEXoN8q1vW18jfYzs81rwRRRvuZ/jpCVCpCcTk9+8w+
RJgx6MD8JqnoVeGkOXlT+DovmRDUjyooTzuX3CBZVxKntRSsB7oeegS7XsL/dBmg
Bz52wh4aEY9H8IcWXREXZOtiKvSE/ncvmpufq6tYUx2LFFz/ppOzAALrA3pQNmwJ
Zr+O32AnuxfzWTXplQPwy+sGcmS8l3uHGVojCksz8GnhAJlSA4YeS5eiY70ek55i
SaC9G7JuldpEqTTwY2xlHbctE8XvPgBsyjzN4N0hjuETek4oLEACfE9lCqLIScCQ
LWYib1zImWPmw2hoqH8A4V/1JD21Y0HS6AWvP391MRC6EGdnBvyUSlzk4aCxB1a7
11M1eT+EbLE+UzupmgFAs14/UMHI71lCaRnDj4OVSCDd26UMOhLCah3OYpAgliTF
+14mwVSWU3FIpCDgGRy8J62TmknjUuTGXAi6o9mYImaeIbmpo705b52O58dBie/P
ehDaWHKiw73djfdfAZxk03ePJKpRtR7d5KHu7I/83WQhoS5GD4II4hqxEVWeAgg6
B3AsHAko0f3eiWPEuPM+T0GnAft4Gk11+NSwiyHAr6FZqTsoN6+o+ujzhNeosg3G
dyJKCFv5aoanakSv2Hw1HhMVqk3rp0LGt9dzrT6CojrkLfxQPiMGeuN/gj0d84AN
tfa7usj2i7cqx0ny47lJY5vI++GNj+LT3bqUbBvsFRCRc0MDWB3RE5G5v38ADNsr
QTq41+gipvDhRh4fwslNrEnhTTqOkY59GcGc2H8zuJo8Xo/NUcN8duCMXUhEr3PI
mnKHVlyXQOcRrgk2YtNgeTgR1yuzp1CHZ6FXYM3Je3HP/oivj6MBfgXv+9PW90wx
PQ0JsrQ6WBQFIJExa3E8S1c90OeTOvPgpBXl/SatZq+dPkp9xeJMHNOSyVKc+xP7
cr8ho4ppXdmfj9lNeHVGMuPXk2yP7wWGnR+qeP3v63vGkSqKqSsg8cy8oYhmvUdW
lsS64t1OJRNOA7eziWcYuWJpZ4hUYyu3BiGSXm0vMOO9NA+TAZqGuk+/rmQEVzUi
ofY+PWlIeIXvLgumQwT4OtvE3cr2Ig7Z/HhghjcBFRXJ5jBtd9y0eDLDjxiPMb7X
Pm6+bBDWL6O9HDyeg1ppgSkmGU2bUgOSDqUFESKvjN7glG4z9YHCREzBeQbGadHU
vgZjhjTNiMS6S7G7hmibHHs/aI1OLZJIfBzAyKK13NfZmKdCPJA5IPL2vSjLwi5i
zgKapX7hUmLEDc56f0a6iZiVNQ/e7hZqkcyjX7G+hsIyj/q41cDXUVycE5/sn8eS
OMJkAMIfcmMVVfZBZH3mvHlIjajpL2AxfWlUAqhqS4JSCQBprrzWCBI3ymK0lBXE
4jqTgdL4LXr3033EwKnQLdMEImjVEVu5GA1DILEYdPYsoQpx24fpdzw1+jNKyRIr
F5gtTq6ZBdGfafGy2baF571iHEl7o6OvY8M1UVEVkXlzY431sYw2eg6Tr8/pjWWu
HaBHU+y4XfD9KggqkLiV5wDiXkbRepvP3WNyCn4UYF5hFz+RhChNb7naA7WYMLWC
qDyV+6bZtLvCoWscGzro0h2T0PDC/O0YOW0j4tUML9UqEYkIHs2ngt7EJkwY0yVu
c8MiJ5PLVr/lkg70j69XK5Fagzgza6U4b6Ybh8uG88O5keKFcP2ke/dE/ChSAgBs
Cq89/WAoRXmI6LvDK0oWCx6irZSdtFJ+gpVnB+5Mns51mQ4SKBWxfP6FEsy4OGjj
qzCmjZO8wVSg3gK9vDemulYUuRpwBoRnwTZlqtp+HHi3hkIsRNZLXg+sX1nrBMi9
GrOu6og0yLpqehNn54a1pjEFQA68qhGgnG9vXhdLwRq5IA51eU8YrR2ryv8fFrdW
b813rZ5wiGVmb6EK+FntuOZd4ay0FNdmfPdBLaGFKLsH14o5smsGU5zTcEUxstlh
zWzJLWdVkd+NDrNUuwoFlUWme87PSg+suEAGTii1w75XP+eTLB288yRQSxYo3BlN
NYFPPgbagehCPAn7Qa+Oa0MstgBD5iTqqwrSKNn//eB6JXWUsSVhnymaMHA8/dSy
GXLBKQhNifLiVWmvIyT9cvegeJLTUq5ML5uwLuhpnjbFsSsaqR7kFYNzKghBGxH1
jTZzX1LaV2VjMpgjMdzZfYS3QSLMldeVMZifudBaxWA+APgKG3sbawWwf4vnznFD
x2Dr5apc1R1LBc/UE1+teHpYVyr0HlpVlKJeOss0iIYghtvOW1qJvQvEC49LJiBf
aIhC5kjxo69cIILfQY3j2p9wImQRGZJCaMFRe8fafZilOR+qsyO57RDGDglz4+Gq
ZCeo0I98GVMvf3SABtnlp5qS3fBSTU4rel7hpcqOz6bGDL7xVJ4zhiOETC4gJOit
FAB6KNoS2mn+y/Q10o9laotfG27Zv/bGfHbOgOBl+az169lLc1oorGVshtUfQIvL
218lp+0XHA81viR80f/ZKp+8wcmq8jQSp9bc59cI398svDsvglRElFvCV/701OFU
13HRgcW+WvvWToyh5vIuvcZa0dxRGieEYAwZq6Wzr9D8uUjUXry9F+zc17LR/5VQ
czj8EHBIox/PBriK7M7+QuAz93VvmUYy9hts72xG6kn6z7+nw8ApOmuKJ/VNoSVF
/fDN0nVivIa6zhbnT1LpNfXLo/SCukJv2UvMPuWAYcTjFfzyo2Y3/4pgTXtbU0+G
JJoWGN5W1tLWPh5TuWFmlOb34OWvcosZEj9ezqktqFht1+/EySFi5kIyoc6AEZGG
n/fGMu4s5aK7u0wwbiZLHfw62KMkSFWl/ZxwKDKb9uLLxr4tw0wEu861qBXHZ/3d
a8Ctiyr8XGyB9xrj3UJj0jFPoK+0BCvyiffB2xO+RdsdnLBTUP8I15TjMtEoQSyk
lNMCdCKPmmtGwRhci305VO4OyUGwkXinfKcEQID54GYiShohiHRrDP4mqnZ7kR/C
fiRkTt+KHiFSYKn67aSZC/7liq36vlqWckXibKvOa440x9eCA4pVUcR0SlzNHaTN
UmlAklIffZM7aV0GYOy9EPl0oEfIy9n0BbzOb/T4O4cMzsG6uoZ9qpjxsmlj2mCD
rJ6ejNdjJKjprs/dTqxTGncPYZI4IkL+SZtHnLtxhOwak7QpHFEvfsRniSm/Vbvn
INMjd2OG0/JGon999w/LZXPfvS+1KBi41a3mLC2c25hSgh8+UHiM+AOcnb5iSAP8
vkhnAivP4cF+HNrrccMgDfBb66MABO7ZNYoWqzh2NMlyqzPcRzKOG1r5SljdmFwj
lrkbXjU/g2Nam8G/UJbJgu5bt0lTKBC2csezpHAT+TkEV88JuRZeeoXFpmNL0pLF
VgXvA5++3ldqMSda4p0BjuZPE9Ix/yxbRc2Q3NLQViqzoUFTC/dgy+DpK+jXv+gz
UDHOirqjdDdagwdje1EnZUVRM8Za3Dd047hGiaPiehqQRmrMMNlBiz0bkEU4zBD+
zSDp0XuGIJF/LwSO+KULhkTp+hdrYnMGizMr3PE787NS5SL64+RMtfMk0AAy8vQd
n8trnzC/NeCniWNdFqkuveGJR+49gFlRAGSC9dxl56KbHnfc/AQAgFcM/ArEBz9h
6ci2TgZeptOxU3v2MLYRrY8MuX0koeQnvafJO1vhn/Srelprk9iCONfpqhpb1FLe
5WBrxRG2d5RIYTBzsNq1jBqiInyom1mvNCABuk10Tvkdxi4+KnnH7oQ+rMm6Fihm
PE7MqnwyP8STjcofh7DLD7BWBVhpaEIZmv8Q9oeiEi5F7tjtAjKxD61fw4xJZ4lF
ojpoSFQIC0ycrWjUEfOwvb7W8rn96Gkv5yRBpW5Q3yibZVoc1i0z1n0oQ2Ku/1Pn
QGYp+GRYM3XPHQ1VgJk/yBpZ39lx4B2TFMWG3T4KDBXtj7t6x8/Wv2rFrA5HZ5/E
z7l5TqwCQFbi8/GU/3J1eDC5qj2/hhRrACZmeymGrB6gLxB9b3O/y6VHREyQ9b9X
U/y/fw0kG6PAEF1C3kNEGCF2aMoh6qvlI4xeahOImlNzVLcQO2/JHkp3AjjO1wMI
wvS9FtnI/tG5olDcBNhrqnHqfraX1iREVP/zL8BfhRmwTV2ufwMbHJ49HuwdruB0
s3y5wvn2TzijqqYhJOheKK3azW+L/VwK7co63nsbCJysoucNCs2ddTM3vU35/vw3
vIMICoiGrjUnlQPG8FvW+1xLwW6XE3/6v4S7UuEdFHqLmH4f4S6WbezffRzjIkm4
RmwC3Tgj62VoYW+O10cEvtYKF/iKSAVTCohmaeULIKJXoiQt+SMGNLOGypPYnV6K
9bqfojgdDYtdoa1Cx/5a7nXhaKzCQOpUZ+lVR0lNEvOi9rcow+YiKw3y/IkdbQ0G
g1h++p1WsCyrSlsJHVo06umYxUPHEA/6WDLcF3SiLRHA7o76NM702b0qRFzkrqgU
U35UFnXieFMGE+6SyUP9lj/mxBqWFxrmuCh9IIDzozsunpd6CRlH4n6VFUJ54BJL
OHyJgzLDDynBorhGlsPI9i4oVpFrlhrPsOsIKs2Q+HGmMiqEJgCnVceWMPDcC/PS
BwlcanMqgupAEan0+B2dJ45uYXjwYQt0qWGZ879nZYvsb5WxX3EekvGqnsRWFLtQ
yooKi1OqaBnhkRIXUEn26n0qAKs7jlzcWP+cmxoZUeiXy77R8/7bKNHSUHa0aLFf
q7/l++Ysp7FJuTwE2yB4gZKKKOgEno5i6xZTYeicIG3Rvs+QNZCNv9zt0Wz2D/PF
Unj/DBwaYEwtBwbIeS7UQ7d79NHYZ63Dh2kJmqk7sdavA+6+PvoCmcB/Cuj2eejN
1DcdXEyWRS0V3TEsmezuFznvI2NvytzE2WjlTsk0VoURoaqcpXbQIXK1XHkQwnG2
VtD7s8ypTUKlqjMInqF0Hck8QNDVEQ+aJp8DfZjxVNO/+1tbfuI6nOvmeYoU7fT4
5fPuTJQKkKCU3CFq91PH33juBkBhGpOlqGQ0QZRYKw/lqFPOxO6Fw4gLj64p/7sO
50dYlsvBSt/cmZ+167qk3xatfvVuJ/ie2aDC6PGunQV/W1g/qBBCDGh84w0d2a/k
BHaFozQbisOOrfgJQkd/XWwrWYZmrSzKB5PEf0w8mm86KtxRujTjIsaHk7MMF1QH
Z34HkqTJHVqnNyfePs/7JmXjVS8UI4HPlQnpMs+0p36VYVBHV2pQgvmkxZYerMVH
QgRJKSj144q5yGCr9Uw/rn4OFxX8iAcFUp4t8d1+A32roIZRGtAMZpIpKPyWlnK9
viZayU7XRtkEvXxfzk51ofOhpz5Gr1j8yvDLkNncR82SS9a7Vg0JDhJivXCBvnmd
pV2OZEr2M/LUioWb4cDjRFZZ/qWW+zOCaK+bUV9k8N0Wd/PZ9cp8ixzfCXmFgBH5
nzegy/g7JsFu792oVwhkKwd47lLeGJM7TFNHFyHmCt7UdMABYug8dfc6lJIy5qwO
zb7Uk+aBGBxxcxcmwpUQwRTYMNvmvvAnzqRbnmFodJGPb80eozCF3bi5zwKTiYxi
tuJ56lX3lPYsun15cUYYmFX5KzJoi5H9ybkz2IPFpO6qnM8Vtzwj2AxOoZKJTeUU
94KS/FmE9LSYd8R/0OVDjjrvlxguzuKOgGt1oYSxHvwtlySV1vnF3xUP9n5AJfz1
9GsXuxSLDKaqeyA3fGTQtDWiF14SmItbOq0i5cGc6e2ZYd6eke3P+bB8XGuOH+pJ
afyTI6P7JkFyUbl759H//Zu5phPfJoBNhbhubFaTyZpLZeU+hee87po1Rf0OhkbB
bwosyIpTCRmI4kZnGl7/MpuAhfP6aUhBiwGihX9GJOq14XAARnCTq7DgQPGhoWE6
9x6zVMf/B98eZKFBhg0ah+4L8Dqx6E/VNTK45DyR04Md38mPEUOViXdze9YQhqC7
X42ZGxor64r7fBEGJhXn43FixULsRnNUa1DGA5LFYN846/+B3F0UesZUPCNlEww5
Op0Fp6z7t9H1zWV9g7eZJFL1Qe3IvBKsiVSkqp6SFlYZJsaMIwgTZsS2wcbi+g1V
2EFgzF4M0I4u57zNmkwTU10bV51yYK1RNn5jI0LNuAH8wtCqHX9W+oEl4vBpb16b
vrt2wCVub86eccaV3t1i3jMoOaGYejzoWq+UEc0p6ggrbvGzWVjq6uWOT+tVhUwJ
kDDe/vcg/iQ10xOi6ZqwSk440ZZV6sFJJkLo2cepgPCkoVhqdzAURBCfTmEVSj51
/kiRPGPLtvGeKM3fuPRrq4q7uro2CnVaFQATd2u5+H7qPQiMaDR1G+dRQZlYmbpC
5ve2Oc4h+GIlemnnk1nYM9siCC5WxRZr47ShzNJpgDaJO4sFTEObRqWKtqtX8FCH
WH6ga8bRagpOaovsX4Kf3BxR0EJZhEvOnzHPwB+GWFqJQyLzT93xF6aFpXjD8lOZ
p6CPztBLs/HynlBRCPGMitKZNa/mqG6P0N5VyhVUAJVeVsXF6OLxpOGAVcvyG+Qu
uAzdC3KGS6E+cLQyVYhEUZIMcCGw0nl4FKAJC8hbcf+KoTgn4zpMvxqxroLwQVep
pBTLk+EHpiK+1OMRwUpGHeeQNbV8wVR/pVK5XNTtc0ty0Ra+f/uVQPmgnYeN0HWD
aE3+cAwnmMn0QCfUyDNgXx+GOgSMYME0gA1JhV+tEW3nI3S4vgViNYIwtu14r+va
iKUONekAQ/xIRv8VV69wS8At53+mmJRXoYuei6IJ9sHJuPgswk+ZWHFfFkbEg7Rh
Mh9lwazRYAyrde7hqWvAnxPMLZg4jqXZuDt68BHdjMG+I4oshdk5JCf4Artey7Zj
2tAfw4k4WeFELDSYezFcUI6n2OsyTafJ608WjXOBAbVXC47heR9RRDFwewceVPD3
ZpvVo3g77a8c/Gub9bXGx4ESQur546f5I03pMX0YfIvlvalYC3pEPZ7OyBZ7VncN
saYryQfr2SFVyVz/AOPqC8xK/x5eHoHfFXre+yJK8CltHdKUAKE44No+8Acw6iRb
nybvgQUD+O+nLHVlJRSe/j7hOC3gKyGOXUl0V63MxfCj5+mj9yADcSXAqaXAulyh
yr+7xGkmyQVzroc+5iCrNaTcLReRTE2tRK7pPDFjAT/HLftQa/nmSmDMyL/ILnHW
AdRCDOaY4q3gtuZUhwzhCyMrYSJ5JOiB3pFhU1Y/IEHz7OVvfMgfub7ffuOu0+H+
+mE0UYa0M88VTEJtDdiRqjbEPB7xZqDiY7T+ECLzlpXW21iplDxdvvFzc/y6Idkv
ZVWa/mGw6GvsFipm464XCaSyBYyFiGY4CRq6wog34AsMutS/5PyUVFUhntu3+KVI
fdBWt6XnCkwZNhlyRLhlX42/kqZmAifhezkb44slyA94Ox0Mfnd0/jUCeWm+cCmd
7a8YRzEi8bR3rRGaSgScn6ckunmWdkYrg5D9O9EbvCaYIYspFbOcPPBcmk7YQ8NU
Ifdv03FCvmIufKhqe3cOQcSLa9P8pqo5uzbgT/fTvSmZLZXSaEPm9h79pedRGeFN
ZmO46bb8RQPSugh3chxC47Nzo59UBPAqOWd9+IwrHW7lP3yyP/S9d205C8WzKnUQ
tM/19lqahlB2kzIacClT73PSlKI6u8s1b4cJuzD/8+Rt2mzSSggzFdSxg7hzyOGu
VfBSKEYwOMwfQ+Mpbzmjz/USD+nKhWgqeaE2D072a3WrHfEyEYntecw1rzNl9iHP
Wk0j5ujymQDWcFtU31LNKOB1ygVbZlbXKXQliiOoXnfvZHjpLYXs9uydxZKnJUQJ
a37Xj43yl7JafVuM0KAJsjqtlMFcZJI4dwne45ZiCw3S072YJtwAvfzkVxfue0Zb
m5OsXTWo/xz9/Ri5U7WglvVE/fqNd9icXhGbv9Sqmfsd8xdN+hIutC8fKwhVBt2k
tXsP23g7g/wPlZIajuMXcDaqcKxvq2WFqRXveIyHk3nY8U15o4yb2y3snZb9LVhd
qIQIxQVyGjHCz19iBWLxUSIVtCVdW/oBHGnP450ktF+bOqgYh26u/dSqypri5Q+j
XoimcprYF7i/uAhErBYZ66aJJRoVRoC2lsZOHtlJ3OegpnMqGcOzfsXPxxI0Ch4R
Z1TbhvkZtXdYWlMTX9V3GV4PiLPRvL48E6//hVCTljM5gUDg3mvDIYPW9cyE1Rq5
LjPu1Mf4KicPrVok0uST9BuXOp2uByAB4r+XPEmMjUcA444iNd8yYSY87S4kGn8C
jUa2BLEmNfLU0u/DFQ6Lf35Pu7VFogV2l3FUDvkAEJSrlXYTM8rk0AOnd3gNeCl/
OMsMClg5T3nSNhYInWAcfTWiGVSmKQa3dOiLKRPU1uY51Qbb6KDRXOFLE5FWwOBB
DfrZiTJ2eaxDSTPQ+fcnmR4X2V0rv31ThopLO8dp7oIYhbvZcNxu6fLmXrWZYyWj
jzxT0iAljUVfGbLe2QoOqDUL+CFciNXplyJxzUf+qhF2sfZrrpTrje5n9DhY6wCj
Oio3Mvuc3q4jz+RdotAP0yQ8VO0hfu9zuFTs1sw7ATT+gcgFjWJnMTLpQuM/olcd
88vLEI7dY1VgtJpFcEOtPuvSH67F3/EgncFxI3Y9tAv4KeBOl3ImRI6HSf9NGADW
OlUzwO5XLP4r7+Ssp9Xgq1yxeqJn6djLXwwXP5DJGeL9e7X/pKI5cGiOhPfxRFnj
VsX0FKu+C8lcCQCjU+ncr47+PNo2S8Mfj1N/r3QUGfidgvmVNDXQKRWw5hwSRr+7
ocFLNh83BQ0ORj+e2OdGUc4gFMIiNYVaZFHwEcK5FbgOQZgB0Ac72ef07QU6z6nL
QBSbibmATz/pKfPqzbUHhCkUcx3KMsX6WI7ksYdv9Vro0fhktup4I0C9mgfhUBf+
ddJQGWdkZ1zev7Mhai4aLfxwUpPhU0U1nntCdsAgtIBxbFKPZ+DHFx5+P6frsHWL
OT9Si9tYUt0XfBCFEL7O2ShHxBbzC2ssRSp5Y5jhH2DaxcWNZo5g1qOhfoReb/ft
Ln8D4IbtjjVqkCet/CPG5dpfkfk9SCMQv5yoZOADgSUe35aiLRdaVhz8d3KBrYgD
Jb8y9A15tYqfMrNgX+eTD+bY/VmIZ0tOK8RzJ5i5Q0zvWCfGgztBM/053Dq0plNp
FV5JQBPM2TTRbMEpVtF57gNVlmlrUM1HmIV+dtsnqwxDzqYJgHX+RuKdKNq1TlfI
rM+hrr7YF/SibekDOMNkV1dA2m4qA/hgo0oXlJucNEQJw5O5Tdh3OXtcJkqfGA/1
c/QmDHVwJk8P2TleShNQY2yLizXgftSIndZHGnZXYu7PQFzjMhBjOGXrcaQYHf57
kkNLgKCZ5pbf0IupwP4C69s64kx09bCvVVEVDNoizK5Rz7gQV71lzMyg0YK8HAun
uA827LNePoOOluHpxzhgmFc2lZy3ATBsZf6sOpwWOsg9jwWGHqc/ye+dBw1FO1bb
Ff7Sd/XfuNepJM2qBsgL+O5BNa4s4Kzq6J756ACjorE8dFR/Bl6+CsU/Ja/H5Pia
vRXJIy73oSLUgzJ/DqvD7er260qAM11DMXIFB/ro9AT5SeTrnm8OZl9vexRuQnZf
HtBhm/PcK7MhrRYEJZF3o9cYyQ7ZYy/Jz9HQub3WRPLFXfYbytqqSz7m96CwOgHc
66udBuYJU29Zflo6DvhuC90By+q5k8GF1/cL+1ZlR5TkzporJ0RTGoAchR1YS2bH
2I5j/hWIInjtGXoTZpnNUBb7bKbycCcoMRn8i7dFF/RkKlfMpY5CEXZKzoN12ruE
7ppBfuUP/CvfgaCVBDdZXeONYjm7VKd0DOwQC3Fb/sL6tpQhfC3gTq4emJyLXUrf
9p4md7ncQ0WF/7uJX6Pijq+cVvCxLmTYl1bm/3Gyy7C2HcB7def/7M7EpGounsbE
2ef5ycEnz5GTY1lA5vQqXXbR+weGNGcUB+bbtMtRNSZH1qegTQFYFV5H0LVa3aVn
AmEAjn84yVF7c2r3J2EzvE+EKmM3nxseo3qnCRCkLlnu/9pThYmVDTNjsYF/8BAG
gXQTCTT4/uXTaQ3SA4v0/FSm1WsstyI8LYp7YZlSNUXug7SSRPzA8GAqzjiCo6Pu
US48iR5nlEKL/eM3YaIRraDrSsPmVFGaAZbpsWQkpVQwF/sYfg41d+PFM9jP480o
oBnop2znJ0jVXwP6dA6r67Me3iv3395Jqb1ipWJuZ1lbq7eGsF5p8OtNE7vgH7P2
rhzRAlsz0kVtiCQJfUNgHNgo8qPGPOl8fE79Jb/0EF1YZd3LPDGuirfjicwJbwdw
G/5EfZ77Arr80eRRz5YefSMIklnFkEIGx7cb/zTYkK5cCRMRU5/mQDA4QPAvngAY
vUii+m52JUYuqiI1YVDzaV7cxGAljuAFtKj+UFLAoTgSo3tig0YYbRN4dwkGuz8P
QsWj6NpH261xxXWisAdpTN2kw5P9AAjD3/jFbIyCde6q+8dbrqjaaVvHC8z9yhNU
Virz14I+tbVqnw371axpv7qoHurFCq0BDSX5gDzUNbNJqDV22C0pys/RddJ/Yg4g
z1tfNCrdoeCKOMg8gqU07XflafIJBnbZCFDKbofYzZPHrQ3D87sgru5AT3svAweE
3OIP8GSpCzavn6P0zRi7B/QnzHO/TaAOTffXdYBq+JAZGe8umuvizo7//rDRTpvh
Vf44jZdY6CG8ljEl9IUs1dCK6N2VLf7YhnoiBySN5/5zHRXSd9BcHwuKMt7u0aNK
n+CjjgaHECNvuPn8EdEKyPaZx+avFYYDZICWZ/qtphZ9hEgDI2IVg2hRjUuStbW/
hHi78lgVmMpiJh1SFsOJD/4mhnQFTsxXLgrHeWyVyiHttjFnX+yNbvb749yti1WO
JQl6kx0vlMJLfKChwpZml32TJKXIcX4mq5lExVLSq7YP5jKzdc2zCtxjPa1Nco2M
CESsO+tgMMHL4+ZgH8J2i62L5OypdoJbZZihjSjJs7M0JPQ8tPUADsHQlHVi5ym4
wcAG3kpChLM969mXlb3UnTvgE3XX7hjv0XWb2pTtFwE5moSQ0J15HSKCC+GA2yWT
HEUkiAoXTVAKCyE7WDvJLBgDG/VyJOTDqxTGeh/nW9R7ru5U47IBjensCoPuKUZ+
xN4xSyqq7fEhh+OXaaqijEmBAB3YFASoH//uf74ZXW2iYy9OXEgVGKhMV/HBbr08
R8Ue5PY+Wq+zAtCukdAo7jTm4IT5EAeTKrFIYCPdmeXvvvbv0inDM2Sp6Kt1or5w
DzG7LQt6L0Hlng77+XZQMJU3SVOKwbzacNkpPL9gQWtgBYbEVmuNvJcS59O3mUGW
DaEKf70LtwT6RjI1qcKMhi/2X1ej+CvIwhzWD0CXywQRJ4L3Zcp7Vs69f4G5ZGlP
R9NZgNuxyQcTQElRPsjYzg2Z6Q1uSi8L3Uy9svjL6OMGReeovLjWlxE/cu9vwiev
xMEmTofDrHyfGBcWnWspupFBKOPm8+OU2ZzejJJqntmBrXC3KfaOHyGy8rSWomos
e1WQZaN38SDSJRrDupJICAoKEuo75y4p9ZvYMZ+HX1YGB79CcP0tfYfjEf3YlSba
LxVZVv4ALaACnVuKMEiQk3aQu5zu43Cf03vStj7Z/4FvpykdEb1cwoWYc0BxjhC1
sVOrbBnf9cZYMH6E9cg3i/O4abLi2owwigUI5jEdqAhRw4HNdZpe8zgoLRgaGVsT
uSAEE9hG19dx5Jwltc/ntiWNxbGgDI0U002G9m4JmEi6W2JSs1l6autG2o4LAVVF
Eqa1vlFYSo0vRkrQM7Wvpt2kOiaba5pObLrwPDLoWQEu4DYzQtKM8Ce/O98A7esW
Qt4lqzz3qJrgJ5+JDMlvZQ+EbbA/R6yLRYDgUaR+iKmfA1lZA5ofLFlo+qfZFjT8
fzAwz3KDKSXAfFQEWAJQqCa0JpLtr03OhTAIlIEdp19XXw0miOY9saZfCoETuBCJ
V73vWim3ioL7x+AMMVdPrw11FQKSVCjtxIVlMX63wyQDmoAw4cvr9urmUsVoGQ3b
rSivNKbnj6/radOMeGxk0KJRHROOvQwqKTnwI4YrNjc+P8X7+pD+uvnfFZmy3ZLP
9afqfJW9Iuq96bznua2geZSPqnyuspKjK44sOdPd6L8fcz2X+3N6iZWtutO602Yg
Gt7NRiszh6/lCP4JtOqcu5/JtPIiEoN+Co2/EvJvCBrCKSfY/DUW3UdNeMvThelh
hzrvXDIU4iqRUxq5KWeYsbr5xSEB4oz90iGMP2xHahgq8+ZIEo1Hi0/WWeNvgOBa
mQFJ/kV1dK9KpUBcfWS3JGYDXrqGybmrmaupbIBu8d9HDle+45zXbg+nre13kfsD
KS21tDUY/b16rzzZuM0zpdaWXZtWPtCQkpBAe4FdZun+cuenEAlTH1Wjt7Kj/Bko
ajFbDcEHv+YiGt/sBDyFsCM6wHSfeSqr9L6xNF1KQS+quR4ERDDz2/Gt3cafufq2
rDyaigbNGGm2Nf1Y8n2VkjR6XMb+c9ML4NzukCVL5HlYSSCZoCSqXW8GbvxR+Jos
46IPs58SijbgJ+nnW4arpA7G2O21lQ9ZCD85XkVCVg8Z5LqbJQFPrsI+1ptCABqV
mgQfulENJgsfKKw02dhCfi31arqWWVexfr3jK4rqgF1VsWU81eMtKWD7pi30KMx4
h7UsMdb0AFQLSa6TdLegLOGIcDB+X6Ohug1FM9bUC8FXv4urtAp0R8LTj2AuIcM4
vcKNRw6eJsNIIP0pT6FDsNzf6wvUCI5un74UCHS5/UVUjvFUqXz5dcFNwTGUm7HN
U79AgAemBznp0L7cwRqMW3J0emKljoL4mBiu9Ryq9NCFCdODKTq/yPNG61Y2n/dt
nwS8eAPcoE9Om5GmhfhZ1XsHdwroEsAXmcRL814SMITOUt7iB4zpOQEra8i1Jzb8
pxAdj8eQpDke/br+QUUryLia6Q/B6YR+fCsegul1sd17AKxz8AF73NjKZFEs5NRL
V/yTa7Ssue1W4Rjmtql0+dVavBuwdyAUgixW0YLmKAqMBNCWUHGtPmaKpGzQmQiX
9hBnikJKzoKFm72mllLYLWZIDWleDnYHMUgpPZNqP8EgVVyj2eNKtWc6ufzlGgYb
nyvyXIhb3rm0j5tcSCWcHuax9rUQLgq/9kMc+OIkKC/OAvoZPEGffga9L2W8WTpT
+AukrTDke6uLPsOhSOGaPuBJ0ra8Wk8GONnnsoT45qOA6VYdE2aYCNmCkdzuKRck
ty+iuijOGW4O1kB043ixNuR7+axRGJTQyBjvb2qdiA7t9BA7X51UkVYInh1ZEEjb
RCaXe2b0519hoObQ9xg8eThhgixiQDCQCCuFGZxzXXf7bwoddJ+BpAhjSj7X9UXL
VTCN1k2x07EFSmi936AE6Ph5mv/teO7JAEMwOw/8LGBQk/NrpqDQ8WGD77MqnN3w
Ub78+iXhpI8EYtUxPgGBM5Lesi+GicVdYGFGuvlPyxzWK1nA6YlCtLpw5tr2fD+R
YF85u0X8uYYc7Wwm5QG2pyLxq9pdakO1kuKOWF1TSjmJUG43+KgqGY05KtXTIzp9
J8E+sHIJyJjCMGzhfr/4Ee5PkKzN9cUhDlf3f862HSsiZ688qphlPVexRy3HGy70
/w8GcTBYka3JUo1x3ddEz4NEDO2TOe7i6jAOa0GDREVgLC4a3dMz/HIXc7v8VY7P
1rmkhnJbe76d0WqAbmqkVhJbiCdCR7nujNMk5vi/gcIyjHt0jhY+6MX6lnm5dCV6
tCaFMIn5bO2LG4/tEGJYXWF91wM6Hn0oaQ7eZ2IW+ooWpBck/WtvQ1Nov95s1bCj
1ZVSCTIgM+C2Xdae++7Em6D0X5/pP7HcbgeDOi6CJucQ04Jv7fYb7vK9s+jGgUIj
JBVKi2KgGgWwJVkbYI8bLwOAiV09uTEGPmzjbzYBfOVH9iYNdrT5rUc8h61Xw3Ri
ryPMks9a5z1CFdYqsYEgMm6701hRpKtvEqF5aJLygl0poaSxchiopRkubtfcbhNY
d6QTxb2k0qv2SwKAeRQiN+jbguPiL5wkxLK/DyHZy6g8jJsgbXnbwiazQQSKMvuu
IBBo7cozjMoJgQ89A0GzHI2xFugS05C1DNMKUBvgI347yBoOFNQ61dbo87W42cka
y5RG3uuVMaG7K+pvKwVQlArtxAeCZto1dJsZKCokL5iZbbtmERgCCZI5YxiMTEZZ
yu9V6usCQQjFsmfRZPCv5R5m+tE45F3M7cJxkfMUlGSrmIvwmgmZx3PreCYSBAfI
ZW2S8AngClAvvL0pMXCkUmBYR/Ntrw9mxWwkGUb7VGOHDktmtD3HUDdo+3314t0J
+PBBLNoWV2c+sS0WAiKtTQVpD7zF8F8TVNGmFQHynWSnmkqaI4KjpOkFCps5h0z4
BK6zw3wygmcd0ajufu1dIpi47V8tczDZ5lQM88Tp6RCCaqDQC96GeF74FFJcmATH
rsJS9BVMWTYUn6TSnPz2bSJehnV9ajAwnyq7vptZdFVXbrlPc3Eofmx+I7tszCdB
R1gMpxqaEKOljYcyKEho+QxFeBTnPGrdWA5pOCjBCMBCI5JwGw6UKtz0DCtuzEEX
cMQSdVyKYruzyJ8ezoevJbXmm+vV2KSbTnEMJU7Ucxfl0D6Hw/JdBJ4SJvdC2Cly
sfXbdNQvm0Ye7YRygszu0w1TYbHPECyQewqhHxUhOZaA9xC9myi70VOZuK9QtFQo
LtyPnOSjRPcdiQoEdbrI9vRf8LPivDtCK/xoIlE5HXD3kQPqVcAHMeka7DOtBRq0
PFQ6n++Pld1dBF+xfvzKMv9etzfHbkRVW/+upKRpkNwyLZJvf8g+AG04KGOm3fgx
D1lo2ybyQ9p32fAuaO38dbw0qLIogGCBI+vDvTxLsJOd95NQi4oEndG/I3VXZYXi
CG6tzISWtZnpRCpBm1mrrAfp9wucgKMayz4yfdp1wZGWa2E4iqheCCbKuAHpkKcx
7R5wVl5fVG9HzVPIc/8MrEsFmOQaZ86xZd54ok+e9IPsr+eZwSTcvhBmSC4N9CBg
RNxOVc7PcYuBKeB44ldMqPTmhdF/yiD8egrOkPdCaeukwBFvNxJ0nxjJiYhCKnTE
nILbXautIvWwCjXLYdDhec+sEB1FODjHWkl5tLdWZxC4VDhvpCyh5KV4j62S8wB5
4bRLXXL+leRjrgRuRLXKTIEv+rPMJsIReSXPimzBU0txTCxmy+f5T8zZU0HbBlL9
OnFtfmq2wtDkXmpf2hvg/UDeS9A8Zddk7VRi9xn1Bs43iy4G3cRTmrmK4pyEaFNG
fq/T8Blv7m7xcx8BJtKD0W6e+gPRNToOJCRoxFYNzVqT4ggdYTZI6KMugknLHjOm
qNM2G+Zl9P8bOeDoSg6dXwZ1gQRcWFTeZEW721uyaxi/Z6e0A7rF7c2kSUJ5UAXB
S1MMDJ4aOI62KGs2LC+uIOptkRFTQpzZRN8ik/X0E3b/7yRF+NR8+J1EqeTDq72H
+K4P191FfWhtMW7f/13KJ+HyDp5rB8f2JDwkrtroe2VG45OtkIZLbKeg7xgao9ca
sqQPWtVF/g1fA6LPhLFuHmpKTFL5hSO53kuk6hYpzw3j4a6jvCAs+tup7LCQycWD
FH69jJEap5/3NYbMMPJBko/CH+kevO2o/NJwwypDb3WgOFwsvve38jBSKeY15ckW
Ixbn5WXQMZ2OFrGmeSGQojSnh2p8yiwux5wWtBRc74CrFmKHaWIMOYyY1f8GgMAv
fGtgDDANxU/N5usOKJFNFOOe342r/5avQHj3ZPPTqq1TOd00JVz7QnF0XTeYsZRA
7wHcKmDn7Dnqw9bIlqmYnlluhuignPhxGU65/8x8eVGnPV9NQ822X88F+WBGBO82
eTGE+zhG2o9vUARq34A1M4/znPuTXaPWoWVXEFXE8xFEkEUH2+gTDDHEUET1Afap
3wkdYcD1axI8WiXnVbb/BfXLf/noqtmkYjG8N0wpUPrdz1t+am0Sm+rma00fZdKw
3dhccnolfzFbqHfJXmU2rFP7WpCS/RrjQrPtVEWq3nGcAeuQDmcJX7OYkQzGOHdv
UEFmSNrM4UNPHWn3g/v1or3heEXNvV8sf75wiTCZyf0RfJVbCvS63schf+IrYwNJ
jnpT1DEhT7kFswfZ1RzgUULhx8KnNDRmQ6GPLmrMCBWK8Awb/J06wF93ER1qGuwT
yKZM8yZFx0kJu59646iCxPLng12b+DEWnj7t5OKs6j0PngoGHIdy9T5llpziICZs
HeTu4bfzex7FFXRfP01KTWpEhZes8Wz5DtSPP/EZ+jHXueAWiUTAPfJzapChFpv9
G0085Lb1FEtT/BA292d5VO3cgl/a8qgRcTWp3dSpQTYN+BTpFw2TQl+2thtE1M83
LIa+UvQCY/5fENU7mpPWbMQrCNK3MdernKYGbVDE/nGuqFnZZIvnNrYzB+voOsQE
StIxs/RdSLPE3exRA5YsaZLDo7zt3jpL8PrhBNPibtVbdnfbralMR+0XXJRIwmBw
6l+5pPVd2G3f4dVrIQEAqI3NJ4bAdn3qEdX/UhqyfkOowfBeBjsCLYMlAeA58IDJ
mrIr2EQ/dhQdvZuyBU4c/uBC3nD11jadgfbWs79UKtd7Glh63dSdZN5T0C8JM4qG
u67DmKHuJQAvZnraDPYGk9OqWRG/JMdzSNZXHNNikwxn1fvF5THvGz07R+8CUcd9
8ozFuJEniDumW7f895nqNZtOReeAD6FTp2QN74IXOqsLPJ+uiScUnXkiudb92FHG
nWKnjRTMsF3SGFwHFJn1rW3VYnoJsj3lvguiDtNnltvAXMgL0ya+LYgXrse3ES2f
TGD8p7QpKznZtafQLDR4wY4zpz13mfI1tM/2urqJ0J28gK0w2VZKZWVJp85KFadm
2SQmLSCKbQJ2oES7SBNvVARJpdj3KPE92ysgCBTQXo0Fp0q1ZulixI3sFvTZI9s9
U/xKC1JsGauGLHEZy0Xf1n9NUt/MfKF9cDuax/goCa6fDVgFcEcfa5bnt16f/Pdn
4AQ+RwDoo6DTc2pvXpGSxXjhJSoe3aRphTYdjnewi9AwVTtJMG8FVofx8ZDI5YYc
uF4s0uOL4nrM7yXGnfD269H/kxhGpq+wKx5DPP+P2lh8hEQI15wxvK3fdzcKJy4x
n8oOLFJ8M1ktGSkE9FK3deQvdS2gALnM1h+RR9wFXbt4jol2r9aO3lBUuq89r/H3
XsP7triFqRBUtcO2O0flrbsl6z2gEpd09D6eVN/DOlD6ZNvb5+geg44mIXOQqEQz
0E9WFdoFnyNuQVGFWfsccHfWEje1VvWuV1y1yaq0BBc6VDrx+zq/rFP1JYPj9WZK
HX/dVZOKdKl7uHEWNyr0zsEoDfM8MnE1zOUq9d2cJ8cIGuTBH1GcVJxZG/Bv1eKv
iK5+/zLSr73+qazXC9IFMXKj4zMXayDa6YsitLfKGsmrcNwfIsTR53wQb7UDFjSd
VcuG7n1xIc0Nd5p2gY3uftQnUfh3xyWLjIIuQcT533ECBt3g4saddOO28coLvwfr
29ncvn/xwYGyLqTXoJe9C0BQpHZbD9XnhjY4kRmmZB9JnZRa2qFJTW4F4E1V+shA
PEk8CRA3HPMJNaupUSExWvMKoMCHTBWNezuHTMvkDwlP8VHNd5ybiJr5bOSk9DNB
uQSi6PTisKKdDGejg2BAA797Ws/6nuwKTeSnIUEPQ24uHwmXVj94n61n9mEbgSBt
gbSUhap7/zFG099WaLWkz8WvsUbUTSHcKJnw+ExC7iXIxxbs7U7lnn36F62woiQA
7AnUHkpJxS3GEHToFqmnTqea0Rl7e+ZXmLDdCPtrzETVV1Hbq8CX3Bwh9hTw12oy
2o5f2C3ukztr1gD0yT6m/9pEBfoAjYxCCPnHDGLn4VcoXFQTUljsF4MZkVyWK5qE
d9lY4zdwmkZGqeWz7zLKgL972bktR7tcHbs5hE1fMW62GBoe6YLsm1HsXQBqWzqg
BP1RrvaISR9sWw/BQBiNN2dRRVqNS0UlaWt5l4xp5gzEeMIuJGE2Vhsld4qjuKOE
Iq92qz9DhYP5tcw6ee+zy4xLDJ5HfQIo0L7Oze+CRZ30FwhVW8/T43Z60H0g9y8x
41JhCUx7Kq4xbqUoSXJK8LVEGvzk6d7SdRIp/+u4o9YsTBuJWYpbtn+GfvMw1PLs
lN7TyAI2fjou8zVi7s97D6VsdYoGIt8sttw+zsGGD8wjkJusdtA3in9RXD/wvdbP
exmqtfkeuvtksGYuqnDBBmemPcAeWCuLqQMclv643Z6YBk19vwlYrzrcFyqbshSS
OFmZIxqtmFAMez1+am+Pwtwe35LD7Cl9skexwIjlZDlC970WRXYHgFWzkT875Muz
CHR6cXDndNzg3e9ZxYHrTURATfnawhy92pGe3eM52X994H9Y9gxnlWUD+IKVyS18
BML4edg4xGzEU6XEDoWY6drjcdZqE3zzoD/JG4yQlDHaKz+YUssroyx1eHAh3g73
vo5aDSsw42lOYeJvT1fqE6p6fIzcntAyohaez/NgeRFcPZ/jiXe3QT17GBwz0WJ9
OlgN1f4SzARVjazD4pspx0KTrqJa8JwSeE2BX3BcckRRq7JsHYO/4MdAsrJdF3O8
GIR5fml1fKGxh0Rp3PaCpui+1oECNDqtGPBJw2ztnK98fsNaGRbxc5wHBEuBD7E/
szQKligM3P20keyKgngKRu+Em1MrjjjDstho7T9ZQ+ZzhuN6uO84gcD/kwBm3Q3A
CHSVYv3+Tw2mCGuMna9bxRsfk0bBWc1Mw6f/v8KrTKGVn/u0U1o7sYpjmchcOWtb
Y7MrPsnWb5xdMRMkR3YEI+lvTOB9//iD/iHtt+WY3W81oLP3SS2Y3sGm+gVL55/6
DvjM+YIJxQCN5rx9r4+uTI8OGCyqdK9DNfYXuD4dx6GA1ZV2p2qnZ/38iRoaF1nD
Ra10Etv+d365gnoPsZY9uAXA9t0F9POCNxMk4bx2ujppQttkLHDuq/2yIJd7mttM
KcLerU9k1Ju5qXqRN0RbfMHWM7XAvx/KI7PxZc6cI/cHSCeSVi2NeO7B4OBkBgKH
rfO0+nVejkzYYFanxvkt8pw6Q722lRBGdQNvwC5qqs2NJODdgwe2T7BmdZYstre/
c9F0lCciFr+M+TYP4jUu1+nnwkY8F1EC41fo2M6zuWv1pqF5xkefNUvCMdQO67Pf
HInyUXss1dEzXrPOE7zUsQM/HKdQA/WNag+zUkQn/LIfnuAIf1PQk/tSYCouGh6C
3/H+UkoNKRZoeenEwFuCSyeTQYig4GHxjJXT1mtwiw0UXOAqTP8sX4c53WrsIRiO
wf9KMm9oAtaX0nJz1HT1gQS4k+sKrA1SqpThnOh/Xp4vwteWOOfhXj09TwZKZfMx
wASS6yzZKuPWC+sQNf+UoylPM7KQL4khdSlk5i0UzipuZr0Ko4u8HSl7g+AZIFER
q0YnDaIX20zrkjG/KKw7o238z7FW3suA/xsMo48Iht45k6xzZ7mpPod48Uq2Mg3a
lM/7RyndTJ6V8JSvfBoFm0Acau1TVHFUVXqFUXjyhzP0j15inj8DY1dDAt9s2sct
nbaJytZR6LC1XPusPqMvVc08AzjOuZqtTFNjKENmvkK3w/4ApBc45fNCALu6tlW1
8qMl/i1pOc5Tybdx46pIUEHnHZeoOsLsM79jCmnRaHKttv/lBw+zKSz2B1rju4W9
u1r14JiTQetCATIxemkx2i9va/cq0mmITFcLBlMF/GX3SLkMeHYvDCwEcND5O49/
H0g74iSiU3AT2yhz9uWD+6vnyFC4HCi1dPvlhFfslJnoMWXZQ8GgfTVCuK5mf6vN
oqMULCA+OzVkAxdp2b5FW3OZtKuvowI/SKIHwPh9LavSDjrxNBsA9/gT+syrsHt9
7ohUyCRyTCgzykNJGrOyfkzKOgfUR9tvsd940nfZEPRX4jD9lMMoANjZjBWlIR7z
e0xj3ABy7KECBH8dLBCvim/RHQk95LnTANHMzYceLz4fHkwI1K6+JJ6d6QK0kYbB
okTmb8a555+5O5+j0Dwj84EuV79AvnvD18dWOBoysDiV8iXIoAIxOYk4qVZcUcJk
J9Ap8uP9siSLgZ3qmUCB9HsIkW7IHAn0uVG4AQppbZ7B0OpeWu/MoE6mEtZNtERV
t/LCO69gnmJMPX7fKAji7ofQwgBNIHag+plyfsAu/TIekvcXJA+U47cGdO1vT17U
5dLxjflgGcja4VxCS5nG87I7GLo8DDYUtxGPHw1IwteW7RsdFtKbS6v4ZSZBm7nJ
EokwEBQmN+g+JPrRbuhhtlwg//MjAjaip+WfB5TJZFtHE1AQSqsVGGLET80MQr/I
VEePo/Xrgt7mjSN42knaIDVHGud012+WD8T25jdIPPZH4kSHgB2ulNbdItupIr3q
6l4mo5OeEMjNUtIvtCpW44m35J9e8cnQXHIqp0uo0g/e9ZiJLvDyh5v6DAd5dUPH
eF5xrP86BK1JmuB8XmRHEfE/h/VDuNRMNjcff7DwAhues+5dX2ozNDo6r+pwBsbe
D6hUWaddoZgNIdOzdi6LEI6qpmYWb0qV6nTjC2FGnq0izy+pjDpDgzO9NedGabmx
Tj+4dKcEC2QEjRuat7n2qOxH0kNQExmf2TvQX40sY73KUY/f86+8SFX7v/tQNHJH
xQ6jZq6fIRX3oBL8dqLvkGHazdX8vSUjuyD0kCKVLInwwrSEvg6pK15fkki/Z8xt
fva16QMZ0hBC5luY8nP2dZ4QnRJhXdNRAzPiBlNaAAvPrN/whdjFD1KlRHm/vNTJ
RjhHwO9wI6yumereHyJFPhBOZKRzkuPu0BZliqlqgVHkqYdNLofysVr24AublgO+
oKo9LDsLeMIvpnRGdKDfwLb/m8ZEmHuUhRHIaWWdA/KNzyYahNckK/ZAfsRnaFM0
IUEaUdquS/h4BhgvA0U5CBM45X/RfIhq7SV7yauVVDCeTs+yzpRfHWPmUQCPoM6y
IRpAq61fOHIy2NSjGEkx+krP7RSNqslAqEhbZ107/8Rpc8YY1QpxIEaa/b+PyKGf
5XcRZ92SXQt0cju9/d65dwhOQj2lTdapIhdJX7ufFhLXpj+RWsyuXBDCfXHtzuIN
PrXX4tVLRurvuMxFHXWQ4ENC1hlVu976rYP6d35BNR2ed7HCrhfdhjuMqaKhckMx
PWce1IoNdXi76aGd5MzJ8jMoVKERFwP1wXY1c3F9Vpb8C+XvWa+B9aAza1I+KHGw
rkFhAA31g/fhJ1TuJcaYFybTEp49dtK8Ppvk9qBMtPzeB0iO6Il525B44eyk5my9
RFTmTz7Jsr+rNLgBiP6TOarRoFFDTOX4F8Eq5NU0RaQXyzxSMxolPdpO1djnKWhW
X8LQYQwCeaWFhVYmX1BOabT25QOXUS1CnJ7I0e76xw95grLBDdrnlr92uMXxYwQy
ckqNIVKZ0i5nzyp3WuyaLaFr12uODFcxuekNn8zKwy8CdfvF9HrTl2cLZUNRZ1kw
jiq1q1+FE3KM+qcUWS/JlaOhp2XXexkiyqWB+iic6cnanhKLU8QqNlq44C+7b+Bf
cPE6nkBRhXsznXwfrrkVwyRi+QoVOGSrpdRcqEoEj0+Z9dhW2xpkeTD7chrhovLI
u+VaBmmddtt1QoVBMBCqY9cJL2ZDaCiEHpGpNyw9AyZV7Y6ngonCNi66Uc7T6d9J
mQcaawskirY4SYejayA8afgw+9fiqNAg9XeYeaAZmT7dyFiEi5zlrOnLwdL7Us9T
zbHYReRTJJcM7jqifBSEVKW+WG7G4W36EoelJejDHVETRuAD6mRjNtO3mJl+vG/C
NwFz9W33CEBaIvJ0pRbiZXN596HpSjHJ83eeaXYgtmhlpKShNNbCY3NI68nEIeQi
+vbjyizCsy8tX8ygYHAeGVITjPewjYQIbnXhEOPOL+a2DG/IauzmbgzJ0UFg7ldU
BaG+PRjVJrm8SHhOanhV9e07FoDYqMRRGnaPgK73IZlRot79yWWptVd/03qm6ODs
x4QI6q+feEIPBldmJiOXFWZEln7fWnfK2kuflx0Nuzi4dpLI0ZnNjYfgp9PT2Kzs
Qt1BSXHb/cLYo/OyCgCTaO2MWowYaqgHy9YQU0xcmYkfZEJTdVB62fTsbp1mxHmb
QcPdi6/L9sU1XdXw33ZOswaerXmJj2OMoAMlWT8qjSicj+febSYMLzTtlRqrDVFm
kVEUVc9KZbH/3Mz4FbltzjEdLOV9iu/vOfmkQJCxKhq3wlkzE8lz9K7DPJGzkLel
HgQsbXmv0TEQap0CAQQIto9aw1ox5Hmzu3IzRGWzuLcEjjOlFnD5/6+aM4blACSY
6LoI7C5CxcLyKkguV71aiO2n6b0EH1DneLkyTCaU90O2Y29Ss+MtVBaCi28awoYb
QQAlZEK+wGaxje09X4RVToD0Ls7Wwybqo5Z+dkB1Wsrw8vufzfyXT4/m9QQz51tA
qcDO1zEEBcuToC0Cre/X4ppJd4EvyK+VTIL59jTlYBuoyHaDCEdat9mOrcIiJMgt
MUtQOBMVlAjqjmslUYYbMJUVCqhShcyuBsU32iORCSFqzUEzfgGFxqt+L7frQb2K
btoav9TReIVi9ejyhne/TP+x+Mw8UwrUy/v4VHvSIdZfaCUTGvybe7UcFcgGsN17
fjQ2rqb364NP3xNhw1SR3pxAdUylcIfQ9CaT3Cv7G9tt6NPLQH+IRgOtET5N42u1
MYiowdpQx49LI4TQun4x/gYG9dkM+Xa1XHLyZ3T0ODACYK79zLz5+KppIiTNK3Js
LMDBVO/HAxDIb5o+lV7LGTG5nu6QkCKLUl8yHC5ZfAmWEq+/eMCDIICTJPmYxlbO
GRfo14PxpQKApvpE6b1BKjrSuZbEilO4yMZ0b7QPlmz2YX4TDk9aqISoepq9U4Hy
w+gVFBXpDYnWpBuuB0gCdpVaAARQDV4M229lqHCiaJSWhBvHNKa0ggBWqu4Jk0Z5
M6ICirHuB4yCmv8Fs7JzF2Wltruml8U7paZDn3Q++XEa0u9apC8ZwSTz5q7sR/mI
ZPLCuFVwlozkPtWqvbZKCWNNLidQhDJqMOv5jtoBxnoBsJVAKh0joN5/qnY6v1GO
E/utQmCePdNNf9hZ9piTvvbqOUOLptO1ws4tYWHc8LV1DtoSEpJ9E78t6ilkuQXJ
Q64pH7wzIfXKj7Ob1brPWhUj92VeboqdCtr9dRLn2cdc/TC6Drp4baLJ66534Sfk
sHCd2Wpwh/sQq6rZq13QiYTTCwSSiXo1HWYlTrC7vIJGVjSTm0i1sj2OkS7R5LuA
sCkhSrF7Mno/yHMgOsCsqyEXqqtKWfY7sCQuK7ds6bFpkXX2/c908PFZfgHZO7DY
9jACp+M62LqHZUU3gTAmyGRObGxVoM10/ztkUB5lidaCcJXevKEWjNYIGqbt72Qe
lOD8OzAX7IorDI8Q8Mbm+PJwF4iWIPNBcq0e5w6R83ybnPY635AL5qlrI2z5Ehp9
/iVqXKB4rqFvt9ynDJTHox6zuhJe+VeuGpNWYULBwOa6V1VWYWawgafh2yEu1Zjt
D2AxcPMRNcJwxpxeJJTSBXdFP5vlJwHD9/zG8useBtZ9av2b9V5Q13mBD5g9X3/a
ZeXjq17dQMcQfT965obFuYlgwCh8p/o/rYJlh5nUlVbi1U7icefals4dvdpkz9gb
32M48dDUkLl9PrEYEI26Pftjo1infL1g4xZxGlnk0ZsavC7W7S32SWU+7D7e8JrU
5/CE7NTszP5PKJeQfcYKbILTRmF67vPxQpzK5ywy9Smc6dw2vknAmurgbv5u7Ra0
y4/h++XjDXGPNbWd5/M4twj8xR1lrhLjWpoqSrdh0DB7yKvcnCCnvOVuxZX9+xt7
Z8+RgRuITYLZp57vyZdLVqShBwH0iOjGZALyvjrqIp/MlrvAx5ae0Q8RjdunymHZ
ZyO508A5QUnt4qnLZBoLIzFzzJXF7ddkhQWe19GdEZ5LVM7QM/GV8QES+KKb/LGv
HHj+0DfEfgn5T6MNN0+taXF0uL5FLd+3mRIrPybD6l4XbTYhAmjlnQr5EDfH342z
UwkYCVPsy9uZ6+70uzDVP1bSfB6y5dGFtTV9siRAI4vsUHdVx6JjGxuNjIlUnL2C
djpn2LMNjdjtxliA32Ean66BRN88qgW8H8hz/G2uRhY+VJViarbBTPp1AuVmZIAq
5tYE+3MIDJVyDgVFt/xO4m3oVfM1JflLpaP5UG7KV12ABYiG67SWTR86fUQNigtO
Yb/hRRaGIr6j+j6Okdf85WhBK8dziYDjUytJwR8IQDE+iXfPGDKEmjw+Y9p3UBdH
wZoXj6Fbxw0EqR+sRGbhKYY7GZ298ssxWIwkinp/pX14aGXUVKO+/CFtIbfr3OW7
xIQfoJ5OFwI8oGE1U9PibpuTJRaVj7br/ns9OEXNA9iEylCeKAPTZtdzuqIwVHvg
/L8U1Pc1Bp2sCYAEMuaISJuVEyuS6uese4sLNATYdLiw8RoGd50e0gNEbCFiKfUr
5Ixe/dxDyIUucvFPrK9jG3KISYTc6PsF2Dvs1MzWv1H6byunaw2wXZmGtnILQ3AQ
ro2j6bNdmEbnYkEIuNdIJlJM/dQRZqEGRvAbIKzf1ips2u/x4ysGK4eqDiU0qVVu
4nFjFr/alAuGAhH2YjhRVXOa12+kRZ46bdw2B1FDd+hU3sDAkZJhnb8KMJrnc3IZ
dLohAyuW+HpjGEGeDKFkqRduSoSsu0+55QwAzDKbEF/ACF/kAI+HqP7tDOsPEIjz
HIa/X83mqDAAS5By9/E9Pzjb4vGqhja3NwkMZMRolb1HBNWK0hZqrnjXo33yQgVn
QkEeNH5LdK6stTRg4XiXgqTP2IxDBJy1PX7wnB5lNsG50uImORLxys6MYLPKzRBx
d32ihLfucMsgWjBRys6HsOMRah3c4PZZtYjkXobSeSKP/9eviPIJ+5V95/RO+DZP
o8jZ6trwJA8QzmOlbERBAcXr0JbLCACjCDXIDa2TAKb+tZB8GfS0Jz9yxOEwi6L2
v2f8+sprDpA7F+SakUfs84mOGndED8uV4BenZ0jJuERupB/vXDIuUCON+9SdXqMf
xHTLmda3rv8AkSgVGeNuiiH+88H87sA2+KL6PhnfL4PKdOyoZsWehP2NMMMdBA1V
x3q3O1uVjhkRdgte28x6PNoU+Dgfv7HBoD+QIU8Fx5VjseWQ/83BLlTmRjUTimsI
Pd4GKo3pRWb9LHEiWpnYFlprD17cnLPGPJzDZVPxRSjvNhVsJXGqKrXpPTiM27nX
B/GyTOIcKsy+b5EgRu8IIwMwlcPGYL3ISRDxczzk9hTg0x8I7RKdsAUJ/1gP8H7n
+CRMNPanqLrL5RMYMWeNqDq+Y0chCTYz65Fj/8NkL678P5BY2O+teHJJZLRBP4rn
vNgy+D1jh+Ive/szqR1IMhAIysdXLUsqnYeUK5trq3nY7UDOX0cvIjyHo1aveiIz
cKm0HngfgXDjjVri45pzNeeE7T8Kcjpy1uHTDKgiqd4OAOAYGh3NW9lAfpFrYc86
YZ3myMLRMG3MmtvRBJpbjwCmhZ4wpCTtEOm39vHQRzAUFnzToI8SnmPGeconLFhg
+UbgNm0ryNo8OXWHWj/4Ivz3B7dfcuOnoAjdBqwiNZW7jWGt2VrqSapv3EiEUquy
btIYLhR4c4dyT7yGPGw7M994ILbc8PMuoJOqPZ51UcP15sNBfATWmXMxFwyLNNqF
WMOzyGaPPyBqiVbrmJcWbxxKK9qi1c8kfmuOxM9ecw+Cj6fM7yP7xc25o0mgC21c
gY+6hkavFSxfX59KRReGujiEZeW/+8yakVkCLfmdN1KHzu0NwY/TdkzaOr+xMKf+
fKfrJFbex97Sffc/iMXZVAnlwtDRqcoZfkxXpM/bfd+/sRlVbFpt3SoCgt0YuT+L
8QkDljSbRcn2DU2Ht0LGGU3PNRL+Wx5l+gaS5s0L6ZBgMvbrn7l4VWFcF/e6EE40
wM9846ID3IQwDJBdE4sMLCA9Uh5BgQwQw9Ix+y2I1atFr2MjCB5abZFag9tK0gGs
xXkSS/LoaNCZA+eCr1Tjx61YJY3CyGXgOGYWYIDuMFv+gdHuCzYDCeioDepxfnmA
XWN5scWaFwt6IzBkJAhmEKEWPiuXX0NhQZU0SVX9UdI9WpaCGTtB9qsDRwnFdj9l
xxCAogiUc6HSAa2aumRlOFrC0MmHS9+/YPBnNJiGRpwS1JUU9UMQg46VsNWAG58/
AYKyQBc3nAeNXaO/UlC59b1FJkcO7nx3SOPvK4mOXreOytXeopTZKLoZ9+d8yr0K
KH/vJ0tN1C4R0KnierT4F6S5E3WVjkDaWpffJ1iIgdmIcPtY/AohPaZ3vBj2UwqC
SRjsQTPSox9XwN8sx+491bVE6pOq6Agd4GNPR/6IaTfjOpnI0QAOI0DN6TJizTC4
7/dYGPyo3ztB1zeHDuOuPiyn9E0Qq9L6ki1B07qa6nfBmElUUt2F23wXW3lclXim
NEhxZfKThRnWJelRkibzwDBe92x+UXI+BZUiSdMhMoK6XnqIPgt37APeFPBVaLbs
EmZO5VxhY+W7Ca9qL0ourpLGvUepOXq1kRzyL1gttR9Fg4EjTuYYLmgvhDv3RMVG
tJ3JTC1UH/AfJbWu3hYpDtDrLhNtNkieD88JjHJ9qbevKIXITAEMoWE8/hyomsIc
hUXhTBTSYw9p5ZCzwRCygM7eF0KwMyHGcJsknLxTYQCMeKSSpfq7IoR+OtxuMlQM
c9RXszx3npS+NToz1DehpBdZs6WWgFKGPPES8EHjySVgWoOVQX29Rd79aBcUBjDH
gCx/W9p9yYq61AIi0nvKY2SrB0768veQcF78RAiB8fx40wtQFxs9CcXqyueJkIII
5hTE47LO4CRwF1IrB17h+8By3ZDV7Do0kTYhcz7itrshNCjiL560+moowQz0jihe
b+rHKgMQIcikgHp2pwjYtwUj+yCJBpTv4SjU7t8pDs22GMzg1d1lo7wCUoZ0N2tB
2fozQIjfxBiHVqX4J3tMNmoHaL73+CEmMqSFbFwZfexQ9bgyicLbG3U/V6MJeU0X
LVD5EOetJAzUsHeYw96ouA7CH9yYCsnwFXdvUAHkTPRoYY2SJAQxnBltv7zysgwF
rj0uI9vr8I51s9/juTGF82FeeVJuaWH6nTy+VFeJhW6MGoPmOKEHPTMM//ijLhxb
NY7lnbFc84faFlhABddkq3o/4pIFI0L2/8f9rBu8qPkMQNoFFMiBf/9T5Acrjjio
0ZhxFSSgjnVUbRWZNKDyPKEs9klqySUp08bw0NolFeFsvULuuq3X05beDOP4VCN7
59K1EBF4WP5RdC3+MBXcleuoCouCzrWpxiO8qtunnmcN7k/9Az4O3JeAGDDNHrma
ld102G6FrBoB4OY3FTV76R4DN5Lm3nE4iBomiz8HU8XOygITP1JaefLwRbBlLZ7p
jR+raROc8OaOWAwMYMgbFXqSRETQ5pU6q3+vyNzhllIXdoS6zrSj7cuDRTYks0V8
q8cRVG+C8yS111cW87Fqaru7gmwBFt3P2hF2hViNRBYM2RE9ORBr/icP2yz2hITW
ILQyEjpWcxVp++Q2icRSMDIR+oPwfXMdNqoSGcxPYlISNTDBREBOx3NqjmM8xYoS
IWdNoxrMeAODOPLTq0wNa2N+ThPnzWA0IOUFqchM9KTVwE84NVAoO2MaYLIJ5vh/
n7kwCUrqS2sXtfLlmTow3oJ1hQyF0dLuS61GeC2OEmSAY4Pb/UJJY9rFTpI7pZle
5lXav0jd0/RF71ZtBNlNoHAzhsvK9QTKwXF7RE2j/8nk3w2oggs81bKxNvE/S8TY
2nbS32ygqbnk/W+j3H469uX3geBuMx3+jSQHD5Q+LqTgTtajyqdmAvC0f3mZTYhP
0tB1GQFD9Rz1Olg1T/MjSV4inrHuxYxkjETVRPHOgcVybOZZPuLN+5nv37dq9lRB
G4qy+mNlEuJ3YtYsAOk7LB+JfhTpONcl5YmQ9VFkVLppFCen4bXKRky7XzON2rrF
/CwKQRbKXcjhcZo/MUB7LfsKr21kNU2KsZBzCbC8cRlRAzGvPvDqKjKB7Hhs6Kgc
32F2JKu7rYxsJkg3BGm+1i49EwJ3TLPuKP+xEP8wrx61PFVRHZjWqNsEJft3ovZ4
yee1/Wkc2CeVpBORB6OtXZ3f9JtK/9sFuf02IlBoaASnOffWYjWoC6SDZNExuwCV
dd0mioiYE9lVXr+sK/xieXfO20GpUuyQRqWVL8fI7uuBt86NZ1PfEUtPHbKhhVcL
sO+XuagayUtgyFu3+sD/FizS0HydSTvj6q1YFN2yo6rHTEoLexOapW0z0//16EH5
aTmWmMHTjcAw50QijjGuygle8P1ikeDUaiCsBebBRypM93sqnSUXeQ6DIQR/jCuG
4cqiUFR2lTyP6Gmie1/2eGxkCFV2/24aBggegDglbJgIY/lJ3t4VyBVrEtRxQw4T
KtcsPfweELh1x76YIOR7xvSFLpKOHQdKWYiDNU/MXMsaFu4goFyvrqMA54VolS3j
nh/EcLcXdG5VahLmFt0wU7bNXURwZmo/XzzZcBaA7pYxwGrJUk1+YCXOduHhdclD
L/qC4LHlcELtbXvEmYiY87z1e/1ZZO9F+qGrrQKnk1RMu8SWhAZwS6wLBHd9n+Uw
fb+gbsYRZ77flOCD0Wd1bh91pjJIuxZMmHCBT9FOTg34PeFB+MwlGa60NIkcL9gT
kWy0AZSAt4k/dQGsJnOmFzvSsz8p+2uAsS4O3Q+/obkC7gxbBT4pEdsRiKv1xMqU
fE5rJuj/uaRBFwIhxrd3jRqcqo0EfEnrXdqjOo2XTOEAY2Ke+gB0oghLMKfVY20B
vcY+PvRhfC4vVPwpywqO5aukTd5jbMnqL9XaFJtRzejxCeIexNck0+BMe1hz/1ge
UnknH6fm/7h7ug87kP7qd3eHXZCGXePJqtAWYZiN2zEEtnsyettvqNYGFR3yuI3U
RK90Wups00itvqOEZe6HyLvkCxm7RWEE1/iYTjD03JKh/iXcA0pA+RktoGqho8K3
ApxRM2iPXXC8tdE895wEE3N7gX+mCOGHSQIedBz5I85bZdrXRvSOvXgOtBzFuM9G
k8wizpJckEWjaE3PlzRjthul/pj06L8dunHlIqg4dahsUNAR2qXK0cYEoQ5/ZlUz
6VH71CmTgxN6CsDf9syO07JHsIl1YwOjJ1kn5M02Nnj9rGp+aa8Z88HVlxblRDsg
hTz3cUoXAtasVRfnVr0horwn244u03uym+wqMj5skFN/DtJ2a90WByLXh7EX7kcQ
jLizFYcGxlGy6QW1+rWJYZCOaEPar8Sl9YUjOs9IvITqf4V8wG04kPm3807Ux9ZH
CP7MgHPoVamCNo41wCey+8MJRSY3Sob7eqvgU7j2rRWTnoE7osODHAPcZQSrzsUx
ELU+J5m8ZsV7lecd+1anxdTx+HYVWc+vqgMapvRZqrCz9BrepvCA+ZrS3kuUBwF9
Pufm6k/tceLM85gxuBLEVVRDQy942B7sOedPKCpFkiJi4eTLh1sZTZjwsuGslXax
Fd49+FyWXWZksPq7Y5Z8gEOxrzn9wDnrRkQMWJhAWxQkm2IQROY1IfiW7ZdnMRRo
D2gkFVoE1ANNTL1beO9PbIsO3Jc7cYvr8j1krV5tK08fCsrIWkTRt69dV2CZJJwX
Dva9C7Gl1mcciKffdL/C6ZXXSG7SxKAo1Wq7yob0QVgCYyzgZzVefWDGvS5xCSVm
C7Nz8KfxwvoKBwjx5Bg0IQTsThs3IJIxDv+6ecDB1jOnAgbviSRrJ8kczRDBSXLt
Rbb8H03ervZ45klgaJnozY+jnRv1Hz8p9rZSnGStabk/5Otm9VNYmkoQvYB9Ckiv
8UrpI05jdSEVQJjSUIZIgSsxFFx4WfQ9O5PHkp2/srtjhagA7kt5geLDLNvFfXYz
Av0og1KG1fCZpUKh9LbPKJHLNV2+jtMkkteEx6N4xpxoleZFYAO1/SZBFTU5bh2B
59ppZwK1YEuYvi1FLufZX7V5vk8zf7eZ67l3gkfzduaKrpUdUxo+JHlwzava/Lqf
YyS6fn5RmGywKV+hH2ak54e+P2eTbAm+5DAmj0atdNFVhwZPxJ4TRP5W5JR5KpJ3
GXb7DiQF+tcs/hfS7KaW66LlnMxXlMcXeRZxtkNf+Pmm1lrbOUC/G4Or7E1B7jdk
XRfLD1psijPM8YIEB+sK1RB8Q9pEWKmaG7Z5gTt/dHIEfdfzMnwrf4PadYWMAVGm
lwtdwK4M9iM3gpi1Yl8WIYs40P23xMxuRbs6verINrKGyXnQfbKwEgswS7GE/DQT
ZlmVdjDbgdAAel28oGDVBwbfNdbUKju8MXpVU1neeuY7RdfSlEGjDmLjQiIp6qta
79FkMej5q02SSwUaEtd0rc+XQOCHZEPoU6ikcxQtEYIfhFRSM/GoqUF/UARWf2zU
6lRXlqWNCEC6KINQUpgl5xj3p1VAwbvPPwuHq2p255GvOn31BYrfz10ovaqp2K+S
IWKfy4Sk5gcKqmbvIFJxVjK44d2QkKYtnadSNVhXi+aSAKXwvXjc67u95hxpzr4B
SDiKqjbF5Vwq6iwBMWO5br6fUMquZ9gYhkPpyy1cx6toYpL+50xicdYgCz64ZPD7
OjLmU/nO6J8vOyfmPA8VAHB87fn9yqxy+xSaYoaFMFPgBBfWAc7CRhqGZV9OKKTv
KfpLI4X9OgiphiWjuE76Q9l5S/T+IsT//UqsQqDw+Bc8NZYa4Ac8afE33/wD2LF2
mCmAptZp1qwUh46NICNnt7E4YUDQ8dXz3GPRspwr00OjWbCPc2yKOaVvBYZUEv7t
4/5qm7Jk9iSuiumYqNPUpFHnd+JDHc4TDJC+om2hBi5Umma7YMnduPwArPwcdgsH
COiuOh6IyiqLMXJfolft21qSxTBRY050U7f7TLuDgGeDJxvTpCLOXLcwSfHUrtOx
TnQMcAC7ZAr3OmGXh/CYhBR6KUYJwBjFRKQRODl1LCOgYAIS4uupW2NPVc3sYyyo
SH4wgqf+VQZ0EzdGbIBltoSzfbjt5AbKSB/u9rl9nIYbwJ4zf5xJcaQwxstbVpTU
GGbI8odnchCa1RLZSt1CFBDyU7vBe7ypx5DtjuxwTI1TQ7su+ocF/1S8VJibdZEG
hE93vDf0Fd2jz3h5NJShdvJTQhtsYnR98HcBEFIREPmrZJDtslKdgtmG6U4IE5XV
pKJfJMDu5AHJ/ef5vsZ+NIccaFZyJu78/tfGakbqzlpvkU2BhyXXZ8JHXaYgBe4g
lrjbkKm/u1ky6pocXCu1A4Qoyynxb0Av+w+PLJ++fIPH+xYavc2Z9DIc5M1Jocpx
GLUz+tVNRMJb+7rBzZ8R+5Whbw00OzQrs81Af8bGlPWocZMWHIOrIExlNpXMCcPM
p5ENnbTHb8i4EOX2aGokaN6sfEwVtCmpr7KmMDjGVPoLzfq/LRkcmbTQIctKOYk/
IhrQfUnTVtadcbpIjkPDsmN8QyNVN+OVNldVsuezw46HvQWt4aLJb4bxWCv7VjhS
sHxSzEFE5LWfZwnQH1Xx1Q89R49sddY4tIGwg+L/N5tt4WKXVNj8sUAobKFsfXRm
ehnCCef63ENicdzUwnvkXVCxYwsV4TjSq86a9mOHw+FQuXxcKG9QQ3g3g99Nv5gd
mkgIxJa3q1a4rVhYo+aae7jjUsk/Vdyj9f1kpXfTVseyy91HOtI1oMPMl+5a18KJ
f7a9XlQGr+HDsvvB9/gNV8osatqP8h54QQAGZlJFPqMwSmNmG3iPcOLjz9mA7KYJ
b/7un9Uihhjl2meGy+dq4IbpKvXt5Z92o7LcMKz8uWfQQZ/KKCd8LvozVMfy5+wz
ow6CuvksoXyM2223QurbiYlY27M0rOy4uDIZ/aRHecgN00M6tc4tK1BwQHC9zzEc
kY7k1wA9fOJ/sKUWz9SVx6L2lx65gis4evXXwP4crQjkjYSvrSfWjO5E93Uf1Ogf
bexkcRSNzuFupW+BISUdYgtI0VnWDKTj9pV7r0HIzRVUNnq/5VHsRLv0fb+UN0V7
BnM5ktXPB3v63EfM8BZZS/MNIiHubr2A0Z8cw8QrkrvTT1kIsw5sLWdc2LJU5QcG
dtTLi2ICdRcYjbziAl4TdaE0CiR4AaT9kp9dSa8U7WGWhhacPcCzNfOUJtvo7dwy
mO/ITDONifI+EPUAsjAaC3nVPJFR6UqXWNM21r2j7FCjIPob8r7y7Ivwy0SnJZ9M
SP0g9JVEcCTrUdC1tALn29g+Jxzj+dVqQbXlYxf2E1wq/j7DoNw4hcjys5LkfbCu
2xxZ20o4rMLbjuYjizGmAYob6oRIzcfKhnxQ3fBsNyPqeZTh3iP9qS7SQ9M/DgSX
oDasgRERU1tMNWZRgLUHUgErKpIAmMOJYMN6swqmc95dBYlFKWu6C/ue6Lj5zN8G
wg3S4ejh4ddgkewZj95dEsX5g6ZiAeX8fhkg9cJM9kl57/zqTOv6i/MtdUotA6f1
Z2M4jWkBicHi1LsYEMYCyIZWWl/qA4I9D2uoha+Ms4wuyAYx7l7/90XaIswinQDF
RUjGcCknAXFCz7BLRy/dYFuqc39h+8U8r66trXaDQIUf927jFRSnp6Oo/XQcAio9
HIAPUPmBDX3Txn1zlKclMcbpRrzvM8wLipfzntKvzcGREZhISVFkqFZ5yGpBb64a
Oku7VQ5NFvdPmNn9xwrhNnqI8RyoXgMgP7zYfokqTNoYtWGevsekvn8++PFexFrk
6VOyZ1j5EMUNONJpPikTOPo3eiGYGCDHs6VDJG2tBTD4830BG2rTZ48xJHt8+pcG
oNxE1N8wVq0bKXdRVXhybe3IxWYagd9qwCux9yY8/mesBdHx1O8SdTNdOLER00rw
GuTmKKk+HE0esc8oB4YBmZyqGPH/KXy80fk9X5Ib01WfLi7ID7G2DrXpogPc5imO
xQvzLCKqgyXAEUUg1w9D/yAH/yps6iOffAXC5wp8r35rPMELRsBPRQ/SFetfBP1Q
rwEIHPF3ezSpRAcOHOVbn9aUm3FUGXkgt+IDdqi2XqAZb0LqLlscCA2GAHUmnZVr
XBKDOzOBtxKK7xbIBJwL9Q7lC3ci3qYgafhliphaysWssc+aR1bVa+mV0XJ95bz+
RxyxIaw21eyTKimY+Cg+vvEoNS+DdiyPSOGYNLYwtmJsPvtjsk34LD4EAb/hPRCd
W6BQ9hbY/SyK0eMp+wO8tqCLbs/WXT4FObAx6B12pqDQYzDlV2JMAyqgNWSe+QT/
c8QNFb0cCx+73Av4ENnACbz6weLos0BfK1qvaLs8+LWxSInT9hVNrkBPD/mEuaz/
hflbqGba8QLeUFS9Nf0vDZjF8ecI01vPbDnyHj6ICY9lx7dwBM+UBaGBR2I2S1yj
ReLs07FgTLY704vGNnROD2PQneB2GdWlGfaelcouJKoqKvZDLsyAE72YlXl8HWzD
YQ3J+WtNokeMYkf5fRw+gEWGAkqUuYuY6ZzZlzWerhUpJphhPelQhFGifn0DrtiJ
t86Lbw2cowbotx6awUh/rVDaEBzduMQaGd4FTVUrX59UtGfey2FiHG4GDt6BtB9T
NTgKpPdWaVtcESsIz+I7qXV1+DSgT5LaGmjRWtjnGs+rK5xDk9YvrCqihi/k0O72
2F3lyFSthmKyjtv8xDvrI5Eq56IygAGh/9beV9tVc2dQioavcjVlw8p6V97Qlpec
qcD9Ugr4WSitl+P6FPpeCPvNbg/8WRQ7L9oa3Ak72/e/pbwRBnVu02MARUhP0fk1
72H/Byx12DNOGYWemejxKWhwv8HQ35vpp+HeQl5TVEiiZjeq189L4qnfBevR8wIi
x+uWwGgZJqg6RqR+BCu6ufVvDBMqvVKhplZLcFPJarZG6A+xEurc672QIv8uLLo8
mB7T89mwoP6jEdDPvZaeH/XW9wHJhKn5la6k0O10TSQgrTx5e/55vggCBoNbvA24
TZTB4TfHaMJwWTO3Sscs+2jrvvFmokygif4/vNDzbND745F/7Vn2Hj4l2IdMDDAs
J6+WcxQiqBes3CMf9dPo01AQudr4lIBfEW0b6LnwO8WQIzw2ju8lX42PjT7vcjDD
KAoC+FR76LkmhzL0B58G2CNsuE3f6kklRq7sKXRaGR4ZAB6jXIn46ietwVxQ70nS
2lWX36q5KeVQQZfii9kOsDMXpI05YTX3pd8XKO+7hI0ntOdcY4YoMvUCR3WZhyKz
hYJUK4VM+0gFTteN3sOGEHwQLJMj4uE/AQxgv4On7kjN/7QeiWphyfwK0kOBdrq2
AQMZTm37HHe3klYvV9GwtSZE5XJbKZ4VfbqFT35e8c1r8iZZdMyqjE/rgsyAioMb
3U1zgRJ2vwYPFmLV2BTb+bEbPouut0261ufBNqJ/dqkfNTR6A2nRqAaumkenhhLQ
xcQKfdF6QtTX1jIJ0QQB3oZzv8yMHD3NXVgPCjYr5TiW1Hsl49VYjmnfMqqIZn4m
KelV2mlRlNXVpcVQeNC9VxIKRT5Y8MX0bGKrND0dcEL21YrIcK4ZqT8eIuGuHUlA
PcG/PjlVHfp24bdMEZJET7sasmHwwS0cZWtXbZ7lSuJwjPJ7O3NssO9gF4XlHQ5m
M+8EevFG3XGt3cBok5R3+vXiXt6qFmbBWzS7VWknERox6HQ1In1db7qksFfmqt05
sPs88Cmx1ocGqsyljDAShP3hvAlsOFnLT3vzwxQkArxrbY86dpfhpeIPKgy/SWQy
1Wt3HVzJHsO99ppbodObDR9CuZ3ABjvPd6ZQQiymnuP1WMjIcXeuoG4BvLCjHQdt
EAf/hEvhKSXqPjz1muhhOrhnrwFrsvjtrxxoy3mKc+SnlWJ4N1Rz0SiCi0nl3Fha
n/N989lmlc4JN4KdnBeV5llT4ViWgZ8sTtr6fHkQ4f/OXVcr2fS7B24d1HXvEJYU
FjTSZreIWa6ZMCAJlh1js3hp2ORBj5gVyU4+XuCxSp21KLVLaIWOaxAD6P0DJoqg
Y8NIlSEk83/yQkdiEQnwqlW+BcUAJ2J2qOWAPND383HbYlURCS/bW0eSGDl5vkCR
FymF6KeqFD1oOqfxwKKb7qDTdYG3Xyz2KsqyIUY9RByWfnNCnoNNnBq3LJ41f3dM
w+7Arc0Q56kDdXkE7HBTDUfihCgCJlpmfTC/CAxmrB/y/eRfAqFLQqTgu6xZWkuK
FsMG453mqm3cgNDFWGBJQz/myxezvVwe3m0bvM9sgYr/iW7G5jtyZtZXDLoXK5ol
r0VgINo9CMqyCVQJcNx+AVc8DsqdGfZX73jpKPDbTwhSoj6kF97prH2TKZ9UiQaY
joMgbuv19IugmwBNBx7N+w6US0DztBJWT+Dn6qU3rRZEgWXFEpTzPpU7n+/p9inT
Hma8OfqTvMQ7t35ejCGRETUQ1u7FlzI63rrfQFoqtw/6WYN/BndTnmmdIdq0EDmD
ivm0CeznwqX8OO/9g51ncSQU6sYuzT0X3CaLvPp71svOavovXo1PjS8AUzttFnKz
YiDBqKLE3T4Z/v5AJ1SlKktaaGkJdjSVRcqCHIrwLjlVB7KVvYcyZ4hgHsfqQiZ6
35c/GICIIWiSYXJxYMRMi60fFy7EWioRlTNtg+CCj6FssrcyfFzFEVaW9z+sx5Wm
/+4csudikiSiTvr3hnxyg7dlTKJobsQzqWLmp4ZBNKG+4WVobhykqRx6EmO35jBo
EBOrJjChSNtwnmmx0uDr8NV70vmY9bO7kGCTFQoT2ph/YgKnV5tFqzPdf7SlwWkI
uFp0DCCrnC8uKlsmcygVyQZtDvQvp8j3gq0RL31RQOaD+SNVo4OqVsic7s013c1Y
BaXSqyelENW3JWjL+nV++elDMhaZ8Bj3LaqHruGlNITyCAh1yoWfYkkVZDPcooiX
sIRc4OCsrLZUA8JHlC3xiru6RFF8Q2Tl3AUix7kzAPhtjcW73MBpV3zU4p/6DtGZ
yG6ysXl/FdDwIFLnxSu+xxenhdDKvO6gbxpY6S1PdZGBFJ+UjsXojb+Jp/P6PuPr
mEH4rOpLuMVNburNd+blLQDodH9o5Xa4GF3/feu0LgdvJtthO8NUNfg6KkKXZJek
VsktiX/BqRckiMknsuC+Njretyw9iditii5S5XkXhaJK9kd3Pl/h2wWZ1L6pruqW
yViKwItn80YvPOPfl7NF9eTpok1/iIvJtDrf60SSjZPtuHjBJFY1dhFkvKbP9cYp
x9FXRg6awAGcsIbbAynuOb3dGr98Y9bt5AKYYrelmWtYG4+ahEaGLCHWFsp8a3bE
evQyEIcLkLZvXe+RSvMJQhedTbJU2m7jV/DHcN2hpJj1SSPLquOFZ5sudA4ZLw4l
HWilSvgQpDBsIYsgDw8kK1rfRjgWsGko8YSymZUHbtZ/2eEkmfsIWbXWruTJrrH+
r8VPRlZStcC/mWzyhwDL0ZebtPEh3pFLh/mcs4Ot1FDqZN0OsXZQI6kkMxWt2ckO
oRcajTkgpbk90ejZSNYqlIA9Gh9DEI4Syaz4B+gkdv3fh3ZaiJYhnAhEjYzCMkPp
ybVTYAtVWulWQwpDgPENSZyUt2aHVkF2VbVt4kKiZDYFz5tO4G/UFTpis/QKqGKh
IfG2SDew68ThNJIAX+ImuKR/aV5H/+0FmMw8soVrXLvDgzXBxSpqniNnHkhQVD1+
H4i/BmI7FgMRla+NJrOH55F0aAwaWDs+xeMZ+03/mwnCiq2zAwZa9NJD99LPhZaV
HCSEUo/jjqHzHr39cs9idNav0rv0V5ev1KcDR+aIkPchRkQBz7rPwvpHtP3gty0u
ZD5uSd0wsobmWyiA5eRamTeDMEHHUMDycYNA0GgPscNA8xlUsfExwAr6itCneFGi
YP7STLe2XlHwFr8lQSYNv3nVdnAgyE7FP2gxRb4HyoMPxpUJEHZiRj4qNQBCHpSt
jOlelpaaVKw7lO11vBE/bLFwPPJukuGMwI9zO8I9yEtLEOL/dtnQbHmsZjVqlwCa
glI8tb+ezVGBwt2RaE2QEh+tNNlWy90SQb4NY6VWx2pZ3P24khgqKxYYtY+PZq48
W/TG6bhfRprGKMRgf4oFUoAyGWF4emonIce45JFcpQ2xKJAUZJBhJQlnIJPSLJk2
ZCRJqdkRDTlnfgMYs1enez+MUy9n5Tc+KBEoFqyrLExE1/NoKX3+dqxOUL5EJ1eg
vnbPTcLrNmdbqSyCBX5EmKqwRGsHgw7XjeuZQJLGj5AMBLc9cqC77LhfRQYGDPps
3qhQ5kumz9nLlyyEpSMoDox/rW0SIZlTdglnv+6DDqHWckHLpi7mCequzQj3h1N4
EJPpn/WGYNe8OCbORNTmLQsP8NXb3GgygUhvtlKB2ZG5vFgMxb5E38gbi+EdfZA2
lSp/CTvBes1msnJzRw1hwolfWuJaCmNbnKdAh3ebjjIxS1RPWGYpy/8KymI+PQg4
emGsXLuMy13DU4DttFhfljmZET1/hou7czJTBhwuwPBbKT3tEy800vOjz44roh5L
eIRVU7f6Rtov8zH/0aopkfBcR0eodgN0bXevXZCL9oKZxdzha2hJ3F9NNNQo/EAq
7Xgo0vZJERTHnR9oauH1/Lfmo7X2mCvHGpjJoFf/S4dDmvEI0mnUPLk+E2gQTZll
7DArj6Xw52mFmioI92EhQG2TbcXGZJtW8gp2BGDoOlyS6XM9/2IAiVvNLUh89eet
oraY3dDW+SgGBVCB8aAELvjUJ6teC2V839S0it4t0NjgN52bz7gZT86CetxmZGID
xhgTliX3oR2EjX2NkmtU0a1g+UzcCknAE4bLdLhKcfmjD6d//xxzfCn66LOYaIlr
DHA7k8AhjNlfEFqaz79ud7tQaJdT8NOS9wt3H6vFlYml6193fmoSfrWsyEzaYO82
HtC41RaobTGT/8Jof2cx+4rf4e0Okmv490yOO3TAPlzS7VaLfAcQUAKWv3cLdc0Q
Thkc9kNe4tiDs3pW3P8pUautntRVMIDjKoGsCkWPup3t0ZOOffcYJfEkhHDPNBEO
CUIqg21Z6SZ1kozIluG+sGF0F65WWO1jJeMYLuoUtMIJwXJ6lig4ZfZuCenf0vlt
8+YFUP8vf/HDo1qFEyRCLRxV6l5XTl+qAcEyH6/eeyMqspmuAmmhu+rtkm/iBF0x
YTUTY526wE7+GwfXlZdNIUcGa8DRwzipjSYJh59A2XeNRMGJJ8q5ZluYlO1E4s2I
00jwEM86Seb+xO4osjjIzWQCPbisALiw9lmYldfHxw/6/HoDzBKfp6E/+/NT27qS
Q/dc8qj+fi0btcgtdgN4IGejIz60gfX744HfmJ1SDmvarFbmt8cAv2+wuxqasdCg
7xzAO3sBlyNYerCFSEJ6M3O3mJDQHia3DUVsfW32H00PTcJPZDQB4L8d8+H49Tc7
RGLEIgG7+jMUIBgp8Rp3nMKrPkhr3gz3JcqiBW3ThdRcN6CE2wpzQgEU/sO/lNTV
AW6aTq+y5+MfIYP7tKEF0CP4TdzSYrYaP0n3s7t3viI6Z8560lb13TcCktBqH3xF
QDF5f5Z/Q7pOeJmN9Jr5KbEy6O5qMTLMp8fzRxpetOc3hnFjaIj/qN2SI3aKitC9
wQsWZ4e8d/vFOVuFQPU8c3ycftl4N7AyDRFItx69PajFyt0g2o3KZ7rxm1tuOomD
BUZdUvfb5/Xbguq3WFGm1gFmVr3xFEC9f5VqSoEXxmbUZ2PIRrHsvPVw1TpTm6nK
GeB+Wwh3IBiKuQOyZDuG59pZfBphIp7zCVXwtcKVkbldh6dgTVplZgQYB405BlQP
wMUsMm3JxPG6eZWYZCoCCso/vg1sFkQTZZ3ENPECJZxzm9kcEbIW68MhS1z0LUN1
XHwKns/Dh4qkJecj3ZgHkFbcukdzJxhh3veT0gk3+UdF0Cin39qnFVv/eJ/5uTqY
u5K9VTCKvx3peDYdutyM9QL1lt2jaFepuWDAp5Ps3ohvK3ngk8gkzNFHWUrE8r7/
AP0nx1bmnf64TRRS4hSTiQmS/WQxDK35SHti9gG2cT8kTYtBUZPzrr69T+aOrKX3
EbdiF75cIOfLSyPyDyldXvfvz1KkfAwscBWzlzpagg1CI0bsPnVWiigMc5oJjgtD
URgSVghlVx6PJpsBfbkjVQT1WOW5SdP1iyfe72jizTuc95O3HU3s12Ti85iRji+e
lj83U5uMLV3O65MBL8bB/dlqGbX6OfH2snwePZuGRGR76LswczEi0dyMIqUC56N7
FeUHO+HSRiiqM1jCVutRMMB5MI8FiWSiYr2neRA6EoJeR8NRG0rz8r2fqdb/VAoY
WFwO3qlY/pUpFKYfHpIa/qCin6DlRTBKtm22gy5Hzgp+icEKxTU/vcRap6Pvlzmg
a4Bs6CuKdwejdMcNjlZbVG8olgK4AquSSXaUNNFT+1EKAW+xWrmG2Z2g16DS8zUQ
nZgX6WfdoHjjgIZMM287I1UuqoO1FwVypyhbccqhBSp8hcscYxEUJyCK9exEdGaa
LWufJcFP8nOQ2ib1nQM7OV4u60fxEq4gsosjYWu31g2S1WxKBvyGWvi1t27AUnZy
uSmkdFrh3oxHKmqFpw7+dVgvLSshbKdyWbKxYpXl/BgT1qCBovPnQDiGcPCVRpaU
XI4/W99uFutGkwGhilFHvMBI7LOEYEbhVGtY3SFHrPAci+7qrPvwvKSCkN58Uar0
aPHqvTfeHucuF478yZz8T8DoxSOxPBkgnLwOX4oPeQKI7AE67cipsUmP4h0TcAUm
86capSVOa4DfDpez23/rWM4vClh4CjIpU5pPreJN5m0zTIp3BADpx3EElWkwqSB9
P2Ja5e8243wk0fPs5ojbWrqDoZ86cDHxLwebpBr6sA+u3Ibhwx12nBpLuW3/D8p6
Vm+y7k/7nGo5ID8Rz0z+2dn5YQaRLqS9fsAT37wbYzij/4VxAbKT7D/d6Ehfhxo/
Zx5bJxJTzZadMJWJPkKJmNZWaebHN3U3QTJRpvsygfJkFmtHW+6049DV1zEHHS08
W7lYxySk2om65W2nyi4fJkeD2rBvbrv8w96j//RmTp/zrYA6oBabRwNVrr86r9pB
5mQ5O4dEPAwi/1Kc5a9UrL/mXbji3PU1WKaQ588AIQVT+krj7KtIZZU3gYto+VM5
f5SqMHIHgbgI+4snXBIJDOYrbY3/dNlXugDCJqVCperJXwY/uZ52Qm5ds2V2YlFM
z3fJKkLf5KyPfzse/6vXThFGSCCU96C4IcsIYETqEs+5/znD1R9Kp2QY2/O1x0Wx
7KaRSVnNRE/etllbrEEuuhZ4H5zlGjcj1RZj/YEALEPwKmHHl4VcCZPPDZLeAQwh
wdRrXGo12WvWAup316Gi4jgLLBrPqe7fiIqtxyziLPYuL3A2Je/bb3emaBFvgZRm
DHTHqMZ5blZWib2iWLtbkThmOj8mx6agGywAF9X0pQMYX8PQxHjTJW3B3tYTf2gj
imffuiHczZ3rc2cfDMdx1G+g6uCzCEPRdwCfCGdz4ECalLNuhVbr89wSp7K1PhIp
bs50Pu1IB3A6B3pLSzC7+nAYMRZTBh3SmBAQDlebryGa21vztFWdz3v8LiyRwUE+
PtOShGyDN///svHoZGolgUHhjMaOKVjcPCOqdg6eMTS1GjdHj1MVJvDocQmgCx7f
lRhaE5vpKbrNysv3RDrK3ZYdio6hGqhPc46eIuFGbW7liSi3Mq+a1vYQarokjoCq
RQ37ZDkqEPkXXoFzAujcyQzdcEFcc04lKlMtNcqceVNhHlmEkY5LKRqyVOX1sVgU
Zx8Jf1AHT1Oq2Vs21QS0DOv858ijWuTYryePFDATBL66uWMo/ILbIdn4ggU9pQYO
IM/S350qpdBo9miZow1tajmRy107BHsG0FKOmOj8Z/xLqKtud5+eePM7TYTyX8RM
/crkqzxSxYjc+d/JFEjlxNnolmHpwNRRYDEN5gBVDc9KFA5lJcgEVLrd6JciYhA9
VsIOd+rI8bKuy0FKcyTJ9z2nCR1hH6Cthr+woWpF7Tch+G5lzUxFJ3DEPOYjcad9
HkMJxlIerdKM4T8n5ycCOci8m0Xj+j3Gye02SA1TiOFm+LsMvIFopbCFwSsjIV+t
Lg8YUSIcMudkrZ+BzeCrO1oEyqb2q+fblzZaZw/k2iu2r+ll7/b8WQ+bZQBns7ME
sFnpu1MT9o36Ks980ZsJVLMAEWv91dFwHIox82NjL/l8/L/nsDdHH6LWA5E6z/uG
N5766JBP0grA0b6XBRKBnHNXv2vpbtcJNLm/keNw9nhrbnq7MjJhjMZxbGB3WrnD
ibQDo0Rf3jHrsWp6WZW+j0hfr74W6b5ChLomYQLi1VbBSaz8+Ha8CZ+1T4Eq3rf1
q/WbkCOGB3TTr5n2OH3xmcIzfKS8Ka7cWgHQ9pyIRat6Q2bA2ZvZCGtsV6FSJptW
aHVR9N7hJCuUqc3w0LlLASq1jxgnUH+gHQ9SX6yf6M89+U4a9CMnC5sP06KnYgIP
xiZLuHIsQGuixiCnRRhYKOKILIMC0ZkLjZNiTAIHJYqpKCHDS9SLYbEZpvR+psHW
zZRDOaUNtQvDYoPDXpydI3u/tD/VVrjFQRG91CJGGR8q2jUCQjw0rOMAe8ViQj67
zXy71Rlakk83YHdyxPYYjVg8rhkB2ezxOVBimHo40bHwgHsJKgqghANDCro+BLwq
xYtrpmZ4rvriFLcgimlT71D1TyGrHhL1kTS0civIyBnutlZNskdFvv+8zoJ8Elqv
Nwl6V6v3qoQIO8NCyKF3W1RhmED3MC0d7h8DJvVzyjU9NiWfyPZtM9Y13Lt/73bt
W63jaoB1pBSFQmEuCpE3vVUyG1ZiYpuNujNeXYe8daTTa0obKw4wMiP39xD0pf5B
Cljcl/P+Q8gdZIG7wvUk2HboiB+Rk9IGp1sx36Hb/Q9rC73PC+4IrSTotlrvDSPN
ghw63Fw8jsfpHJ4TUKjH/gNQGy+L4lpN0L8ZERcoxqicNcKLQngIyc+xDecg4lwv
7vHHmYD3qxP2n9XpNxHYI5qb3mddCVs3ICZbgUxSvYlc1ksqMd7iimlil7RZKXSl
jMxvfDEPMElszCjv/BURxtFuaEHSgM0hsGF3APD7Umh3lcQW7PgrpcuN9m/J8kVh
enHRXz4Hi0VGEXDvQgXGqqqNyfzBUHg5uxka+xE48zV2NwviMfhwb27PHR2i8lmv
DAhuf2UOCKSM2CnLH+QmLmkMkgC10uZ2jTeP+Koo0ue+tXMZWR1UaMf7vWHzqzPo
jAlszMc9cskqr0ACZcA3nqzlCVA/HEbwPFu61mls7L8PDhpVcWCFJ96r698y80w1
HSxYqCe4rt6tziGyC+XyVXV8/5XEf0LOXgUrH1J0seTMUlGktt9GN+x87PY+2B7y
C80WWSuN3xLjI/H3LwzuLWPvlpNsoCKH6WNlETrEVPgiBkmvL0MMmjmUaaJgp5CC
fCHqd5WdKy1CXdj/gqChCzMRpqAOWzvX5XyfXnhQuG6WXKntnzl+CrPabHQOU6oe
bMxW3HQ2sJLajLIMDjfSRenSjmd1HalDrzzKL+4pJ6IvX3MWyJOOP7kkPbRdA1Rg
YrsE9ioDDhLnqRPYMp7ipQGjDB2b3WPwMhF/HOYKZ5OL1BWJrqfXA+eOgMmNO+sb
S0FfrGW3iqGfsbW4mj3PIOXy1rzWInEPxFlC0TwkLwNlJc3rhRpCzTqS6u+lXo/2
4Tvh/L/3J489emMo0MS1mHUVYgbPTxKMuBGjB/ArAx2KC8+OvmGtyAkpfM88bZ4F
pYHJcl5MGDX8r2IpkONBAl/FprvcxRf5y+8IeZYgEQGnk+zfjxAvjsdKUoYJwxjM
2dVJa3oYvMIi1cmwWwkKdeiXGNArsKw1MriTlUh9i/8XUvzxZkE3vBjzlF3S0guT
ZdQtAURJtKRNMXxQCdd/SBeG/mQ9lOIEuPsDLtSMXIkCXi1t0SqtvmEVnH+Sdy3N
OtT+5ObOhLNxlNUB4EBuvGXTJECe0UJ854xyNWR97CwvHEXTfcpXqIzVCFK2wHyW
qexCxx8oQ4PkIlv/OmxoC2g9qb9BPkwEpn84682lOFJa1eX0Q31+4NihSvOe2IXM
C9SQ0YQxtzjXOteUQtLyxjxUvqlO+OB3MgExg0CPPQQecrNpRYFTJp4jjE8GSQAT
km/HRR5Yp79EaOjQ5JX7BRzecPcosHyUOfqfk95bEdkjQof86Yi7C0DIG9Eb7ka6
xUUSdKcsO5W0t+A7LHFXkeVbSM+8qeW6ic/uTGOL1Kpma07gtIU8yMRtns5FGuq/
dHY8ZkQzqa61SgYJQ4uZHFBWKd8ylHS5zp4b3STR+WXg2ymlYH3oEjGDElR3zBlk
vdjrY8nSic2q53Vv7IHeaAaUGRmB8iV5kCE9PyS+CWOJhANQ075DjAyCTxHvzsJ9
cvO3MYAI/pdLLcJUYzRe80ehZaLOzzAJNZvhNQlV6DdH13kfI6kRk3oNYyS2FZt4
3pK8+l98O8p++nq+hcPnrogXf90zuI9aK9v2287eFA7vwiVKs+qRkomh0osYJhlX
G3u6pFLea4Js9a7/hjB2mUidH96/MP3HA1ipQJOBoLyfzL183upta+K+m4GOnegy
VUM7mV6EbLepClFobEKoWmVlPRGlvofuKepih9exMOCGu6w0iHrt6rHx4WjRmIFr
KQ5A8DGuEJSPWf7d87GrGHMKhlPhvI6PBocUqwty4jQmro71+Vkj3+RfrZj3/eej
N9L3dVzGJhX3qC886MY3Vy7KCCWvzzfSH7zyWWG94iGs0ykg1OXL64E56cBNWOUw
XIpVFCLSXIUNFMpN6wpTTiTkpwsIgKRTVg6mTcXML9REBx0mduc/48no4FdDGCEP
y1S7+4T7wF2P/iRC0TfJvC9Q5MCPcsTkAZ1ygHzZGOcwNwZltspa9MgJFuCknAHE
gSzSQmbpdh/g12PXuyha7MK6PiUO5D0xc5YvR+CbihohEyd7YOLZ8/d6sN9WD10O
pQDZBk8z+qxUz5otcNhD/dACGqnlXb9JP/R20sNhZVM0q7M65byMhAt1hw6mUjnP
nNu/DYgEQskAfXwT2An39uhJ2QmsUYpoW8BxqskFFUAwkUSSrsgp3l+iqfbljwkb
Z1tNzUcPVj/TTPK4I10E0+CGtrNhkM3jDhooEhD+ahlW/DqMnieM+zq5NQ+Dc6dJ
lK/d6VQbkBg/J2z+lV81/sd3LrkkX4OI8KLIHBBJsXBb4YvMW1I1H+JxtzSv7R6/
g4+W2aT2TSwKsh+CQScP7wTWt2QqpsptCB6BKK9zj1SNb9Uw1VQHB3W4EiIgJ96T
nDzKJ2R7eAgM2Y02jNrdq9N+GS9mMlIW9jnP+6cwXRQpnEHf1o1Jp6VR2xQkIjGT
jYvyhiFM1TMZcsuFEqlEaTWYWpvOh548DO70RVvtj/u8yJOlYhgiUgZ9GMYwM+4K
GGhK08Fs8Ixkd6MW23aNSy/5Huh2Jm6+GO9qyiyBft+8VRTbK8dIqLvZpxRhAk+8
F9crq+egjdtElavMzczBW3VmGybvCwutOVOixS/GtCWYWuiNL+RwvJIkOgLWlQMm
adDqm06BxVRlxOlB6swVmjw4c2D1aeuIDHiZucLi/IxnSEu2Aec69v2o4G3CIKb0
m24A9LsLBNjTaV31+6bgYzppDFPAqEohBb7KaAA7OXi9QndtL0lO9zUcNEsQe+2u
UoQ9nRfqNorpyP8B3rGyiscc5uXUsAzpEXYv1x2IhHs3bl+fauJGirMQ4w+mOKQl
nOTwLbuvNoATwucjuHfoNz7U86GXiscgpBY02wOb8ihghbzfg5mjgOR3q/m4HpgN
q1kVCj44cJ7BIxcNbeGwVYbyJnzmGOtyIfILWjVD6T4QXM6w2ybHsfsf5sirWzoz
jWg0/K9BRyHaIG+V/EsfDE3r3PcPaYpnCOUan9UhVCF/HiBYhXwHIY8KjuBdkj7p
bZiqCerOGpEs3pwpZ9P+61I34h0ico4ykf7ZESMSAmY+LP/L66biat9imwhLr2PH
TIn54xHdYg8rjnI1WbR5JmfS+WffWaFo03unq1EEcCeLLzBf8GordT0pKarDzKg+
3Z2DKNMkt0M9NXbxiWWbsAliU5O5QS3VF0leGi7LgIwJzaoNH/TF2xDuXTzkILvj
awhVEU6Ns95Sci+4+60gOzOE1dWNAX6WuBaWCBANA7eEyv7mLMOYF9FSAgcU2yOG
qH4AvDKD9YfcMq+/Nqa40u1aARLtPPeW8QfVgRLaRSU9nwop7ilPllxrSUi9MSVg
faKMD0FniGNKpPv6GC7vH733LbnAuV/qg3fftLNlHRkaKpYkXyhkQnGtL/dMDPl9
ssKz9SAb6As6tFqQ32N88Jsu0aZGWXJoZA8I+GXv9xmot1bFhFd5EQdRoNGARtJb
vJouIijU9r5XDjE23aZ2HFBd0Vd8wPKWtLf2eCSbjatQ6aIw80eYSHzFmeOXQGaA
Rl9qh0P7O2TQYQB5nEYCp7PuK9EwuJDfjtbEh5A0j+VnU4CFfYraZdtiLMplEN2E
lhoEdtK8lNDHztKkWjnJHtdRyqzv1PLhLKohokrKb5OcMPOUliWGAjWPZ35iOiPC
Pt0xFFIGZoAf0nVm4SbMQmPtWaeoHayN6yRnouNBO8kQXc+Q++dPPa04UN1vboIO
qQWUyH9ORhzIQm5iAidqDG5CKvNpDQ8U8sTj1mvs75iW1YSZimRnIUt7kR1GyNck
PuKvsEVTYATuW0ezB0WXtAGUzVQ6IW9kKXd/5TO7kVBCtUjynjJ83rJyEYGV042K
hjLUQfjqOFx4BAsO5osjmqPllO2NOlbpgZ2zfYRkayzE5YBBXVIbjvotkqxD8r2m
kNA5GwbwlJUpx3858b8VnVieX9uN4v2Cn8gy9pnzlTXr2PFy6fapEATYLJY0gh7A
nzB+IjKlbHS/kqpIUJ+ODr86CCWgHK/ZbWkGRYIljG2usxUROpK2OPZGoN1vMoLl
/TYxO3Wu8JTudairapCLohHlKP56airCBKGfyIKLneCGjqzhUxNB6ij0467GXHhV
tZg0ckppX63n3soZ5zDn4C0RFHP10UjpYVW9kgozXaQrgnLZFmageaH6KvpH8JpG
8WvZCYMBqTXZ14ILRrZFcJhNku6sop/iKVNzHMIq5peAuQgvC2sogCK0AjCPwjRE
nHsYzHNXW7bM6V9iHaOuKg4p0WI7Ong5Xdg0FxF1fxg9oK3ja5Hojlq6BnbppJhr
5699S04y8uXJGNXaP+DjfhW23M8RHxd6xFJv0hDug+1arIvKkDuR/JD8Ts5VjUXi
NfKGRgHaOnkCy6YY22+69f3O5RdjEGPb4boW2Ig4AS/gYY2jMETTilBMbg+XseT5
cs261hHzGXhiYQBNeqAQ/9Az2X4htq4Ke9Kw6rumQIGK2hhaDxcq32Um1TuafJ1T
lCmxym0zq09wZ/C36PSi0g06s6RFdGuSmfRkPGuTZdJqfvralkFX4Oer/FPID8Rs
4ieCpWaT/OVGZtT2Ca9JdaqLMyvtn1DHMVUEHuCpfpva2koGBLn53nIrM9uWnvvo
/BhGrBTbmxtu7HlF20jiugZUkFaNaMfBMrwzfrzsmSPse+QfJG2c9zi6x4c60N2p
TK/74disdVEAiwTfqEu5pOYrBS2v3TpDpTcAhDMwB3cDgLi1u73hQ8TfFT1akt/U
VigdsX5PVpUCtoRWRNqXzFjDm5lnEOMS21Pj1SSXa8lOcKLJuM1JA8xTRbtQ77YR
kjDFF9BvBEGQglIC87EtqGjlPLQ64e3U06hUDS7ZWTT3aPIQVDIii00fNmkW52IN
b9He2rv2+Fs0DPlyBDo22uUAfVMy6bk5ftxxNaiRYq/lvC/piD011qnZeP5nz0U8
7JN0jWK7pZOSjeQ1e2htl8/LSL2GDPk48yN/OTL4qOb/p1sjez5LkHxwOyomSSo6
I9yV5fxhUcuwfh+eR66lg59yETybXSXqJtIkNHUjyy76Ouw/AjmrBAznl0lyT1sY
auC9hXZJsb7ciwirkVT81j+JO/wfoodIbm/frGUAZFNU/FBjLz73bZDalRYY982X
17OVWTVbg66qjS8IELbXHp8ifedtFXgZAA/jH6421JSPIadO0JlE/iUpTCbrV0xG
bbGZWhQ+Stea0k/ufqRFNzIu/rxeYk6BxPnnmRPta1OMCN9l7Gkt0sKxbJoGvGCU
Our3OnDUhfkyfCNNbIf2CerY/9JFICr7PpkkjPJet6CiOenHRARVnNYzz9qENxI9
xxy1kuo5S096Em+k0Gh1cEN/BezCCEcJl8Fwc7fHNUH9hJWcGcWKOgbP3DNNLnNi
Me3W3XCP66IFPJ5JLNxv4edCEiAOV7hYd8Sy2UtJNfCQ4GiO/tDxXAg38TChKU3u
uE9NjzZtV/7oW8QwN17bY4Kivd9ONL3Y5BjfEWVmpfKeihP8ONJSzDVq5OQsnaKb
ttkfTMfaKFS9OTo5PKzvUyyHerx+fE4wV+fNqjMZbjCVloGychtSFGMKx6hnTIs0
Jz1SJuXt37LagXY7ZWAw5MWfrWDMIU4KhAicr9GajfdPK5aHQQpstkJK9mTwF1Ef
A4/NzlcIIcE7W5d1RHWqyCQ7UibyszJe57b/swWKCIjwD57o7PSkoUFa5yvWIsQO
e0gaxwCrZUUKAHmEZWCPRgW+5UQvGr277TLSz7NCuDLYeRzFRXikp4rBn4GhOMn8
qvFZFdfR91TuUPH2u3UvYyD2BhhQGnpnAycyewTm9SFz3ftLyqegWBTLKq8A6eA7
KkCSlCMOsoc3VpnPHsWx6XV8lSmwG2rH+vrnZJPcKn0r1TD10Ut1auhoIz6V1ewT
BWDFD3rMOlT+9+8xzlySl0x4m8EPabbvUqeltgA2CVNS8DrCR+p4TSjmm14zDcTs
lxSiRaVMPo0HjBnwAA+m3++Qusco4ig3J5E7YdqRYA4MRxw80aJk/VSAWLp1YVZ3
BpAmFSvbauB+awYC5Uxk7WgS/VTXchh1i5CxCG/dwgdEpLBFF4KcalQPrw0Exjtv
3E8qs3YibLQMsjTkAQcZ2edkfPxjFG9yBEFPtiUaRpBFdu2bPvawmZRTb8050eKs
g93jMqDyAepbUIlWB97cdci2t0mclEI5H0KTmMoMevUa6NZqgOB9pjJ3ew2ajq8d
kJz1rJOCgPfBiQfwnvFbqeXvNnjrVB0h7PsQz4EzmefT+6dIMPAkKGGke3y3L9ec
F9VWOtQeXaTu3c7Rs0bwnHuQSclCR8hGthfthskMHiKq3rzbDH7DkHVKeptmEKOz
Ep5c6h490Q/5nbDP0md87P+va2Rsu1AAeSzf4ZsysAZck492OpZyCtVrs585qYkn
4U6YKciVJ9UEDRkOF81eKc+TmMRUjnhNkjJT8iuIoBFVoZhVANI2jBji5dcNeESU
/D/0b80NJrt8AGmX6YR8kdqyXBSVwtAkcKukqf4Gpi1B2PHWe3uNyZxHNSGs9UdZ
Nc1rpPy7mLSxsI71J/WsilGtGqmTXzy7oALF2zOkqz7bUW/ZsDQPgruUX0QBn4A4
OQzi7Kr3Mf5uznfm0cC2kGVA2Agi70eNirWg+c2Dt0zCi1gAbWOWeOvEdDTuM5oy
7KsHPOh44wwl3Gl8SxIIF57wnvORDw5h8gvIeMmcR5ezD2Om0AR+J69ppY+zUyw0
ibpcFQeOS2uFhJEiEf61qwOFlCtKPCv+sLe1IBpAcSHFVHvwbW+oCCRpCLJmVzOp
RzIu5sBPtHdClP9WaUEDLlAeVDIR3sL9khGK+d3A5s5c4vEv0F7KxtloHVjKjP8k
P88yxYnQowZC66yePX4EykhZvvDe0benrfLvRoE+AZJcNeENeuy/AIcxbYdHzNKO
TcqHI3l4a6P7Qt1Zb1tXp8T4I0R65ct4xm15a2WsS0CBwhK/1FMZf4AY+WJrZxUy
61tIZYm2OH+3gRB2MWqnM/Ny8ONaThqMMuiRGv04X8/lJLW+meB38tpNWBLEdlr+
8YkxCMwcVHIwK5s9qwHY+uWI0Q0E2jxK4qh5Yhbp1qjYOFWjobYOmts9xIb3VhMP
03VBYBH8HWPdVHDMsJE+YPkSu2cRhzgnJklYqq/GmQ+nWE67GrvvUZycRPeTARnN
EFo0Qf2buz7WrkGUFXdZHi/qeY3gB/1dnRRpo6Qf4xS/qYCi4cKaNZ9k/eyxrjT/
KxgfPNulSNDQ75ZffJJq5iDHG0fU744w/tO2q7DpZZCqHtuf8XnvVdO4SDUKFKWO
fTI4tS5I0YHePEVhgjyOsvwZi5aXVLeC9wdI4/GfO7k+d5KRizk6SBIE+YrzhphE
slnMns0eXb7Lm1jMQwAn0KqAI859MH7fSntjlPnHzylWHfLbAJbS10D9hb0HUtDC
eUpIvW0IZq2m02W+C1ZJlcDJdD6mSHGzOdsVv4bQLbvsIRs4ddwANXSke4zvSo/S
xsCX+TohUiEihAeNJN/sj64psjLKlJxhBCHOn5Mk6kQ0xPE1CQ/QX26inOK3llLf
04Pz4KCLPRlLkGQoPkP3RXOGJ2YnWy1LHhJssCfaKeFVg0THLA1dVsKk6uhLstOf
lqS9KDK9o1AOFhAR9XWfUxhExlBIqBXFdkxfpknU/a6oDt/03BSHk85KyStFnpUS
7dlzk7TFD+C0jHHPtJ7J0PKUxQWkDSZkcu7TBjfVrwhTzdaYiVwp+olDfNKPNvDS
th8toBSsr9RGWmGVcMke+A2xs8Si9y0U/rtpzB+B7VrIWNkWvrUUmy4f/z15pEtN
Aqzxavb5SQ/64IErZI50dCFbr1FPAqpGLGL7MFpOLrtmNWn0L5Y7jL/0Rb84QoTS
slNQH8MLsXxKWbBJU2wU3p7mJFgz6tJOSGthUJ1W0zbe+00Yorfjlm7TBfiBs2HX
ZAbDrFKzlqtMi3Wj3h5tkF8EbsnvJ0le+Cnq+HVZTCdsAYdKkfvr5r2tM4Wer2Aj
36Ee0lo1qVfWaerfXkk4eeAa2Wk2DMKX2wfLKu2s9I/ACKVlTa/n+XjuQ0AlfCrK
5AFJxxIkRpHxsyxZymRtfOisJiHl//bBh3hIlmO8ZoG5eQW4aGNG/aQLHynpiuAp
idQEKPFpKrVtdf+/H2QIIFBHN/+EaqAqbGBILId9qwSK+U/dWQ/Q8GnxxtaqZl3g
rF71rYJsbdxHMS6QbAQbBO6aGsVvvItay3qtBRXHLpxNj2OVMDuA562hW0yZjRhk
ziAaqhwLqQZzKFmGsmV+/R+Hzd9BYi3q7t92mUaeeJ3K/d75Kf60zD+MMzHJZdXg
yviexIDPWdoyTUbb5QzCh26mhydeFf1Zx/5mHZzoMEV1uo31eO+zy9+FkyDNQuEJ
/5+1rXszjNKuQqBsux6A3r1PKS1pEsSlsGeauv7uWuJIodI4dBu11EsxL9VRXxxY
q6IjW6qUW/ssHgjfKvo5AivCLwatOuF9X75+wZdBJ0WHnUxA6efL6jlxFfvYwHZb
NAfUB5b/jiOao4Mms0RK78+x5pmy8DElPgictWGz1xLSW1iriQ1KixX31Dozyps/
SBxU4h6++I1JMf2qzXOh5jXOwoy3s/50MlwJcaOYU2lwp51/5eWx0O/nBWINbYHV
kqXvAsTrNNY/0MjROM289q/UDxaJU2nIGyxjk4gpbHBAdzeEiF4j3Y3OIqzwtjx0
FEC7I9MjGDBi3/o+z8+F9JzI7+c6E97Sc2tbb6AtsuAV86HXW7t9y86aCmhWwq4K
4rla4Q9Pc6XGzKzO3kds5/8ux2M9X2G/RgUQoC43oTHRBs5gH1IYjmwgDKrxParu
9W1OqREDVX7YFFyO8kxbax0K9/05GEiRNDRbB8ZB80UeX7fGVemQBRJdcasZy0eK
DBaIEr8fbE3cc5MeAhg5szxI0uzjjI11gk++Bfhqzhn9ltnYLJvVw6pMTxUPGmRv
9dfc+X6fnY4TZE4OB3Zq/IYW/Lt+k8BItcaxw1SZnSAn/ZpofqArvf+WCKqYTdI8
/0LqiABH3kt9fvcZtGa4Dz0mYqM5emmCg7dA+3wwkk42U8LdLgSfayk5Lfd2Llri
xx9/Q/a1dMrhGRBB7tdUf646yKmU9UnWGc+XTvNm+ar+KkeXjhf2zBy2tgV1+AG7
s0fm9Lh2dbWWXwq5Lesumj6Np1qJV+o+Tc+fSfNCctbGL/3+gjCAs2HCHIQs9OU1
4VStHioSXOLXO4JL5H5sqpN/tnZWuhjwe1FdHBRlaaj+9t+9KKn3oDnuC3RWs9VX
uXVyR0Pj/7lRivjaL1T2N1O+Fsvmx+Ogoey0xn7n0nYi8yiJP/2B+WXDbnIE6SwG
5kiUqoTd5gYsolu9GTUQhjWY2uH0rPjJ2sr1r0v94vPYeZt8I9tLAxs/fzEyopPk
x/btqsadDVJ9fr0sj8NdbVAKdnU0+5ZIY80fW++eEnpMsahL39peBDgrAYQ5/L1S
wllSHeVurcYjdf7kq1vH+nYBcu/ZVLqO17+7xsW5V+x9ZI0udUtfKZRp5yAb45FC
NHJMKR1UPtqI21bqtqgqkZimHN379ykUJdY/lvlY4op88IdZlYhvC9+HJoeL7Vaj
VKbRYGvTk3/YFW3b9uLeNDwzWSJaBQWnyoTJgxIA/bcjfGOHAC3uw2ENQqNW83g4
Q52vgD+7fXXfGwK3z5CxudiDqgRLAj/u+aClrtx7NgN7GXRkPao9Ta52IN4D5kdf
lGkpV4cXEOrj6VbvTNmfjjG01xpUNNxvoYS9O88GSxEoz+mU39+vkuZGGEPEdGUI
LJo0I6TmBn6ygud2aaaUxAQ2s7yxi+d3pxWI9Lv8H3LHTTdOSYV5SRyreyRc0fYu
nHyXXVL5eisfa68FhNb6JWlTkPwhx0e2fjhguUNdBNH006Fvg50zD7paKuP3azKd
nsrI6f7wUF5QK0+l8WSMtHd6m50GGKaK/MyFFYj1tRBFkaoD+kZ9UHOFyPNTAsuU
Vn3zTsH9Ou+zf8J4qPriAHUDzvcKymfCLV7Tv63E0XtzDJZ6HkhbdcMMdBY7qPxv
Sy/GBnSuCnYPcfX4bQgCohFe7lelhFv3CGC/YGT3ZYbliBhvJMGv+Ub1vB3BvZKl
VfUzReDYfTQwQLhKqySQ11Pxc9VfE986ajsA2E00rJNZfaFnDDib4siDzqVokZE7
0H3fAUlJQwjeglpjFf7vbkT0+2LMe1Kk+FWtAw6fy2/2ymCLal7Gt0rGuy/SOqTK
R4IJo3BVulx/avUe5xPaTTdUwlroxNgkm8dweqlBnrwFEdTiDfD2YnnV8mgobm/+
THNZ2SZKoPvK3KttA50i5G/xn/ByiMf+FLwmeVCnC9YUqSKNjveqC21ZWoLSQZ0c
mmNuPDdOWXfGDgxeqbof8Qfmw4iHGjy8Nbk1Rre6ANkjVbrIEU9uVRfdi7RfHNjX
qkdKQJ583oeqHEwrFqOyBWD09Hd8uDseBrqgq2NgPJLgNcUhjEnrOn4dVvV7dK6r
sbFlDCgF4XlYZCvwxYjuZGt64o/YkTABdXC/xhreigCT3uZewUbyDxsCnKsPRqom
z3ucvsWZJARB4rqLDJJvhuT9tMjwFHTeB9sL1TgIVsaPgIXF8TLYRnq6Hz4HYInY
BMuffH2nqlX3XS5MNl9lazEJqSi8uM3hz9P336evTIqTvQUnQ4jf989FFn/A5RUp
VhAXGgSNXml02fWWntS6iQhxil81HKqYM/oiewkzEsvMLK6CJsCiB9ajpjAn4wVQ
DMZ0YhgEUwVLfUonFmmhKKPH4a9SkDpRIeA7vlS2Y+0Ovb5/CwBPwZoHh9xyDSH9
/aGFi3yN1TQ6aTmOX0XUg7I1ObcwRCx2npGwcem5idQ4drY7twk7MASNrgLQG6KB
m4/usi/piZinRk5xpo7ALSC+f5usyQRkFHtIw5I+ICp6aMuH/ksKl83wpDRoBh4q
cva5R8rq5D0AAaL7OXfX/cnDuR5S7Ew8lL04U5Skxy1ASWmWd2ROpwmSshqmE6bS
bCw1wvQdZjGJyUxi6Sz7eCP7GljNxruDxjhPX3FYoLMn512FQ1iZl+bi/CaNlZ/R
7M3vdSTZx7NtatUY4Jt1jbDQTjiK5Wo7AA2LV14W7Ge5cQEsR3/l3i/AtcE/f+qG
We129Ha7Bcryi8K0ML3AlGDLEyUJZuj7nVzMJTD8N7jL0V221qQxKI+grHlPV8Uu
BAfvAH5dAavxWfksk89tQSVNPYIcSGGeg+flABkjp/eTRQPqeApS7OoKczCqQlMD
0YgMkoIrjDsxBiG9v7yW3A3wr4AvouEqdna/kzrQcu2GhpBhksbTMYBp5npKTp0V
cDlwNqUBjc/43rCvSQhMHVIpg2yMrwQ1KvgJ7ougg0pfZsnszrg+rTpfu5V37CBK
e4w2Mvmmaj+xJsDiBsZwPv65ovLi80NFh6G6/w2Ebw7yVsRJlhao6141lVU/sr8p
6H+/SDwOf1UhucaX7BPJwcfKUro++a4bq+MRChUl4ROZHQn9vBvsMokMdkiD8Znm
3UF7aSeKtwp74d+2oqk2XkShLa4r/7E0yDb0kCEwoP6t95f0oBc53KKDKEO/OmC9
KTjnUgHY45gqs01ZNPyYwHr5aP1rQNtr9Iim80hPJtb8s7p7hqFdLE7/WYGQraeY
72JdNMX8iY5bCgSinVnqA3nNR9QRKMpzRa6MdBShFmJTM1ZZnbqvgznIlMc29k0w
/ubvubbD2f5dGwlK3QnbfQbOF9KOCNM0VXze0RAV3vBN5pk2ntMiDcR3j56gC05O
jGTEKxCvodm7TXhXyIHb0+UcPxmxeVxuFdfIz+ZQUgCaF6DxSBZv1hElTVaEwH3s
nozFw5C+GzBgWCZ/s3DGiUOe2nNkNbOnlMlAYs4Bcl8JdkSiKeSivhVo/A0cZdz4
4gPjIia//N3eFNdSF7y9ezzSr9RACg6Zr2v0xuGLO9cQpAOB2OtB+MOBg/Dehckr
l7GIqxEa+48+bCGF+Zn+9j36/iuoMaeIj59AnLLIRlZfIER0nqMWtEQpx2Ba3dz7
r5gODKSfqbNkJHKMkaz1Gx6ZGZhc6kMluiCnaHuIFFRYtNaQxSuwfhVs6w0nkJ/K
G8y40psYBChRF7Av3zgFRjNser60MtN6qYLCaCT/UL0X36E3M/YJrVZIdZatDUnF
zprQKEWT2i0Fr+8Wstjgn/fQ6lZZ8SH55d9c5cRrFORUq2hGZSZmRYoFQjlm0Iao
LDyBUpHdYhdqxnBBKgCkuqgJn+fi9JxN9UI1siGt5puMCwCuzOs8pDftFV4mGMV5
cvV6iDrJlenkbJdctKTQMa7tyVOC+uZh3clsWKW8H2w8r7ynbwQc/qLtVs83WT86
UbSIHehZM2+2j2I5Te7yDbGbHODMvYlSLYnahvFroysC7CQk2iOt+B6XZpVt5PWI
JOMWI5en7DOV/bwSBsCY5g/+ugA2I7nbR2B2Uzh+04qK+lj//EVrJ2xe49mP12Bx
E9l7L54b6VG3CvAkLHuj1xkkivEMPYQtu8/Crx0K8AQfPM12tQuhv/+Z5wx/xfrc
2QqhnCV/5Pjld6ay+iIgcFzi249Jw4q5B0A0W6dtKAiJZR0qhpAMLFYKy/veOLv9
drmcRLz0Xr0jOruOY6NO0a3IgFlb+mhQ4yINAFxlIBNfMWfMzoaMz3QXRrlErEVa
t/2fcPcSR8Ie4Th5AHv9TddjLeUdjwN/3LssgUPHQ8jqWiWyqjEKDsnBMEihdvY6
WUCsVnP/iJxY2JPEYrJ5fgeBtbqcvEoXQi7/Tc9TzhsULTgIx7poV46ON/ML6gO/
uAg07R/aeIRBtrYtAZo5GNs8Rcx5dRq7GI3npYU4JQ2f1T6G1Q7KjCmpCs+TMwLF
ykq0p+mPg0QiVPy7XMdLRVG3KNnqWObV/WdTz6RJqkeFuGz5B4EeBPnt3mb4HZEb
Mmc97SnX5wrwRdlgpV49eHyuCcZtwO/uCl5kfOQBAT9JZXbdRqM1G4AcUJbCXJqI
tw9QYLRGn8hLV2D1QRnOM5HdMGZJ7uiTt0c6txFaff6vsry+3jeNpKRb1tQdvGzE
4JDoaIhx1szbAenS4stXY1JnwRQWj0W38UBseheHAl0ZiA0cZ1V2jNRatwTz9IOc
jR+xGUWh/vhKdWKRA+wTsxJthgcPkEBEmdgqdTnOz+rmBo928cWrTGF/OupudeEJ
eeSLgNVtiqdb6A5F8niJQ8hVTAam0fsT5SNa79qIQroeUIhDmTMJxNmwQFx0I1lP
/tOEY671lW6Tup0vkE2Eva8ucySEFMcCSj21+6EVas7wDJsbVwtZp9lUkIfW9wIB
PvbDj5/QRkEZ93ZkZ11FmU3JqWv2ITnx7CD48XeGTUuWeoQDCH7pUa0PmNRJr/08
EocRIO/w4Mr9Axmy5YxWB8O2KC2ZgFKisfRpb51OAtr+GDMGXn2ZpoFKs87q7ExK
z7EEmEIn9yY8tHi5HUYEPnwgBexKxY6MJV2v9prx1A8qbZBZ2Hs2HzqQPmaKeN7i
7HmN6d5wUJeZOOxq2xo/7HmZLrJObxVRddPJa7FqAwlPWeOgi+R8URi76F0VaWZ8
wZq5uGsakGLfBZkn5BiDghC+PteWTxLNbMeSRNuXl+MWWtm9Hii2DG372qM/x/Vt
N8SCxa0BSnFgapH0Ppk70uAnqkspSxVRzuC+ERmFoHj9PU5ytQ5aRG+h3cQ3RuuM
r/9AWpjvTE53BliGjEd3ZH4gd+CdZhodIdv8kIrX63pthb6d8evrnzFijfdCBRP5
jWNj6rQEzlm2KTctZq6dgXVfKFt2VlIehVegvm/8gYd/Xn4n5O0mZrLg5GCHar+l
oUxIGg4BBLcVTA+b0eP1/j5WwyuASWwDD6mu0UvUeW+uYuF1EXDZYJvr7z9FH3aY
Kgqiw/oQWN18E9rpvy99xucwIt6lt/qRDh4eyFu0Aqvbho+i7GqRVe1AC0sknPpo
LUVcaz9ucgtH6XAAbCqXG7lOdNAh1sEUFZRyPcxmUXKV1CjogXINGKUA8XcMjLfY
e8EDsXjjPvj2SJDdi6URc2UgovWA0Fuqp7oTv+1shkTa3v3bzG5YHpf4LgOxiZI8
AKfCGcOWcCCQCRwOlPpup+CuRO8oVZiR1cro7QCz4bycfyZAMdFdhdmyuPhJe/WP
el1GgrZ2eqW7xp3tk0QlDMbsSghPAEsAVM5i46+zaEU9Nyybk3FxcBE6xgk+zBJW
DVH5gZ0r4vhkXzSpZh5n/WOPTAY8IxjUKNz98jvf1c1A2GC0hUhfcb4qCMamRp7h
0AMG8f2LOI7iy1qIs+FC8x3FKKM+DonPePF87E6kGcXf4mfLfR4+1zo1tsmO2+Cw
EjPRBHlt/SBkxF4QIwg6PlgahKjQmnQ44//GRL859Z6RYYuQBllxipuOd4lZ/FmD
klqMo7+uD9mTmp2RRaVvDpUlOVOzBlbThI8leKB7SIiHJAcNwDXWY2PRPlNizqsO
QfsETPsymy7w1vlSj4MTEzhoouLrjOWy2QJccwqm+9hjEWEU5FucohrZcdqucWEP
Ehusrd+HnfbLgq3WfUlS5HcKzm0wGmSedmyPQZ3voEU0jpdUDOL6lcoXl93RJMjR
m/6m/NTWRUYwlw0/HB1f9z/05YCmjSOqzLVnK9mAV+zFFFOAvs43S3Y0uW+8CPsg
xBAXx3CtcHJaGdLDfDyQJOEKm37gd2oV6kfuuvz+l3Y1A+Fyb+6XqdbcbxG8HGz+
ARQ+UOseG+O92giE6rkCvGezieegz2dBqA9T8/l33VL+yQowoqMUxIKH9OcpUQUn
e5yGqqgcb2z5JCYQjVHisRZH0rQQ7psSCdXwI0oFl9Pi7BWvIRNIj2aUa94TI5m5
ikjaPMZcpZnC+eTO8p6qijkJilFzp0Wg8blcDsKufg+npEsiGdnvyPbkFmCRFjMO
Nwhk1mLgOmwRoaSpSdutESzdkj3Hu4GP6MPsGCFfYkMiSKmxYBpoHbFcKx3GSK1c
iTV6JKLBd+SHlX9x0JM7o/EAEG+ISZi0PMiaskWEuURr0Y+0XINHfWHqfGYgSdB/
/RLn6EPKoyaHlOUIGokhbcHtRbpEvzMFk4SmbP69SJX1aotVWQh6Wqrcr96XHc3P
tlwTGXMafhUSsj9dA8PWQ5s+PKEInZPZaQvq5iu8Tw0yX8S7s5EAvAljvl8hS1bs
bWLkFSGcmjth8Ke+kpR1o+uOEE4NY4L9qe92m/8l2rqy0qp2ALtfTj1p24x3hsww
N68Go977pnmuyRUVWhz6fk+YdOM/lJ4Wl7Qw6BXZ9iht9MLi/OjX/hBBfXFe2DEF
YLoSlzI2jEblMM04xFgGO6fWY7Kaifz5aUTkx7iT4tASJXjIy5LiQmLhTu5juHfl
qh+N4/t3nBr37s9+DocygOkzCUAbKGxZYQWS7bPsuLmgRzScimVq7hUEu4y25bUX
pX+YdDgGvKfHBzoArzxtOZhuZK8VPjekv+RZrEf3nDPmp4Bv/GwTHS/1OwOBruAI
n3UvrsxLLZL8fWVQG0IheEoXexZBLCC/gLqu5yA8b/RDgXIhbClWunQUYAOkNwm/
EhwpgNBtEbOMdFrjFmEbQCiH8IERe03tcqx6AuSjusW/TT8orkjOMU/+R30tX/nH
xcuUazauPj68okxfd50W39VDv17lJHqY8KbQwzAwRQg5kfoxZqXXoZbWh5QZQ8q3
KDICwHPLp6pfvYHTK/PsGeLQE99eivUwwWc9uls6Ms2wCryZMvogTKU/rHosMy+z
2x2PgUs8vzSRrKdAZpmCzX66N3mna6K+tqrGqypiikPZRndBvs4wX3s2RXGH2amm
koUf6TZUxOna/78EM0C0B3nVUgWeoJVBumMxADHaUuINEu3thjE7FvdhyxGKn3ua
Ved1mciToq3jbny6FB8aq55/P39seCxmnD6oEL3ehIOQtI9touiS7NbJJyVhErVr
aC5WIAsKArqAsoC65SUR9WhzDTF3ephhxdKLbGkisMPKWLyu4LTKIYYKP7+ALAZu
ZR4prQaVvabj78fx2tM/S8+QZatuBGzMT9wA1ag1FfaxhLYMFe/SE6gAqb27hXZX
n1e4UH3uOW+bbdgo2bJCYRXeG9cGYeOX9jfAvF14P6nbvET+p4H8/apeZgRk/fxZ
P+uFFp7cA2nplZdJpllvc6exFL/LbyJglQVEh+QKZZhHlNEljoYtZ1TFbiwWVW9Y
z2R0sK4xZXx573WKGyS9U3Z3+2qkdf51+lvDdvxuf1TqrJXk+DjMGp9rDjWyvpXu
SSx5+v6EGDknbBdnzz5HZ8IHpNjT7dsby4KZ/By/Pf71FCSgtmaNAYbzdSwYnF2T
Sxe1Gpc43N0BZ86XYcJi/CO8sBxHOFl2vpJYWIcqdunqOBwpl+KcvsIXYGcsOsB8
jFAVU7+pkDMVqsypmwwDYzCrP77meaTy3Y5lKMlvEiL+wx0Dd3ZHRUBch/60wyWN
IyzAZoADRyIDYmrgC2dPTt1yPT/tiQxJ9uxE11Q6zUwFd0G/T/JrpdyOZF9MpTR8
zWriQexmFigXDpZglrQuYp4dQNB6Stuj6FHfboqrURhNnR5VQIDv0k4qVL6XDrLY
7008J40gx/wfWu5FG6O8O8gn3DPAitS94hN0LLOtOsPshFR3Y1uiz9K04txqSW02
0qXIo/tivDFdl36brycTS6kLLSrQNYryycmx5+yK8kSvjnbcaa29YXyXllZrZk2s
syUMbvM4c9lCvM/2OdBf3TJrRM27XcnqI42wxFHmV9KrcjKk1m7scuXxwAsk9JMf
cWsTQdA3u29r1T949ZFBOkQjT1wqdeZG+ffvY+WTJEiaYn/HRQjOCmmVUhdxHBW/
fEKt/jaz5JbQznimH798GxFSMGll1uepLyZ/tbvu6T24j0l1pNvGePKFg4+/e1Mq
kjKTC9OFmXHZoxr0fTLvUbP48pZZeZm1OiXygi6a669xK7q/nQYhCJb3KS3Zd4y7
CL2KFcgiUgvKUAUg8pRFcpkMpicuUZii7oWq1MJjQDDpYbF32Azk/0XMR93rxmWG
IojuoHODUX6ENW+Ts1PuihKGrZhy5F6K387K4X4rCeyTVRPfNu1tgpGppzeLW8y/
R2ijtchlata/K4aeA991X/JE/LComTu/J5Go7/CR0sfz5vwpcQ4nCjPL+wpT/Tlh
cpG3okXuNR0eiSbunZDLc1oSVIlLFPGUZRjZB77sqsLTH8ri4J+dwH612ZxV17bl
4NJqBilFj2oz3+YQ9euKjzgxAr93605qFzst8BIRyz9D523+YW4Qzo3rzFttufpB
87H7AZRotQaQMVB9Miwm94nEwhAPIMWKQC6XKyBEOgy6ifr1z7lfl9mbGmpbHdjJ
VJuORL/FA6u7mfDIaYfedr8FbyOtGJQOAs6Cerxt5F5E65wDoQxH6lygvBRfQSZQ
y3/ZNesVIF275c62kgETEiyB4gd/I/sAaqF/lEthxFZaM6wR6J2S84fy6/rcNN9/
DS/2MMZm4Mtyb0gUpKL2DEHHwsE0t/2lMpre2f/gK11H3QSBbVMQ6nU6j3nfFyBq
nrvhMRXgINghrinDj9V9mXHmuLUNOH6L/+TERPThYcrja3gtZsUHiweh0MK+un75
lTfdhJaDOZjmKkPEmXiMvqlKzIYAjPMeD+ZYVUsyYx/fpanIHzIocMKs5ISpsz+O
SRuU5pI9hAf6oXdike7o6L7K6Gfb+HTCnC825GzJBh7sftL4se+UtJ5+BWSM+/Ix
PCeYUSpqffsf0dPVGdzgbepqCBO9hBIEGjyo+F7JEDuXcWD6zzRz0jziwyuPze3b
OEULAPRtGabvskeMlA6PtjBBxheSuTpSrmnLVTk4zCo/too2miHzz3GVRLBXlCkT
s13TWvb6NtJQNqCEvYvNtBp7GbLfk0JZL7VEuhsSVMWjXXO8I6Jr5zUVitKI8WZy
0VXq2VMB+fE56YHVwyr+DzTBp0pXgMFqX/TyL3Eimw3H295MnPx/m0oTfXykPdlv
8bbR6GM+w4NXE/dt+a2Zuy/eqtjEM5JCUqk9SNdlUTlW+NDxYNNXpdnNityQbiJw
s0y48+zFnB1Hv8s8iDu2T0pESJGiL4Qn7uTT4nQx8n0fXaz7uACHY0gnG0dxWTj7
etvVWU9ZGadxPLeNPtKbq+U2fb/w4LUiBFk7F2MEiMHxAXyPiVII02/PJ01uVR6/
gL2h7GeJuJznivj2sJ7OgvF5L7gl13xbrp6Dysitgq4xx1jQs6KOc8G7zVj9SsX0
RJdrJ9ujgpRpvnCNxh2gKm2p955mdri87sZdB6691U2LXLj4lD+SmmHhkqKwsEJ0
ZYaa+V9XT5+Un0m4dVSdBkg7mtB9AMKgZoot528KFTCocBWvT6ytejTz3xckSyDp
hWnFPNwiusKuUpGyxlF/YQ6vhbvAEtgHvvpqc3n/cnYitAKzCZw74TUlU4PAAPIb
1YGqucLcXq8l9LbPMoU2lzzuKoSS3nb4GIc9Y/3wNeihf8NSIrUYpJXPPQUGx+lD
KilmCiRK34o+dIZZ2aeE6far0I1SCh5f6MoPKgj3aJLTcLRLOKwbWQnbB4hixPQb
U1OFCDrVyAN21GcCw/De12t/hUWJF0xTkv2IHsPuoiN4wPiXkYkPISThXi2kusHw
rVby3mbHEdPd9V/dMOAUZAMqFV7l8NW/tYFMpYke/hMKO9Dbw/8wlyH1PYMJsf3/
74B7FOokRfxnTD/yC4zXpOsd1yHEmsha1SbYItu5skPh8fYxXyNS4bDxoqjg+i4h
Iay4OkUw6v5exsemgbJXOZINDp+m9lwigzGuzq4mA9so18iLWI0MHDQvbF8PVmmC
hqjzQ619U4s0BVDpClOBhhGz8CpIoRCBuoXsHKOu2426ANHc/IUDyzRlyuyqLmHc
1vtNfHZC42ynXW5hNGaWHkTi0bEN9Z+JlxwG5IsHFfvCTu1dSM/TTC6K4iXqFW4n
f47MrFA+HmIZEa79IrnwThO+KFbg63hdMNYxvoNA36SiLgZOWorSlrjZlN5JubzR
oisPBrkl+q199wi0k0puZo7m0DxBQgmpC2BUSH4hyDSs7GU6ZBq2BGRR8ff9dnzc
NWy/abPO4CxOLvRqi57TKtKBHPSQOuKXrSh2fgRposTrpngTeh7vBymctw16AO2V
IlLt+BMiRazWk9oARFsbTEM1YNVuOIhWtbCgHtt4LPmfKrv87iZ/Ayfsrt7p7FMU
WOVVq+/paRQtwRnFhcarBk6zsTfFPigiXK6OFBvGrQfSPz37K4AMTU/t3dM6Nntb
MB9jaqGhjRfeRhnZSlad9OwEXMrOD54Cgs9rEVsInAxYfL8HmTWX2TEqFBK1HPt+
ZWlXUmKEncnipmTVqr9EAgE1Vad5QZQNIile6WnwtHqDIm+RVTlXbjimdivUZxX/
ohj3aHcMa2eeOyq7+EVWSxEUGJ7V5HmJp45vP00U3az43mbWZseUiHRtDaUk1ELU
XWLyOjBYiKgvqnxHjivNSCDBYyW5JzmIZXWAVjdsRPRgnGZjFVmXnrlKACBNpuzd
/0CXJCp+M6bsfETCOu6qViEEGRmnBdSwUS8ocBlvenz4BR0JoFJqnXuGUSccxFe6
GCz4V0DURg77/iHpwoK14tZZorUm4ybb13Q4SOyiAwbsipgyjih9tKEd/pT59QVw
mSP3n/p5VJ/99N4b3Wh0ZY6tNnCs2Dq7Cjrh0VMTstsMZxWogqL5ZdLh5oPF+fzO
qczoH6xP92gJBbp05Ak0WJTlaQVvX/727U/rAj5DxBl/jakoLQ1azqkIMx1ADSui
Zj9tMbU/RE33/qRWEfxvFA05Qqna0s4NniZFb4zfr6rJD6MncdhNjZCdHUNkFFGP
8e8vw+CDcjmsXY+T00huBfgtYLAgk8OK1g274Mrb4Z4z5Xz1o/EJ1lZjkzQ/8yC/
+byaHocYALaJZz2TfA9BQCMyh1xdIvHkif7MO9dpDuOR1y+narL+1ZQHJuST9wHn
/O58MX56EVW46UapasPv7BgjhZmv0thOoO7uRtvTm6RmxPOqPYfG8Jdr06VndROb
jbvz0iow7z0ejjihO/d0vKjkijjiPkUOSQwcStKHPrfTNS29ej+jecRgxXuim69l
d7uqGdazI101k2P6mwDVx48IRAbz5Jw9odLBbC8G5tMkHHJOKMGzq9vA6J4+rBJR
9bGmcMK3UPbAMPPQ2iwF9pucVFoxTk8D60gdUdZ8Rd1rvZrWYEF9xJmD5pRLKEUc
fupoQ7HB/Ny+5xN9TrJof+7f69lP8saI3UvYQobrJelrugCKLjc6Up66Sc1A28vx
fBKemdHuyu1igeLhYBLiRDRQUEOz0BlRzMGB+0s0YGhcjH7lX2vpNRLcUxtXOuzy
+87iQK48cnLMqaEvLB82orMQVBGT1H6dE9JXThz4r/A8id1WQyBr67U17EG+5NA1
qm3b8TZYxQnuxydyuJNPPw4vug4IT1H26UkBhYuU8bygXb30z5cXqz+Xcr8dw4aK
Q978q0F+Iww5ibiE3vrM0QGDXURixi/0zzyml2k9DZbMIxorZh8ooa3kr95LnPBz
e2vYQ0UhmfXCaVlSeZJ1b3I97yYGFfpzdVpJNfpSPKbP2Iz0Cd8T82oeevdH/0C4
UQ8WrcXXTEWEXDXB+0hyhQ150ZRRQ8ngG4EIaz8cXhm/bXLLW3wDtATu7NXpLn6A
S2O8vBrMsOnZaLiyzzzAWKOOQ4fvMCQwBydNp/TmJgfYDPlR0v5df4P80NFlk7SW
mxpH76AiPzBhkV8lkIjx7GjLo4Nxzs9St0gegAZY3rHKXeslsW6ucZDdg3ymuCW9
v5QsurwTCRSkB+3IsJ+boIIUL7GtOejs+GJGjpOtKAKJ2rmHTz/M6NCPQ8r3bw/n
d4ZCvda3GJcO8WyD3+8VQRZkuJxRh95YgNJXwDMpsau1WMp8QaC1utM5slsJIdp9
CfQegTuOGhlFwUl0zhZATV/Ta+qyo+53qXMwKui9P2syQrw/Hp9pM8BZezmTfDq4
JY6wTz95gk0QjmGiX07aS5qSaZAC3AqBpw9Qttxcweo0wMcg9yJMqacGzZMWg8KE
sg1oTDCqIqwLFzeQf+gTpxVDIyOa9Z5dBf0Q+dxwRAE2lVZN+v6zkPNYb2ve8Mgo
Cvx9YuzRA+Obg+9vQ+mFDX85sidhuNSAK76QAPkUCMX8fRonOtxJeVXkexuvlC9b
XNiVi/WFMa0Z7pT56OtViHIajgHca9ZZ/jW9u0qxQ8It2SbYxI3ee7IpT132RvOJ
fZL+Eq7vE1a75gP/uYt93mQd/V80qGd9ar2k52B7ZKpWHirE9PuHc8o7CMTsbCdB
09hpQgubdYIfOFOt8V7E6kGBA/qTL8IRulqjUOrOrR6lCTYXRsHibFL3vc2xASDd
m86UirMzuL6YO2TyfjaUTEXdutGBA8Mj5zptUONvmUImEFGP6Jwm2G0UFqgFegaf
I5grt4Q8YVh0WMFbdvg5Dn64Gv5FJOlMp35gxxBth0+wC0PxB9bAY1JDaO0iOLzf
+cfPpOT4alWWDTonh61QJg5zkw/ZsJZQrC6vhUK92SAAN8bAPjPIRAV77LActR8W
IFTBkEkX8N7j3+W0x7Mwvr7V7axYoQ+kO68IQ9VzP95wP0nyn87cUzvLffP2dyc0
dPwUGoP6Z6ttKLOI3i0k2bqNXc/Qiw67248wFWbZQixZdYHTiksNwtbmWc/VZvJU
PEkrHZChk/DGaUm+im4HzjX3YDhkPqE6pLekw+TAmAAEkTd1qz0oDLsmae3qQl48
zdDO8DUh68m1Hzn00VzY9jC3wghCTJQkCrzjiHQfA+jxcxlCFlH2JIC9NFkyWsV8
XZ9vhHuFaUcqfM6S86oranINFzQXwGnpOWrn68GOh09a85AMbP1YUyARymtLoo9e
m9SQ1+KdFeAjgb8n7H9IzSlyYeNtjoGzvyvvUM+icWWM2qNinkSDFxle646U3c2Q
2GN+4mfbbo1uDSZDYz8K1wnX5fT/glFi+A6ugAIVeCR792xreOM+cRQyKlgcCO9V
r97SePz6V8ss2VH41wFGPonBCm/QNP/zYwxlJfeqrpzbsX5S+Gj+nY65ygu6g4D4
mgTEHzBUvZH4JBcZW6X9HCDDO81x3jJIfv9OxigfLJ/LEzkdATP96jisdrac85Lp
YbiJhd6YOlf5wwGis8AWuEVfefoiTGHHNuzVY4Wjm2cne5sWoKboBENdl71ASneE
52GzqItJWmOasd7kstQY4EnXB05bdSmhUZYUgeFU/yj5kJmBUJljci/bpu3iey8S
TKInJrh4cKfCuW9R27SGYFXz3eO2C+lapUKEpPkcbhscu2Caj6HS9SRxvPkFx7b4
kCyd8lO+s5aPid52iOSksV8g21cO8X4GZcG4yiqF1xfN7WoLe1VxsA7LwolVDCZm
nGryjZTI2LcwVy0E9Jj9RsOL1UGaY6c58YcerrtAvcr0mhWGtL1/SM2lTaHy601N
hQk4P2eprACEk3GkLmegfLIjmEBvUmTg1sxnQF62cR2qKCoO9YDwKQBvkh5upwYy
g5e55kvbxAMoxRwNDnOwdfJtu0yHGT1KUXHfGSkhrdAwTOscF7LgthLp3RD9tA8/
SHaeIdH58efKp875I3CEwKnhfJktCw18z3vwipCV1f7/8n9R3wL326gYNnx9ZaUg
kvyBgTy/ubTMhiZtsk44OhMqRs1ofqvZtf9LCMhx5dlkDv2Z8Kk0Vlrz+mcPIR5f
GkSV2J0R8DAPtzyXVcBIv5XWiXaLvC/inTpMXOxQi2KqeUGbDG6ao0yDcew9PIKT
+xhgamZvOLaUdSNiWAjFQsvrdgpVTnGfRhijhk/m0UvspL7U7GsPKjexzEAeaZ0e
YMGhEF5HhkUocY8V3IkZ99M0oSiRARAo2X/JkKi2u+b2ccSmHvcEd8qzr08akhfW
McHTe92LllDisQyiPwCFb/9JlY54JYonX43OIoLrgC0zgBvPsFwRKlvfVIKSsDW9
fE9LE2gyGfTvMbViaJHhKOYlh8mI71M8nnbe14AnLG70F31031PJmHuSmZcyawx3
wtaNrSgC6+ve8CI2isYaNTisDmYCpRLze1xjzHlP7OwI/vCWkZZhndhLIF3lDWMG
0f5Tqn+hFUfyq0hYgTVr/yu0HpFQ2+qk2qPKZ172gdGSQ/+vMmv7nwlX/Kw7vpH0
0Xga8VL2SqSGiPquyCliAkO9GJ5+weuhwyd1qe4bfSZB9mDb61pzGCPs1OTPi1Wu
T/a5tjDFLaqLSkReK+6F+c/hjvQvYt5DMD57ghoBqd023rGR0mtzUAAAItlft3Qa
+gyhx0CeQyxkb8Kjk6vSbQyEMEjWacInm2A+fCshEiHZDx6BhmpCdgTp6bnJZQFx
04pQjSFQ5Ygk0mB1jMvZvDWGlF08zewEMiKMXEE9RzCyEdzriHDFoBhVYvTRpqeJ
pSTyLhBrGGvyDxw0u62+xDjMycgRNV0xjTty+fmBBObD+6cRE++ddgoJ0iZnIexB
gH9O2pIIdydZLp3Shb5cAP93/N9bVAWiL/5wfupMWBx0o3tFXq5OR3DBjrXKJheT
55amfBVdOmjw7O1qKwhhib8G6/Bx5zZG4BFDrP14NrclJ0xDzmnMReIHoNY9sZDl
T9Lb63mNg520jRMaS8p9vgRTwuZwpu0zvBEntlvGpdqI85Jng/9I9wCb7rFiFLMx
7k81fkv9bHvXB7PZjOYCJCPAuZfFfUMgA94HH/PEYkY8MEDQdnTDcpNBSayg/oYh
rQHadVpBfjz8HMGOcTiiWyFArs+bjyVFxNJZPRxFWYoesVyh8eWcH8tnoWrcjS8d
Ucb+lmq+WOpOMJu548JDdk681xtB0Ma4fo6dbdBK5uF2vZ7YgzmxN8imfHFiwWWc
ssZERv2JZrQtG3YWeNGPU/Lus7WgN/o5/LG/Ql5cl9oNsPz7M4nWqPBQFd4TJ9+m
8QGiv08n/j2lr14d8hfqEIC62+IauN/Ax0tPTNELwin3MouPXhs3zkk6sFf/4iud
Cz/5bEEsmNwJqehvXpBk1JOYnSm68s6euYeYnzBwUlIzs6QkUIA/mbaiYK7fVSrB
8xUc2/cQCuZA+xbxNa2Jv9nygLvFFeG9C78Bp+ywJWjUxqrmurBgRa/Oe+8d9h8z
wt1t/wwR0j9jSBlcSxGBbzSvicKM8vkU6jJw3vntJPkFJbQ7hrsX2bLfi/meCrbc
NWj9kU9HqqS1+s8k1oaLL9HqLYOxcXVzwakx/Dh9/9p4Wu9EMeC4WRty0MlECqF9
xFzShLkf8J3ibV2rRq7NS1P9+hoYAHkujqMzN6n8+yZt8xAeT4Tw6TvAErBpxxXQ
aLp2P2VH3dOn63PvFZ8OfMtIT3z/6H5uzPEAuZYH/yw11poagzas6rMflZx6yjJn
Xwol9368OuQmDo7iI2NUxhLBF0sGXbLQXx40MSfmOilJlgB/DplH0M7LTO5qDafa
PFcPb+dty23w+FRW19vLBZ+bhxxx/4Yqt7ntmeCi0XwIvhadZz8xAY2ASoJxmwjg
a/8sgcYNoDplc4Y7MoWaiFzE5dup7zgj0fqNHhnOl151wnFb32rOwBppTc7bnPZZ
g6QPh/aGkxwnXSepkt6NTbvFNv2XC/R2k0t7unVoCibGuc6aXnx8uyK1DBUWNQmw
Uzy8Ap6yO7B+ZIWf+t/Xx4NT7YT/IWE37mbAEx+Q6UfHHEYohPMG16U2DvoTS1BH
AXg6yHFf/zIdfCW1yoQqpk3ACE+Hs0oSUpn5eQxBa8si5kRnUL02YpdCTXKaShif
CRD1ZcWp1mAPYKcDwDMOthOFXP2FsUno52Wg6CEQ8qa1bQaT53Dtxkeu2iGoNr1C
Tl1d5caqsTutnZuLAVy7NnFLZbFV2C+ShW1XqAeXMkjXdQ9H+KIAOlAh2R/e3d4l
kCPCoiL/k8tyUOJY2+Wxn9nzKaNMoGxVAnRU67ODyEIRxiDSaVHFe+OMPAhmi4na
Zf+qLnkiOsEjQExI/eiWIsUjEIus2pZZnc4Z5L8LHo4DrQJYZdQr5zJkx0YMXvm4
szHbN45CVaNpI7h4RbITmat42ElF6/de4MfWyAVtxyFGDqEh/zYSpcVOiybBtM73
uGlaF8GcGw9Bcsbg8R8PecAx/Y0XDGLT59jnB/l2G+cNzkc1hfBFFXuvSsjN7rwx
hVGMBGWprTsctqO5gYV0B5VyNHSxFq9UwELzqux2SliMWiDdLVbKQgxe6rbhNYNK
K1jPAbTtYIbi/dA8nA1pcYzhqzy66aGGQjBh7YKrEXJnDw3ULh53VxSxWx/a3AbR
4w35JDxfrObGz/QQIjZBTT3R7uDgrJDLUSCQSUuHrFOpVwIt62xu0YUtUxI08Y5M
urxKg9DhHVycVhjVEyHUHxPbfLpFaj99KTcgSJwYh6ProE3XIPZ3vl2cEZNYthrs
Yfzp7lPt/FviImQrHPeI/uAMpMP/R4skB7vCQnJT6cXT+L+IeE0bJaATaEdZYtZ6
poMQQ47wXESirgjl5O87LWwx+9WhV1c8bPZLITB/KBNI690XfsmeFhPpGThCdoBU
iiYbDUoJs6R+ldfkS3PEQc/tm5MfQ+xPEE11KjROHQSOAo3RZoBkOdlOTBf3z5mt
KmGRH7+XfM5FLiCrmqi5nbriTMYQrbVDhkh7hORRdBs9hklybpqDxccXANblPAYm
Iqd6kqdu3p9d1sPiaSG8m0Lhttvv3RvgicqTn0nc56zOH/PpDPLSPFflnwC5emjD
1Fh/Dc4ZsZuH+CIhSr47OQ4N/GQZpAsidsOBXoYu5xLTjNwPRPauFdRVU61AhLQa
KnliEoYv2XinOTmki9kGgNRSFsMAnEQNEHCqzP7g5+iKdy+t6wBPK1/mXpvxsN6z
4k1u+vdQND/tJNdeyBJkzlDrF01nrlf0AflI+m+cr1FI2arl3QVxFqR8SztThEx5
U7980kgy8XBvaEr6F7UPvEwjBKlWQGIVWyNOBOl0DWr4TN9L00b0UzMftgdQGFKp
vQZDS1OTDfhSrXPmvhHXGQ99IzuBC2qqfIq5vkaT3ATGIbTv1pqYZ0CXZPnJa+7h
lgSK3+aXUon/8z+XWwhD7k2xl8PeGa39pK2yb3/Omxvpr5qH7zDG7QRnyAKaNMMx
BB2PHLEEjheH4+TTWFfL4Cyr9898WOirWrHeiyy9VVMw4h+mxYdxAvDdc9Lwm23d
lNueNluqry13zTT4CPkERjTwfJNA7yCgyCXtkCajATsOBcqrAXNiZqlRnySvT+Of
P5IybQYWFAU2cHZi4qwKgKNx+KBcl4ydiCwx6nVoImYslT3DS5dR2Y7Sv+R7Vmhq
fz1/mmJjkN6uvoO/EegkiOqZYlt5tPpRJbPBCiMaMgtEqrDMbAO7MdeWw74j1t+F
r3BNutc3p6r+tT0kwzFVS8l/UVnIgnCJ5ls+xK/t1ZrKlq+BsSAGVEGB4C1OMMMK
/jmjCV3ocEQrIjIldEyzeb0kmzhZstr8pX61Q7o64l9XnAL2uaLISzi7DrZyfrwt
aLcnepq1T/apv6xs4Lpzo/M/G39du1VN2Gu8ZkL77hcKgpX+dyHyM9WIAuZGIqo9
WqzjM7PnWS/kxs3PlYdUrPjdFH7zoSapqI1HHP0Z07DMYJLwnkgjT8jTbbJVMuDR
lFpMPb6GvP4TZVtZaDeUvqqwngB53dnBx1tvPLOmEu4S7vtYGb05XZDki8g/Ni6Y

--pragma protect end_data_block
--pragma protect digest_block
E5R8AcnvnmmL/Gh2TYDCKAqc8CU=
--pragma protect end_digest_block
--pragma protect end_protected
