-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
cDzDRSvJqcOvx0/u91VUDGc3+Nj+5WUBcBCtRoGP6wP3ryivqWFTpB+6zsZ0KQIq
DSjGf+xP9Y2Ogf708BYsYvESfpgHDEHptLP1Ark3iNkAlFLL/SEn+sD3Cq2/PCZq
BVRKvu3c4F5607gMntUv3xBpAlDKrxbE1BK8ktdQdEc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6448)
`protect data_block
yudI68T0G98Uo2dYWNe8OilZ6eldTYghLNFH1kNCKnCOMw2SRUtYf7ZNHMIymAu8
nr9iipNyu36V/y4l/VmRFgGN1C4iMTxGqMpEEop5C6MU/slz9Fos6GAuIjCe0eZ1
5uI18gwAvJG+YzEgnrkc4bkJN60zzmk7TfR/XiieBBsJ5QZh5ulWdHN5tRRbc4zK
/9PeaOI3WkU5gsBd2N3kKrU787T6gh7yPKsyrzGZuO8nlK8UWmf0TjzJcO47dcVz
QleYl+0zzlteEugzG6GaMRtP2LvFjTXZsy4QdnzXdb6wJ/ot4eHpj2FVEyiehJIv
/pue/RDsSUbClaSo6xIXuvSNqBlF4OvArdfikOoZqpw60h1J127mfhsX3eQVKpjn
0fWQwpE8x/+kLYjxH/8Sh2/r3QUXjTDay7NDuA7tndl5U31bE41duWT7Z/0hD3Zm
JpZVKu7jDq3dZsBQLJUanOIJIoLdyOJxIJ3dGoXxx3N+bqn0bJADaYzq8rS7Ws+S
/ThWVmXR8gKYEahEJDwDQfMrSPNhIlm4tbthqlVCW1rrlzu321DfH+fdmuDcok7c
ZyYovxJTsbU1s5ozGSudtA1T/LIiEwJ5vLBjHJG7aRFEPjyTVA7qbmDAIk2vNKzF
M/odNHRz2wbcu2bDrKN+TZxU/oJe62OMcIdJNrRyKpb1fW132NzYKZiyzp/ifAqJ
y2VgfEnwgBA7sjWWCj+TMrm/IJUSBy7lk10oE9uYl1ZVwl3/Hlgkw9yzaZMk9Apk
QAprj6QqazUN+edH3VGwPUWmy+f22Rrgc7JdJw2aIfuCdp3/an7tsrlZxQlT6BNO
z1C1+CMMYf8i7VXCvcARLytExMeBDCOTTJRXzUi15TTN++lmxnVxKaloA+SK0aLx
lxANf9ARRqxNJnYAhqIJ6WhijyLDywl1Jks6e4gdY+NjSnwf5f2T5EhNfJghoYPk
5uYrIZ7Fss0JTh2000GsrSuZz+qC8hCcvEf8PYcGxfXW4nbqhXTpqUVt1xgvaRE1
Z7v5Gxj1tgtNPPf9enQU38WdaW1mWNWGzgF0EEYl50eLBlFlt92xJ402UVGPwjr1
ErwVLXnwVpgotAGcmfaKTyiJO8lpq3Daz0PfVBghbese/ABSusqfmjWdWFoNPM0d
ks4vecj2aoAwoYBKCCJcR7m3ECNuPX9gyVanMPTH2usvFybtdL5DXkZ09vd3l60+
fzRBVm0+6D/FPEgg8Ot6WsbKB4HbYIqyaZPcQYGpXgzslUJl+eBE3LrbdKSxULUD
arvIsRcSKkFTralxwJtcL4jaIbWXY5myYD0n+hmFqQuAt2CCxvkH+Ge30jIrmEtF
igW6p3qIgW+jHoB9mTlv3LD3SCrtsxdYUIlXYCCXxCFc6Xgi8pEH6xDnJHRGnS8W
n1IWdQY8Lqe7EvhKSdF0oBHobR75UA+1E2TNA5LJBlxiFL2qgmfDnk+RwJSP8Oos
uXGKjm7qhPuEBxygMJMitcyHfbaxLl+UYfSsvfZ52nQw9AtFTKaRo+Fpw6Z3skvm
bFNnL9qp69dd+KobyDTanpS2h2cGGMEknKlmODJPtV2x5NafCqcqJwkp9tsQATbh
+Yg9IklN88WcQC1ekVUODcWf42DpvjvM2seCKwvRN/UxU8Owxb/yDhCOftx/ExTS
d4MO3cL7lW2lSqNb8srl3vO3uzIeCm2ZuIG0ZxloU+ksRAdycuSxyzYBlLYUsgrt
tgpkMhGgy/SeioKvZkgYCmyLqUnq6muuVJpvkPMhm9Ps3A0N6g2DFYkapN8/O3Bg
r7ncRcOJ745wup340aZzVXWdrsD/uAV6BF2Fl/kYcOmMG/9N8olcvDgbFLMbdHa5
waoiuuiIvGHJf2DT40OyJTN4G77+pgYbplFLA1Hw4X1HQTpaiBrFQvVA3QxoEnQ8
0BjX+U+wjXOBRXcwcdNC4ehcENh0xxEZMzfB+bITFaz6VU8gDugY5kwcRPspfElZ
BwqWeQtpOqgqtmvOs9R65VIhZ8teGizmkQg33wR+3D3ZxDVCzNey7hYhxDMYOF2i
RsbybA4Wo8KsIMTHDKsDRW5ndUfQFT8A92QCyFPBchHqCuvsvlocwB4Rr9yU22Ke
dPJqVipSyVlUZXITq2OOQGlR574VrQYCMhw/oBXSjvD0Y529FW0dALHTAX5JIowH
mVi+pQqoeVHVTteEy2mzesNyB/0prooHPF1CithF1lyYAR+2Fh6H+ZOjedShaIsM
uPhiHdzySZSLl8JyMIf9B0N02ifXIryjSFKO3+fbKg7xF9lZT/6DM7d3HLd8q+Pn
w5JTV+6S1UbIInqNOjUNLgJsz+eSamZN8tqiw48LKJBizYroAJXHywtHC3XjMqwR
04pm+O+Ol1/Logt2vhgV7M2RNFRrfLpNDuuYpX0SVakAH6mQSGgutdautdVXUanz
AAaQGBLM+aRY6EnTVWaMMkjpsPotPjstuMcBuD8C2GdxayBbgRiius350N7K0W3b
LcMThgxoEVAUA+l9r2T0AY31eMcO/AyQM+/JFP0v7ejDKGN4cNv6BHSU2qQ0lQ0N
fdmgmE33HA6jInZepsy5xApc4HxIz0UuyhC9bdVYUrL49m/KIf/G2ZyihoI6qTbv
ETqXc9PdFHDADKJ/YmrHxX8SftAy60BI+j0i7lT35Ytm9cj2FznVUOLrueJc6XoJ
VAc9KV1z6SiJ0hRODt4jXH7YKBQuUnPCYspmxR4PCVdmDKhi9olABhiaheSyZCC+
xJE6GbXGBz2CJhf2VyOltCFNsEcBFNkFNP/RYsdifBh5Rjc4V8fhYrS/pFgdPftf
wIvaiupP7JBVPe9gBX4lfcS/JcKLeqW/nzkBZZZdseGTVUKCRCaPC3buKwGGx9ks
tFWKxAfu7sQsDPdqRnKYzW2FaGGUtXpMEZ68eGJh7vv87sPknnDb77WqKqIikvMi
hVEGfIhUOgjjRjmFX40hgkj0/jOoGyRLPz1jCobB8d3c50eGzD7anzhEg4LnWfKn
3Pe498EUPMsjYGhc1PiFRot7gupbo45nFb7eNv3og5GQoztmVhxOWICDUM9P01Pq
35LanI5TwgGY0uWxjhzPaqBaT3KctzI46Y/vg8AosVy6d9nobkwPIlJ9ohmCoXCS
I7Bydaufo/qcEnjyn9f4ZT0qrwbc1gWzsguUw5vxQcF9K7cX+py+42rRZgmF5+1B
KwkngZ05jIT+puP6/tKrl2bw7sDMFUkFAhBlYi13xwHMpnf55IR7BB7g8lSufGVR
T+BOWzai+dMPIxK6gbdn/k3a0A7JYW/rUXxS6pwjA48s4YhgiGUUPzrd4NQeOPhU
dVo5tIKO47fy9DQrJTkJimRt2dnDnok9dQB7hND+DoADsKUiafhL+atJh13jSeiW
LXkNRx+MAzy4SPviC4WJbvgQhw/n0kX8MFDlgkE2cMsQQJTmmA8mZNDFxe92zqDa
jff9UsvIlQaQyG+M/JQsi5jM40GJ4HDr1Z0dOQuT/UkJpDJ7smil1RwRp0Z00Qnf
nWy3qq2yrUNDVY2lS8xVWVjLUN4qHkeELdh9iWSfr/X3br9C/0nOmTncpsEszn6x
AgEllobjmMvNy3pWAaGj+LNH604g++V4Dw1qE+r8qwiPaBWMa8AnHS7mv7Q6p0Ij
3EPD5tPMhsQmEcwTiVDdV8q0Xq7mJxpqxVVEXwYOUxx3GV821Qywdal3OAENMDEg
58rEVzfOcL8z9H6TXkc5of1bxWGLphjabgXuRES/ouPV3ub6VfNPgckSt5OxLUGk
wWCZJ1U4dwQdNVxffxx8I1JZ1wIzGaFUSrv4QpDLsX1chSD6UdEWfcxN1lek3bW7
sLNPv4sij/DW1WcHSb/Oea97ZKmGjsySbQgyQ/gIHRnYY5Y+6i+VAjfZ7DZ9p71k
qqRdOK0DhGHWJ8kUPNXaeupMTZUQExJokaOKkLwMSIAYA44P7Cf15mK9gKQXdUjp
XYdJL279yp38UMwla65v+cr7K8Q9bxCnLO/4Yed0HBnnsWBdpHlN1GN6ze92RARx
1oZX6eceITSoM4Mci5uidiyIGpwZuOrpY1/HkdRiLZNkmywL1mtTV13HXJbwyS0H
Fq7D90Ab98ysgIGMoFMSIPwu8Z5Ge1/wj63QzGXByQ+LM5kCqGXjXgrqiDz36qFl
4hfDqROUtZYIjpP1Xr+s5pSj2fDnGiIdK2XOE3W2eGbHu8daWCs96tN7dycuTLL0
yXf/unjTUZNp9fWN0OwLtdT4L7b9VEKvMsZgrDDiXxFYbR0vF0psaUx2B1ofY6fB
5bVr+jkMsWzO4GvZjhDftJji8peR/hkvduq/QFX06OYjkHztH/pkSnGDo/u8mFyE
wtd8wuE0D6jWwfmFT4iu7bkVzD0c7WgENgsUEyiNtTita3Lps9aAWhUqWqFZe6Gi
r9BJpzJCbIueE9pW1aYKdfPO/4hjr4JVtHgPmFTdfieyY05wHEF26UP5kbH6sOBK
hfKDFgyng58TW1/h3HKvRnvYWgCwLl0xvAb97rE7ayitkyMwo7R+yhC14nTAzXYG
XHs9fWsrKaxXNkJES52vR1KfyHKQQXch36LQRUoSvtzqpjcZGLpvUWWo+AFgU3wN
eyHNT94VuSQ7GIRAB8SoFClBv+R+R0eo+YGV8iCDvOK/Mtk+kBPXG5vsQPK5jnJW
9lvuLFpxozvmaOtHG5N2askFZasSTNVPbaC0KonHp8cxxirJ5ceSFMb/Iabpdv7y
TP3WxekrZntEyT59v0Fy6Gl/2GJJoOyn0PmUJBF8g21U0pbOg99rUsd0V0rh67+/
zIla7b1n/AgduoshhXkEeqFD3sn2+UZiQGxoHMoeH3EARlM6UbkBcwwLZ5Cfn10r
q/zBwusMZ0WnPAU64wabMTn2ZKI+IF7FTdUi3sUwui9suEIcbH3sowEbgUBBdccQ
+ng03S42xquvCXKhEIA1dxSibVda6ccR5lhTYhV9Es4FrPtZMI9wpBU/7m7bV9yf
uV728nKxTQYghmH9JHCLvuSy505CQgIDo27kNJfE5mwNx/pJjEu1eOS93GHxkpvX
kG3b1JkkujDHuw4uL6KIXzrCOKg3+p/Vkoq/i0sZS5kOq0yQKiIQQ4CWPqc0fA7y
z3kvj66BN+BlD0I+2ZzGo7qV1/H1R7mjxpJ8hEfGrKl2HCbbym1pVDbwYl2RVlHU
VANYt0HZbybAhRrheIvt68wnvk8NZN3x8+mbkwXuwWK3apyp7Ct+QoumgatAwxgh
BRHOYsD7M1POxSwsl8xjyc/fFGWgPieQkB47PK7vhvd4D17/rbDT7tNFrQuQzE6K
qKDjal8oizuBWj6rCIMjXGqYveXFoNwyEMwAqM8+1S/m9NetdcaH0xgj0CVoD0Rg
DgaFlStUIm3Y3o5vFdDLzuyT2KieAIVFJx6bOjvdsRWjWEPfZdsXwFWu49jfKB/C
LhntUqCnhbXN5YjipS5eey7HMKo9SUFhjqiFZrWuDfQyWmr+aH94vPMoRl1uV7KE
jdNtg/M70uhY02AlqIUM94mML+P0/hjgVLEX7yTSEtcQZIM9Bm6vkyTscOxsxBRO
T8tbJHZZOj8S4tQ3YGafeFNJtXxZzUu8Ro4yriJcd3NjhyW8NFKJIXAE/u30ODmH
e3o8gNUasq/O7fhedbVRCaedr70JoFao2cB/aza4SXYHkyUp5I6f7J57Fqhf+GbV
C+Wh3/T4rimvGR/xELhYu1S9UMDlsvUJj/yDZhVfGbUiDueR3P2k0i/NfJrp1lyh
5mOoFKsXRQUxeedEftyH4VufAV8kjoZ1Zlbzyarz89AvTUkU/lsl+veu2hAAv4NZ
gFXDUg3h0QmusRDeY9692ujlWBxfm6TtlhBRBA31T4KmKfazcvWwPhTkL1dRT9fF
54+mhG7dv2MbcgCZEAEpalU9TQbCTEQt5QWMQgwk5olWN07VBv39HTNnZkeJGwdM
TWGEdFiND97fSwZ3edhZOqBr69lAYedsyvdJNfPlO3ReQrWTwTsLluTK1y8xzrIP
7mU2/tlgNKgkP8h4c2obilSsv8NtyzKW+TW3Li7Jx0iVM80emZAQf6olcvZndisH
NU6a1EzaREdZYWED3B5woRIzGjr9n8ioemlZRfQNcE6/HJPFW/OpNO3LdQ5oQvRn
HUQj0YQqf/TNGLIvk57oIqKdlIIJR43zbYmGZNo+a6cKNnVPUShnmHfoT8J6GvKV
FTKwIKwBZ+AlAP/OkUjCKJ/lI3ypB9Y3VdZaWRWtD2+I9YEjrgG73tqc5YJm3fvS
u46fnYQ3wlANI205KliOyXZuI5ukoPmnNSzxhYUVH/oP41iOCLFLfJIlv4FrGgwb
FmQz5e77Ybe4DJl644+Br7+xH5TFus0zSgX1GCQIxXmI9k6G5nQUbi3lCkH30d0J
d0mNYyHcnPVmVwED7Gyyw1c5CreHqfbUI+g2LHT/Jq8uStji1WWQ3Kb6FGbCdtni
PmZUt470A6Vfo+WTKnR5ruU6Jpc9rmMSrQYWkq/NWUaNZMV0C5LWAxX0ocRP45Z2
TuojlfP7Y+56S0Tq3RcrYI5P0WTQYgejs5HppB1Ufe1NZwHzxV5FYcRHiqH0WjUN
0pBjgEZpM9S9x1oXOhVgyXn6SIndyhiNAur6GWGT2ruzYw/uUo/emp7aFBDZaT7v
7NwC0/YiKC/sl6wkLEFEPpKPRq+6GWdgxA9ygRs6gca/j0l8joW4jIh34iH7bxwE
WVRAkWzD4BVUxjNS6EgzMoZhbZ5a4stkhiUPxKuD/vVnmkqVuOi8lPXsC0Zd/W6l
9YPQKErSqdy3Io4WOgHndoRqtBTRMKLn/3lYIxKlu9ie66NgfqwoRvRoFOEhnY/w
rM7B67RVLiIfle60W9br4UNBB8u91DXfMD8v6gDQHdivL72/Tg6fPZ3clxyBe2ql
R/eWd+NGWeS8YvR9Hpaa3k4ftsWtwqwaL6vlbX4h21sMbXd+eqZsXkEoEGchoUXg
47lVkOSR/X+h+WufGmSariVxmN+SbrDUFFIGV2Y502VI8jFWbpFewE+QkLsIm0Ap
Q3Qu053jVz5IgACvO8bFXjdzV7f9vvV3JOc+pgtE1ga+ZTEJnAAV7pqT3qNukWBy
1eROVadSqsUTA6pWOvDSym9Y7CUNLDkmqr0tAevtu3rYMi8uiM95h7OYofDiT700
LGcfnIZ4wXhkCv0Lonwv44vn0mC1Zj9R7xcZ/ugWc1d2e0/2XzvhgTCaDoAFLm+u
XGMVJx/IQO7WGg4DFOsCcTPyB7jZ40oy8zGIK4cP/xiYe/bVfSS1M9oaCP1Tz0iQ
6s0zc4CUT8eO9M9OVhXg7X2V9d5zx8WtQRMFUMfQEkVkA92Hb6/Jh6P1/lZjmtOr
ZZEJVD/E4VjMIVXPf0PUAEzVdEtdckpfPtcCc3vCfOE3oSth9mwj+WGsoB/vHTyE
Iw4JHXNpLusC5uXrJGocR77rhtWuoE+mjlsI6Gjjb6/dvsWEUfbflXuAEI8p7AEl
Spm6n9vz9JfSKD3+HQ2TWdvnehc/0S7z/7JkB49TDEQZIWaa0pqB/EKE/zsSBfS9
lO5sa8IaXVoi54JRD8A7yVkvadsI5Kn0mAlVAE9yg9QxqezjoOQeUmUtV4onz0SZ
3bwGVOWsCcPiz3f4Qokyb9Vsh2Jgg1cVkLWz7DGSk7NDyHGGue+lJD9JO1oJYiT4
ooFP+zeklidqyoH4LZquiHgmk/33rh004PB3cQk9MAKPCLbo88Vnqs02kuJJzbXm
jaM5b06PhZEOM/6TlvBFhzJWDoXoKj6+0c+9oBMshN1akea2CX9Mzm+KsSSNiO+d
vanfLVJZ3+aqb5ElZhddPElEa+e8nHJ87EsZawuhirmNari/KoAiMobC/G7Qu7NC
37rnwqLU9xYQ5nEvN9oTKi6L9OiMxlS6EQOKToSe9wFQrRb8uU5gm7scaIZlZnD9
k2w38HnbGLUdGNiaUeIUMlKxginfVsC8qTzAJhbWaQVoJjyxzamt7WvHSTosdVF6
8hbKR3VeGJtVTo5iE83Ls6Hx7EiGIPUzqtPHqJfbzKBX2TZLbAj5+MYLrX9gUwWR
SI4u9Kdx2cDgTJ/VRmcwB+XPV0mqd0MiG91WI3fm40/vaxZ1etCb+o2fDh2fFGMK
XJ2g5x0+hUopIxhxmnAJCnJ9iJTBv8TS38dGEckqAbfdGNihY5JHly9/E16kled8
SRsju46D7lG3LYF6vrE/2dGEVzYaUynErNk5xUwQgh8B5uEG8Xu1apDx2yeQex1+
R0kweayvkvOKdbvs13V93w75ghpm177kYgE0AC3VFomA2Z7oV4c77deqpmJHytzW
epxaYkPGiZNSL1RpRdHA8CVoRshEkr7G2dZSO7OJPuuR4CBynOLHmBQUAfD2RmES
Yf7WGiBaF0fUkG287uSlc33S1s+7rnUao4nJWvE0mry3zirERncQH2Vsl/nDWFUP
5mmax59ua0RWIZhwljJP42aegrf6OjAlBcMc74YfwqWYvmCcrl3V25jXObnBFpAf
j7dwcAlpFHjHm+1O0LJvrBmrwvR3qBnWLyEawQGTMfy6DWb00izfeJ+q5Yeq/iuK
Nx1LePFdwy8/bfW9q3T/6w==
`protect end_protected
