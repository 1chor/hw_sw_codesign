-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ulOx+7z00RmL5Kqk4shbaMqTFK4x+AOogmGWXgQRNksOkhroHAtKX63hhwwxiz7XmUwX21d5edXo
ZB30E7ZeG+8oUE0/z+63heDNqatpVYbYsV3akka7ki8AfMpvQf2bI9ls3jTe3xDD1uBD5z0m7guM
STXev+H5dt01LdnqbmSvePdcagTLJFFsEuEsFhVoXR8Q2xQ1Fnd2Jgq/+VK4JK59kt0Qm9t/zZ7g
ovY1CfY28iIbtReiPKKBBUjnG94iSOGRZYRS01WLwZFeoLv/AB3W+IwpoFj7jSmcRn3URRY3OcID
884qhUzwaYe9IhOZv1ngBDaiOwRR5/SHnNP5TA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 190112)
`protect data_block
kR7E/HmocHA88OzhV6YbIuxa9pJ1d0BKFLz+L/ngZH2x+e3qSKfLB2HLbQV5JnUEIPg96bLNihxd
YnIBrVhR2k9qGXHyYyybSG5FTHSAQvlH/DLB8ZvSKjPs2HnF7/TZjbNdl0a3npuCspwr3fB/imOK
x6YSSXFtNvjH+SuqOQfkrPNslg9QhS0bwmyErmPzIKa+/KMSfdk6xRqTSlkPfuwaEFqjGjoRQXHZ
+17kbUAwIE2eJ7C20XoFsrjMsPgKN31vP1BhhRj6Q3GxmRYhUXfnx417f5p6/KRlaHu05PTFNOPO
IZOMAgfGV4yUWMmaJrw/upV4R5tDtOJnsGEJ6Q83NZdmsPchx4+XyjruqTofm5mw1QTVCV46Rt+N
VVqxhG2gZEoUwNjRZxURgGIzWjj/+Q4GEOFa7eAZtFzvqyjCpNKMbwdkdyuHUsoCo8txx/dypYE+
oxghSvyPHCWe8JAAUFXA5GrseEa3aio22dRWRiRM3MPT+NvRIMrwVfFR0k/o83CCG1kxwnRLTfoW
SntG11uyUTusCsV8tDO4Cq+EkyMZ4aDz9STHBxofPeOe5U9DllYZPyKbRSOoSNCFJeFnN2sDWzJ7
eYwULnSbgB24LA1INTb0cQPYYLzuCiWEzUPYmY2mMk8XB4lBNfy9mLraQbkYKPfI5zEXIBLXr9c0
oYCkuLHA3qNYa8f42dLew0mSDEuBpjIPf456nSKKurr9ky2HOZLLxRM6OHZEjlZYZVYIsH7bpZFZ
pKIpIRFSf7r+GrMO+LG2639JiOIXo5s/sG1bFreW1DCzRjgdHJTyrA+8mnhBq8nOB9oFiZ4+Rr9h
ajdg++34N5v0gl9sphJmQbFPIceqzDyU58ikmu++oUQty9zu5GYXyNus+CyZxlI/VKDZzrqNWTdZ
Lk36D7/v8GNcsrvyuDOxnuker6jQyLbFqp7YLEI2yoHZqWKxcSCjtmMnSpPfqUUg8eq1X8+2wfYX
9kmx475DT2vsbDwJvK0Ve+cc4XZP23j/CctXKorkYsLQaXYVKQXNMdJY4P74ohuU8y0pM6dM8SCl
Vv/JaBetWnRd5wZDlV7a/T91LAv0pNmB9X+6Y97uRWdwnCstPD/tpj+HqOcHxfGQGX0bRgrw2nKc
opThnwMWA9BdSzAmGZi+uha9SYQOwv3ueKFI2A5fs+oF33zhRUhVOZQJSFcHX2EEdGf2VRZf8g7P
2R3hPoMFSA8m3e90w3VyfoS0T1IzD4gSqrdBGu786TZOiJwvDeLD3TJhpBzOBIaQbs6/RJTRth2X
V3XrUa0r/M6JTes9LNAPWv3mgI/8DibAriMWnndXB/Cj/Iv4WRq12fAR2a22UShno2IlHg9vt0aV
O6baksBkkXYHee67ymvsgKrD9cOwN7PDiKjR7IIGI04NNQYun7HyASJWs312VIXRwG0bfpH+E1Lf
KXPz7PnfvC//pQR1B9az0Awwnhvtg4XEr/5qSWnNGVN2Lb89x5MT0js04OwbMSHbCKBQ5iQVO4Iv
wR6aJ5SZZ9EqoLH/vwtalJj34JQw+FA9te0t2jeddM3XF0YAI2xAuGOeUZPxAWkfdVD/olb3g5/z
cykKUPs2x0l4KMnhAyZAbqp8VcqgzAxWTeNS+0Yi+neNOW2mEEI24OzB7b+1WCwlbKv4U7k8zHRk
oE/BcT0vgfPOnSm7P24q7dEu764ILuQWLWJqow8s1iV+zGTYhI8F9Fp45BAIJHhMjw11l04dlKg/
VW/ntZHoEO2zy6F7a9+tjIk1KCqw+q696G9z2wDKDf+ikaPXQRs4CFUxdw0GUYMf/UvhmWtnt3PJ
kJKWaxHIBXeahNuOqqhwqrzpR3IkmNAApgKSXUTdtt67NNc3KQZeal+6ApQmXiUbH5Ym0/yjrZzL
+SiKE6AuQ7iw5b+jMBSiU1KW8ep6Ii4+nx/vZCNxNw5+t/JS2j9GPTuSr7rQGlMleXIxhZjrTNf9
ZlLSlnalkwFZSTW3mMgHGY+KxXYBPklvlJ3ARz1fiIHxnrJc96a6DNiXa/2+UYjhoOTT85Y85U5e
y5U38sK3NuGh8EvbH9MGSYePmM3d+5XSmAl4Hbu20LD5MT7kz9+LWmf4lO+jJCg269t5djUd9VfU
CbxJM0CVuidCynPY8Q7qfHKXE/l9hBDb1Fu2waMAWq5AzlzdgbMvOQvBDkANEUVf8g8p0gjigIuZ
t/YufQZK82p2F9kWxGeJUOvtSEMojJLICvK2t1QP8JawwAx2paSxdJvYObEK7DZBOquRdpm3LiJ+
cWNfJ2YrJkSuwj7/ise/G5QkATh4Vn2zBetxw6E9VBSHG//9AN+VdULCNsC5NX+cN2UGGA+DWIp6
uX7lgKVlAm4v5Mduo6QZC75/klV9VWLiJBF1j6ktqUht5Vy6d6dNIOcd6nP3dyJnKUDHPXRItMfE
aobsXFSVyKnWcLMFCxl3Kr8tpQa0L/unEeNNaRFlu1vfp5WIVGlLD027HEzbpACYeu9HsIDG+kTs
bC5Zzibyx/v9yCvlbohcEwJAs60mWmazK3qpQt3kOk94f9qy3YiopxsfOSAlgmyiqelsnDfPmdJU
Jaqx6PQ1M+BlnKRiTUW2kLVpU9Iqi3gY/rRM7FkT00AQdZs36OrSbcNtpSkbxh5d65HUOtqI0lhF
/ToLc0Cm2VyjVmUMBevNMhE5MwuC34rc+Xzo3IXDx2oOBLaf3VaHVvm3z1/vzHED+dB9yEVEyUMt
anZYtolka1KRPAF+oxXc81HnVM11g1rZs2e2tfT7EcehdyhKuKuPAfvm+QYUEvIIaU8nWgPQzrJN
58qx98ANhCmTbqjy3Zw2LZXfOryS0rqaQHpvOYs+VjtGZp+l6de1U9OyG3o0gZ2z2dtu3i2z8DSj
KpXioAXZM869VFuhjJn8aM+c5kfBceeZuso6xfjxG+Fp8U9eC1qZTm39WXtt2EbVS9xp6ohmCKOa
acToGGP8A/CrRUGKcZ6XBi1lTq+wL4XGKCaCjC7fNxataxX6GWDrwnDfzmXUDyTXE40C+dL480CY
qSTKNL11pOHEpf2D3ReeDO9oFnQVF5BH6/+W6lDmpGvT1ZHd1oCpmjnJSDaN4KjpF1K2hqk+wGzy
oy5YOfJOclvRsQYmyNg/e0rqmoTbx58IBvwEchmUNOBT+jrOolwZ8FXwml9xi8C/1jBcMopAqzMk
XjztPEfZsewAVKnxEEPi4XzZu5puqJpHF5q9r+ab4Qf8qADA54SeEAy6Ix+WRVXjOraFawvJ+SGj
8bjh5SUjaADjzhxRIrGoRgQl2ePEkP7sK5FHL6RzyXPFQZv+lnjcU/pbkIHwpRibw6pIMh5iyjsx
SRoJ/iQb0FkK8Dsi40xWuqyuvYDmYh/vDadqKezO8Wz73GYkTeDerXz9+vqo3n1ze9YJ96QVWyvG
2DetcKfPeafaYbzeklhmlkzjvGTd//sMipIrCzCEx8vNuCBbhbk5ZL9zgM/lyMe8WfSZLrBLBg9l
hqgm9skJSqexx2QBZv6vV8N6jxOiwzVy0dRCKzd6NMZkBieCPFoehOhHu4Mo4TVdM6oqPgJsEa02
e/2Eh2ERFgHwNBRoEgXlQEMrzMhi0WBfVMFufWTDrCq9duMtixh897dAk0THY1y2itiKqlBkrANY
owytMXWevn6pZQWD7HTWANTRbvIbCsIc7wSMix3ozd5OUSzm8WHIsXGdg9VztLSUIG/T1HeL5YKa
Bo64cT7hUj3oy/6mzMXCvPNkHykDg8pFQX6QrxGcHn327vOT7yiKPVSE0kIfxy4BbhozVilISBbB
y0GpbN2rfjJHqAYXmiLpTzyjkp3wHOTHz2DTFkaW0tKMD1UVjtvQ5775fi7ZDo06GpJZBP6z1qf5
W6HCBnBaaH3UXqX1GhnrnPZrMro9m3+sYzTAb67WKeGcvDeUaqFa+C+h9xb0fzACCJGwlQFfCVlh
MxoQY8dECU6Eg/VMMl22qppR+qrAqDaY6SayFJ15fKPxHO0w73dWtkR8I3N/qiU6z8UO/sGSI9+K
PgF07j6Jqpt7m74qX5JFXaJDx2HNSD/68iVliUd82w61hWD4SkXbWL/2Ceemq2AuTk9FvwerClov
F2uYKQmqf3PDM6C9rgbzYtRIJmc+Xgc7AxeGtB2/h6No41NHZQno4vpiGSiuYWUBD8KcNOcaegQK
RKIKMwyLD8EurREJqbuzbr/RGpyAVdhG78iEg4LxYAtVSVPOKrqG03PxjMHzVuh3kuYClxPcgDbY
5T1ZrQghLmF1Grx0fI1caZvC0nuO/f8FStNh95GNonrRjpFwBtJE0qIhjYBbWrHkUltqKdEJR1Vv
Db/E39FxwvKM7n8F496DqfhE75qpRCEL4XaBCyk1fUle22e04ykw6cp28bScFJfr/tV98n0EGUR3
6sF9KOG3MPgrPU1pXFhKHLisnHr8dEXmX01GedeNa/p6ZRcuITNuKjakTZA7YBSBuhfq3uYB6hvu
yslyGzkf0QJrA5iCwZUAeDB62rEHFNWXSFwpuLA5U4yjCNG5kSVXkZPUOeYy90I3fRyd9Obq77Zx
IW90QC3NRxkX9c1nknJOkzXeMPBOsD+7Eqp6rIoUmXkk71VPFbsDxJwnml5Lp6McQk9zZsWGfFwb
zbj2bhXq5lUmP7R+etykz5wFBVljuPRwrFug4A4ZkngBf7hoZS9p9HxsL0ev8GZOM4vNMaBwoZv9
63P51RC1SrvChIb7wiEq+6aV2mU/mXGJTVmxKanoKZXud1ElQqUV7BwwnxG9xai1P/52r6cJMdTX
q2ITEiiVwEC9ew27BwhPFiW+Q/Rl6l1xc5eeyQrFxZnLN4KZwgLx38/utQk8yo/ASBp4WUm/8DnP
WCTXN7iSgRh+od/ArUGwlOpmkFwKcyB50eGwAvGTL+he5JFQlDkD2bcReXEsyaO4rb6BDqzpkFrX
J8oNno//IcnZOFpLHzrJ9c+2QcyLsA6FSGJeDNs5lDIEfxK1Teyn7WNBREj4//HCIgf16hs0naTS
9K2GXChq/Q9QEcoJFZz1CXVIThDENne9zMfXRN2ha0mmNEv40HwoIJWGBknRTXV4PayH5ST42yNj
thDqi2Jz+6+5I4ioPPF/zLfaR1/ZxW9CiaEtigaISsm+DuaRJGI6QwtiWwL6rH+4vL+MHs6nt3Pc
JMxXz6X+WkPc13+pHgTbfTK/mBsLjIHCApRtKbo276FFFuwW8vFszonBDYbSFgCPP/HLEOU0PaZH
LQQYWTEU5JcPtMXJp0tDfY4VHDQwYJsJLyTU+gS5/UNlI6JcgUTrK42K9ilM+ZOidfjnP9NoTxvB
6K1VAIQCPYmeNb1NBGqirFX0dgX4UwdVB/7aGRp0wy14Xav2GIcE0bj/8roHg0/xdqF74wvXcWz8
2ia4ge7BbUNZPGnERjEMWOLLFXl73qVrzqBt9eukt0S0/9eKiRND3h/2PQu/1o/FVAxUXuiUPBeY
l6iFH5+EnPG1Tq3xpgBdugxLjTsG3USALR51Ls9kXv0Q5TxHzd7drucy/dTE192j2x0Ky1jxGize
0cFJ6+0fMKcyD4xkSTPRX6kCR5tcAquRUL4t/OXgyC9C4pbf/7InA44KGAhCy3Gugh5lPQquiQDA
T991MCCgp31+Fq9kYizipOSbve/sX3FdcGiSc6wnV1boJCUFsZf5XQ2bL/DPkBoB51DmiekkLDLk
5RUwRAs0WwjtOo53MkpBjJsGNerVj3zrJcpAMRc2n2Gcjw5OU7AZqLn5IQ3DrDIGRWsFbUltrrog
NOMjHQhZ4WFRsqQEO/XNcjW+/ji4H3iXPEOAQt75jv/4OHzVZg8MNmPMmgjiLRzhM62pwktWtc3r
sHBVhTYfhzEI5CcV17pD0+wrq553KcPH51xpnZDdZm5aC7eT5bW+JWaNTmkb9kk1z+YBFP6kNeR2
Bh+pcUzLtHesod3AHjWX1AwYnx8E/sg4x9uu8O5EwoYU7sUomJnRtCApKYExxIi/2tHMoxfPvD4I
61zxaNkTmhpvgyg07dYRKMSDWdg5Qpg4/tc5KIQND7/2GIhbnot6vfxAqRbz8GFJedafWim6RCWk
XIAD07uQjeWMGpo2eNlWnBByU+BFWIFClWR2U7ZgqBJmguXrhHlT7K+Hhp9u0EdAtlWJNDBpac4e
cvkE9AHilW1psnlh8BBsT8rIu3pGUVMWaqaHcTJ1zv+h2lyStVTfz9NgkE1yk6/JZH1nANSEAAVF
I31lXIys2oWhJMHaaegd5aXVTsTuM+nFygZ9SzK9U/sxi04h/XOLZWoSATpNZk4ekm8yKV2lxdy+
insFY2FkzX6Q+34HHzskLFwUNg3dghrwN71947lNZAB3iRWoKJM8sZLJ1DB651h7ob562kffv97m
BP7AYf7U69Y8XXkYC2av+zjgoGr/qpn8Hqf4/Em/U3Aszi0KJ+P5vZikMWYtTtW1biXAkHbRk0aU
hafL04fya+RneKUKqecsKM75kQTaw/MSfUIAqL/msfahTOqZoZBwEB8f2Xo7C5ylAexSwIQdK/Zf
GoXE3RC/6n20xb2cJY3U3GVVirYRVP6LClGJFIxABa7VzPghkuvMEKJfNrOF6UxMBIko2MxHyeCs
6PtWu7HASeg1z27GKwrtXYBCKmddic1Duq9nnI20E7id526larhFJd0fV53y1maArPO6GcFuP/FE
VpU2Phn9o6+aBN9r5G6hGFajD5U5pn69XuHhGcnk4YzyniAdsAra24ilG3EOPhwHa3BXuK+Ic2lN
scg6mjdpGTgt/ry5cxYuTYPQ8lzJ6j/0QHsFKq/POCQiXZDhh+WzBcEKwXiplKZtPZ95FVk/cKOe
dwIJ5YLJjvSWy4ycH2bTieLwNh8p1Hfok/1fd0yEeTMPI17rotngU/4GJ++nn5wUuXM26z+uhOYJ
PBIa8vvFPboe8Q1cNACJa+wgEg82GdcGHG7sTtdawl8evb75HiEi3unz8Dj6bJUQOrjrqKtUJQO2
1WRYc4SL42SBTwJXIavSC5B9GVO2nweEMUJsmrSq2cvvnfX7YpYWf+XvhQLEiZ1z6ekUHnllNPjS
E2J085uGfpESvlz7VzDwxg6rGMBguRcOz/Vy1lbUuyxnL/QlNsGupSsObZ1fA6DF6RUJSU4B/Gxh
vDO2tDf9c6pQo4XGHEW4OGL4rlyhTg5ETbDlTbt/JOIcEyLoiNmUjabRr9s09mAOdp8jHUkjWxAj
8bQAQb9Z3Hm2qTQbnHYXMsr8zomNU2HqiTLT/fJokRRABdnG5doGuJ7GyQKS6OGQMuI4gntRs1Ib
TtFEF2yYnKTDfewXHMDTf96Vpm8Xdrny/sMMd664JyOa6sg4YpEL8qD03TtLtuXsOL1/aikV7BJQ
SsCI1kuHAEh/zzlFEQzCgjEUbhLuy2wibFo2E6QEMCwpghDSUvM3g/hK0SZYrA8ydG4Jtlbrl302
PVG0Tb9C7EYPAFVFXFLT/thxdEGaQTMGX6Os6kYCa0aF31v6TgR3S811R4Z3HNAqn1NSIddo3CDu
t7vAFM0REbaw6rjLrzJyFHSfivHc7Y6ndXkmjvZQDp+bMV8cO3PoibLVaF2UOqIThwplpaYoMBzx
YyxJjJEyWRsv/8eSk2MToxv8ACnN2cPrUz2SZgEJWmhFWUuOmkn3up4SDYkG8AXXgWpboJmoZqhl
60Z+cdvItMn47JVru8PcMUYE+5+HMDsahzwlvr0+ljhSMyHUY6RmJpp7Qte7N6a0AYcnVNf5b+X+
bfJVaUkmje8NS9We4f2mB5wNwUPrXHMzEj617NUPb1Yd+6DngCD2It4WMVDzuohhuONTDjhgjn8m
Tx8/5b7ZX6pVHv677lYOlsjE3Khe5cboRAp97zjCXF5XFx2aP7nHNy45MUom4B4jYrBds/Dj1UsS
qT7hfHyE2U8Pw+7hIiNzGQnYCD7PUsFwXIpaYMwAsk8mf3UnHajNcBFNAgVeu9iIi12OfhIZwGa2
IxZL4ASK0BdX+I1p253oKkKB2GJO4TRs7lSpUZA9i+hGDeV4dQb6XYgp0WAcJ23xixFmfI4HjEqr
07gVEKfBR8ETWN8gwrIoqA38krsBjrWNSGOguGiRs3GIeMzpkylivjTa78KROKOGIvbT/Gus2qgO
5qhy/Vn0DX4tUo8KfeiLO+4IxQ2jbmL0J1VyMyjHvVZioyfqkauT/j1lPL61ZLcM5u89kmYD1pM0
BurybciPrIkakftGcOPPGiM2QCVmFwFAoHBT7kPmrR7sziyAM/YprNX4t234JpxEBn+svQYuFhKB
Dlv/rQkCQkl/kzVsrsqEu945C5aS4ZfUgjg88O+H/hL8I9Zj/KnsIU4FDiZkZ5HOy5bSbAGU+QnN
b5YCFVP0WJ0nCNUKZKJ8fnL6dGBhvQ+GuVBa3UNd2hL6B4uqfn0tybYMtZm7Jl/KxR2qAiAlHwmk
5KlnuGGI9FyFjLNycKtVSQR+949CZqEyGzY7GmQd0GYWeTUJqZyYgE38UBSiC1RO9G/hKTzYw+Rg
i9J2AaQ8m9K3sSaVLoxkg+v4lILjYLnajXoArKgqi4Z672LSIJIWbP874JquG7p/Hg85+D+gsrxJ
ScxQnId9lPUCKbCypY0XmAenh3ID3Rbfx0CX5nRAoNtIbhp2b0sb+/tdILLEXqV0TfCC3nQKTyZk
sFdoHZDwWlxLksR1IiCtQjDn1VM64Q8gAEwXs+kG79gQHjcLBhN/EnW9rgvYyKoN7zEwSGA/y/L0
GJG4MijGsmH8cZwXIsyDCGTD1RmQNO5JDke25JWRnV/2H0AYU6+9u4b521hJE2HukMf1N7Wr7v3u
UiYYOd4Ky3DncY4fTew2HL9Mz5ROhbGm+BZDvPYBfSQeFk6TnR8JuvvJQN1rGWt3GakxLSjFEFXa
0yYe+7gC33hZorAzNDvLyAidObR3GuSCWx6jLpPLVBIqyAyDAXbuQ8Xa5iOyNi44lFPxFwzXJsVH
w9/yT7w9Xgoy0apm96YCr1Q0oYiyNo6K34Wm4zk/4+LD61B9AyD5oNDgq+/Apb+ENdGoGc9Ur+Rg
iS5vFyxPbJQDF0/hdghnDrK+0pS56YQhnzfputD+YNsWxWax7TV04JRmGBXL7enjd2z8bOv6raCC
c4MBBRCp/oH2fF/RwzDl0nykc2hmcll0YheLhU2D37w10+WZaaI3yz/6BOIfajeD9YITNeazGr/B
R3KrWsx6Hmvcsigvda2YZFmB9NefQYgXews1tzfY1lmBZLq6muZ6RrXaorEI7j2t/yVA3K6JKLhI
JEFLR6lKvOV4pSy4ZzrL8kp0IWh8rvE5dOQxdPAlwUA0IIEK8P6FnKfrpaOWDrJ5lDRvYDfn3ZhE
iHVtTUJWjZiX4BuamsF7bGAE8ybg0SMTdgIQzcaC03pQDKFa6Bl0rLlVSH7gIHrfPkNJKdFyF/7L
cYfXUYg1IglXTTiCuGWH9SSD8fmeGpKNsoQnfkKT0pc4CeOYRBova3taqlsdphQF7PPxhn7seSnO
UOPvsFczGe7jgNXSdqH1HCOlryUVnaBUkdE7q8H+kBuynjFx/vBmcgieqjWweh4HqMNgMV0TPt6O
cp4/MlTA/+dVq3SgvKMB/+c41TramtORQFLn/pffFgCwFIINhiMLEP26wPxA+4gAUymNJyV86vFW
wI3xi01Pwry5bV2YM4F2p2WA7a27bFgeSzj2fDEokR+OpJFHl9m1InTTN0/TMMee/Ldb5Se7dl2x
AB1aSP7dBBaduR5kW3+ckbi+XJgsxXOTvsyNfIYsExg50hBC0G+FnpcQSQIlHUT2EW5NlUq6DzVL
8iFyvqpMuozRDAh9RBuWjsuXQu3rZL3wkm0F5nF6/dkNYtqdWHNCA8QtKNvqg5O9TmzbfCrh/UcK
Idj8w5fskkpwx22DjrPYntUobvBxzm6BFOH5KwreKw5B/0tQUbPGexfCZU/59BOug1aaWc8C4iFt
6IPIrBlpH97pRhTbXBvv6ZICwUDL5y+GMFOzgVhAIWnLREW/PFzlK4K7e5xMiRhTN+Aixaaay4xN
ebw30fD+brwkGhGa0SxnMSRXsQ4Ax58NUOSwmJM5i66IC8Dr/f6VTn3poT3T1TDc463TLsY0OVXy
4iDPbNmA6E92FlZtmB3ieLhiX8QCuKk5Gj3VnWRZlHG0skCcZ+krXUFEZ88ia+egZ3AzrUBn3F05
X1jwLaD8ZujweLwrs/1jQD13snziAZ+3x8++JEycdzQJVK63JCyjUohAGSfih8Wq9g6xqDnuoP+u
KlPDo7+lNJStJvxlHhlaWR/6N7GN8jiApqIe1ih+VpJAIEY1VAbhQrpVt/5d1WROimRar2nHdXPI
fbekqQH7vKSpcams3uT5BhnqdzzThwm0a+ozNLDtE2T0OHYWtO2YX+B67F+s82PpvaBLzIPVf3Tb
EpRBNEWMO+1G0xHuzTsF2bcsz735d53uTqKbi3SlnkUxsE4rp0auW5qA2qpMgg4iGaWN2DOx2N8f
xYLno6XRYVK+MqaVrN/cHNqbeljRSk1Pg9f5/NLJPKxn1upSuRvTQLGE9H6D30NGapwzroVXvfUz
eH1MUeuS4WavFhaD4fd5V2m1vja9Blzt70RycchHSJ0spr2p6fIpKAaldpqjjRn2z84Qm1yewMOT
SusEaPe7wNCD97W/mj190tMByHAtNbk60hpYJqLU+gWfpY6QIRFY8fOiZKnuS04dy8d4stwnrnQN
YoF6U3nTVLjRC7uUDnoR9WPtJwjJrHq8K+MCNogqRE8+3m7ycPidDRWLQjbXIzd0oDu20+oJPXdv
wvsBYK/+CQiz9QnCXE92wdGwt8wiQ1cGHBwxRvsXvScme5QxLIyIPv7E67m1M8OBBFZotQc+u8UW
H4/dBzqz2cGwrwabeBSNWPpFUMyth0pTTagV+w+aXSsb+ZEk1UKBY7D5j4ttSgZjlfi2zB9aC1BB
lULHkvWPDYuC6ljPdQ/cKF2zWuQW3ZFEn35EwqN2lX3VMcu+rxaFcVYP6GKvPbtZsx15PJszQeQg
Ap+DFjfHYsggxy3SlufeKyZahVPdRJp/lFU1OU7HwV2o5dyWg3IKZkUVx1NHQBmRVVlRfCn+ZFpD
wnPebx9cj4ic7BZ1cyT2zx4sRC27bDaPMGiyRCLv3aKBIhWj2CYVj0ZcT0xX4gmGWSU51ZVxEkOP
FzPC2IO2afL2R3b/i7fya/jlEyRwEwaf4rwTlSfsi2IPMqOeGG8ZPpKCVkE1QEVnUv5ECsV7PMl6
OX2RvNoaWh8OVeHbIc6asL0k8dFaa/Qv6aBAE/2WpItwrH5fephWxpL6vjPLh7azZ2vQ21KiYeUm
0Nh5Rk5iU1fyWFTbyCBYrfyPgZsNEiXOBukjDyETLy79EqK+jT/SvuyDI0YZVe5Zcr7FEr6q6ntA
1U1OMXCqGHvzcXfdgPJ8kxUYmyXixRBkk8UefgfEaPL7wECoDh9B021mg8pQX7IrgLdHIl2c+vUT
cVWaEXoa48mOhfDB15HnoBsFX2wNEunsEehnRaPjZFuUckxbVuUoK77NU3d8dDKCR3wehWNT5QDO
tthXHSK0FdiEAnjmo+rmbBZkw7axyuWNeIvjQvoqS2Y2EVYtTOZx4frs56jYHoDhdQbFcPoqu5Lt
2PtV3KYDFAbHuLLxGiyW23pmqycxnvcqKmrfy2Il0orm//lltMFVroWqMTPs3qrv34syPr1mVXu6
p+fkvNyep3eoh44r9HpJx9yymZFd1PwaKoFCca93i0KTK9LU38Pv/6NFXmAw8Vegwe8XbQqOKeVi
M+JjaoqPbposWwr2Q/Lh7Ob+0yui2pB42RgCR2dUv9CsKimz6ZXyL1GfMxef6zT7E1y+i82Kl6do
3UhfFnfjdEmYUjylg5pTPmTrw0vajEINJXzrrhJSsx3OM/xLc2Vn0wGqAzv6g4QA8JKlMvLeKeNs
6a59exXDVkWiAuNxhe1yU3Zd/4+CmsPmNltJvTE6zTiLYmwyMmJ1LHggc0u8g7laRRy2DOvQzu8C
QO63en5G1LaGLgZtIx/2RpXxojauKwTm2q2xMrx2Ryp/d0VqKr8J8OJl4pRpgc7gRTpepXEyTq7W
ofKBZviwvZZ1YNDDUkjxYR7PIaeCoyyL3EIY3z8aYiVzI92VT2WIIo8FnPDaJEVtu8qipZo2Z73J
fuG9v6FXcqWdhSu/Ok2Hqwm5sI42daAh2VvD6o/DvQcMp0Xr/Vs76lq1ccbTxSTOtrTJb8Z8/fys
3sdD7V6q9W1RniB5PqKwTXI4WfZXy5nJQkmF77iKysxEvqp4N4P9p62RXCZxMTVgM6DaC5VQXArF
32teBbSu7yM1qyX2YthO72WEubbey2t38PtahbLAHY4xaafSJVTAWhmf3T2hONZayBKhMx9m2lzD
LGCXr5/rAbTZgbiyMV0vqcTkHs9L5CwAtr6WZvXY4cUljTA7tjlz1Fzd3B05qKOWcob3YE6hwKyX
VerSqxg0UMz9SNGJI+Ts8jfUpaKXDDwkVYQyxr4lu7PWtWao3aPXmJhgpN2hk110AIPF23XbwN9r
d/vxaRiss+sHCcNNSKOt9R/tvfTurDpJCoUJUysoXny0rwNifV62L9bCWrKy3wd5A1ubctMyb5zp
L2DB9d9YIN3k3eWf9oGNZCVod8DJp4ONVTuBZ950xyAKZ/fiM5m3LDoak8DvacmwuFBtqlWNXczo
0R6f9F/ZQ7MnzaaUap3tZissGxTN9m718eVqVAX0KDkPgWGcYFB4QmCmIUuv1JO88ob6FQD4PqfG
LGOWqTpiwGXKDsv0ZRmi3H1+NUE8QpOMox43XeOxjQW+i++nCrTUDmNJHfo5sERsSJqt8Kn4TSSb
nfe0TvGlE+0kSameleVdIT7RkMCrU2zTzDn81lDtMskvbVElCIAw5HstfKUrXdtYZpYaTJ84LRV0
vyPHHL2htZvXRyZ2W6ExIAdjr/yBHPisv/M6LTqyG5TSoerknWgCj6lh42H2zZI3V68JJwIQx49J
4kKpdzHK63hN/2yjevJti529NDKEOIrQASSHjLwlRAjGLyKGYNJ7qTWwi+psMnLDbn9hbEWS71FV
tSfPcfYhNF6Cg7Obr7c528ffKIEqC4wWXb2O4huAiYW1wfQ8aVlvajCEs5wG0iVZDZyQb5znzed/
fP0gX1DkZ7PV7q9sG4mkYhN+eQWJ12eCmpcfbcZBiaigx0XqHFiCQ2lwMmRu8CMy6l/IlVFiEqj3
PVaDUSu3vZ6E7po8ZLwVZ+f/XdnzOp1M0+aFcDkOJodm4dIPD4NPwvuS8zHjzOue54XuqVLYHlJJ
eTRa9OU8AEoDWRcsz324QbLsWGbPh1Q/F3SaLRA5Niy0wngowWboVlshZ58b7AxmQAX/E1yqjnev
UPJKC2eT99dIE0Vr+UxEM/LNk7MTngLwROyNtb8ZXAIOa5VqJgwjw6PdRcxfm2AcK8dQFpXPLktD
sb+1WIJ+ip6O071VKI5WIXCf+MfUcshGqX/lls3N1TFcw7+gj1VbOqBQsi1pxMGdtFxLtqbthRs6
uZyfuw0M5zI5apY9VHnNFNKQQHQqBkP86nQ6ZOPkdmsEyR8qu4oRfmtsaJhLwXWJB6E2yg/Aj/oi
eMLalfq9hhHXQCPNpcHyOAZOVCkMkgl+LJR5CZwJNOQrIM3vhCWtZfr782hkvCozHRr/cubDDeAG
ubVlmerBAJBds6kOvjKw65mqBRdqZ9tMR1K7wBhSOJqN6IfITHBzeD8r52TO3fMxusFgppuw3JZS
h1JUht+CNRUVjcPDkNxTNu2L762DUE/MvSlQevYvcX017L5J/zTsKM81pv88RKUssyJZZi27ML07
IsFPD6g4r221MbK3ItYqNXT5z/TWBzPEw7TadwOGxyuEA/7Djec63vt/n0uXVRmr3oy+k2OkXSyU
zarN3p1hOmiMqsl361QNq4qAab/zvv3DY9QVUrhdmFf5PMLNcffhIVBR1foZvX0qe2zuue42LFO2
uhW80g75w90ZPvZc4dmgTNskVjm5MZcBaXCkpK+ax2PkdmOuU9qy6HSu5xd7gtSZ16y1AhIO6kpM
sy01gcdpCrAxUHv2eTB6gyNgJtPCooSDsDTrEwa2BcWm5O837kZAeqAO0/fRNfbCDxn/VuKAIFx+
8wPVq3Zhu0BZDhZ1kh97i2JBL6XVNhRtl5syBsFravNjuxYh2NM8/CTprTIlV60nj1SMp7rsN1JE
VdJKIm6Z9BjDFH6l3VUUWy5FI1X5r+WqYliqehFwIhalhDKAeg7oGsjmbR3SRSLiTikZrdpNa1YZ
M1zTDP12s4MeBlWPGLerRlXev9DzXDQNevnvxIHqdcnZ075pF4XXPNcnzL0NReg4HyMdneQzK6Pz
L3bG/mkhexj//rRue0oCeX5vMzPGmEbeyhddwhqXskOvWQVaVT2EAjNg4pu5jNT+jnEKiXI+Y4Uk
W99CNMmbGZFpOlaJ1FeHG/WNs6XG9Db7sVN6cN2vFrR7P3sHcp1Y1lKuv5JOhWs0Auts7Uw3LcLJ
GIEvIn1HCroBfCJz1hf0DPC8Xtr3sJ5x1/6ThSX9QrmGKmuMOCtgPRnXesoN2bI1BJQp8nEg8NKe
k79FQr+ns53wGdqOgQMk6jK/f/f1VEsziG6wPFXu/NZ+kqWjZ9jssLbuJigLCPpvd7wZWGLjvTUm
rA6qPZdkT8lTaHX9zMXFdzuUXlAgs2HY2Mge0d91SsuA1QEOml3xX+5a24Bd+b8Z3LOXAlEqGphI
rCbCb6Iqh2LYGVLvyFdXKpuOvirv6h3Ce0Yr52jANt5zJ2zmS36Fy1px3tnAUyvhY8GUs6Ka0dIp
WXxu9MZYYlO5P6PkbV2T3BhVyXzVbcuhDe3Tc4GrxsDV6uzRK+u5wwkrbPabfrxlbFWhlbDp4gaV
ZeQduE4TQ4dNTSM+l0oz2LZ59HAZp11e/C/cNbbgfxzQudf9zu4/EWmLhWiwI/Re9Y4vzq7tCW0N
HkIabkF97RAvwM84ReNqO1pVaQfimwt9DUISku4Nl9CdDD9/fqmIGrduDf/cKSZxAm5CZ7GQphpt
wtuTeqWO5W5bmLuTHj5Yblw+x3tTHydawVNUpUAMejoDePvI52DmMeB7p85QXtRhze24SL6PTHFG
9AK9NgJoiJ22BQg1RdYowKxkUdalkaMbGE3TxSSNC+0aH+C3nyB7zmoD51EdqLc32z7fe3hJ8Zqw
/0iDm2622cSL1XxlvKPkppiM8Imm6/PjVTK6BsBjPXukqFEn1OKeK8nMhCNX2LHUjkSDJhhmeckt
tcsdj/h9nvqJvyKernnoGcwpzSWSJsKCV+UaPdcmon+Um4SvOCQH0uHLa301BdLi4HHXtrKV9ykG
bC7JmD81rFQ7LvXBeag4LN12FWZkqWJvx7KOVZ+bDwiKFV8VadRPSrS+cWQZoXt9JQjZQ1bDX+eb
KeotQEFJkhhrIh7nrqpt5yRA8SD5HEdDD5YvJr4vdNyBLCWvBHmD/IIRUgMluH6xmMsbTpOS8jrC
eQxeZ/H+SrwVkG1tNVBoLu7cucX/nIHXnMa6rWjjLV5tqnsyAW4a04YBaFfAK2Bm09MlmYN12qde
ZJoy/rFXaMKIW6jcc8+eAXyNiEfjONiMkCZ1HmB7I4eDnHLKE6IJ7728tr8Q2QWsXHLjMRHA7v9z
W5HsRPfLGLRvqsHkVrp5wKDGAzKWSF9atN31+evIYNXYjGMMtBmZhu/9e/Cu8iA1h3eqnndnoMbE
dWm1ADjAaEglvF6/06/EJwcMYVRmEv+1zm9fPIR1VhzMkaZlHUY0XRN6PvPGS/rAbZpn822hd0jt
IGC1rhz6HXUpplb4R/IpZHKTzJEkZ7Z85Fzuy9I0FCMyEIAMJsdUirNGYw+8uqM72adTkisV9tVG
+T7ot5rCjWgezOGPFs7aMMF2P64w7M9d3seMlMPbcj3kpiz8m08VHWLLJ8hFq1E0jHIQ00u/XPy2
Pw5kIMausDhTc7kN0AM7KBAOJ0RZ3jkJOVcAJ+0kv3qSpkWMdgzJSSH6sydf5GOPm7jwDmCNspxP
S+p2aEfDT1s1ENzSLmiKWKjc2EScfFqkFoxudsfd3G5mMICaMRd4wumhmbgAOQ6I8MeFpFYPx7OW
gR7rpr1vWiWWPnKW0SXJv433w5nyYhESYD2JOkVCwG69WKt3e2Vp//SDPpWxTWSz95YEd7gWsveX
iZ+aDmS/GZi/aUuR9uww6OJeZyiod21NZT8MGw+zLH9afgJJykEXpoOjCYW5PXJONW7yhh0Buazd
3gxNWwpmVPTZgqELO02dZhls35R+7ptUHo7mHe/hBExrjFwIOikBlfm99DHnp6/SHGu02PjpEdpF
Xi+GN4/VzzegkGLM1zIdGIy0wUgOK35VldfQaGOzzwCbOb9kF6H/q/9Ty/9GgGVwMhE0UyXPcYLS
D2mSrFx1muq9TQ2yLNfCm9Z9Q5BWOxvIbW8VcAtNry+7PfUmy9/zIJDxInRijbt0Qcr+mpe2gNhN
+b+tk9jDFJu9ZPNmDOulmflioX5jpOwFjqV+S9R52Oy/fDRW5Tp+/qS2/Oa2MENTfGCfGKq0yAQ5
uZh5NQcN45eNLtswh7P5NRVuOUdxi4H16HRjNzCCtYAUIbiGDaO7lC3ml7++2LJJv7xS+OS7aNq+
X/DAcFhmYFBWKxQwmc3xzJisuzU4VOaXQgTaWvp8dHsWh6hc/oLezcDc/Y+HK6AOyo6guMhXcxMu
YCXNzeMJJMzXiIVMJ1o03PqgyArEGkIJ8MrrYBZrgNVYfiDOt9pfIRK0p2wt+H2QCZRXJX82nVnC
YBn3aW/ZArx3neEYBQvo7omSGMaZs5F3C/3oCG7xg8yYqZzR1BUItDne98fcFvpCBrp1ifQj91Mr
/Oci+gAoSuqGl9/CbPDHAv9133LJQgsokYaFfRXhmWbKRA9bu+9joy5vhQGfKRhhrZ2iG24rgdGS
foFA4NiIXAI6kQnUb1oc3S2rp5JQmFaEJ5+JdB8ImsyCfnBDrbQ2yRp3qumTlOm/7BqVLvmLnGim
j6PsYiMhc7WEGmymkUxOtoO05KYI7bLOkY7aYtzU/wmPFLZLuT/BdQ078k5Whxjsnr4ZoKzmPRNk
+qcpuVe2ARQ0nB4RasR6An5eBQAsJHYr0hd3vz0ZO/iA0ra0MGcjoMe6ipOWt3O6FP/4YU0qkLSZ
E2o/8wXa9oW0yCSpqd2H/cPe8d+4K9Sa0sVFPXzu2cDx3e5JY9mV+bUhRJ2GyBnBzqqZY3EHv2H0
yqYVA33GZ7nZlRihcn4ZEqGwXstvdmAGzk50qf6x4TXh63brkierDRkwx4oakIa5yHbMQ7+fXE+5
CZP2b804XyV8DZy6muYVWj4q187r92CSrl9lmW0yNpTXa5dZWTW9aruacuMRPrDvzeJFiHnr170K
RBRXAk5/W0SZ1CGEss1zkawwfPvR3FFJj8xjoWqHY95nh0ToFBxmAAjNB1dJh1sJKd4DkKfptwwT
xY/pONs7cCFL2a0WWGItiq2FAvZjuovuSPJSgvG0pvOkY4PNB/NnRlCHrtJkdQEBC3gsmkGu0jSY
aZzIftgjF/qUNRnX3Pe/fbGtxTblrchxaruz6mt+8HRHpLH8ufbIDgK2Ni20NiLlajNTe99hrGmZ
B21qsuFqrBqQN9s9/jIWcZaGIgD0UaGoW5zy1p7AKm77YwS4Ff/n3T/sGy0OQo3GsyFBFSpo5PUq
xKLdeZ4Di4i0bqPNDLqrC8VONi9qJWNy19Y7U2v1nPGDjh/wasdw2S0bnInMFn9CK2xWwVNJvl8z
FGI+fZQkaF2TSBztogf4rw2cZUkUCC0xNKPseSJJ9YSGy0kD6KEhvUnYLau8Wp7RZdMPPr2ZpxoW
OZB9yvuaHBVjqE0OruTKjSivoRG4YhCxC/QpSD4dglaigF02uD9qZi1g/3wnACuTq7kDzgDNfOsh
VbmHO+yQWRIf1xS6csrc2JsK1SXG7VOW46HGidOXvl5WETFqjW1C83zDrFEaxIFXXCLJ93SWkrnB
anwEYMxuyXPwpyli7tclBg8Hy1XsT4JQsW3z5gk16xhZYA9QITLUBHE5qmjcFSA3rS3D6nlB8wr1
7POS8d6GGIS50AblkBW7rEyGmyCsYUeKir2wMe9G6qz/7+CO4hWQjufZ/Z6vKLi0GODHFf20Wd95
wn7T8BezOfOXsfZ9b7jVqsDNkt3uCsJIfG3kDM3xKQea5q26ZPeS9dFXLLsplfCwtz1mmMioz68h
d1K+aRthedo+pGhESxghkcmiD9xb94XegZa2Al8+Z+zPvwxBkAleIeQCz3Dy5eBunAKVr+AqrqBu
ln2Gh0jktXVaJWcI8ly7HBO7qBecEMsMfm1DtgChuvaxCEp3GSdJ9VUOZCa5AH8JiliU/Gh1Tuc9
JGUzk31VLr04bE2HyZzyqwSn+1AbBaGpTiyBPJhBPh5TQuDt/zuRHxdcEwIPlZH4sxwfyah7+J9H
TxFIH34bUfrfYsCunHtAmnaUujh7eWsUKt97AeLYvMjCJTuBqPs6aEXKURZ7Am3ADwjqINK35tzP
1O26mOSZlEYc5KWbSSG5uxkbsTxUDl4RJU1TtdB6iUzyFsxG+InFd4dV5QZsHEJ2wS+L0XcLZ5pA
SVizNnydZ7QXbXTZNQMYZ55jexN9miX+9gd7cr99QpMG5usxLmKToW5u2rwZYfzBdfIgVdCV0wYx
wDxeZ7eeCUcDnUcDY5cQ0MLW/LBBdNqxa3JJE23aL56gqNVhhSiQ7XjbmKULiSWAKp6PryGiO/07
4aehNsN1xaudecsx0SxLb11dMwnf9rJ8H3YB9FI0Mz7cG5NMtuoaDV6PpUAAUwODeouTEq4ysJ7A
4TbFf8R/vPec/yteOMifPlKJspQaNsCrdzBX2Yuy2G4mZ9oWBYSgJRcEGr36kZPyQHeHxHqGi5Cl
s93DAeq1JqGNRtLo7mOuLjHzdY5DnoYBVyRJ9Dl5kflAFrs+oTh2rDunPCINHvCt+ZcF8NYRWEXi
UVaGjJdI9VEae7TMGo30tN/ZwC0AAgLZPUFVqUCiAi8GD8ozUNGz2dLtrmpzuGboaQdx7HOBCBfn
7Y38EtNA0lTf3nRDu4vGoUAQTPnR6kPbI8CK6vSMbPnTHgDR3sDo00OLNbnGJi3zz52JNyzl1TyF
RlYeA1z0XN5qGxWyHXjgVKjiR/STyoiCGfr4E1hTCek1/rlfet/0RF4bWlTozwH3ztcIpWyhS9RP
nN9tp33sGFCX81gzVrPGifh5l/PEbuXhjWff39c5WBJFUd7iNzt09ZWUUcKtMkqd7crXZMKEA9RS
Y5dXU5t1/wsawba9KLeRW/b+mF2W4SwEZaPvyjvrkpqYhCjNCOP/UqNhAP3Rbuyq7BUJnbIpaKG7
9pgTbfjT0/Kpp6iYb6VCtKq8PHh+V79nYLl6DCB4quAu0sKf6eSpOHQesu8jLt1zZyeHCbaSrQNX
svFKZPgVL/9X9T8wrgsYWOvrMxLDAGl/LCsNqIIiJXKuYll4+bGbiefE6ZlxdSZj4EZZ1ybFnu7W
N1cVwd95BUnTQ0Oc6DFRFV7HT6y/n2uUCSQMo12EQoVCLLxr1ZF8KUjjzi7JgHo4Z0Ve/q+Ug6I5
f61mBO3rNBsc+4R7ZCpth4gkTkEewwG5iK0caQ71HYpKSYMm8bHJD0YdJuYJIhRBumDeSz30QdFT
q1SzYYa741kz3ntKqUrSePBmQFHD5SGcEfYq0XUPLzxmPSEmL0z0uIEB3yD+sjgBnpCo7YyCeayX
Bgcj0sMcJjUKRjUtmTPnA/G4RrMS8cH+ZZHCfk1XDAVZfOu/jy44IX4uV2JeTllLJxCPj6dkewWX
cHZ/SP2PWu6HhrnXy6BGDwOYq8e3FzYlEmGh6kN1VnQed9ipQWoFzKVjCpYvn4psy53NfSj6DXT2
VDrQyQFtpBZCM1eGUkVlIVoEnienpZLGmlESxnsDjJqAfcLGiHDtbNiHx/LsNy7+KWCkqfShwMuG
IyRmHBBK3kVZmXNLV0CovNBbDeaMnvWJ60P+fFeRwOpYD9LuPvOilECeh3rhuUTTQ0qSgzZ9eK0X
8PS+FBiwCsqW2MtWnYQsdBeS8c9b/Uz3f4iNz1mV5gpjqybSax17HAz5pyTiHkvYQl2Hzwt0kCcF
XbGyq1pLDGmg1Tv5Pm95foMp9P3R5RG9i+JxV8I24U5DLdGtqjSI/+rGYP9jkP/zRukstJIUUj4H
xQfZBOYtTY01c9gCF3+s6nITFqdrsijMvdzA/2pVryZTlwuI9asgYMymR6XOVZF5m4gl66toMuwi
w5lNnNlkXavjhHmAVsaTGfyohib5PNMXiGPiDQkictE1+7QemFnTzCuhDzEUE6uMHdVYRBRUat57
EM//1uzeIE88dTrY//mAzUFMwsUX/ONbXWwe9Os1xuWVuVnOKWPHpIi6gx7qSfEp4HNLPuVuhy/E
dhBlrGb7Cba+tsIn9KUa+vnxb/CHkt1lEJchKvNIsx5DE19jxfAhbhrEL8dtwi9HIZYOf2cMArVk
w8B5pq0xVtKJbpST7p14i6yCQcRUU99YZpD+OA4z9SUFBs7wSdW5TddYDWBxjh5Rtqk7ICRtZ8Rf
JCe7eQn1gFujJ4PmSFriEks/BVrRoESDhXj7lsKX2zV3JJQT1ASHXrnG+Or9HHXA35Qiy64AXf1Y
pzhMl2+G5NGuyvIOFsEfOuM7BloXFl0AI9XK2UR3g26+xMMDZhGta8T8ilaJ41jWq30fJLraIfq8
H7qzC9eyPdroEpjUgh4Vx3RCOtQay1EKKPidOw4FHHIM8VAfhY53AmcHg/sIbzWw+oUJ3fcNUeaW
wCE0DsPalKJ2cBztPnShtWqu+B3w7EvbJtRlTeYVZvJovNWMeaZekp17zw0C1hw5JLq268Pplr9w
sgwriO2eK1F8NRjLoM1S6r8aF1GFnG6banhhk1QPLjOAs7NxcICslejHzzE6W17ng5z3rcxI7vBd
ZgBy52JFYiAcoyFb8RDyX2psAOuirrnXLq7CM1ocqiRNq2hLBbMh3DGDpbIMo+ljKLUCRHebonBZ
z3bAcQrV0G2UanVnxhGZAzgmzM7ULPMmtA8Ao9PjmlxHIO/9yzxT4QKtKa3vrDI1501Gsr911cM/
M8922Ysx2zbhZ5blzODmKnKoNrRIapc8zLQzrGD4AzdXJJM6lMHDjqqNsjhOt49OUDcCjA7SYJAR
lmE9evdMsiOIcV30F3yvRvDqspLMFzsEV1x4aNpmPzusKWnHk413EaI0Si5hLJXAvyi6K+XQtiph
XQ2BGynw9vmu8hbsQLg8wBl0JQvSbIH23insB/cPrOsmKZqSYiQ/q0DjWeRAO+7DdgpANlgNFZFq
czP8nFjh4wLPNAp5/BWpOzT7OVobm47ArGXZ8nImUEUvq269o7xZwkNPc9/LxGfZE5qTdUdxqans
rtqNo6x75dF6sFSC3lJHo7w6JOgPBL3mGNCz/vhri92+tJzSFFM5s+vEjCLXEPqUmG0r8vqwrReD
d2bxkcceeDsNaQUN2usPqbVow6doLlwAa6atzD2DUIBqkSTD/cDy/zvHUzJbXyLCDtRob+LoWY8U
45LaRHsteFSYWCnrS5b6h0HwIvXLkrrw1L8WFhhGGsmMeFnZ+drdauPCz2yI2K9/s2EGFngXnGtg
ZOX2hDwqeehCbP1MT7XoLmFTzJcnXJ0eZKP1/jXE5XYP+DaR+R3sIeVRacbGcgVERV070sYyhO+R
UUtnuNLwzPOvDFS2Lxtp+ZwYoYN1Gq2uAaXeHY9eeH2w92F0dK/gbf7Y3RieW3RxLZZz0/lymr1l
vf+gV410MdJPGu/1mVNRBCnXQrstm8ta+6jBHTjpdhJVPA1yE2QRyQ0rtQ2v5L1paA0vWvlDaC9p
VkyioqQYK7mv975ez8MJYCHW1XeyDyPLFFp4tssAwDHiPMbLdIVm55qBSznR4Z9F9eYr1Q1/XTr/
9sJQfPhqILlFe3wwpAAVEzNMKabcktBkrcHhUuYUJFLfxK+wngUQp9k14Igk0N8RhGeAeWOlbakv
PQpwinOWzGTSRI05elfveTJP9Nn96p+YUvLHaNtKlRQWzR/NcNoFOxB83bJZ+6ZLHO7qqOUpBOrT
KRr4aL2QRdTHsjb84I+linxaeAj54EV9fMP00SjIvqF9DslJNnsLpFBFDkvDhGVYPuw8md7YcfDZ
eK4ND6YzdI2GyMvrVGDYkUSdbL58CdA5i5VYRG7HH2vlwYWrXpe8XB7r0C6oc+z++EYptPOsk2P5
8WrJjH9QHtI4OjoIrLP58rO8/rPI0G8BmdkbL1YIauZz/OS4jhRkxuR2HoHIp+B/5cbQ3B5qElUT
zmjjzWvP1cLa6Yp7Woj1JVPT4nGW3M0rwypebqJXfIi7sZeFUEGzXJ0b97sp4JsVuet1fe0dauxM
bwsdcmX5aAm+aXt8EYaeN85dAYRWydflnWktInTrKnkRm/5H1XJuGY4JRaMWfCD2BHQY7PH7857i
Qhp4hH8chHXCFX4/+gXNhKTbSsDGoyxTdAr/h/UvcsvnnqgRfNjyzdTLexJ+iE8DhBawVbxlPDIi
GS5O/C1e8oQeM6thzLocnYKCKHaermDMvenaslXvWsc9TZyWeHY2Po5YmZD1U77jBqcFvsYg/ZZ6
xgRqmJDDcJhjOhHAOds5+Q/M0MQmOgH8ctIm18LwzsIkMJ+n/8PFfNECFj/xXYC9eQ85hWvcbM81
JCD/GOyWuFGNrjTGq7CjAqG9xeMtQNRNyhb9lXac5klfcGebwTfDopVCDYCPFW3Z9KTrf1hfg594
vjojknTL2i1Mg1OirJXyQ59W3PYd/v8XJ+Kppk5jhXjD0H3UE3S4r9Yjilz5RmtG6n9fcgKaLaex
s9U7AZMHRv+0O6lAwdkaEKsuCKMUzPRIdvb6CCEl/AOMvua8NS4DYK8j0nrnjrPiDC3mpFQxsNKp
vEBpWvGDY0d3kdHh3vKm9Hf4dqpZJ8IIbf7kYu/+vhlWimRGke5JT39yNjY7UujGgV07AiNe4Rwk
Kc0EIzNOtMDsa+KYgonriYRtfAeLFidkxCwvZOu5/c/YrUj3ohiXwWWRg+iAIMT9qfYzYg8V2PWj
SQwJ6tOEu03IsOXHCRltdZ2IpztpL8DWcGqZQMXbVkYaThg4Oir9WmWiN0ZMO/tH9li0xkkt0hiH
dMFYFcETnCkoX9yaKPvbM96cysd264SmAwekz4x0YsmWR16S9pC0mgaGX8h5bg0i39TD/2oaJLbo
ZUJt6HOdZ9s4+RcH8oRaaTzFWZAV3rAGfsq5g2UHFmmcq5ISQztAh0AQP2cGAPzeiygNGsaiAcjB
WB+CqVB9shEIySY6wix3nZEjxeUeuDk2zkvSCZMRqGpYt3sDZAXcXs/9e0D83SKtUqmGaorEVrm/
665Z+MgFgSf3oIrqkmTKa7Z9bwO74GLJR2k3o4MkMNgTrr2+ku6TbN0zjtEFuCbVKRKz10ab+Qra
dWcqOPemqtFcS4Fx/yKf4bI931nVwE/HMbj8U+UdvTKRbRPOTMH7sjyWfbN1iN2/kv4naXFCK4G8
YloKHi2f9MkRhF3grp4ZIlDj/3DTKqB7WgK+qU1KkiIFz9YyYEf+cKv1E+A7QoneINdpBl1fmp8E
ybDNVxpdaHRfT0BmRnRXvQKFks6YdGpMuycjsB05FNkSyszUtV4+wwivfycaWitrRV3+JkqCMaNG
GeyODWjbdwt8SiCeKjMu30ncS8+05S/tqzxuv9WNCzKuQiYOi2RoFOQVywwTSqgCyYJLST69u6lz
EXzMCDzucerVyiaXmynDd2C6TguV/w7eJ0E+7OgxIn2wlool7etD6yTk/r7Mv+ZlPfIxi5eXiMrM
/Ui3KUFaY0rrgeTk7OpNSnqTkA/jjpNTirjqnbgqpCkpPWFppkO2mi3mNWme/WNBVmuKwiYOol5Y
YKFSaUIu3lFhyoVXdQ5ZFRiMW58ecYVpsCSFkEDpHkZSUBYe9EP7aJXdEJxdu6pJE1/BO4w331O+
XNr5atOohoV0x3PEg1QG9Ww3h7VplUqg6jB7JPAgtonYIY6iCpnoSt0xmr5oOmSI3tFH5W6usseF
CS9kld/9eQAxaAYju3dVYQsJ6VQdwrZC0gFhEBl8kcSfnoj9Rvx83lTl5mxOLz5DvPcpI4UziElH
QAntqDaquY9ka+1S0fcMDHhMFVQdxkAEmILi4ZZV3W2LVhgFHtHmZQgRMSYvQpIeZ9D0ouhlLw/N
lJZSptt4cSJnHO1RBXQBC/C5ss0XXXCaUlcwDQD7AKnDnyeU63V3D7HzEm3ehg0oaVr+2fQ2clly
sh8hrz7EDK3a6v0GoeUarBeqTdm+J2logWXouPLWWl9Et5d+pHpVFvq27vJpme6kGSRqrGbpqC8M
rn5n+97dbJjezUaborQ2sA4AnCIUIDa7zT4XEEnoVy/ksALLkv6LqGlbX6DlIdoqI+1NICuX0sY1
94V6VmkgI9QKaqeHxZvfqkNOOMhNcuMJkzFCbyNXEU4hzFC2KRRsHQhg8CKl4bOBmTOQuudnvVmJ
24Ie7PTiqUVxooWKmaqu2r2+knA8eZL02cER83NXWT+BNZAJOLSruzY4K2xAKBCZ8li1pb5zpP2V
2mZ8yVv9LupXjOuul2LNskl76wf5SSTZwIISvgTyxAMRJBoYdI3gmaFxqp1BZ4GI0DZg56KEZDUY
FLZSQt/BGohFTdoi+ZP8kEixazqpcX2V9v7jJh/MVgBE2nMZp9nakYCjzYIO5dxtfn91Yk6M6KoZ
dFbQ+dKAe5ytYUw3wHzQdYh8mJlVe2yaW4whUn497LdIslR1Sp5YXUEnno5YriMQ+KGapaszO9GK
zegcW6xX7ZS2Y968osThS/OKY3qF0sG5o2Og0uhDMEDqqaFx0/R8fv7LdC74UOO7FCnLSdPAtHei
iR6DNe7wpGELx83iyc4Z2HYDI/WZ9WOzJO385TR8sLHi/57b0eovg5knHKM5o3oYDUDFlf0oARLp
SYHjpOPMpt+ZcZXI2mtDWkxhBKTBrXRWCC6SXPkyAcpMfezp0sJIk975w1EHn3QcIkjUAnL8a7w6
wbNcKlFDhiUljcJKQGkaiCCWJ8WgNxl4nDUFx/CeK1MJss0NSxd4lgmhDaSht7z1+n3fu//HOCw9
Ch43IccfPKlQxRZEjsLZI7aAswn4mjutfY7ocAzFdmoX94sDf2LpAjnVtNQU6VSA4co5U6hVTefj
zjuVtxHxxL+22Zv2aEbzDdxFNojNlQb+DjaQLHv4lHohZF0wkYVSJcxcOs8fj+VZVNHrH9LR1oma
PS/7Gicr/lCbAhOGmvlDyoC76UI/uuW08lcQQwXh7G4kdhyvCKcKdwYURX0Yq17j89xMSjPSNJ0q
XztM9kagx5BHA7XsL+X+bzOaj1JUb2weOh998uaWxCokjLfL3J6+PZiXM5JlpKmRGvRWq+RKm2MA
J1UaZsvV+PsJrU09dz69ndtOgme6CGbhb5nB2+ZaVU2Rqnv7/e/FcpQq6eI4QvNXYT+73Ui+A4PV
KqHeF6sqOJkCXPrgSm2X34yLrczR6s5T9YV4QeT0n/kLJgQYU/e7fvDafX3ovvx+v/lc63TLHMCN
T4a550My/dZXdWVMg7et2hZEkONyvXW6w32dfoxb3KpzRNGCfBJqMECGAv7ktiKfLuaXuY9kvGc+
GoMbAr++zZ2O7A0+34Tzyy2vhkiI6VUNbq5Z1Wy2UnCMA3AAz7aCJ76GmZZj6fh89TOtZtkW9uM2
C1KskRl8gkbMgFG6PKoJpdDup6XSUvrmT+kL9TJOg7K9u7JVqh7LITxB1MLLOagFhnfa1Ss/UVqi
d+Fue72njDOJZ7psKn+fyd0Q2wiVThZVxZqo5iFS7bUGhqjH5ruJ774r0YMLY+Gub1LHO7AIUID/
wMQuSAyaMpWymuzTNZWPSEIHdjQjXNlaQubpYVq0nH7QsDBjrJ1UHL4JvDXotyKDyPL8W6BNFLqJ
+YIcgm5m9iaaAloAETxiBYGhAQwk4tvN3nYzLFss0+m4Efh/mV9O//HrpgFhfFkROfwGaYukEn6b
kPfuC1JqZ0wsZF21K1788Vm/uM4yAtMk1lG/y4s0LS22j7VVsnAhhZX8+hCUGiXjbkiijGG/a4RQ
dXBPxJFcLOXcyXAH0okyLa+tesJG5DA4FwHYSymV3ChSmSAl2aX1GYlsCQ2HyBe/1DGGz6ww49b7
aSJUTCA+R5YI/vvZP56FaQJ521r4T9D6JFxKqoU+dKhvD+5X+zKLv9MPhfRkugX2EQM531pJwrUC
FCtgnCnca+A5l02B615JKzJio60SHPPaEW6fJnj9/AFZGiwOUubFvL5RK+v5aYtcBUu5An2iBDNP
RWNb5B7xaGW4prGDodjTwQFSWAbIqDw0QZzWPPuooTmGE1uyKASYbyVtf023uM/XUiwiMm9O9jsD
7GkvZZ7kgHrVCfwK2TntvWF0ODyboXFCS4BrOzkxzXPL88aXUaZHKVEdkZIsZ49aW9HCw3Pt3m4p
0p5vnsNoXIFF6QqcbUwyY7a2JJ2MueGNmvMAR/cRgcNc9Hv3Bp55KGx0tWBKrWQMRd0DHT64wupV
HR8MyoEhpW+u14ekpeGf93OzEnKttWavjrTXdXsbkUTHc9tXyc6U+KeN51Kf/rl7heQHSelC+seq
wcOfI4mQnhQAo08C4Vw1YVHRqL6vQyjQq5qKPWPkf+JYgY0lfczqbObSbHz7Yit7ZBEXTdMUmJPs
8wpdJ1SxYPbovFZqjyTe56rq9mtLEkgs5ScyeZF7vA/IMBEAztEcOo/calELkYskBJ2n6BqX2RqB
yISSLRipNsIHqKCG7ObTDnwSTTs3Ip/56U8Li0USfbiU7x+idjNY8ex1ncAEdh8P1pcjqBDOSlZE
Bf50QcnAy6l0180avHYndwWeP1G36u3X7MtfYJFUKDaOhgyocAs3AGnBSj74P16SLEtaILACzmL/
vOw6v2HqMUpGQDrX9GCYg+calax3NIffy9JNYEByDitX5fnwdImLQAKGlriHOAziMPBRLIl2gSm+
9cbJ31z+jirUaKlf6Boe4CQ+i+Yk0Q6mc+omUE06wzfHgu821Y4JAgsjVHA95ylFSrzwtyqJ4GXQ
0Iwbcl0brIqSw0LofOETsmPguyh1bQhOqJfaqW9jkZRad+5ZIzHjqFmDjO2vDHL2DweF3dARdSEi
uTwZ+L1ZGB/44eXwzpcjAjswSlyf/dVfR5X1EmtzBo5fmg7scSssN9KTrKiVooTFnjkBuXq7Mix2
nnfrPUMkZ/Az5NSfIApyIvtJ1/asgDCP5XYfO6q+cm1a4/dNNRQ4MPrpabaXecNt8e1MbVkHMRjn
BoYv82/qfJTrmICyygzBH1ra2SYxmd6DNwgMPrh15oHFG7AwanEe19rjrt09G6o2fj4Cj/IZWiTD
7igvnBdaBln0uHvL1RrFv/ZS6NhZZ3myanjLUxvPsa8UTcZvR/a6dWs+RwmxQiBFyxzGuJYkIuHT
Z0Be/aqxshGC/1qqCoMjbItpQaaeRPEZ57S37Y1Un1blJ5XX2T3vHhPB+j76rvFggHw6yNTJpdf1
fGXMA37mEi44EMWda+smK3nEXaYK1bNPB/aTlIgjOZuZrhzdpvphEUljvVWpZHopxSadXmZHKGdz
LGWj9SNgGmikGrurRxh/tHWkPy+92LbjHewM9L3Ptj8n6uwMfoWOgIdBw9l3T7uYzuJemMI5ecBj
n/zkQTKOumYeKvIcaaNQTtRQ/lAE2iwz5RVnZlZTxfwNAXfG+csl0LT5O1iXD1xlYKj2ku6z08r9
X0npUmMoh3zXa+GgdAbEngHVsqnx0XRzLew6N74oNNL1Z8RaFPBzqRIGo95UPEtxAC/VMOA18dkQ
Zh5jwsgOf8b4oDhh/io5o1enHAqcS4MOihatwLzEGNetH7PUV4oQtg57l4HnX1SedTZgsRBlQBX2
DEcIEG4oFhjbYcfJVvR8zEGT0c+HfhoBuQTO6D8OnjNR+lwCL1p6ao0Js+MW4LDubrR3+cCwbeOl
g0dkulpBcTITG/kvQkDYcsDiaWFTtMhHCdK5iU26NUzudpzdzsflqGhxzVp+oeNza32rz3bjUOnV
D0HPoDHEJmE8zPEOQlAqxV07CKakbBoZh+RqZ6bvfC4odlliH1JBojiJMFsavCiRvoUVX2gyGwXI
nwotYMVpACGHBb1VaeUj8IdHEUNdopYXQtOXyQXumZO9hS0JwMVqEO4I8N+EdQCGEHmWQH21p/FV
UiSyg5wbNr+TajSrvWzpZBWuRaVButF5OQF5suaHuV+isOOSQiK1Jq4eMO8OmQbSHOS1tJ/Svzhf
h1zwAZTltZn8Pj2afBd0w8sfqFfn4PgNW5j4PIPyOiHd1l1Tht+b98fPTHY/z2uYjCuismcFWuyF
LdZ3fuV83m8IPg/jY+7A9Yy30ywHIUbyLMTC6EEfnIa6toizlQGziLzhr2FPpopYOeNqNcWm0w8N
6jpszjPfI5UJ/vQWa8XE9gNjOYeFucV+0syv+Lx5avgEJ6ARGoKwe/ebPzmqZ3/TAUkL3PcgbsI5
KSzXJ4/9HIhm9i8im/MtBhgfWtr5BZh5vnU/lw6np00WaNTY37CWSCAeyOQ6hkZY/9heQK4jadZU
ph3mArVNsA6T1u1Gq5mn+QZX19ZMiuY7voaJ9GZkggwlZ9ftn923l3MbbuGrEuRCAlUowButyOyG
98mIy+WeC6/AV9oXPgsFd/NX+Cew8mpQWKo38o47NzLgweqee9aUjDjV9h+c4ZfPuGp6u2JGjX/k
RLVLne+K0ofPHkGukkBY01TDfEuiR/HulqU6zl31MChcIUHrCN28lAbVk24gUATHsCIHXTjAUZhz
PmLZOI25kjscWy2KpByH1RMooO/Fj8Xfpo7xEkgfST/gVRjSiO5z6VSGq5Y8RQA7YMYGWQkRFOo7
IZ9vtuZCUUHqPLdEMkOyUMVl6y4VtQdZWky1qJcIjVf9Y5vKbCn4e+B96AoN86mWKVC1MKdClSiw
IxRKl+HxxNEtBPr0FVzaB/jGLZfV+9kai5QaAyzXt2Uk7a6r2ZY7ByAxfsBKM5HSJqcGPoKKaBRK
EfjgLpSb9O1uwuDRYt5RijhvbpZhlNTkvAMHUB4HfK5/n90nK4Umya7x3tJJ1yEgKItEh+ts+due
RQ3ZOjwI1gdIgArRThNq2LfO6QfL3/2SRXdn7pogrSAqsEhi81CXcTZrs19xvamk6WM956oyvmhW
5EFh+F2LPCutqIAPWEn6IkS6dI2jiS4OalLRhuhtrUZwFxC2qbu+m8IkCFQyhTL3QvTZjzgc+0X6
orE6XawPcwlus5VusSNyknq9OWxhZqk+bbQVt5hmKLhXIYp5vNRqm2qfhikZchnxkACAOaJIHBWv
1M6GZGHTGTJld/mBNAOkeAWh5SoVA3qMFjjYoCvqaosbMbR8vuYzkZW18tJeUOrfdANnzWZB+Cp5
ksGp1B8oYpxNRjcWQ3zXqMIcbUwZrFG0pUdnOLdKWmkD6S09yFMjB85xcd84zm9DGKcvPri81IP7
UC7OvjiDRehBaO4h4CMR5m/NrXqJ+POD2G45/FUv7901MYHLNbUpU2jtEYHMXzTI+Z+M/mbejILS
c4MLh8rcSCM7Pivu1TluYV9IHQ2yfwD1nshf7qlTZqNG8BZDA0nNnaxQdbKf0HzTgnK1u8J812n1
OJ/pQCI3LhrXBCda615Arv3k+712y5HTZmhKW1iMPbBiUcO7y2GdQHujHINS1p+1Svt6DZw2fBSk
T0Ot3MWTseq52IATMa+KP/stUuBhAPxbFDGBcJ+OSulxAp3F+iV9j/tfXQmxNB7x4uVfs19McCNK
uqlRrH8UnsPVmGHx/LQCkJTPuLOr1WP/GhIw9DoVQbCP1zniXgPc0qQG4IdKkI98hN5sEXPMUZWG
OgAMpM3vthXeFbSEnTBhY5kD4bpmUeZ4xcKbneOJe0TWc6PAhjZZ6sDOFsUSq74b/1knYM3V6djp
sdgXbB/xv/15pNcxnCCxrzwYy0tHo/qN3Pj5VrcZhjGchqJJpmhniwrLUXB/OEeKiVUGavFrWf4P
TKoPNiaR6h8LvHe2OHwRFqf+mivGV0OFMz0gNru2h4IBQXhEfU/uV7LtE4pklMWHtA5iXr1pI20h
QIDUFkRLgkDUKIwwcwpoB23/t110Sd8iykN+9nXSTIVO+9QbjFXPukX57bgg7xS4WB/6nqr4D3mh
FNvSJLYmLlndQdo37Tx09PHKTYt9bmp4LiwfZXrIhWh9nRTTycPeGOKQBvmx+OLgJJqQYpTpF8Bp
MSRnFNO7Sn+PIg7K8z/Jm6IFKeE54obu3h8zFEDMD9YdgxAYGLKgLYY2nJk7vac6+my4zK845qLA
sNUEMh8f11rl5OYno77wZ31yZ651/BLZ/Gqsz6xWhs/415URp+0fdZqLSNgzHujV6T2Za2N/Bj1d
HzEOnKiKGEFOQk0DO1LgaiA3xPIuGH31nqyweK/8Mi1A/99wNCrCZGjc4oGygyfUfKeVUy9S8028
HPfhM0my+AUd1S/iPetZMG4nnm3Ah93s60S7Ob1yPYIfXixTGmGawMhV7QJL7MvaxXpto7MQmCoU
SXIrEJVzfyFG1CgzXXRN6q2u60dJLyk1/D7Y6I+sgwUzbnHTQFd1cVWDGk3mjONZoN/TQBsxDyot
/NeLWj2njvvU1SoWDKtP6ZBwrO/2kyhxLLKw4KzLQO3rNqSSTxQkSJuNUuNfUgNwP8IwBVZu9AZa
YGEi0I3xGRzBdAs54AGNFvKXhWJQCDkQR9w6+Idi0u/ZCwVyvKPQ47YjsKk3kpCrfjUzsOoLgAfZ
g3Wsh1e1ak1tOJn8FDSehxDS7FzEzwpoBgj5Bma1t80UZtQ7tHLfFn32wphfxdROr5d8p7oSJamN
2Fx7bZS+XaGUNMOJDyMdqrJJNeSBlhXpScdNaNycfcFcm4ne9Z5RtdNhvrBZ2adxLBz2WBU4Bu8M
IymEK8hDcG1MQPOjb+yhlSZXBLPgH5CiUC5xNhDVi9eelkJ1LaP+DqXC1S5JG/yE8RmJgga5uMH0
lKbud797AE2EduWCetilB+KoJHTV02Tqggdn9t0bbRveshgcfalotjulPvbdtJrUNweDMGzJtDHM
t8aorSAsL2pag6vZaF60UuMa+uFAmwxARlaFyAs8nsMSzFpk6SxQskfRex9sjTqDJad2otjF1UIb
t1kTT5Tal3rCONIyF7JVMFIUNj3P8iYy0VyloyblqiXVZ3dWuuSeZYtjroIFggeDO3+77zFjvrIB
YY0HMq9q3Mv1KnvAqUGEhPWmB3psqU0ObMzBxdNWUR0HqzgRhsCGbTYgtgoXvvGub6dfnsIki1Ty
OmAIkktfv/+YCqwn62EtwmZKMta090ov/PYeU7oRzPVuMX103Ijx7O9hZQ8WHiRf4p42r39pqxWa
Qv14EiczYHi6nNIhsnNM9Is1th2FCOEHyjVHjOJzNn09Ph2m7l/z/o0taKIFwxqqHf7LAvkgn6OA
GHeDdnIeC0hETOBJU63zjL66c6IkxSYDj6mimFbknF3gk/IDUyZ2xhKGQ1eOg4Z6RhtCVjDglIeF
VL3KCiy1gqu2HZo9zI4JgwsFB6noNxbC5pCkJZqvQLFTZaaTJIQQX/C7w5A48DZytAIRyR+dpg5g
MnCKn1aTec959aDh4arDXQKodx+L+t+YZw9zUXbkTLdjqH457mzDBY3adVbdrptajgDUkQ9z4Pt0
kFMSqQS85fIi8ubmLoCt3DwbpxSmQYEw/wtnWeIZnuy0e96QjubKV1NesOuykuBZXb/uOVW3x00Z
fuo9xH2Juw8B0jAgbDIcPTLmCKbSJ55WjY5NQeaI40SL9xEELtz/aIZhX0uvFrrWeMk5YSF77kJi
Y4zhTmTLdMkCM708QKwJK8iKKW5AIURl881BIR0Ngyj8W0WNPb1xf1DlrByyMF8Yt0OdHEJGrEtU
joDvLpuelNVelD8uBZzcASrSxPT13odHfXBXGfaIb0U8NW7rKJOx++5n58DgHj2JKP15mdfkVxxb
SnMF+SRaG2XzRPdj1o1v6pSfaY0U2v8ciXCjse+QmPjb8+KcTy8ftfeaTgT8aSVObt3+7/LQjb8W
+Ay4Yl1Q16iQxJ01Eb7jD7NBzVfLxcG8uvsJdMhLzUGcTYOJt3oqXJ0vyifQFdORHJBQuagDUZ9R
rrwrLX1e2ZgF1f0imVD/HLi/6wRiIhU/SyKyu9tJxzo08awKD162DlvH6Kpo3713Klh1oX9nmZIg
Jhg8NS7ucBYRxKKROYqVuELLnW//l+e2eeMOib/5TPKlw+y+2JBS/2aU4TOxsjcGyC2/sqzrPhWN
jPQLSb0flwZlKMLa+KElDy2ndzYdI/qHOIVqPJ0khWS1tShH8ocy8whaGbcn5tTTf7sBDIIFXksl
dKeVgh0t8/msZam3sCGZDARU6W/UZuNTgOEjIaqEr82wL00SDbvJNUSKe5cvPeQN2fpJdJR532TX
DbzBpA1cDbpOTIfoDubGZ1xaXOnENwrSeubEWlqJexvaSwgnDhvDZf7piR4VdAImdCqx2ZCp08ih
X8A8vQ76ANGPNY2aIkInFCwuK6uMvUmL8GPo7eNtdAMN8+A5S+qhmvl0CpVPueJ4ddVH8I7lg4SJ
+gTpNk6rk+0aQte9fns8CQjXYT9XqEw7/DHobk6e0VHjdiG9QYmC/bMEnZkFbPhJgP1Yr8bLW3zC
DXhhPP7jE19hmlGmgp2LaTUGDzrW8MsZeP13BRXCN6E+1mOT4qI4/3JZMYRru+ovOhnQNO0uP8on
2AgUrYKQIZEgYe95z/7Rk+VUQ2Q6FQt4D0JVGmSgCplsVBmcDLx3r23YeYUab9oSzEUoKYrSD4xx
5GfuxfsvBx8ZnAbv+6FtN2RfjwtCABHVHx1rIzA7ZDt3DtwCIEf+tP3wyhS/PVL7yVZ+gumIJxsq
so4QHD3mnRkNjHjQ0+aE93vvxvDGVe9HTflmRJI8sJah9RyKT3w2MR30K+u3MOEHOteqLH6ZXZ6H
e1/GdFXwghslJXRIkK2MKz/vLC8PIgnz9geSwiyBL9AZ6ggMM188eOBA61Dloo0uFSdkpOl+uso9
pHEBJsxHqc/B+NC4RWqG372Dg5gnZ+RFy97jtaOmMdXwhr1H7bLbewd93pb12YuTfFvwdcbuV6/Y
Q0PqBKCjyfuUwnJUdXvRrLF5HlFJqAPQxoSwS31YWCy8Fhv3VXGPsynVu7+Dmap8z3S45WNbiP+h
znkMLcZVYcHWiPYZIV7/hakVKe1avBL8/4XYJbyMTUoEglKxzEE1XK4Ojhh0Jb0HcVZBLOefaJDM
Htdqpt4UhHBXyJicDKmfTnCv+75N75tg//HRl4DHdE+X8ac0DM6NTDzU0tJKmbasEtWtRB8tHato
GxedUHd2qKB1BwbFjKKadaEjGJPGb8fYdQSz8AFnMCV0bZS7WB9NA1LLIRr536FDa5nJwR0UP5dn
2YqDt7bslPNgbTNrlxV4s7sviYuZIMIxU7efahKKD0H2RwVAe3wLDRp3aVOczY9h1BHH3qt8uJ3u
oAGulPI3AOmqojBrz0MqQXktPjPUfY0dmp8UQUGAfXAmwwwn5T/Uf82c8t2vXXkU2dwl+t1sZPpB
kZpH9B1jcw0barUvI0kMREWmLP2pb1eRe5rLR6WPumDD8gWc+OyWQY6l52oRY61GrKbQuAzMJdPs
PWgzqz8Ihshl3OS38uSdMM7fsaiQYHa1+OLLPftihJVEZREK2NAoEoQoFvBSUeNWQqV5jr1ArGS2
m1nNY3BqrE6BjRXmiggBkySwObN1LDmHo0viiUkMFjUqfA9LetmSgB0c+7FG5skfB+bMypqoYzoq
N7ERnQY1ldsO+MV4G9SsNOWUJruoWB4kei7Bw7+G08Cvt4GN5q3hXUGwfETz2sAsA72D3XHY3pSf
hMEagMO46Wck+vxxKy89yTVE0yaietI3uzbY6ax/9+DEYTFEwpx0Er2/wSXYKK5U+E/Z9KJSPTnx
pQqB7uVUY3QryK+/LWu1G8pBKIX3WKh9HiWpQ4LsKmurjSWRl9ODCaobPIdDMpVbzSWVn7v1HZCl
yCxB9RyxLKiQWWI34CjQqOl7d+mlLT5f1DSIyQ8VFqhaTpRhzLh4+hvwS8QheabD45QsWSJ8aJg3
D7CAeZy4Jcfl622jaDgTQx40Dxnm77udlauTI3SV49skj/NdIql/RHOn1qogpcduowQ7ExFBnZpV
p5PnCfdSQkT2KK+oQqJkVfmj1+1thx5SKUPPbwrNADq6bB+ra5J5qZU6l17opjI4P5y02Eb4ejv5
e5szlhqWxkFDcqi9gU+Qq941Y8WVoKPnx7VCGQNqAdiUp548CWjKzAtfqSdCmFqJgRffh8vMHU7F
LJuVKAUH1SBso6eXMg6q8jnEI6Uo3yJycnY2CnvvC5GNWWlMMcA76VPSXsgy7NpL6HaDwMe+yIjP
B+OCLw32JKsZbV0VZ4WLp/JhsLpXDKGJCvOy39FvNtRz1DT5429SMKzI2r7M4fdgaSOKziZAWxFT
KI0IM8YBs5LkZxzjN/D5g3JvKO206gFs6kZhoLbjTkVokHmREa7+Y6rzm8M+vnnsBrbR26WZseAZ
WAsX8Nv4eJjnK8rYP4a6oMj8MOsRAGpcmkPcz22MGFhdmexkhN2ZXyc40sO/4lKBZRmsd8zEjirA
qMcNjbayF2c6PyEyRfpqx+OSjn/feO9ufKcMnkugw76kGsmhamJoTmiwk0veotBCTtFBQNO3SmMp
5ncGW7QNXp+ZnEC1Gh6jM9+ri80lpXLl9g4AnV4x/X608zBu6sdqHof3w5wTMY/Vd26JLXLWjEn7
yyE54KI6xIEyzBr6gDxTK8RgA0nXUKfHye1BHiRbYp3W4eWGtTWyXkBUdvq+cx25v5bwmOjRIohO
VxKRJ0Xvu8YZGzn2aGXInYAQvX+6riAYL/pMqGztZoZTn4SKtLfHS3IRd3q8xvwzCExw7CJyvU5I
V9ORqonGkll9iREW3s12ew1MjbHB74p8wx+naHBbyayyfrkc3rln9p/LFHIyjnllFI1PviN+cTfE
T+qWggMlBS58OFpEoGpx3pBHRPX3eY7d1ewaLk8GPHp2uhhkcS+y+l9j0pPaD2ZMW1TSNZP2ZSBg
Fl0Hm6od9B5mU4wJt1zJbXayDq/ceM4mEE4rHAbrMLFtg0Duito7yrgHiTXKu9OIH0I2rBT67Q8m
kPNhbBhiyUYcrooHXIj1QxUrdTL6+N9tPR1B1XiW16w7BYrjNRkETOhyE6MU+qLXR1Td+DSARye+
XA5seOsR/HGD6jDUQ3hpJIsQAJXevohpNh1GNwzZq4X5QuNVy5iBxNbFMxBoWcwf5VTyWtuWOwvl
oOU7jkr4VMChziG9bMoY/I4zgz//zj9B3mM+Y2x11ydAvMN+Ya8XzR7xvjIrLMQy7lvQeMvjsHxL
52c6XKlUhPaZ9Mal96gYSDVgD/Z46t4JHjsMrpt7pD/VtcvUrei0ZUG3Pe7X2pKQgvcSzB892xfB
EY5y+lV1IArAyaWGK94vEa4/VNkdzjrEYE1sOE+o8xh7Cg1QJuCHEbUVN5TAnxkxUJsMX24/Bc3V
F6i2wxF1rAvvvBFOkjsV3dP6wMazW+gIlV976VAn/YlBMFzhcxFEOzDTdbklDJ3I4cA0nb6p7YxF
mknv0abpBWFshSsS/GFKFo3ywQoEME1vysilprC/gh+uyTJ7VbGZHmcKPE+xNKHjuDUynLEt23Bh
axOlRA7DAQyxxLadxZNq9AJUL940t0oI9WBmpSR8FyileHB9QqHiYCZc9A67FRS2TxfR0Mkw8FDH
7VEUvcuSVDPiohLVSzvgnKpkX2htGgE1zAECWkXjPQQ0o/iF8dcUwxiiz92d50wUygw06Y164TFV
/AKOp1Mqw/8gY1uzElEzYYvyhsYM//pAIkhrZcH95JQhZs8jiumn7cJoN5EpH6SvH/9FbfSPO0BK
u4UUFdXrjXpCvTfFQtv214ZMkBME+ebXX1dIwZJL3B6sesmZVFpN9HGLGH7gFBB03CMWVKceNYoJ
8Q8yugf537GD9FRXzaNBJ2QKGIpBm/q9DToY18DlN1NillsLg8LyY9baLwU+XFTt655vIH4cYFFT
u8R6oLmMY9MGIp72V5d8M5Z6BpdaeCdzeAXwBJklNSt/wj7lXW5yJ7nOyGDnWjLhWu5YXz/aXFvC
iSeG/4+3CjjsbMIWlMGzBVSMAmfmT+oi5rskOpAEeKhT9nBxuHa1e4JpDmAsxhfCdpt6x1z9EnkJ
cBPlzJL1XQ6ONuzoE48rG25wH4Ysv4if5DkHvBY6auNU9VhrPJHUK0k3BvLVHwG4vKKTIOCiii1r
foOoyvL1cRHX9miowfkFHvuw74DuS6x+TK3fxPmin80o6E5xw56KMi+zLFdj+hLYEHjaJtk8dTrx
FhfzxXvvVPQrgFk1gUEvMVRFe98628oDV6nmpaSgFVynxt8FRoxHX5l1Un+iS2DNvmtmO1ZYkBms
oxKAnU1VwuNGDx6F7BNBtYOO0PEYwqOvLKXiJagqnso03zGCzQjcW13Sq8g+68+PeJsXqoXBmp9U
N/XBgZPFrpH67UBKQ0Got52rD7f7ivE7RZEBzEsLpWzASCO3epVQSXtg2nqRiuvEpBWSHm7ndwej
zxg3Fs2YndP5jABZaaXPKSamcl8wXbnriDVuukVRFkdCUPzKKs3M3DTOLEx6xed90ltYZFKZ52II
kOnZSV+z5CiW06eYumKF9M9n8wRcKOZklrFQREbJO421lvMS2cJx1RHHfJ4Qgsh8dP7czOeF21oE
Tzg2/ccwyHMG3Qr9xaY1wcD9B6QAcyiuI7QE8XnASKoNouui3fsWaphOx9Zw8bp1Mdndx6rWjeJW
TiXPC6TF68vAFBBDLqDLxMQoM0y36b6cgtvuYxYVZNKzNTkauc+vAWmLtfqgMr6CN/ZleFbSAsT0
NTro3q/5tO4+TeI+dv7FgS4F4suBFOUFyZCdFIk1RffkLW1s5wx+H+6c4nAwK6jgSlOPvXjkuSLY
6CGU0BiLda6v30pMuIG6DRYiSYUetuw2QWtRxDFHbx9/Lhw7gLM7GdwbyG3cbff8l5mLFJ3sLhXL
YZqgwdUoPFg50mW4JaqevxNTSNSi7Jfkk/4qNEbZXEStwUswU3km2rbOTDOxPnG+3ZqdK+zoyRwR
A3iiMFB/S6ulgmyH3zbcgHn1VkmougTD8VQ4EuEbW0X68X0AxeBa+mqHdwlmnDBffSvHUWuub8KC
S2z5gFePgU2fw0QhghIDyMCuHny8ZJ+xW7Nc5MWFDFmOVXM0stCZxh50ROJ9OvwCjfGVHwOdtVye
0N/UuM8yqo5BSDs7Pv1LDWvymiEsMrUeUwl53vgBMWZhK1gmZ5QA9VBaAw9wN/ZafpimpAmuZYz5
tsgmS7wqvkUN0Ez/VslemJmwg3miPzxRTraEXXUyYo9e3C/k7VFvokQkXtVYgpgtTONArNkiW44C
+Gyu2AvygD672lKpcXsMV3uV/f3adpYzowwDsVMQy/yyTtGXD4iCgJ8zd3/r+cLE5IUa9/5CWpeD
5Cao3JZKNGhRAyQjUxwZvXFgd7wPi+DI1o12Q5ffTQ0iYNrsv97tqqGkMuyS23pkDaGj2Zths3UN
btacNK+fHZCnhLTK52We6hvNNfquZVvHWkxuIX6Af4thu0WgoZUWfA8sB9ev5+lwYfxxGJdVbau3
QP0zAE02DRYoSuo5emj1alyZlK+YjRPT07sKfA3att5SP1FcsOnppC5Fzb6g5HhPhptID9J8CwMI
AMr6IlYZoWPqROg4pFEdqrTEprC8S3kKpA8k40/Cehm1mZqQk4JdwT0i9DrdDvF2vkKCigeV4RKL
jWdjkLTRFf5P9ZbbW6Q4MK/Zd5tI7Qhj1vIfd7u1hNUW3RD+J8JkBWXqZ+NmhI3pZa0RIWTyDGlG
fQmFv2ZvP+m/+AODTOK7hv8IwR4H/O6P4VsDIBRtV9lw+GkiB/56gQ26r0CGiNCbPe97Le6eE/+I
SBuahvkaBX7fE2hXB7O/pzHrFQT/8p/7XjS7gNyyA/5Fr5+F8HMsBg1c7/ReVfg7EnTTOY5qkY1Y
PRJObRJ5MUagOtqNv+iTVMlagrwQz3w+u4G6D+Rc0vv2+/YUuV8+s2acTV9bXQxiHrRNkmtkKFmJ
y0IhGAItwz/8THJA0pYBL4hAnxYV9Zc1CPiEwRE9soSmnt+xV3MY08LA0+uuxp0q8i11V6GHFyjm
fVb+EjMuGeadfEn3gOu6m5ya6tkhxqIsfTXHNVNcdouj3krk7teDLKxhkxnEHeA9ILS99Vz/02aK
UceO0vjJNvf4Rc/DpKa74dxDCMoZjik96KV1uMZISeLVH4UP5OBmG/RAQMsfrvaXuI5EOfM89+HM
cLma6c7cY64WYbn43X6Q2sPOXJPit4EPXUrSa0hbbfZ0wu+WgJprvCrWBYImX5UU4IL8h5RgpFE1
FkL8Vu85Ty2XMh5bIK8INEOXob7kiPscdwN3KSozLauggn4nfQWU2LM87bka5uGR7szX9MKwUymB
9yIv6N77oDTA4pWcPzUJ6utVunzyOY2HJ/tGTKPcmlHfj+HC6t2Afokb6dvwhxJmtADLn/cFplv7
vjrRcnjjV2LkaYIxoMkSlP6kqh4A7JZlS9Qq21lfza0+RxTeybSFpW5ZqcEk3f/6zno35DOz4xcx
DYqz53b5zfB8qSrHasMgYNBlhzREzSlz9o3RLhiaw23XYYnodSdlUr18OLS5jm+7Q3P7SBKYRqdj
19lKVwwcnAXqnxtva5hsptDF+GyIpQoLCD0kMB41Pzk+MGaQId7LoYwAjsjGFWVMz3HNN4fs7lOP
sY3FolmD8FNWMXERdRljDIyYl+nFR5XiivT3LM7oe//An5y02ZD5yDqyylAqhQ7Y983kS3DArTFJ
RxBhZFJzZspl/M68zxvZEE6O/WRkGBvmJgUATJ3/GW166cwGJq8BlhFbNan0TZ4GlVulte+lL0Nd
338ithGcuRy/3zfuaEBnqKbS3VQZtDD5wFG02mIyn2Mg6dBgEYBVfsyvO3jfyW1zNgUwQdz8uwWZ
bmfmzFOVSr2538AfkQPEFu39q0iHhH/FNWva/v2lw5ere4qmqLkgiZRXKp73cCj24ygQH9E9m1p4
EJS5Ls4OC9PHr/EuY+YFScExTVroI4DiiQfCgnkF6YMeMT1yLXTOhReZWH2JQly2o+3q+gTK/cvV
m+OCcbH04aBNkeXUMgjh/W40cduXO/10DSDR0Vzr/q6s7jqGquWYjmOBnOeQzUmmrvTD2IMJ/GLa
wgDgWasYndpEMW6/UAX0qGtnnHD6NuGFH5WkOeBTcvHRwqzA8/fd8YlqaAkgKzmgbTGVN3M/GMWx
BvKSwvHSrSyWQlee7WGtkbL3bcTRwKTY1WnKIY3KZZqp058jOh2qvPG8FkOlN1Szt4Q/KHhhbiUd
zgLmJB3IFEMP2vd0pQp2tT37GBlQHya5XDBKHIgfuULwTUdEBiybJW626hj0OdKdvWUPwnVuF7bw
iPDHFTqf0xmNdaDKMRHjy2hXVB+P5VXcOI7ROIzI/YaU/nqjDcvcT96E+Ki8vKJOjnSlfG4+bz6G
VIhRcmVBt+kVhDZE8F1Cw1I79mpSR4TLTYvVriujBBuN5cKBorgynEFGw3b+yLLpeeEKEgx6DMhr
3oeJ1DLDEhsEEZpwSdXOtKh9wShpBSkXe5dKY+U2ej6m2boA5lLrDmyhcnDtZxBuaUcqJGdFknwP
9bn8Wz6aTOeBFISmMh3oSkFqZ1yIgvLGHObNJwCGFqsBD5b+mChrLMOgBqpTuQJqJGXT/19Qj/Fp
OkZtERBTh/AdGqPhwFyrmFvptrpgrzEcrBrthmVCyxAkB3JmmzhdAyNR1jEVXCePyAZScewcdDGF
qcVfNqq10uDucM95dEGdSaIYf0ul595bU1lz1ka3nEfswXPzat9ZAPqIfiFOEAqn3sZpAYmRgdW/
zXYWu13GHkNTb96KCrey+R5Hh/JBCM6u7sXQCLEycsatdQJSZTY4tTwBR5usOKWFc2Lj1iwTTuiO
8P88bKlvURCG9ab6MYPwi3C4PncdtKCu7W/eLwhYutWJEd7N8gZYPGH7N+Aitrw/JD0uMKfUTBq8
YVyX/z8tgTpJlX7PjavDBSBv3qcYWRSdlN7RrRvh++cMTuirXC7DIgtzHIOvoDxinrA7rJ8/qj9q
RoC5Sqru7uMWzw68pJ07iWzmHppW5QBJDRE1GURB+Ciam6cJspUGjbrek8s5SNsADN7A9R3sjHBu
DV0DCtA2m/hCZj2wYdwCr6L/l4UvwvVSqKGJfpXKcioBUIUR3tnE0kPFJqxrwLr3Uqv0alpIys/z
DKqqbHeh5ThRDKpAo2GCAwGbOWtHihERpYowwmKBfKoddjW9gnub16L+Y01XwZ+Ol8G387dlH09G
FUeaN/SBSM2l9FZw9/kqTvBpFX1Z8NXi2X+UzA3chkd5mEQZ+TyfJyzIJgaE7UIl8JYByOfkvuaX
AV1WdjgfJrU6X/IlChdYX/htGufTBP6bjGmQbDFFeTPrQkvaIB4P78JYmzAQbO0Q02Rhd/OhaEO1
3flT4Y8w4c7Q6WZ4IOSDrpeFMb4x6cNgjc3WwAdrdXEUKsbwx11Z98MH+1rwySMjLpRVMAH50cSo
3pbJ0zCU96QWHHaJfvN4tzGGJhCU3fweCFGYP3A+WGCe9jQVJ/PBRM4qyocxTjTi5XqA3QK2WyZi
qPxNhghyRJzeNbbGrPgutzFrLCoSnnMNYmTj5DLxUSrnWcC7ODT5L/NExjsBxpUq1j8YJigQf9x+
Np+AAVuRDbh0Qoh/qssQI986P5g8GBVdXXdYLO8OyrPAUHs/p0EhnVfGc5QTLhsH4A+AIOEXtkO1
kzTgm9lXxOUxRUHiwq9yDOHTGLv3JMhcAHVLzfFPUo45RmH2le3iWtJeqqmYhaGCUxV9NsyFkbzF
Rk81UlpuIwuFp4QrDmE1iIcaUXCYTy6OvzxSczx8m9Xye6hC/E5GJtuSpzj4u4jH4OSWPt/jYzhk
KhbrkMj76OmZHkaaB40cC9KWnu/AZsQ67aJBlu8t96/dIWAJ50ALvVJBRlTPiDkREmQU3T1A4Iow
/5coHCdYcfK4BKgd5f+3xtpT3la24QDMkXZk3usAKxoNhU8PEdy11b5CZBn3UnP+8OR3cBp3sQjj
Ngt0/xt255c9TA9iFGtgbW0h4sjfIs6oCOZJmCV0sEr3Trb2k+KlbWCIlhwXmFVkrwtHQr7iL40O
TgwsIa7IIUk59G7X0uYB8oFUAUasyHDrOc6VcVa8Nvr8aY73QqJntjj/dk1jt6UZkutFUh3Z2pCI
F5gcI8FxV/6EdNVXbKz8lER7Sliy2oPx+A8aGVF855RFTfTTzxRsAzTIAn/ghAj6z0Za+hlmzXVr
Jm9S0yzGDOghdSJxAf5MULxFZpuEOi/RvwNeGtojUDypr0xrjPBO0ZF/VuFH16HqC3RlbaCPYFWU
RUximrXm/Lc9w8pTzA9BE9Ld5+kCsnHs4rO32t5PKckyhvIS7t1TPoZNRMw24lGEZLmkREOCFuFa
2SfMgTBxTYmChLhkprdeG8wFNaFguWwQefSo+MrvmOFa3dg19o/38ynsqwGU0eOR43nDlFgSpLvY
IeLY2Awq4Dd7j6U+dvcSCJ5ULEA3bA8eT+4AOOqOP8xbFsCK8JvmT0L2mGfb15fYV9NJ4+rq+zwZ
47KNsKRqWFwg2FHGn+YruSYcy6Pk09KgTd1nSAs1tURpN72TtNf99dwvutzDPPmFMfP+5JKubJ/o
xKuy1Q2qc93D52wrrtN96KF3AHPrNT1LWOksoKnyyvkgCAp1OEhYdH6uScRKGGwEeGkMPq+1Ysbb
q6C9Lq6fI6951DkkkXV8+P38YA8WjUUwzMoOAHCenCBLlPRkjD4GOOFr4aNLca/nLjrSmwuKHekW
MLKsf9r5Of6VLuDvGtL8mRXezbs/qHch2IHnx1ed1/b9IdizsX9G2qvAiVF9eUjXwecnw+XMZK3y
ID2FtLWW0aY1bFxHAxZjA+bgGkUkcnd324pGi4kuBRShnwzSjtThqCwlqFnmj7nePAm3gD7eldUA
jTJpgx2tO3EZR2mdxRER6nJUnzHofP3h+Boz0yfg2j48e/gEy8TCkaXtO6FR4TzSrK7SJxsqy+Qc
NIdj3ROLJ6I7L8/R5ixGbGQDxs618FEXaUjy+vyCyPiX0DIY8aLDrLTCtGEhn8MQqBnzOf/BeG5U
pz8QldPXh0hK1He0Rx3k8UwwfEpKWUnA9ACDm0MXee4Cl+7AxF2RfFL6BQjxClS7R2DrBtHuT/Cn
0VGdBPck2Jdy0PcVxBME2xCudmFFHgLvMGk1q80Au8wuudewrgNXszBhz3ENS4422KJ99sox3Pmq
FGBDbeTdsrZevXKKI1BUwwgoA3EwzsemJCUPewOPhGk0c+7IqjNG++ZTKS8+bSMnwDMKOwwMTJxt
nnHvwgXyFIsotJ+2lChL5CMpB/Nl1eYJ0kUPEfN9XpxaQ9AbXiGro+SpHKSI/IhuP2GP/UXieMWQ
3kVs2YWnS1Hbx1DFvqpk+oK2irgm4vpz/hqN2Q4ZijRkUtHxVmfxIedvo9xFlN3up/y6dAbqMFVW
VuIMl3xuc99M1m3pnskSjaLB/uCnVSkugdWs5RwguIDAj/2KNaNbLWKHObzKZU4W3eAvQqbOGddH
u6BIG0zzYeNwbWS4iTArLsXCnlIIfkwYMeJeBqvWyP7KZQZ6vT2CNeA7b0uucyOlLlMlzEN8NEqh
IisaCu24SWGf4CPoNh2T5VCNHyc3TaZ0QLpmrN59cDhmOBBlA1qfXt40+AzP4vmFb/xb+F3QZkPV
yACtC+BzA+MDG9D+NTKLXqxZhkHPihfxx9gpMk4lUhsO0JzIsZrC1p0bvajUT+EGrC6vrlabE/GV
majxcXIGBvLfE9+jrCiGjbfUMMnTdAmmWKfME6CYzSOnaTdeunZ+5AeDgZSzgXKxucFS1uw5cxaz
tck/a+4Zenp0JYwud4L6zmWPrrvUNgNenm2yJZYKPIzQ4YMnvJ/K/GmlsdVczlCUzEZqTzicxncP
FTgylTmMd13Ajln7LTlWhxjamQ7ey5UoDMI+uD1U6DqUtpMyq92xk1F0mB1uzzbiWlF8tvfy8dLf
0FiAFcZVsl996O/RdFm7p1BKyxDJ6Bx/o4TqzKXxMTbZ1Zu691VJmZiNpBcnfSTP1/k4XPj2WanI
K6F7jxmAebz0Xqvltva9bY2aRCqLgI6KmJibZlYR5vBcaTVFxuSukuxVeYZ9DWTqEdgtiO4WJudu
D0sm5z5TdOxd5JtqhQn8qtGCIMJECWkXqldLp4clddG7nuDqqpDYajmSPvcoErGEP70y7BJneyTQ
4v0cBchsEBpjUa8LeeOVip/EWy8CLYEvctVLsUoiPO5In8gvsSfvZD46sl1tFEtk/tqUE7xC0Pix
PmxBLQ92IPPI1thE2VStCUahZeW+OBkkPGx8PZrHD76uZiBkSnR2qkaIeIlZrjvet+t9oKCBnjTp
6NrSJn4KsBVQmIRvVO4L2DhScAlf0QNAl7AW1DtVnABcRFbUzw6b2tRHiwlGjSJMH2ruCKCThtLi
Wvrn9N3V8cDMJZXnkW548D+0MGjaZuGBWRMA3UJ257f909eqV5eadMG8R1YcaoGhI/brsdubbZok
cm/eUSFXJilWAF7MFyKSmaOwBQ5BhG5XLsnKeI+iRAIcE4HLDKds9uYLQ8Gd2d1VxkXa7Na3wx0Q
rbbq654hmIVET9cz+MuqNCfGssdeHaWfpJjU2nFGDNa7tWaUHDpN7iEcvnrQdr0JIgZGyOXETQOe
+m+9KmAIE3qdS7cohAoi/9jvjWFSLSiSDF+iWnCkpbb9hbfxD2E/KzeNQ5qgcW0n4kO/O2cNMsVA
mAcSVvinCyQAVJJa4LqxwEjD1M3LZxOnnDherVWEmF5Bzcd6h1ny1tJSnGY8WcgKneD/i9z8qnxT
0lOehW6dyp7R23RAk4PXyl6P/jkolSz5c0ZXFyYYfR5WpfhygyN8d3PPVvfkWqn6ehkGYlFd3Ehb
ddoMIrCCJm1iw/ntQ0vM6MyLygEkMy+IZS7Kbq7jLjWVCPaVUDJwKCrI5mPvlOFyhY3rBEXLTIyi
GRJMLoZ4XyEu7P1AXey1EW4PwYVD62D7BpLtWN/U8VkhLDeordULj4DloUqb9v7Xqjt+0ddmohYo
xqL7SqapuhlFeJHAASAOwvwpnFpuCaGEobm4+v6CZHnUXPad9FGEu6FE6JA6mx66hBl4LAPmjy+f
Bf5NEpqwhFn6I8WBfwPUVV/DhQIY/OtUInSmhf7XZ8HzV6t1exABV3yT+sHgmq3pHPls6PMuQpWZ
nuwXQWcrklpQn1CLzoJt9r26C6A1qXRsDm1IlJVRDuiT2+FPipy2cTmgrPEF3ob4kfxqrGeH6rWQ
6I0UBZ2zllVGBvFCZxf9iNqg03wbJ/rO/sTH28Jbc1uUA0VNArIxIXvfhkJr5eVsUgecgWLpNCWS
8DwOY3FOyKupT96x51G42BJrtRptnLqJzcUH7gWQjqgGKBsJv6L80Pgg7sfQAOflB8M8WTezo/Fn
gam++fRfb1kcYzqXrGVSh5T8B/+WCSxsjl+5raY/Sfkdy0Qz0J6sx8MRvxV7S3vg0bMzDCzsGD6J
yVv1be3EGvilv6/47uxX4Ok4PSr9WG/fW499QueC6njVp6P82rGwnGFwriuVcaBtWuZGS6uFg7F3
7Le6JxYJt70kzb+mfY72xcHhUyWAf036rg62klbqmfILQpGepKjTgCxM87dyrIDiT3UJH+2mGd+2
W4B9Xdv1VeBuuDLZTpe1v9EwdSd7Sn30+t9CreU3FMjab6c8krlQEjKJ3ycQlkb5K67f+nxI1qeB
37zFnNWfhl/m28/K7YQUoEV3GSKfgPK2MyQOrq4xHAsxgTLopLBBv8OoKw2o9CF2LM2zwD6ZMdKu
A9sawR2RTDILzUQbGuMNFG1CCfhIlpll5WyhcYN82gg5cbf9kq3LTuyV0keveCba8/0GsUgkamRw
gnaJP6+BritP6j5Cb93LCwnjglzvcVgNf/VKlWeI4NQZ8PafGRihQcf5kcpO+lzXKq4tAdNbdyCM
Emw+RcRnGpD7p+FKrPxA92bYBlV7VftnXZ7uFSEB6oRlayTBB/cQ5gVIpdKN1vMI/hxK/CqS2ycc
rj/Z6PFrBR2TO/fjVW1Az+EP1K1EPf5BZMByTe4nHRye9VqetrNZC8+oeLAR+z5XViggsNucOk90
VQPWp3KbUJgUl0f3nkSsP0sUJk4+yx7ePX4ZuNZazt4DbYBx0hv4DNAiSZfw+JGx5id6cthTw8v4
KQTUuIq0cUQiTa6aBFXpxy4vg2oYhd9+GDTok/BEeDSW+HSf5W/SSrcFTRWuPJD4ivVSn8weGPJe
l7xpKm+9zw4ux1f5IXjnXYoWZdH7aaF4NRA/lEqOIWm/KUQbE4zIJcEF3CGZFOtbdlT/tXhq5hFp
9S/vTuVbJs7D2m3lUiM0ppCs0apbK5ccjZKeo/iI9b9lsvPb1AhQoYoI2RT3lz0aor3/sQSF5H73
H6kPs0N+yW93HL+xwlCDUSvPu3XLjnU1920UmKXMdSVB5FtqmCsfcoqOkCrzEoQkYR7vf9N/zLKN
4rpiO8Mav4HZdc8NAnGrBFd6OCiBJxxruicPAyzl6DHrubm7dc5PYn21rVLOBpZF2cK6LdjXWUq6
sks2PZLWWyjlq5SIdGaStEgG5jon+lrswxygaj2rqcWhI0XNPyed3s7DnT7tCj55rTxCt+3C3sc6
Ek+7NCT7qLrClxu0fApWAgU0Q1t5kocDOzbzxSUknR4beoakEgzwPI2HkuOiEpWMtJ1rfh58cZZN
ULRbHbiT9P6ANRwoZTWO2dbibBM2PgO5tCAHlG6f8oiw9je2AvqqVPvTTdhHmel1uIjg9Uv8wgti
nM7WTCIJajnRc5M6Rff0PJORtm0ft3Whd0xQosGEkB3Wdv04yaQ1VVtpsDPUDm83O3CYCojIQ+Wg
xJtfNNJAtVEOsr342atl4o97ghYv3CGe7hKHHmAiSozK5NZTVmbvjvApbT1ACuo+6QyPxCbziv82
mwnNkl2SH1pTjK40SsmhTDYLffsdxAkWOHznMBTG3nnXYVo4XVHxZPA702Mx+lP/DA7bIgjfiMYD
yODgKXmLqpI1o11JshfDA4wc+2F2Vt2Ms+tofKgb+sxSVjT3Q4j6TQWCk5a8DVj9TX9I2XG/tMMR
ZCdyULy+gxQfhPIIy37vKJa1x5f8k5+fu2EZ14Sbuku8rcuVPB52aw51PTyp3Qjs3t3T9pbZqhys
emIuBTSRbD/CKf40ZaUPlXkyobU//W6XB9365qmbOHn3PYJc38XTrQbWHl3P+IPAZ01Syf9pPQp/
RuZVwUJbXcXllCp1L5WCOuBhWuM5pygmP4Kl9fSh3UEDRukdAUerd5SEheambf/P6d238GPBYcAf
c5kgHCjcKD/O7nRe6zXokgb0ufAWkoB3zq6lnQZyTvdSeL4Zs9HIG6y1lHPoNkt+nHm4Ph2HH/Yg
kVXOhlJG3gBRLHodSOgGpcNulAX/VeZ/ZJ8M/d6qRFpovcDlQuhZitK3kjJs49uHByCnYQqIohgu
PT3FgpfCW5xFObVLVrCBvd5OrFE0+sjkUqoAshw7yDfsByFJCzamwvteVa7gskrigEgnedxuulfk
q36FIzQ8HfINnusm8/62AY0oQaQz2koA9iXamT3Z0t/DPJfl5OlHAm+GEYTxTU5KbrrMdE8YEu/g
Xge41SRAfsY5y+iRfr4dgSqCt4m1YiwTxEKWiZYKuHcMrfBruCH8BvsoqFtB3pUlWcL5OewUpnV1
omNqBtB0pIj+q3dx6/1kyUkNHpuCH7U6Ze8Z04smU4WGR9Jn6hSx8QGSohJTx+3tz/34P2SRy5tj
30UsvPvkrdyVkKxdcg8mLBcMD9LTF3ZNiEBGM6g2eX2UV/RrSyA79SzBbFR95FSZWB9+0/wQPPFQ
ZsEF2TTq/FQAOwpTIi5DvLjvZ3ruyJIo9f4WyaPC3i29lRiaLJpPY9w2fd4yujzOOdPi1JB0ujOr
1lvaAB7b55x3nqrIh6W2+7t5biOUTNuTn/87bHedK/WHznN7RO2dXyQeBOKJ8RxTS1EQO6HJHYsk
eSLNgO8s2ZGWSw8RPDSvnnco1OnlJHv/FUH0KlPCSzFJKyeXyGLuGpumW5jIHhk7d4TYYzN8rhka
6d541Yh7ClDEbN18EjifnBSdW0bSy/UJZyIZLeJTCD1u8AcKfgkw7AbolxJ3q92t7T2koh55AlaZ
5N1Eeq9edcY7esjMWHoA7Et7nubwyp0QS7+xadis91+oLW+zGPPkfPSK9SIqfGLwSUsXr5Vn2v7R
ULp/bKTF0EIIQVqT/4F7R376kZut6xtC1GjUulitm5x7dJtaeZBqfSIK40pMykWeO9f2UJg06bxV
eAFsmDUXrq6G5fqShb5bY9JbwjTv/UbPhZO56F1WVrhRp1eusqZtItZfxispt4+J/Acn2121zrP7
snqqugeZGQ3Uo5C7nV/ytAr5xRaj/ja/JD5fZow3K800vvY9jWJ3O7t2Fy3d1tUUNbAuZ0lm5ZYp
yTmoENSm6vfrbEk2LsKr1NyN1zQgsJ2mO3kduFKDkrvP2fey7cnsp/KfTZFjSvQmzUHo8TO0l88Q
imo+C9Jb33H7pGuqdewwhT3jTz1tPi2usCxtcZfWRybtKieir8pddKpygI8NyWp7TO3fgTU1oGxG
o3Osk9oBeW0Puy2tvFtzU8J4kIQAEEBssf6N4l0BcgpklrmGSDgZTMJ+nwQJmak3fss9+YbvtXGR
nsgGXfq/9rfLGZoLXkC2WALrJLvOm6FWmXd+5n7WybQqk+4AwWPF/DkW5roCI7MUoVRiGxpMOOLL
SPtGxahnFfsjGjk44T/TXGAU1IkXWviiwO+9gPaRr5grK+Bluc3AIscXzi8wgCZvIqdQTVxvKiIU
tHk/DI7BYbYTitNht23jabBLmuAxf5msfuJlAbXOWLnI/Db4Oxq3RsTzCWgJGyXjtSVBBER8BCwm
Z2V63pjWXoEuHurfIqR6QXqgqixiBHvPAmAQSNr6B62lQdC7T4ZWjMxon6rKiTSRuRc6Th1mG7V2
8HK1sVmFOBttiCq42lY3rkwY85G4xhnFcwyZgPbOIkBe8xQfJ+I49rPWtc64akLsvcpAoGIhK0uF
nomi5uRm9shA8ZAlwlyRiGhyGQf1Q6fQ9nTpaymWB9lp8NzJn5qa3iqfJAmZgzy1+SXJFYxCpr9X
PgKVtblUbB8WqXZxigSUGR7/zG28qQQND4k49WMIMdas/zL9reqbEYGbdGSLTHXwp+VvSuzcye1K
kCHFqQqtB+D4pOuAFYbzufyQF0z0fEaN6RmS3O4kUTN7Izkb8S8zWaUJhLbt+Arylvd1x0r7IlPT
Nbsbnti8szS00JSptckiPR4t2YHNKZaZZjskESDlhybw8bwtKeK5gKt/0NPWq6G/zTZPR1fKZoUB
2ipPsk+CUUSK/4J6+9JeODmGKAbXtSt3Imq7trY/XNMZ44aFD3YvQ+85E0SHQAU7HbPuFY2g7xM1
wJh8eJrM0nTYNZcEeORn8f0iEAPr9YOyA0MdPn7/uChGie3l8KAz3U6V+xRPUMrVsbi6hu5OxTeE
ArNO7OtFDZC97nV5kqjhFrk6apO71i/lInX2a2SHZcTZ30ibhzh2MjA9ES30eN2gZD9Iv49q9VkK
fcg0miWkOsAxwu5nX7+5Aj41As7hpT9stWW2gyvKL93HOjobHsNeBUwj6siWDYN4o9CYfwTPrk0V
bMv8MveBTRN+we/wzqJZ5A47wnsjmATDXSalChLRr1KXyRnfn7VUiEtuenSCtxSiwcve6G7McESk
X3P4b2aUn4/OzG64Ddr+NywavUb2qnyPYKz3lFEnM4yjqk8ktf6YGkob404jkU9cw7+mdtU1Jha7
j4aIg+NWXv8DTQOLp52Xz99qICfVB0R0VcW+f3xMrtb0iN7QdaPjn1pjmLF+fzP65lYT2DGfALt8
OMlLrRx9S85SIdqrhRSPYBoy23Tdp3s2/gNVuat2kPh/HlvzqV3+VOtBI/lu3EIlxyL3sTORBDbg
jcHStot+YSoK+i5HT49B2uCo5I4qhayJt/TeEJxljvMBXsux7zYTpMQe5x+2lpfpiGg29IWxRrwA
wzkL+axk1sMNNLqW5ZkhRjH/Xx99VbTs8cd7K4KC3vycxowC5H+nN1CD8yBLLFS9z9zF7CaHXYip
aQxQVYeGJmIEwoaMrr3fkSsmc4UYQlJAW7aiCqxOggk+iKHpzm6cHAhdqjQxmlbRuuJP2WDGhh7u
wiDDPGigCOUJbDFNXzjh+qlfqo7YCbVrhsY2YF5WOuVJbgbSYQllIStVLcEpZJYFLz17eyAdP14A
vQAdUpX0cuNkVfsiJMU7asWTlC4hhT2vSSoLHyg7ttM+bb/mfOXjBZ6ZsZi8UrDxH022Y8Xs5oRv
PUaiUzzzPQxb3rKepLKsFM1ALkv+yWHv+gNmiPoLthP6JUfEd2rW4SyTn7bpXjQ0Hzln8KeLUZRB
2qdHzfqLi1PBwQmGQgCvfBrN5gb1OwoMOijpQY5h+NXsWWgzkzL0jIgmfFNvEMh2s/0Uv7djHiYn
mdEWH2cWa5l6z8iaDZ8G+1OKDcOM4De8CzwB7pdLuaUwTdhoubnVMAjMzryVf11AFTfZIwdP1fE1
DJt+fhGhvo1lnM6kOF4pvMq9KnPYC+pxfBcuMKeU2d9XG0c173u1dJUNYASvT1Wfa2PPOTRWzyBi
8DklHjSFLfMAhoZahl58Sul0ngkrAQYc+mXcvjkHsokRhWNZPaIOjAgmcKdFkHsdwDoZ9QxFm/GV
mEsIwlPowhbbuiYQKlOBxGGpZpOBtmJMAD7pMr0QVtc0GsKLVBgKW3PLNhFn2SMpHXbofipfZEzT
fRUAjBJ9njRTnkfkPRXOzKnN1aijFRVUBiYGwDbVOs/FX7d0Zg+vCm66qQU8K78Hv7L96jgWCoXQ
izGJpjafKY3Xe6pDGEcxMROqfgJDISbCm1dsE8A/2mHHQko6i5DDkjYULduRUmb9J+htq6cOxXQh
nibKSSAkI/1Pi0miRSmj9DZqXWSa3GwV1z0oLbSX5aMQxi4hfSB9I48sFhBMiT4GIKT2MN65ikK6
PetCvhzi07rjjxczo/1SHNxZRH96RFNrO2iWO1AXsnm36n+7uDyYJ+u50bjza7M84ZkkMzxkhZF5
OXJTAFyeHCAmW2q7oxVICiL00UYCQSxrRSARZkIzOQdaoywgZDwNPDNsMUX0NleTksEEXC8CDcSL
pibhuaRtqfgPFr+l3uQHFdBBI8Zwq/k1jMMXhXnc//o+ao3wZsP0zzqVSAG7OczH/wSyF/FwJNm8
oXiJtkGrNwAONSf8DMHctCLmqDS0vomLYKkILXh+96BC3T0oV1JH+wxGOZMRFTAtS1jiJeunPoSI
H9wyMTrNYOkRMIEjaRJY5+SXfkJVzjfVsDsOSipBAUhL4r8vuAd8WowBZf8N3qlVMTofoT9deoRx
EGPIL/e83emDMko00PA1HsV/PyWFJKu/8YQtvN5ppwlRwHWoNS+UFN/tIsoKNjUW1AZDYYPoFBH8
3tDAPGA3xcmdyLMsX6VRTCkcn/AVTr3nuiERhc0xq/ZiZ64paURbxpVkLRr4pYMtHnOPz4m04ugM
qpbzVlNdJvErV4eTQC+pRna7pkrBnH62/JEOSB2A8Ff9tPyWmG1Fg4itxdrd7CVJZ5WHcH9V0Glb
buVPL+14VZVgmJLU0dUKeXkBrlx9UxXxwnyO74a+Pv4sr0/aby7xuHihzMkz5iIlX1lnDlPK+fx9
I6YWKx6JwXbJ4exrNUYYQOdh1cu2D2LHI7KG0bpupNeBXJlawBpcS7EUkKWRrmSLDOxJr742juzI
/UGBKia3ftdV/QIzO7rEEd047nesVwu5fKfTpmiBGqcIoPUjgSO/kIX/qw539+4x1W0ntGcqCuBO
PAurooOE9tD6veYU7A1V8JLjIKqo1BxvessPLMD7sO83C0dWV0FeMmYOagyawppQ2cyUZ+/oAO+Y
1nHPxHvCjT4WUDB/rtf+kfP5gbvGsCh+CPksayhDhHHycVD3fNMUPNcalEfyKwYFPDjvOandUP+K
24UMmkToEt9UUhQu9joHuUOQjvkghB1V6SrHJBlFF4IBCsfbtcGeAmibWIvcG/2gcA00PrkM1BQK
STKsjcye+Fu/t3vW/QHK4yz831ZYC735L3g5v/I/TBkuoBtPFqrtcM/laVyPD/2xvAGKJ/Tbk5CL
Y0sqSF/qgEcqsvph6W8KhI1eDPzmm8zmSe479IJruoHkAnkZdKPNWLZK6YUmYRBO5f87gwIUeo+n
03r79h4AvSofTDgJXA/c9GH1IDMOwYE9PrdQtIfNjeed4FznPC4zi9TUNNyL9cRMdYymp9GR+vVq
36EYbq4eMb89iMNWN4O9Rdmgo9BbcVUlxyKN+84sTwCNtMs9h9yxpgoEhhTEF0MyiaUdxQPGRq2k
CqnsXJJEjxkfUqoxLLX5jHwkM92rK0++g9fHI5JD78Ko5HlAui86Qq+XicBYKi+koWBD12q6pZKZ
kth3CC7jTURsWj2y7IP1KYvvLCdthLIWGMTgHiFWLrGPDhf2WgtOZ3YnlhNkk+WGrS0ciB6ht9Q+
krHIgHDIcCPnTCXo+N/ddEn7QUOfOHQhi20mYsNnDvT/KIjASTI3N6DBz6LkcO/vk8o1bxYTAqQg
a1mtr2KIO3Lbf0BnUU6cfgyajMwNY3wIAihvrLY370Vg86z6wizABvZfGORKjbYgj4e6Pc+KNSiM
wtPuYuFTQCQcpIraG89zA7Vg2FbK+XyY88UO0uSjiuk68PNjroM4KL8isyN5K/tvsR4Kmwzd4/pS
SJ0x72yTIfpdgWGZA7rD6kyTyr76vvEyL7xivY6i2Js7zDopGxds7lSRJd0U9Tj0ZO8LQ5pcyOlg
0UMWaTP4GIa7OLvyveXl+sv9f4rkCk+yyqu/0XIbzwe+8PknYDx+Y/c2+P735h3zWAZ5g5y14RCl
vyxX8e+hBiCEIeUPs2w2VRLrc14ErDyLKW0i1Qm1VXV1r8IAIr2K+Xsbsl8JzWJgtsd7fFRMk/0q
NUe2cAjG9ZXLjxGdAhtgDDJdptv3dcf0R8lw+8eFTuvUKzgM631YE+2NgSdf9d7ND1Tc1i/GXD+E
BBJI2/4hTfUXhs6aXvYkrfyhHOqOrpLwcNPv+T+We0+tL1iEewho2eF+j0kUDAx1Vl/Lmes1Y1L1
/7m/d5NH7IUdZ+tPiYxjzocctCd9K5qosY1b98hps5nTbGWDkKope2GzH1R4wYn3EJmjfw+bJsF2
Z+3RgI4AkIX93stQV2vG0+Hvb1ZDP1xflXnw6i7g6lf6u45RdrVYBW276jmhkAYw5a0+7Tc1hPBt
nqAu6FuReWmej52b4I0BK7zr2Qx7jBj5+IKR/CiNcDNWiABLq1F83UYQl/eD6sXfVDVaYfvy0b6t
+ClmuGSSfJnn6y1VXE78H25zRtz+YzKQ5Z/ixg+8QXXvcR41lsCijxaX1/S1Ax7O1+m4GRZFTWjO
WpO8jCa2pNYa16MKDbuABpdjvCUSiB0WKsji4jxtuwch9PBCf+c8/xoeBti3E67iUhCL7PzM4JWk
PqVkZEvnp+yBjoh/Y5Kw67qFzKEC6odf46x45lJLQ+wkzj3YnEzwxBuNESiKNidEcVTKbx3rYzb8
bLpJwon161tVkHDm5annx61zERNXR75R9ggxsZSneq3ofulJAD4T43lLT+zbiYoMGBTiwoXwqKSU
/8CMm9Y+FibapfmQ6eLVUMi+IvsCAjrG3siLg1Wz3hrBH4JiRIHS2w4p6+/SrTq+cY60ahp6YHQk
ykshq//IYMM0EmVue8kz0aWrLrAPvxSsXtRfKq1h+rm2gjLvnkgR1Y7y+2VYJb5SlhCOxf9hqQZI
lp7nxd6nqijDYuCbOj19/fsqoFdh4vFZwCg1drAaaFWmI8l2k8r3m4uTAhtN2vki9AaNQVmTes0Z
KCIt3MC2BuCwvnVGnLLIrLKuE8BYZtAlmjtDuyDY/tY0SIjiAsL10DAePObDgcYvO5rM7D1Obe4p
YuEU3DapSzuhReqm325NGBGIFsio+FljpaqjSvIuwE9Z5oxz/rKef2sPZ4fz5IObfm8kZDetalgb
8z3c2UuM74AUq/3pQtcvHXMY9Q8yIrSBogxd0coKOtiKEfaSxWDU/lpF3aFZLG7MOkvc6HR2olAz
3ueXUVrGsg+KMbjUCCNkX2CxFynU113q2dK/I/QAzc1L9xWKOKC1w5gav8MlTaE1ox1NmvWJsi1m
634Qgvm21s2tWYWZMnjOwU32Thi0w3Y+rQWY1ohuHeIKjDD6VNK+S+8xGtsyTyX5h/2Ab6wAK0kH
3NUMIRPI+Hnw8tn3t9UqMzMCl8f96amThv8SRr6QHdY8uAMaVYYcjReYS96rh40kC84Ed2adtgv4
4aghI5iTNWO9CQnayxtLwDwbV1IlFpFszAoj0Mmq7DRESFQ+QjEsDePXAUHaBa3LdK0SEliM0Ab+
zM3AdsgMXI477rjJovDI9tDZUc8mEUZAxPcLd0uqdZolXfikmdy0iDKaPPqOLdts/Arr2qfRI4+J
qGqUZ+cHf0EDeZPlAI+4moJw1fzmNFuX7BlaRXhBtvKTdA20mKQESo1zGBgDVpx/3aorBrM99fKY
pAH+1ZEGeOJZvxfiw0NuPnbSstRuwQ3QZYtC//YDgI3YtOo3hmqfWLNQI8kaq4dG+ocOexNhLG27
XkdbL/FegTCFRQmPVxuQ6YUL3Ym+YwS2BASFF8BFCHXMFtFCV2+H19d8KM3TQYitmt3VR1UeBaMi
OchOA3vgPQ0IQVq6ve+3dL4Xc3KYc2GZsnvY2XNA+QfCAuHjd+FmIwFm9uPjq2ZLXG77AQKX0t1C
FJ9oxHRoGgf0kf2k+ocHLub0O8i//5l9qEOvs0lvjZtapsh2iQNcNE4LJNo/JUQ5Ohe/EQitb5TJ
BTftIK1lWjpwfActo8HoORO8JOzVGciYMce+zvLBXEVWxAqdNFbuRCdkD5DAPUc7ZsgFDzyvNl/y
lhe8Bj6Iyal1hBu0TOVj++Rf6SYzCd8rTBDS89wblTs8do8QQne9vir6i2mXYjRKGMTh9NPdPE6X
t9jEU+wRB9R5lME4wnYzBGbGWrNMuSU+P/YuB/KPW3y7eDS3QHFJLOijX7Jgzp2lkoIPyzKPmp3C
vkSD/mO4OH51oGLr0wHO5KczNcfn2Bs8AI66Wpnooqs3LqcKPfYTGwtmuLGsoIM8HU6RI3BT9jMC
wJdMza+a08W2uYFV6FnxJPO3WVzPEtP2vMAGFdN+cIkMMk6MLwwh2zGvrzBbgcvUYyT2ODYe3hss
NwzeR0Y381PYEpTcIR5sH0WV1DEqmsVLNC3hmgTY/f8H3ydiyuRO5WkUSlRgJV8Hs/mNxiu3s3BH
QEp0LS6HnhvlOthw98SxjDSdr7KcsH2sEDnGD542mUqvsZsa5Du+65+Aw20r/js8i8e0PtAYYicQ
v7kvGmAGqdQvQGEvmIMQvgUUcwFXhWTXBt3BbJXKvDxqLSqf8gcZDjz7pnJXG7A7mXjySPSxqnJI
1xzlV93r3U9yd11+EM+l3AejVLMzry1y3OkW8ApL6qcejsMTUPXv+po269XfQxfG1PbdZLouPcWM
w8d28EH3X24Ed/dH2aTyITdIJGdRbfGX/YcJbUONx6dSpVopHWA+6GPIKzIKHclp+BvOCk+l7pqS
Nh6X6lXHs4BdV8FPHGSuLBbxMfq9Uog7RfZM+FpQ2EFW79r0xe2Y4ipW/nbIWMNSSUXCmauBSug3
VmJv7rmggxU5TCMO8Paio5ey5pUpBSH6rT1fvQmGjf5aAGsQQeiJX69Gi7QnzookrAnS2GY6GlRb
GMtaWQ5k4ryP7EPkdRRScrGlTDzVAXL+wN3QSrP5OEU+vhQWHH68ccZOfpdOTkIPS56u0Uwo7PPl
b73UUmZ2DaYE5LZoJoMA4VZQ+E7tKeqHG9VixQP5RNplQkvzjiIbRdeHT21iRl9MmXkjO1RtuwJD
CPtiqJVyctEY+0XlbbmvYi+0WQzJz6KquvS/EJDx7IiRnCHAc1riDR0Jnl/X3SLjpCJlQYxmePtm
MQ+wNR7xPhdZbclirX67veuDsQp5FZWasw4TKJFFWo0zW0o599Rh6mtIgjT0vH4QoRlacvTRtcWz
p4psee1jTKNTvWxv3PY21fLmv29hWmkgqrIDt+XjmVjohkdWndLlZERNAkNIw8b8+RzOHrjkXg20
9t0vTS1bUU0XVWOkE+FUd5WGFQfrtnxhLrOHfCxXyZ80RwR5wns1E9/EzFZWnLCdYky1bVJUjn/P
W8dUh9EHEK0SlhfEAPbcj6lD2hxjty95rhsu0sE1AixHgRnanahQrvze1pZXMHjoR/q2UvEbKZ0v
4Nhbx+kBfV/mN0ueQvRUSu1HWFQ+M6ejGIrw8c0pHOOf+gcGrhj90mBaiOXTZVBgjNI3kKlcCyUv
jE5+N9MJleM1G0iEIuYbGOacUZKi43EoUBro+sjQndYXschOFa+v4j34dSlyyNQS67WTp4keWVGd
GCA+Edd+Z9jevHISfkJ72JF5fef3sgGghpqfl0mpyCoweEygvbSyyh+99Tkz6sCmycM8S6zWxJev
E8N6fLbOxIckMZU5L8rnERj08iE+bBew8+2U+TTUC9KbIH1H+oz2RWfxk691QtvlS0OkNu73cZoN
0roSV9KOtlW4dGJSHQQ9R5qKCuDxYr79/eIiEYQPRO4UpbbYpuLTziKBC99SHG1sJ3JPyTIGEJbs
0kKEC63+P6dVjPCdoUvyfQy8DpCqcYGK95XpUE4jiGnwANIOqKMNWClNoJOtVziwwe6RGHMC2DSu
ASlvQM+Lv4M2wA2gahic6h1N+odny5DxUUbNHIJI3qz5WSNcLCCnQd/zAhi/eJCXQe4B6N7nNRc/
EbUN1sFO5H6+3LVb7p0+HdOHiHN7JIE7hDCaY0xZMcoJ5JACH3TiDosjEjIP1kUNIRJJTNVzqrpz
5ZOQe6vH3DnZKcUPKtmPhR/mGy25DAkUM7CA8T3oK3aVqVWNUpXkE/fzI2ai3i0JbNf3ib6gZb5U
9mY31nbZQkMFZSm/FIK8VmUZFWD6uBLBtRpb1JrrT7+X8lCsb+plXT+dhSB2Egxhhm7UlnRpoXPr
TiusHF6jqO0JAf90G7whcF8Z2LL/C/2iVVsFZGtZTkpPlSdNvffmK6ndas0nMYYsN0WvceVRRV7J
6WvmQJCCpxriUICzxqNBMDoEoQADzmz2Km4g5VPHCBYfUIDLZMKA21GHUbRzhWanrNv+0XKASN4j
Y/JHEvnSJYYg7rJ+aWjuwX9+lflYhHxS2vIfr9H8Lv5xEqLlKw4HEnl/2Ur0XBu4vqbGPTDabp56
f3ymYUoQI9pH1lT9DE0U8DTkSjDF+Oycii4q/Iq4bDJoUfFwobMqlOu09jTJv8SfYSvbRlxjQEnp
K2EKJk/waeJKvL2WHHralIJuri9+uttd2Jclrt1Y0lihrg0b5rJWbVYzWZKzFQp5Zbxf3wtRRjk0
U3FslBgFji39krULpaNR47YhfEE5HlzGpdJm9/qp7RW0YgiNEm3YK8YwFmUPUg4PqulI0sIYxKdN
hrWnvUv0PNkoPuATDI+Kkbb+eiY7u891fKVG0ivdD2JQEuwqqJqJEhosBbva/dOKbOMlV1+vPmbL
+/Q6DB79zACvveqEKn/gWEE2gzAkQTvRjYDu7p9DmmbzPovTwZbt4PPvVBj3FMs3u8TLQA440Gzs
kuiBriQ+kOZs5X95N0ESk8WhTkmInmEY4gVeZ6gMscjrIL53t2uDgqF9Ro78zfc88Sj2IFeu7FBX
yhZbHbmKAMLLDI4WpTFvP26nVCvClqKhc1aqPKO30vIwdfNYnRWgDEaMfHXc/KGzm9u6ctXNHMBL
S1Gay33uyts/rSWctaiIJjfztXAJPT+RRjH6qx2t0/Kf/SzsaXw967Zz24RlvRFuPuK784RJ9Da+
i5hu707Bu4A0ROt0alTNsrDEfZrekRQfNU9c7EQPwzU9oDJI0t3U7C3USLsDWbZvT/9JMAS/Siiv
CI3ROCqDTuYK+vhRP8mYzgYXefCf1yvylnTusWwRfk/NDRECCUfw1driB/9CYIJna7IOd89fTBw4
GDQwBvc+1WyyUn6CbfpkJAmYS3j98ghUhFXWGsuPxJj94FemQpvNRFIfdMzmoCLVRzn0gCwox73i
2eFC66WPqNi1FDyH+pOJAFQ8FY/j5YheaE60tXrhfcbfdKXcUSvCtEl7fZ/Yah37NL/EwVGCLGK1
jOU1lrNAHepW/ynV4y6D2Wk1ssHNORkD/2BezebtZTXvHlgc01WGptV99K//SV/wcRk7SyX6LOiL
kGRbQ19HTbMuHmlY3slne+Rys1tv0G1lkZZ/9hhn0ZRECKVPZ3Mc+iEB5MyO+GUYyRKnnNXH6lqo
lfI+I2BccBAsj1+2271T4a+lnsb2Cx4Q3oLV6NZTTO+DSGcx3ccIgx3SfQkacHE4UjHfiUhlLk4K
JXNXUe80UlblTYdquIW4IsaA0mU1HEVOEkl7JlwunNcEIOMhaeLKFLshpEUxHXFj1qa7nW5xa4J+
hBzsMzo0P/wVZ9PW20J1szApTbx/EkgdxYs7awr+/QtgDmzpeg3dBqGgBmBE927HJ52UbJ2IHhe6
qL6tuoM33tQY66y6C4wX2TmZhM4bwAt6P88e60EvLuduxaYsdJ8fqbWRownCKhpvX7sox6R3Tr2P
SI5IOj8cdlytZTMmjq8afd3QMdYABovM+psdwwc46qBayKXMqzzrzoRz6ZnPTa79YjPj3w2oj4Q0
u09hdJl70r55Cb4JsLJHPIGcEnNsjvo+zUUAubJzCpBqPMMQjCc7JoVWjFsy2BRKNNHUyfR6V/6c
SvewRx+yosNzOPzBKdJzrTKmMbsGLMv97XC0YfhfwBbWe1jq4E+S3E5Lsxc0c2LLWciB28ceJ+Wa
T5H8HJh9v01yCURF3kFV1Yjf9q+nCxGT6iN49yTGFsCsv56X9xEGM75CCyHeZ24AplZwsd/lhJnu
ubHqYwSLGJFPqvSzqaPXiOKnsGPry2MbmQ7zWetenN+dVQ7uSVIfdcHeCVfZzg6Tretc3MHO/Na+
g/Qfz+xFJVa0sy27gg+TiyJYeGCXnOqvDB5fpkJxM6u8y7K3WtuV4fjtds9jDfWeEb4FdH6THNjB
VrO/EqwUcqo5DrRAuIzhddoWp+qUZtGExKjUQsWUc4Fc5L6dcPlQ8rRK2o+0Eb8YpEddPuyXrrYl
kLfZLtX2nbvZPSc2WFx8XHYOMhTps/zud9rY9TZezpguA15z4dfuzGi58jUC4ML9joRqmmBgb9/J
unulv4+mMnI8xR9vixH522nNqytK6SlyMEwGWoVZXOhnZw8T/UjBlkBOJT7i9m2kQwgWP618CbJV
suW1dbhaHeBGhKw4Nah0yDqkp0xklCjv0LiNgJYbjZo51VZeFB2ugJT3sBe5xx4ygU2GCi8oKWFu
4P9oQKsQZBgPPf9lv9/uR329jF5H/EgmIa5EW4x4dfllIZb74nrRIykAfnux67qSulfmhDkuUK6P
SuRmf+WfzDc1eEsg8WH8dvmJvS5ZqMy3a3hRl4Wz6OpwaAYtjhdhhWTrg3RagoYtUE2jaJk1l5S1
6UGSmve+2zpKUbIAtYJdvUT/N4fiRn+0IBQ39Dqbw0wzy5CSJ53Qytqv8/Z07u1b4W0n5U8fMVUt
GZD/YPaX+IlnQLfESc8bxlYTOmS1OKWbaEZQTdMUF0iiecy39Hye2cLd09z6JPvdMO6BFNSVMRXW
vhnj50hm5/9UHa9Sbh0YNCeXNEfJP03g1L+QUNGXoJPIar6W6pTBiJjuzYfat0ETqvOXPplyzApK
jRFLRKUrWoOdW3dFUKxf3zAQyRNjJ/OnMhMW5sM7WVZ2eFVW+WBS6KXy0B9x51xEpPl3uKkOhURi
Hig1ycxCiT0W/VlMGtT1Dq41vZjX60hXukiItCcOn81fjfyk39kAd538iW61aUYiWb2WdsBr041p
22iIUqYCKPIRgWXE0atGiHUgO0J+JMa2wS1L0XQQ2i1WAYK+2osOl16m31zqE8dqInye9Ds+7Ddn
kTTgCOz6IeeTdxQoqd1rC8sgyinquTolGFv/qVkf6QCD7hDGfcaE5BBZUScgLpZU0TomEtvSxMbT
S/kJyhRpkC+nprkFK9aw5KG5JlB97G7LbIId9yNipRdq1AgP21f/zqxe2rcvQwi7l+/Y5numxHK5
MyjVYxVL5amg9Q9fksqC2sRdbDm/ClfYQJiLs7hLUdqbuTk53JEZYKx/CbM2Lr1CYlIBFnfdXn5G
R+wMV9ItfcA2duQbO/2s9DC7ezwHHQ1XomKXUQo+9msn6aClqMwVjY0BLZqVAKdVHVbN1m/McR/1
4jP25i0u9hQX8rPXImGoAIrffBceFRz7iyA3fnpFlT/Z7BAtbaywNd0g9ovdI+/d3wyVabMyNhU3
HDHrMJiaWWLVSW8sDhuuz3ZEqSqZByb9MC97y3VYCdaRI/Nmj4K3qs+aP9pJZ2W2idgyp2VFeh4O
kD7x+0JbBxixPnqlKAjk2ONGKkgwvKMGb0ha5sDxGp94nWpIpHNXBeAb8sSEl4srr+NfF36V/J28
WhZM18rnwtBofbVu3erOZj47ASP0xzToT/uZLA3JgRATsGK87Z/ziw/TZc9P4kQ+cP17zVE38cWq
9i0lgc7hHPf4T13xo/H4bMWRAQiRCHe8lKOX5w+lBLcEDprHuNJEW4TgH2izHPYKTGRKCvOpgCgE
Iuspj/pbItBkfl0owJdhSbq0ZnZvfggwZU1STcWCwuFsacCI+SCrNaMphXVoOOt/EVVr8BoSZRND
hgRNawmhy0+xAGs8RIAZde89XniayRtDnu+mezSLvwrCO3n3xKZW+TqppLbcEbXNZrTen7eyY/32
4wbOsC7rrG/KhyPhhThrmkfuigBZpBx9Bahp/GOoxg+6pdF8ZXDqF24b7rMEVN9eGfgTJlNisPEJ
WxxvCeQqQSFy1YD1AsE8ZMqdGNYmX3wo5/NobAXyw+5/ugimkHr2VPLNXWhdETMaqfaCb5oJD0Ic
KuilFFYJFXEFu0rk9/yF8dok15qr/k2UehUl04hHZG4jxPkqNQAaqHInQ5F43F5pJ9AVj9T970Og
7u6WWS+4oZCqQ0aue7KkKsMWK5/tAZqEXd/dNFQ2BytdBS0TQw/Fnebc8xidbIivBsxGMk/PugN4
n9XTWcKHLKRZIvTPkbthO/tyD52gQuYCgRwrBUe1juSP1zF9zCwww4f9irvRMBfdmGoxwV2hBGbI
hEJHeJfxHcjczspUORgOlYARRUqxL9i09OZCRvIR8k8vWEwknGYa51UmQDrktuPqZV6tceiNQMNX
iub6BHXYVLH3mLQEfWQowmNuheNgJADxqCQ7jRxzowuwdcEaWYgKfX0IWgFXiRUbDiC24RsU1wZ+
F5FIDNVKWIQ7HGbJ2QaWawamuLs9SLRjnHi6UtGnaQ7BxVSbXBWB1NTWZUkR/iE8lXUpEfDMm6i4
xwmuo3a3QTV8KTeYkpeMcj3qNsX3U2wnqJXrSLdXnrGBUdg4Pi+pUXtRR13bC+oiLWJNnXcqMxD9
cxQmeTkjMgnDFCnAetDsEd1+BLaTPr0CnjRhXyYOYs2dNlyqI//q41IrWZMZlJn9XoN7qXnq1GSN
2CLsSUQy8iWMhJnFxQbs2cmG9zE2GgbMizFyPHTbvXBG797uuqCHWjc2EyHHKUO/GOel+j4hNHhb
MQNNQvtL2vPrEUErtm9WFGYBOcc4yk4Bsf0F+Kp/UZ8GAE63PljbbsomhFyUkSp0RRXIffCbgXer
YTmt7Ur1d+QYCyFGpMfKzivql755a/+1VcPBHIyl6xB/DnI5uBBLcTM6ox1z81QDpz3+ywf6A1F0
Vc6AH+r+gF8fIvRjhadDwAt4vlfnHAWWDsuJTa92UnZsXlcoy9IYiKb+EwRMA0W9OiYJQXM6vgYm
7msd6VVDLK+sNbZ8q1c1KI0JTPBOg9FJMzoQhDdN8VWomveat1l3UOAULOLaBTXuHYRrtn8qMpEh
5ZFnUn7qCSTEf78yD86lmxbfJiAnSAfVw5qZ7Hk2aaSwssPxHCptPwSfLuEI4zpB5pn4HcTgeg+a
HtFFeBH5bjwNlmSjsuIqQNsiBARBKqh4Z5NIF2Cf3wO5enf/jwxuMTCkVDCaEARCOLnBFiAqDjfy
V3iD86dN69nbtCNkYfLgTXqiGJX2sKMdGL2VI+2mdFC5C4bq00rN7gZsfFzS2vq1zqQtID1YJRoh
EGIkOWLvStxwFXnuxfoxs7d1QDZ3K34kpQooK2KcW9zP70ldUrXIUE9t7jFUmK0FP9r5Qk2FtanU
ia6RwMl2hJbSbQds92Qiy9xXdB0s+DckyT5DlTc4Jgpl04g0kFv/QIvTERnwIac1HpfD8Cs8zyMr
6wrMg4khwtvekk7Adi5ShPWWu3hr/icwlOdWi8K+nep9wMVsHnvsXeTvOUGThXCmmT1m9j1b/0l+
do+P0GYgTV+7XtTHf9pZ1wi5Xmq4ZzxrufGTZH4MFAQGxvRm6B3/KikvD+d66Mb0VjuM8vLeQ+cb
WX7I3F55W45Gs79MCuyt+GKaTyoLzgvJpDh7u8iSSZZm8iQMKlH6f+OV6Py65b96wxrWrYqHLtlP
ZwoO821PHULCVniM64Kpf/eHE3J06As24H+wfCj4eLNM0lVPccoCWsWXNgr3f4Vl+WP11mNdzGO7
o2wyIODXwvQjRsdQ76keZokB8mYAyIRiaa9ivlZM8R8idy0UVHDnoKJTM5VEtF7Ohf/hQAzVacce
2jH+EGJNvB6KerKdJpdHVJuKPriqmlmn8d661brnmB7HDy7nWBck85Uo6MYv5D3AOf5gUVT+e4kU
EInj52HX4NNOxFacw5GRd++YC+d3zEpaXsEyD10ouz4FKWfUB7gQ4tJKG3cFEDghAqqc8EDPYuFK
aD8M66ppgdRGzry/E7S7p5mrxtK0aQcPTRX4xX+nep6yO/46+bnDBHPFINq8K3zkR5wjRS4lV0b2
j+HlEQuE95egPbEAhApljMhI0hAeJa+l5rNw92iwxKEUZa+6E3qF8H/dyJ2pdNnw886SYwI2EvSD
fdnnXArSAQkISb8KFgnVt3Wjq9KyaT8T4z2Oa32VPshcO1BXP2nAIG2KDmmgvxpTVZZqlXcAg1lY
f7Dlw7Dp0mBBAGfy/mTS09b/kCQcwGhpLCQzAC6K7Ncj8zRLZ7WJW0nsECZTHhzBxvdzVDLYPw7q
vie7BR7ofjzMdaRgbiCExqMkAj9k3RJjP42YA/tprHHcTNqBcXufztAMruetyzhIqhGRLPCA09Jc
R4jYD6TzbPQ86ofKudg6l3MSDPzywcXtyaoF0zB2cPEnrZtl4xdig8dHIIEvDSKCzrLih0W6lKcq
Xt+wF7XOXpf/Kobx2IwrjXlh10JVmKYrLvbMKmwQdYwmfKC5lf3HFQdFFHS5nmYBXzugS8YfMH6e
q4mv8YHdlpF/5XP8f3K/ncH1LZAh56b1gyaarFMFHlUVcF81vVHsKNnpEMFMp4Gr4o8k38LiVEX6
oMNzo8j2mRCxONfCFWSaU3nKGmDRbK5m6y4SfCA5msgh+EC7matIs/I6aVrmFZ89SPuySG9MeNz9
k5xN+vC51zQ90NepDySyR8ZnPLgjh31pxkl0aY/h4/rhBP5/V6pGncyOabhFQLEhYR5V3+oL+fAA
JaHtAvX3Pu04KwePSurqiIHrNgBWZYXTlGKM4YxOHnk9c5rmiOkE5KIp0Y9zdrZNCZY69LmwOtu7
SJVPelq1OSZlHxaiC+FCL0hmrUQzqF1gsZKr3WSSUu38QsncUWraSSVyBMCELPOCZxG5PR5gOLVe
4lmRppXPtpVabVFDYVKO5pK7a7kqaGQSMuefOF7c0QmCBzOVNPg2bZ6Ohj2gOZMfKxtNryLqOl0Q
DrwA0mUP9CYA7bOu9NkSLySLHqQYMK9M2HQ+LPBqxUZ8P5z99AxA942LFIOavFUlQd16cCL+kb4M
AHE3TC+sxCL1WNsgk3Rn/1Miw5ZrH6QuwG2T8VQggFipoX2HwNkjQR5ubHb91MylLvM4/IjpD8iP
F/hPvN1zH8OTxq5shU63hMBMr9QILKEPzXZOw9UtftvyyvOvhboeS+NhzjEHXRivZPJ7lMcMCw+J
k6xL7M39TsuMMuACsnSyy4CW/kMGoLcNu0L6+qljK0H3GnXAU0xiTWoQVehprZsD8KpOCyCQQcyM
Z85LawSdQe7IzG+9d/d7Yo5A/z1u5eEgJo3ZVVVxD7DPIqvwXSCNr19No+XjelC+4dH1WL/R5N6N
A5+jPBWRQ7st6CBpvwvEMT81uG6HTiwa9ZhhkbXqyqcfuj6gPrLQNqBto79WmcIMTmpLt7smM/J0
BEB0BbLeBeYaT+MR24wv3JfjdE5oazpIrh9S0LQGN8A8dZmbW2p1jW4tNiHNXzPVWcXt7qZK715Z
yNiBDvYWAB7drB42dvv8yYwtw07uTqo911fH8TBsqxsd0GeArzV0JJ8r8tP4MHRpU9V3rwU/2O3v
u+cD04LNXlVHGOp3COYeV4BT9HW7M4ruoL2sYX/zTEstRzNpKFvx8ZVG686du8/SbgqC8NBAa6Vy
FQeoLoSvLNB8FKfrD5x0awOw/07bbDu/otQLLFN6e62upSZDy+72R6xgHXbVbQ9QaqKC+rpDf9gu
oZiIKT5EcPVBSywAWDR/UhrrrvTTM8Ye6RPsFNjc29ohmxO3KfemM1OyLksdECova6zU3E6y4f98
+ZL6tWMJZoNLPhHojzPVhGhIvgJO4IPPAXPXMsgo0/IAzndk6ihACguJ7TtmleKLxeSRiea4AYpn
Mrfu4cZ1C7vt5kP6ag0gNoeD67ljVeajDFNYT+g0ra1m9sZdD+ZBatXnx3tC9+pvx+1kutW2gSDo
qUOQLSSmLZ3Ljc/scMonfclBBfE4Me1JoilSO9rFQ1PHEROrX0MeUg9wOrHYp4163mhdFyTUYbhY
LAfQtH3qLn6FLcH1w2cxHBiL7QruBb6wS11FgfWaDCn2xripFaEhFwqplWsleHoazDYJNj7/Z4eW
6+KA97Y7Jn7gWYV5KLUpBuB9JCt6Tc155Unjzm+MBtMhAvw/hNWfBHQ9GhEEL0/IwjGM2tgONUON
ULa0oa1UwY0QTNLn21oMfHTe6t8y/dHjtQcHvWTrgEe+JDclqOrI+kTl404wnZAncYj59jiJd5Fu
jSWgfsrwBeFttfa2rNl7WN3yYdPLB/Teoi8mmoINIteIJY9MhT4c8fo5G7gA71accp1no+y+2jqP
9Q0TYgHr2+fA0QelU0aymtdARIFSlNVXXcwBcsK0bQMq19HFWIkCwWm1+AYU8pIL9U3qm92u0jN4
weEy8mCYgaBhbgAVlJlLQ+8XFm9MfbbHXWMJn1zuFUjkTTzI8fD2k/K/lcD0x8Cj7Y09OZrTcjJb
OS1UerQIMaw5K8PLJM+k3VRBUEOr7Dkstz6/gVQCNkLK222axTOfSVT1DK8DbtF5u0isrFElORQ8
xEFrsbxpKjB6qHcEVjiM8UtiX+mEof277FLJIoJs3QmxSCJMb8ELe4odHZBNG+4CcQRhChlW8JfQ
3khYwCLTWaGZsepjdRmKhQdc4llbXzwihb0Gm10LKop6+SUIZwJMYeTnSo3ci8cFkBSnGwdymxnk
vH58ZeNKYIVMj1Os7+LOnSfwcUetytq4EQj95/NZlBVDzArnLOsshojIDn1D46D8lefRQq9zuTgI
jJBLWOBh+OKVmiSfQSDhDGhKKOpdLYdCiyg44EOwj2qtWV9UeVNS9LBuIGG8IR153bknAKxIlRps
QjcmwKFwD/im0g/XPWqGN5Wcsp8Yla8bWWo6dRXPTrSLxJ9nD5spNhuLnuUg8AIxzIALFG99krqV
YPFpPuUZ+9n3CG4xkw99zF9ftGHnqA3ZxVWZiZCSYaHRxR2jieeTY1PYRrYQBh1MAwiBX14Tr2pr
NRpEnp8KdPS8FvVuTiVgahB1X+amklKIw12KWe4bLHB5d3cGfNspI8UVlgdc/6fbLZpAWnFu9WoX
pHjtb4tnGrCBpgrPLaaL8Wsxp1EE92UlKfL1bhepyqcJ5ErUtKY1d7dg2GX8MCHAk3ZM/VFENZD7
JPc/uCmgMyP76jFK4/ZJGIELKBZa3cE/v3530cWFJZ3FhLiEDEM0gpLG7WYA82Q6GsD3eQTVdFbX
xFSQUL5bTOEigsMyV5qEy9AHsF0N/c+/+Gaag/d88uTd1NwAmsrmz8yeNMESkvbUCwq3EGeUyHFT
sVhW+bU/BHGAZ/Bf7HbTUyHiO0QXQJRpCg/doPfSfLc8KRxENPl8r81Hjkod4fcXXAGyyb5Ek49x
cehuQUeuN4eNUoXNuqpACH861EZqKtaGD9gUqt9b6NxywFFpumi5zyZ2Eig/hDxu6vPeEzyS4SEt
qkkjAdGqzADGqqHsFE/e1lBAhOb7PQ67zj5varL3DjqsRQAI+jAyBcOQgZsFvC2+UYmlfkia+ZEf
SPbVOkqtk7F+2T/J5sS6anbRktdn05jm79CFMFfP68w2Kd1L0avjPn7XlUrOwTgOHOvfE9fPWP+b
/QcvU1BGSMs+MRv0KkFuou4g8omQIjpJJ6tQJnFOBSXHofKrFuR5hPSX4nHI2RO7lotkTC24DYk+
x/2/0sd8eYi8//i7jF1wwWAHGwva1hNKO/7fyeWNfdApAQtPMseCbBTl2Z7O1GM+Si8JDOyrsPJ+
jDntpgT0r6xG6ZM48+y28L4V7oaE+iDgPNJx5WDGXD+t+Itrgdj2CRFM9kwfqujrg6R+jw0f9Xhk
03A07/y7NdbCnUi7+FGqhgjZaJc5DJUECJq0RDPPd1p9EQiKYbC4GJ/uWanfO1/75XC9plX79RR5
Dgry9bBj4dtNA/gYAEQl+OUlSraJGiB8t3jPKHA3gwVmyUhTRldnPhpQWDLevkW9OQmv/5I5lnYq
0bbZN7LqPGoJA6uXimbj+pULiBLt6NGmOc0HlzdldU4fJf2X6yQFi8iWM3QgC3xw91XhL9oOKllk
dZp81fkeZvvEtDn7cErXjCR8/jcBcag3E/XaMFYQ7MoUDTLxGP6z4yi2aFqqwxPKjCG8LVyB+zJC
fT6TYuJUfj//Ndq7TcMQQsQviJEHm+F5AKGtt0zLHMREXUOKsavelZ7r15IrW1iG5pRQtPCMwIW8
vPofghYu6pfAptwMFirOuOekHxrgAGStGWEh4DZ8aeGKkhl4+vBJ8LmSt1HFJStLE0y3nuDZOXHp
arE7YR/Le2v6gOQIVP13jksbC8+tEFTdN+eTecFSetAGSv099rmWo861fPJhtSG9ZCqCSvgrh+Gh
IQL+R3ASsGplTyA4W2IGUhIYpOKifAMRrFRIy+iojQ+Fw+UNNCVzksyCbyrLhHFofnb9TQctt5Ye
3X+7e7fA7okydtvP+6iqOYgtI6llMlyXcGu5BUDMdGDN62wlOIEU3wvnPKwr49ld6KiBnR1bRxnm
nlOAw5vRUExWtfRsetqn/5jiJJaYqaw62jEOg8nEeaK2RoE2oAxJvYhhFGZWw1vnf0+ce4k/YXVb
tMg5f6E1ult30oqdT9Ehg2NcozUCVOmBA+8fy5DV0pU+EsGtxoMFwzmfe47mwdC48KEWxNrFy9Wd
nDSMeXkAkg6rS7dyPRbo89Hmkg8A1T36EDRD9s0FBaeiGLwWmTC3cvWeCKlVvx6/4lXhFz11VTwU
AtQJAiyht0W3vd4KcQclVXpn2GlGzdxbvrJFWoQVPXn4SJIKZ4vpFA7vaR0jh+yPQiXnMoQH4zVs
F4RJ5dkI1hSiDTKAqO9xC+Ff0qD47jk9Q56ysTP21858944TPAePs+Jj86505JGkKFx5BYoLwpOs
PVOI7au+DlkJpaGbTZvMqyk44QLwH9Kxj/ZD5gPE98Znz+jRRk8isqd6/zYQ4fC9lkFg4QZLYfSE
oqinGLXQxiAlTaWbmu5rkxaHumpXYzD0Ovqe15+MMFWyqK7bEO7bSFEjUXJ+i3PGpnE1Aw6CZaPJ
JcFUn0DUuh77BJadrjiMIkIBK6KmF/fQ24u52a9rwPEtIl3fa5G9Tj5izM/T7reCKts/y4cvOsmr
pp7REW/O+tBKM8O88hNCJnNb7b/FN+txCJGBXPzJzyeXog912BX8zvMG/kpuMkJMegraZa61HIA7
w3w1bOi/X6x1d/gMu6Dc3D16rYvqtXwZUkUJIg4dRWNCJPxsvHlqW6W0KZflOcwlLO+TJUrh27Ls
wm2YdiikLZRPGHgUIvfY/pzdLoE4Y7GSBYBQQeRrZ1S18rjgTKjIZbRO2LAStraHZUjjyUxP0QPv
FY65RoDYzVgIVnPsDL/iD083i17TjX1KwbRg2dKZvzxPGtJE4XvtAZJ/X7rcdvHUTF1LhP+agnea
V3L0pTM+T9j4OEztkAMHy+Y085Orq11wHruNR57o3LTy7WJ0YcTUJFAigXI/Iha9i4on64UOqHoG
waNFkPMTRMa5vQygdPbHpbu+FXT7WHVAQRF57yViXVUkccQVYx+IW2XWkuKIQ494EKXyi5evzB4L
6f+DyTPV7hpBaqbi+fz1Mlu1SHS0uErnjKEhwRpXYxDoHmWeyjaMt+OHQmU2Bm4/Uyv//vvYeQsG
qUfYIJKuA5k8qZ5P53XXYGoW1jFiDOFpLqbBMuUAAAClEjnaWcrskS005B6kBN8SX4wuIUwzrh3d
yz1UQVB5UKsgL1Hlhl8S5My3Ejw3F0hLl2Ji4H/SWJWyKLdPxphMu5bc95O0ikj15a8L0rmN89VM
85a8XIg33cU9e+/oj30fPPWeniMDgWCHmtkkwxxqHDRp+g5OJEhlHc0f0xN3jBXvAM9mu2r69ylM
n7d3gkOVZvDP3zohGrxKgd9briVopmqaKrFEAO2l5Cez3AD7OdlbdBjjz5bAp3Eh9Cr1krxPrLAH
NjiOhS1Ip4KrHrAkP+90QxXA6ddjnbvZvwjwVZRNBBDNi6FJRX0dl4Ry47UpIMAcxfRK7d+YahOe
wnxgHNsyDR/E+oukvucHUuftPqiTb+ctHzg/0fD25daxhjY4udv5Ermz/k8T3AF4ei0yrhTO/w5B
Y+O8FqScjqkTrLZcUHBmkoo+17lf3fD7fpQ9ab5JKYvOMgZOlfsRGlI8kqpVxjPayhZexJzPLe6n
x1xn8JjALtwIrSrWCYMnCYGAEH+zNGmjppQr7gXX7S9kGs3CyQnfR923EeOekA+W9gb/vd5qRfZt
Def31fECuZtu2gBl9TinXITvf+Xfd7H5WCLWKAyW3hlupI6MsQdZ0eWozDxvnPlY2gimMmnHNRtk
6ZZT9D1AkWmOypYVvrfUp8S8EAolvVYffXPk08bLzzzO/wt5ojDDUh51/emS2izOLI16Dmzv0y2J
BAeWnPDZtcNhDllhd/eryTrB88gRlQ1ekIYUvlxPZp1WRlm4PXlslt/ZBWgQ6DgVjhTAC81IQ95y
u6Poex87xViU0aW+a4y4jLbpNZoUQn1z2HikknHdElB9UNqz3Z4SxWmWsZ69VcJh0QJfSfjimz38
xdMZoNwTQ6xmFj+W31NDzNsNwm4X3F+MX9bS/hW7XGymji6Kv5QqMYxSBB3WF/UrYEyyxL1TaAuE
Q/cUKHXvcPWcghceDtdjZxSERUpaFHCKpmV0MS6eM5arMqw+8y3S86b+UyW3FL/MrLKJ4dBEL+WK
yUi4Mi+OonSGAusms9OpxUKt1+ttz8j3c/e7jx67g3oIzbvuI8R4yjLAkoKGr3STdPp/LNrHL372
79RDZynyreetbnXIPrtJ0K8tzJuQc/rNYnkYlucRUa9R71ww8BdkxJvdFMc4fVbKDcEsDW3kaIa+
nHGs5lhGplAHHC9fl0rKkOICmSVWpk2SRXRwe87nESkS+trlykSkM90jacfp/A3k8cH7zc0m3EC8
giY3OLd4vpWIizcCV581Fs59OmtoWV7C+2vBXqHeqEOTrOIF6F1MPI0rvNCSRp7/S6u5RnK/aSHw
LnPjk0nys2zndfN8iLZ5hIiDQaos1IZ/TGwstQ2WvSH1O65j7ptE5b9DyzycyG0Cnw+uxqT6eYDd
YQ55Az6BSJ6NvdTN/n8PNGoO+wTHTzYB+EuWrH3wVLHc9AmXyIIWEALW5ALWlCHE0FcmdzxGn1tJ
JH+4Eb4eEgi2BPAENj7D3WNgvOhXPwjLQegb/3k2bFgsUECcaPKCh8hNVbv0Rs9o8TxeEDaJUE4a
CosGz0CjQgz3dGTWAKg1xNkfx4ic3L2KqGSYEU9Ry+SFU9OCCH84X1ilphijj1ihJrWQ2ZzH6Cc/
KilC42TvhToKNWNh/gCmmqO2jxIqXo/joID+/K045BNgvqTJJEXuNqZgqfr00LE6g7l9pvQMTkP8
T0SixoWkavyyzmIxcsm+hpcPpZsmOdi2go+qJIG3x0IFODnW3SNJGCROBZcS+KSHadWBFAqn5am0
U7deksRWVFBiukxtEWTjpdDSMwbuGz3SizzCCIR/CmwJBDpvCrfBG1Kle5qUUs5iVORTgRv+w0zm
T+owcs+3XHImutg+ghX5h7nyXlGyq+n2jZUBtRjfZav03spz4xVEpKJQrlbG0YJ6yd7H4YKFm65i
Gnzzr8wVbmKe9uSdLEA2vXwggYR/YUzcL2KU98TeNp/c7VuTQUHnv6aU4MXEn090GILTX8Sp1hKR
Z20SF9djYh5t3Bu1efDddyaK7K3RKm5A70b2esDSi4KTf21ZfqW2QG+tziI/mjZsh/yGbzow555g
0z432SWuCTUOHdWcQWAHYNvbp9F7ISman/nZ8b3vl9PCStXusTLD+Sw6gbS4dZT+Ak4VfP/FnRXK
s7Db9QKeKk6T8wNSmqqYL9pPUiH0bHL8prRy2blYv2sMzHIwLVSgBEoBhjo0x1XsGqyrAAUAPWRI
eQ1BMhhCHo3fAdo1c9igXLodwiHrEwux/p4M+KSVCvMcHgpiUNzWAPrvEpsoTOM30fqNpDPf8upN
8UG8VQSZPzdGLICtBaL8oCCBs3F1Me7HRx7T/S5VQ2PDhxBPj/zzOZJgg4APdIMB7z3x508sxsLr
KMQ52RBVS3IniYsyEM/jxokckWb4qfWr8btCxA1hB4kATQjskoZG3IzqAdZ4UZECajFYQDCGAhh7
g/09if+X1tsdHNyxKchPexYyZ0EwDveISANQXeZAweSdmpXTwUMls5QMgMbbCJ9NiIlz85ewzZDM
Kz6iKNZT1/SlFXRjfwvCodhEuOGCJWX3NwGv+VO8iIRsyZyJYESxVbQT5wT6WRIcaPw4TmPNCG+g
BMXpcRyxS1S6Yyhm3jaQscr0xLvLjHuNCdfk3Lxm0w+ieP+iLv84+d15uM1spO4ca4zmu92Ly9HJ
rYQ86R5sm+/N9V2dOfrtXCmw1JJdzfSDu7WtRmxkd+wMOd4hFFbpGwtmH+hjtDIPNJ6bDCTjFmTc
qcb/eWcASHC40QgWs4A3Ic3sD591YCTpJa4qoKoL5lYGNlnQLaK5Kdx+LnNsdwdWoGr4AHJndSRX
BYXmGEcZOgKGUjFgzqbIAVb7XRN35Ewf5VLURsBotS59hbAHCLeSiVvP90JkcWWcxBepnE0Qy9Mb
UR0Ya95BmZ7TfdXGKukWiJ4WwQfnEhXKuxy0J0H6APOEPYDrMgBMU97xq+wygOR2fKK9sLVNhuWa
7RTP1Q8bZIE4Ro5P8mEsFoMUuvMlW0aVhOlmYMNDlxzSuEjc/tljLI0cKy/j9uuiQXcv31xlMHAL
bp4uwNFNYIcUTLRgsGBJ+QS7P/CqsesYahI2g9ua7zzOlQhsY8WvWamS9fZcWQ534wYaglH5PBrf
yN5+RruEjNDFCSSiwQ25vMOOYEILtTg4MhP4OOKjvT8w6JBYPhAExvyhx3mJfc0MRAV1oASy44Aj
n/SEfCOcCM2Rrn2TvTMcry4DN05L/qCcj8GUchMAA1PxCgK3dns+gIOsVftlHCnT1XHFfwjJyV7+
f2BzCGKXAdM+WnY3wRbCY43qJjW9sMgzyAYEB/hX4caham/vyAGkv5JJwOjQRA8naNkymA3XLFSm
QN5eKKHHfd81ILe6qxZpH7BUa7gooUeLgMexAGnZUwKRHpvtrF13b+i+W60vlX2UXN06gi1DRAf6
KlssYpeEL5rETMRPHWYCrjHJeMT1HWBSSItN0r1TcrlF91EteS1Ee0OP8T1f6zyEC0Pjl7ggfJFr
mKllDSjRXGFgmOP/wRGcy9C3ffs7pn+6BI3RQVKiuIG3t4+J8Eld+t4PBmTN4mZSA5bC7XYBhAke
lxwMTBZLKIdsPhptmTik/i/Ce4UIc6hRNW10Gp/KvHIH1FD6AZwilb7sMCnHy5pcQ0IF2U7YTxxt
D3hePYLgmRGY+GfPHdFNIGhWLLXdA0NIwZfVcZn4DTTf8xBOlhtlSO9cgVOnR+ew+eb6YTVtVRiP
NS1bzN7mqE19jSQJbk40Ad5iD5tRuPNRz16gtJtjx4OJR4mi1c8ASgEYz9Qk+oEd1DTR9oSmR0Xd
ZuQlSGHVw3lLo8ww3OIraNOHkdoSmSWk6BVqB4azV6n1gIbq67MBh3guGW1mszHSJg+DHX5Q2GoV
3GVKspv4eU41Wpb42jGUARf90dS8WboSFOBLXhqx+sbZyPKulWuUWpeOXGMnnzpWyqyiVjE+TDMI
i2h7CAgYeh4lDiOusvrccpdgqM8itk/rYcS6hJsfidI0rrNAFvHBm71CTdlQK0aEBDi4sVMZEvv8
KVsOfYYFcYXW/AxxI1xyEV9SgymyenO1P2aslwek3p/0KFwwJGuqf+2BLEh4AZnrsZAUaVcRP0ro
absM5YxPoANjn8bPiPxytD0tmD4DM2WcDgLzZPTP6I2F2hDfkxAP8zLI9RG5q72biSArq9UlZdKM
H2+VPpvf6m9jgej+CXjq2BPl/HXN9CT1z210gQ7xcTc2PGEuM07gJQSJkqpiVuWd1NX2kHXbNWxt
QKYBNLhh+8KCPjWj0d/YP8/Ccd/JT4t4AamCfQ3H6iVb/iz5ADjIJW3xYgkTUJmmCia+ZTCpSVud
MJU6ExmL4wRoP8Xq4UsXaxJzD8G3AeHoEiDXMcb5SOJxwKwN7ujO8Db28ixmGtm94Snduz+Tk95W
1S1FhztZGOzQMbprNnrv8Rfxs8MB9eHvpYcKhGueZoS7Pb18s39iXc5QAzW/S/R8hXVjBEEySk7L
c3nUEgQzqkBnOaoLQcP6JxiLGH1c+MLaVlkulu2u4m3gglzcEp2l0OlIb82FzDMhyJ+Qr0gI4C/U
JzGldihPtEHHj94x5qulz3wj3o3Ay1RmpO7Vc9G7D4k6wG5RvZQ3Gd9xHCa0C9HY3wdlDq9sDuB4
sUnkH6BSx08LCAVqVJr8TfEy+pCfXOg3EiizFkz2Gjl05WZ/gssJXFunDmYQdaKTJUXDPKjTRjOP
2bDD16/ZzcC7pzjhTVTGSrDFcQjzUuMndgIDlwSuGJDkYFLiYeqHjGrgUw5l/NXbjlUlHcwsukQb
+Yk7bR6w4uMT7PouYNxqPEM7Iv3KTS9zvqD9BBFW90YX1TcmBHfcmTPZjDJdetPYVi3r/Mtf9eOT
PJqOHi8za0+sd1ct4B5L8HBFluH4ruRpmvi33/ioF8a6Qf7VT22YQ2fHAx9d4kRd2u1Uu2LwKmlF
9TVmWDaIgvIfkinyfMUzrGLkU4Pv2fZYuCwMZJ2UePOIpzEon8TqUitXA+cVJnWWgVBDm9/sgUIN
L5lP8XqvWVDBw2QAmx+jGbhz1hxBS0aGwQ5IrwDDJSKxoEOYumYzIjZdBoCgQNcwq6Mn8hD7BExI
IusCvJCCWB/3iplAMTm1sbtJlg78PTNnq8y1FvcKCbsFkUDTBqW6L7WejdPCyYXNQSID+zH28uxn
jlmnL91DfOAp3xmnWz5vnkkhdWnkJ/H9R3yJDOi+itEdhPXQPjUvBiTD/S0nx6el85zjCwFX2p2Z
DFwskIv0CY8zxgbReDO74rA45o1cWrIngNMAjK4uncos9O1zXc/KzKhhu3/EBmwVxdxiW5elRpMB
9VQWmJJM6MS2+W7MkghN8VhlXqGUK84YyUVCMTan+rY2uTy7n6jZdDLp+ZOtxTW2i9AzOOnOg+aZ
+eizWLrNymaSEtpPksmyW9qmHPrxPIcgcuTo4Ll62a6xd1Ue29CyywsrR1KSJQ9F+/R+6ex/OHY5
UbQmnVa9GljM2k0nTK6UF1wmdINDMKFneI2JUF2wqUUDlEBdTEAZXw77txq83hZcOE9l9UmFi5FD
YRC3cLGnGpP6bnqSqM5nw4goanH/O6a4Zr5hdtP1oBO0C/CLcgzE2R7BDDtubCS6bDFVqBkWyihi
L7HRFYYvFzTbhvJVZ1L2UvKsAwk7bGsmYI8eZNq6t3kQZwE0UEHcWxhwdxAslk32jRGU0LU7KQbO
B26zqEqehlTSLMq8u9bGbUZ96resGpqBRGjRssGbVtPAh6g2jhkQEEUdWBPDcE3bdOrreXqshqmb
yZhap6/CbVApw9PfyNJtczew+tmbfXPpNvMgQ36L/JLYNVrNaI+iQvM+2L+B7++zdXiRvOttGaPT
4HQ0d0aER2BorpUk7LBmh2NOqsWe69NOSIFjXusTPYG7W06GHpYp6QjoMQMTQEWYtBtvFM9x1qHR
ftYp/Hfu194DlChYwLRiLN1gLAGyHOi/5TELXiUziCZHxNdgiPfyv/r1ChiBFzpx162JZp1WsRQM
Pc24EY2xfIWjtlhxEZ/+i7e26tzxEOVvm5p2qqZa3ryI1f8atONFgREUEva48d9KP0oqNe+dB8Ow
gIQfkPjFLb4FOGR+zRRlpsS8ZxSJe4iJwZ5Lf81wKwAU8JBPvNT3WD715TKQ7YPHQP7lTwSTaoco
UB+adZGPIahzujc0HCl+OECC5SP77MgtKMwGLq6+q8ulOFzEZo5e0hT1al+orl8OO5H10wjGo2Ic
P5isexlzyp6ID58LLP3Ck7BzMiDyZvm/EEOxr5REvAQIUSuelLjrw42v7yBFwmtpB8ZSBQ+roDBd
aOTV1Sj53Nat1uiCXqdy56XRIjdz1WvuLylNnl7B7yDlwkyUIEranx9cQtJTiQwFmrxW/Koeb11x
XXDuJPCRXwCOABu2YOE6RRvqgPfjc0f84GmTMrjLmOR38+vKVTjODq03jOnp/Z86rQXxMDF1plVR
Xfrwp1nA4GpvizFC3SJDram2EziQ8KKZa3n2tHlHEKAab+DGRIwRrrad4/mjg0Xl0Kb9Eu7hfoUz
FwY43BCYIL0GJsFoAoyFBYSIJnwP5btybPJj7f/EqkCzxYLqqexuvaBo4Vj2ACpTqGWCFQGX949x
ob38QzU0ZF9kQprDd930xagPv9DwmjM1RSiWOCERUgVAgB8OfleunQ3ynX/vWaA3TRb6BLlfDW4t
BkgY0I8YG2RZjTxJmWPm8aQKlO3Sphk9W7lb8ToulgC/1tmFFKuhmuXrCbEy7Cdpby/9rqexK75E
qiYeY81Wf6FpihDVNvydEmgcxkew8SMg306o+Nb34mCM69MI2paH1OhSRuKFTeR4rNyT2Hw5jX6s
9vtCK/9g7Yh/4gY58cNnt0/KTksm07YZGZmuO92x1u5N7JDQgAbVaI05OqJB2J1OivMFBxFYeITs
Ec1aD3KLbbTB0oWWa/tgQPx5OptBPJ7ThWJ3eCFq6+OB8LV/oAgftwlcQfVnDYHPTz7JMkL/dWEv
SSRl1lm20gC+kF2/g0YOdmUyQcYBPp3pxDLdgvGpRCmP7TLuiDN1NqB5wfHN1oY9o1063fxSDobG
KPjLzncK++3tjvUPEYiCyIk7gaLLJMOK682rxUpYh2ze6NkT7UNDetkfctr2bLi+zn3UIYiUibbX
4sfKJ2uur90M7BbSio44BAE5hSdLmhGqSAtqoa3gcOPDfBgL42JKWgAKU/GQRX2MAasNvsMTihJK
zecNLCUPlN7p1FrBbZ4uK+1o/UTUJ/CmUU6yGyxV+J0iEn6INppzY01zQ0vvF5ny0Sg2SR6anqm5
omRFDJr1mwbbhLTzJ7XxLJfIS3Nq67I8JiMnwHmkq5eEzB+y3PhTAtEpRy8qcVuD0sN0tFLEfPlj
HfL+MuszmbrGe78S87yvTmHz1o2QmVPebnQEGMIHjOFjxJmn9Wx/8/ryb9K7YRX7axDQFumqni9y
Icw051osHi/cw1Tz/HwC4k16fMCWwur1ai7rxZKDXaR8pWq3pb/BqFHNHBSNIbjkYslkq9ytbMgW
mRXdua7bGXvDqcmJRhkUYuJS0Z1zAseUGzfy2uh0noHWBLy2/TuUIvF4yYa5AnM9ml2L7QKPLIqv
4F6t8lClNp6GnxEpAquEtjPamBWBNwDDjzUgQHDBn3y2wRGkWEw+89FfFG45pZ+LFMdBm47IV6vZ
KqyMBiJzC2ASoG4GyjbDWOyDFjOdH8jcqYOHB7ChKPN8iIwQS4b3I89F4lZe3QlJz+FcA7WmPhjC
B8QGISduT2DWkQmofYyPle3emo0Ria4fwfh42u0oP2BDRT1mWxHmgynNV2ydB91WxDCe4JqVuLW3
U49SEsk+6RZtwGF+8zJ4GX7wgxPSUisYgHiVewtZkEGOUicFuriIpATXaGRs0QCK4k3z1ypb2JVs
WiR/udIl4OnWzZtLHHaeLsOYpLmrlLA0d67SqQ54hJWAWnMOEEV85u8h6fQn8cUhl/1oW59zXtQL
PY0aMgxxamN1W5l6JVIecsrHXHUrEzxaOlWHdDzFSE9jP4EVmUMPGdJTYgrLhabG2Er+lXEw7C6M
GJnvS+svM4RuOOxlUciaSb+mUjr6S7GshQR+UpFO2ofcb4jPnfaFLnUasWlaut+xxu34boL5XmPU
dCW0DPvaQxjEtLAC8jJe19IUrAQ8k8/y9onZ7JnPzjSSAritHBaMU4un7CMURpXfhIUV5j1g6miU
c6haAxz3RNwCkru1zFcwelGKW1px7r2msPQ5vJ3NJZ6PK8sy6td0dS/fN0QcFyfo+y3HSS3cevem
M4lCpmapW5ulp3TK/prZ64PQcVT1stBJbpbVx8y4Ot+0zs2CQKXG9OsrO/nX9mwvH4GPpMkVn1Ub
5rofP2U+n8asIutAgnfma/eY4niwUdrnvAd0prGaZA1H/aw7SKG0hvY7hyxW+5Xe71/0stkGxBPq
VEEkw0Y35hytgj9p47ImHMD6kFDn5PrTuC0g+6W++mYnBcQq1AEumS/1lz9Mum0W3PUlf56TVkhP
/mmI5dH/33zXvDPcx+RG7eGE2tgP7OKJbcKYw/N7iJvNh8bJQKqWpJFZzTTUZQvn59uPZYi50Fjh
1TCMYuYPesVUP1GDMb550RvXKmbLOsd54PKGCAREte/VV8zJn0m93hU71wCgvKkFk53I/POYvrag
ufmJs1yXNIWP9eTU+vDCFkQXe4qPx2bLiFCeQO2JnbQwmD2EvYp+TXLx007WPGjG6bMBF0pOoNvk
Sn2q3/PJjqKzNs6hYO7zmC2CAexa8tqycex9FCRtSiGG6E7ZUZ9IY7ndeZcydxxyL9IaeoF96bKr
FY2KF0BQE4OzoALH4kP+jcGnGLzI0lPPa6KBlZwdBF/unBiPS3L0APtUkN4KSHNpOi97YqNN2xF+
y2gnfTKSoTKkVer12Qp9vJbnFSl4PsBM/KRF8vee2bsAbR3sc0G17bo5MmjKIMuADXwgGQP/AzgE
khTwmsYg5aEHr5Rv1Uq9J0qMLxVyxXlYMjqJVwXIABiyuE6AdjWItWV+SsntmcLNO47MQJgk8QSM
+Omvr7KHTBs53LUL9x5eGhenrerN0bZATje2ZNs6xGMRxASKXJ3EXrrsj98DZPhFdS1vcimk2WYO
jng3OVlKv+K4bwVJmB64NS2sutcN09sQnUyJJkRcZ9E3exzlG+u1Ba9toGCkmaFBljUL+A2yeJC1
JiaqMdpWWZDbZ+4hbT3OunaGcamDxSz9qV3eVliIzdetxejQk30JzMpWW/YXoEToAVS6b7M8dq/d
uW7akT2CGD1pDD3wSvQ16cKs/EBTyEeZHbrc7/55wV2HdeAcU10ylIPbW546z27KFW2sIdxYgrQN
lHXXZOxMuGAef6BBY3D/J3DywytrIq61coSSWuPCUJriwhca6MggnSySOXm/Ru/U+t7Wh+8OoCk9
PuaVdiVFxn66AXvTfPwpPG7soqLyRKWTZUiIYWd2BEP9bQO5nzQQc/QoN8eoETzwbkifUGCc+cbo
WF07vfloN4+O8W4nbEs/koHO9lFqayRGpnNAzkX6XC8eS55vmDyUq20tX0pnD0pi4Yp5djPBHY1c
IyrGQ+/3wCAqsRndG/UKQRypQaNR4oT0uxezp1VuM0GXnbsCSZAwkOUyLDMEgAtazZppY5Is7cct
i+ExCyyhDRRd+7nYz7dqaG3pESsUzN1k86SgVEnPlkgvLZTDuzUbkAMJ4kOcp5IqykdJc0EsIn9e
SoTwZWZme0DyZea/6TxwJjrB+cNvil/nsAITMhw86ihSHNDwX+J3TTh8zJlOzn7eB3lQmuGA+Kpw
UQ+Y5Aar9swvNLnqv/fLpk1gIrFlbNLF3Guwr5xmBWIM552Lp0rbWULmO+O//5zHwxjR4zBGRAqi
dEtqRiiYWlpcUjAh0hzH52tWWQK3L37OS4tXd0FP+5hJ9vLNtFwqRbqqU5tsfoJUzVT7S/hCTllG
5nTa4r8PWWOyjWNQRD9B1b7AB6YZQCTr4t4N4miWRXQe46MrKAW3HyQ4KhSnZZycHwsSGJ3gRTSb
iTaQgw7j73GVrhBexgdDGKcLyTg34lW1ksHnM6Oc7nEhJge4R4S6kgyAssNRgeHUfwonCKmLov9x
pLmCWqkUC4fn8NXFKRh+vwt20aRvGXKe8jzCWTWxtf+XGEJQEPan6Ev1c2VrKTvn318NxAaQmOhr
YwbmCxETVSppEbONxe+lGa2yb8wpDwhDyMsVaxXnvRKBTrqZXsEJ0/8QkjweFGoUtTK9r7/SeiK5
KuqtXxJwQT758uBnNqP1b9CwuEzZxPx4VIu0ejtkTi/B5aJCxf/qp67t14+8dvsvDlqypBhvQHU6
/YvtrRawABMPLAEk1y8BHl9qbyswieov1ty7I4MVezRnIx8BnRjKvGNfx8HGaFuzM2yFZrTbuUMR
4G3/dy3nIL8qLaq93Fe4tZlth4ssQ/+ywVsuz9JoYWVxCIiAcx6A2PdPPPxSFoFnBKUffuNuFwzY
YU9XNdaxi2l3jx5yiYApP7q+qMnYZeB1pXsE3edYpLGNeXfUHgnjyPGgVoVT7ZQkwoDHUVkFhyvI
lEyJ0iK2Ne3Jq8aGsMAtFmgOMzT5qQ+1L06iSu72e+HNwYnKszhLEIQXEcZVkItDBgJK+RPJAPFh
b02tSHWMylAzJgyJPIgATK+sUUh8bTrG4fa472aet6G8pXW6KNQ8EOyIJ1E1REd8oXcDgSGE2jSE
foWVnUd4AkAv1dQReR3rTVdfWjVuxyOorEDO4qIaulqIJqiMbASZ8QV8YxY7TBArIU9BjHndnwwp
bU/hB9QzCgawV9XLsbFP+OU3d1Czd1+IokXv4TUL2aKn96IAUzOgY/V20bAFXUYn4pMn4Ss1/pWK
+33m9hlTA+ZjGwvSlCzJ4YGf44Xo0ryw6YZt0yKZ4thsE6N8mlZ9YH/pq22NOWF/LYvc93dYo1wd
m3KlXR5FTHtoqSgabUTpFRVslF1qA18kMcgaTkxtvjwpXkWlczXzDYhjT0VDvB5Z0WphejgYBJoH
Mhkeekk9oori2IsHUqerDPNsQR7/h9xIw/Ppp+OJGiA6FPGrS8tThfqqplm0PGbBinQQrRdzKMU5
GVmFzz8kTt8yUcHFB/ZHhS3k6lPqwT0A0lP9L359CMjo5yDDjejhtk7HJTbA//oTYxtcr0zguOrE
ooQSwDBqQPOU0nXFrp2r7uXWy17uL0hItpC9/ZY7zXoKFlxVblcUi2/gF2viWIuHfNiugWIe6BBz
9eEWOJ6ruen326dPGtHYXgWmfrZpIfssTEO2pIrCZGXaxXWdmiofrbXQRuZr8dIaaxHDpGYjD9gN
hcx2A7uMjGlQ8xD5kYBYKc4K/w2SVp2zKQ1hXc3MlU19PFRiqUP2xBzy+3XEf0UMScnL1S2IUJP/
UgRga4WOSntWFNhSuyCX1d+hu4/575tGrSDml0clkV5b9CkhiACw+RzQTjcqgfwrTYOXy6YJl1of
ODx2UfoBi7sm/P4IWBYx60f69W7kxhFyTLIDt8nGI7iHJdlPrx/A7iUKjBSdgWftKYKFqjE89SKp
yoVR+VwbjbNDq/oMmLXHg++1iPqfyfpZtvABtZX5gN3Ju7MzagXS1trAPV8kUrPbYvCS08lsmzON
zu4IO9W5jDztEZECvb68A1iBRJ/xxEqPGc7y3s4Gm3oPFNzEyVrhmyO4YjHeRapQl5w54UU+eK3t
1hP5Xb5EbgmeNDy2nCF3euqyeB5krcWr3CQm5Qe1MUByNoxMGVwxww73v8+7w0fj02n92TI2kDt+
udEJAcefNdGYnZuhUNithLaC4X1IOX4b/5C5KSchJ78boWT+ELbVPQ1akdA+1eK8jGpJT8nenES9
7zK7DiDCmZyemQOQNlhv2hoMgbwxIecVoyw6K0DnUhXu9XomPeq8ejM/bURFUqpUQFRrb4pGXZFk
shVT8acraWZJfsgEpvHJx3gqYDW4Qd0IdXhWMDNiidPsVXRk3Rf/0+gfkyH16nQzarTBJvZybE/l
rvxr7V6HiOufw0PqRxy2RLHqQePnchOCDjPVe3h4wc7zHaSH+e3ht0RM5MRlst+mRx5xM3NAlUEb
ao/3G9m0gXVaCNoHG3LfSz1PWjenywOQpFBCp9aPqLV/yCKgRmESKaR05RDSLtC/avBmTg57pETK
K5WO3KdIh9ZqjQqk6SE9dtuELvhKhtLWnOdE8bIgiTVRzQmg6cRMDwNFW7mjVruTDbMVW3bXDVdW
9tg/KRxxfUUUOM0iJnM6uYhTvOGsJRl1wYaOzfTXfBG80R5zxT/eye/es9a6iYBpfxSo0/KIg6Ny
eUuqY/KUIORgD59fucrUuLtVelzHwnKtlVLA4PQWJ8xkKErrvIfwK4QgghvwODzlDWEaPh/ovc/a
IhwCFMCH38t1wQSzUJaWn5kzoyHp4wF63VvvsPLmNPpMbz9LGRZ7Uu1on6QSCPvIaAUYVrWnMwTc
k8D9hZF5a/sKPiv2Mn/rMlSPlpH3Jx7pkfdXqE66muJmv7DoAcJnnFN2lWVZbxK3tk1f3RKyvOBI
Nmrm0ylY1jTs8bySf9Kjkhow6eY/UP8WwSp4Gt0UP1x65lKU6XjKxUhpjYjN0cIQuoOozU1FlRjR
2aU7qSSqkB5oGyzakMRknCi6wY0ndiJvvpWMqdCCnHNhqh54tRaYO62swcsU+G6zKTuIbXMW1dLd
cJv8ArbeAWEVkKJmSc23nvDX4aubqKCYKB94If1fO5Zknt3t18goU7KbW0NYDyF1d+v8Y7xfvt+Q
nPd+4+BofShnUFq8C3U1ZeXkbyXNzquPoKfRRmj6Bc8XikIBwr2nxFsV2nAndn6t4+g9WO8QZz/z
lNF7X1DdFPXNLDkRRwnIpERhQ4K0NL5/Y4mubOrDKwOCpQafj3Z3Mpcm46/Vl7h8L32f7X7VjuFd
piU2STDA16r2sHY1CAknOQ/SD7OKS9bfBU7nCn0Q5Gq4JFzpYCKHOd3SCku8kRn6wxV0XzTAQWhy
SlcpmkkToc7NoRo7k8o3SC+p9sCMvR2IfA144Wy8i/cnkLdyYM6on6bl2mAy5RgjMRZqSv5fZWQg
2c80OPaPvIeuy856k/czcxv1gdA0ogcNaXzE8tE95qwvEQPsewRPCs8CFYPIKG45eZxsQ7HmsV7j
BUeJJuYxoCUTXCjOHgALYsldynAsx4ZLtIObziyD6+HvwwGd9ZLl112rDU6KQHqHfnuNbhL8W0eF
JojAIGugCIUAyVa9/cDdS+okKPL3kUUWg3S5xje7HYQdejD68rdKbj1n7h3MySDIVPXOd/g1FHzT
ntEui+RAiwcto9cm+OtDv6h5RTK3pXDpnn6pZzSfqdWs+v4RqzD5BTI/+q6FpBbW4WpfxvONEyAe
N0tIOj9HT0RNZ0mB+Lxwa9Zj0KT+aMbi1z1X6CPM4dizYXAD6KkYi1tqScSeUVRQdKBOJ6PXeMOm
HtBccJOy0cp81kgq55M70u0ueGfXfBEQ89tmWN74onYKv5fmkNY/WUXPLCz5aUWQVhmiUvlXCCF3
VtXr2OW8PzabaTby2J5puUqTTFY/dG6F+b3pQQcUktc80LURXoIMjFfUAn163Nr+w2aLw3n38Hbl
JKV0ovoNGDjQt5X43Lv3YXyEmYKv1An/8OUWoWntvmlB7gPfA8K7Wepc5xEDVphHFL94VqRmje0W
ZGQuJFcnQ/yGzZET8VYUJrarUW0lHsR3qz8JY9oO7nUGnmAFbWwVnt9/j4SaMTnfgeOdQOoCZPCy
e1qnRHY19QJGCXMSvnogiLFELb8dSd/HihklSqOXFoOVpCgvw7VZwMlD3cnouT/gimDH+kvKUxfa
umVyt7hSTK7TM0gHial4BOhCXMJsT4s+AXBAkOMefJU5pNveftjuiJqFwAceIprAOm/LNM+9CnGd
9SPcq6IcaOxOzcO5NAms/x9bmLtx73AbbO4O6ewKffWE1fcXkOYPKJ6hKGDN5v+zOr4UoUlBvajq
Z92Cjc/QBj7VDfmdsqcaXBHHF7UfjaQwRPf/MzjjC++EhaBfdYTC55rXG+E5EzQPexx40QX38krH
8C/KUZmo8B2VmbQwzcTxnaUyfm7h85MXHrQYkHgMijspB2YWV9d527r6HJt6M8tjLSjzBRIY/gJo
pIhJbZNmBPvpV0sZyK1oQMwH7bcKZKV0ofx5K6cqfxOqdKLlexwkSEfFlNb6cbxokKHwaTOitOc1
qI85Tr+7rGHYld2LO9RBnCDe/EonkAfiRKdQ9illHS2i6pHwrkPQ8QXHtvamdz3bNqKsJ3rgxhxq
8vk0NdIhdxaVOLb22ST2nQPHtoF/hkXqZqDElZQEX9K9w4V0nC0WAlT4711qVGbxpEf6aqc31dbO
Umd5U83qf0Qi3zwb3A86fSn6ssP8bx7ARr1IZcnN+vMZ4uu27qBNYZwojYz8AywvCm5TlTMlAlyQ
RsRjepzkeiVR9tRq5q7l6EaoJlVXPZb7BY92n9JCwp9KYoYxDkPYJYbEJoh5L+47zeDUr1IQQhl/
+jGQAUsWYh9dWixQIwVfS2UkgJCDTiwIPOIHFNVWWCxkZ1HncrlMollZfU609xSHgZgecL4ALCXy
Wqu6lKu4OMp2PzQB7T/W/UrrUTOfzEiFWajDoGV/Wq+Uyeg/TBh4XPaoumXWMY+IREU+elos4jM9
2YapFI+a7yq/aRthWBdYienTVYhLanhl/AfudcbbVAwwB1DXxuxwPrNa0QehxipX8D03LA/zbQgf
xLFd2Tr4ek7MBXv+DoEEFwugHEyvUHq60EBVI6Zbx5dlUH0WBddYZ/MMqEypOdlkf4Ty/836xAdB
DXUN2k2eR/ZuBVY3oraWtTtx4vzpWF1jJMLW9cIxfx+C9RaRCopVJ6im10DONqkWKaeDpBnLwNLm
IN4LK91rbHm1zvSb+XALORVHcjalBIO/uO9FTYRpb6iHqfDiVq9zOce/7hW/BgZTccREuFV4N9U1
78adwPOT5Ow35EdSHE8sY/FNhf3iFf1zTomLeRsw+Jkf3klZ3Ap31OTOVVupU4P4SPTGiCTmX3K8
LUju7uPObfkK/AsB3333/HSetjODhCn5WFhvnCavHdPmDbu0u5dAG6DjGYKTz/N3nZd5kzJfmlLy
0cRdWMoNp+t1RH5AY+qpfFdhJ1WbLLfa4ugEbKOWWIaJcPWu3Gn4vxwpDsuwc3wJFEN3PQXM655u
XQewZId7NkXNQrWa1tN0jC71OrmeZlsOuyQhK4W0JxeH6alGcSGkdWluWC9K7qoZ75NNKApnczax
PSgBmhUMOG7CUfHTtTVxoSZnAw4PAGcsHahwDwg071VsFzto1bFK+eKUoxpQ10RY9iaYd0qOnydb
sKnhZPfcz+jgxkzU3a+rK0BlVlWETX+FlNmdPqj2vQEMsZ8mVzXRdNmYj/D16syzZzJ5ayw1TbYi
Cq+3W/NtKI0GdImYM0scVMXGgoaPuywzLFQ3Q324pxghD0mnmepB+TmTpELHHyDyB7P70u+KvgvP
+B3NGIoroukX+cbIPyx1RvQDX0f6dEcseIz16trIaZsGkWDcwTK2MfczPyTvpqvFiAmU9tbyyXMd
ohxgwT2eNFy0Lz3ws5UzRi9fQRfLXYP2V6cEsPcaSjzgjTxy0a5fcxI1wvEYL/YUKC3l52Ujnla/
fGIIKCeW79f0mJ/LW5f4sgo4bWKmYTvbqO3WPR+/mYVsBbApraJVD/8ez4srCa1xzfWCoWs+iGAo
3DuludX1kRHkoEOjsiqahUmJnUGHByUqtjZWrbAw8ZtgXXt1ZLalYEC+Xu0wK2upvs3nLorh9YtG
6uEBGpKXB3fwPw7wjPKk3OpHAO5s66h5orC0LOtkHUTYeIWukwLZttwx+5WOldYBdG4v5ulK36lh
im+glXdM+F8/vhfBn6+LvHujXG+YpOwLd5iTqtiXW+2Hawru5e26Zaseh9MFckezcbqWxYWuBP+D
usa1cNYrdHzS8m1rAamIxsmrd8guQPJQenbqlA7cRIJGSTCN+mgi8KlXBG/BvwSX8iapojRKa3of
xUKDAG3BG/8KiVxBaXqvOWXX9YlEd0zbT2d7aLgWoyznBVaxXpXnU6ukSwPWoJ3Ba9HdvouEy97w
+k1Efj3R8ag/qkLkx6mFxRB9s0n++At22cBHO05ISrsiY50HifERXIBJhh1EU92aQ87Y6VyvTkN0
45KnuIUdrABHKXuyzwsdwds/3HCdR4GbYYaTHsK31mkSNRqNS3lLCOqjd109KEXJZueAvor/3N4+
HLpoJFtxIS354NG/Iq06NYunZwANEygqJw9Van6dPNQxKA/f4Ebg9K9eEikVt0pxZowDzalJO0u5
+OFbLTdlujBfp5ysa5g9rgryRVxd5CB4Lqn1rRk2NAuNFOlVQNoO+rfGOwRIuLznOJdL5bnMaumW
Np8NUS3wql+S7FV5KFFLJ58tYnD8WJL7dT1bQ9WIRCsCfVmJdbIk75bwSCD01Z2g7yK99CYt5cdu
bVUiFzzzhfnzs1nyUhEya8WNa/81pq3VfE4/DKTHWaiq16VSUE6RBbkOTu5lFccHa6L1SEDfKaP0
9bH3WgGIdOmSInBUriQ6yNhfRGcUgX8AvYbDlJrHPWOX4tuJ980K+3HOTj4h2sa87HAZUdqZKYJN
UrIkNea8DRA0RXVcAzz7ZsblgQaJkzgNtA7j4hx9sXa2+WOCchYzM6lwq+Z6LiiwWcYg+dHWJCqu
VSj/yjkGaxSUdWdVa3LgEueXAzQga57UbGyJde38DlYweFk1ZhVtMh7fgb90RxuoYI9+m1VIng4c
Zepy15aLE6hnTkv8YkjBSTky4uWnjTggl/8MnCehDAWFmneK9H7zx8Tl2GVs6ZOGA1EvTiSeWjA7
0C2FBZyh+aiwMr0z7/Yegd5Kof9U5vf5CJAm6YLGaAob51WBRxhVECsQNKMq9KxIPWT81kJrko8b
vYK9E4kbUoeHiaKgnJpZZKujywXLxcZ2HqA/AMcLfHPzTfDFFoIxJtpsx8wyKp1LsfP7J6YQ0/bo
z2XSIvzNAAMhP24n1U7++Ig90/YLf6jodG+iCg+2ooEwsER/XEIZPp3ApKDj8yv0mtzVwlRD2Tk6
MstHlNAO6J7w9k6Bu51WF1zNy8p1Ap3/jcLYuGBq1puUcIojvGjPxQ3kCjEK5+O3n/QUT3bHZYdV
z2zEmlv7HKdkrfdfVtBFfWISVYod7gKaZXI3jKPiZerFsRkI4wQf628HMLqLWriLsgbORlflUI76
KpZYOBIUdrQCEYp8gO/DLzL2u1Q/QITrZAEd19VjNmLd0EZb7SyI/CVk2B561CX40AFdDyge6mAu
RYL/BtNX61WyJKXWZVUcHLboVcYYCix2sd3QwqikwaWACNag2VjBTOn4ggpQMMim761tWmZj5mNT
7aHdUM0dUpLZlCDUV2ay+Q5aWPMijhj5YnRwQaepiBFPSB7HI10uxr8AlSV4D345J8zsYYSHLsGF
RBKxvEoLPrLIyB6cd6TNoXeuEHeBZPGWg5kAXutVVTxbbDiDvLOzoJh7vu4/oOBaY8A4sbaYJesX
BxsPD+3YdxMj19LuJfIoqLknsMvtBwX+rQH800T0zwF+MA0SriIWBJUh6ms2Lt4l3LaeYFYCmEtV
vvbpr3t8gssl3iNV/JYS709nBRrWHBEwLt1Z5utskXJBVHxanxcdmUqH+gQK3MiJVRyAW86lkdQ+
8omtqZcuVpULAVLEbbC0jxZnPlJN0mmy8AH13394vscVl72jez6rDdcZMqiBojePWrwAaCnwYxRT
49OJUcqlNpZug48Z8bQrtUIzmKmboi2itloONdP2TivaepbxFIsBUxCdzLSxEL/sLyst0qosg6Dj
ekmzzSAzRVZwmbRnlsQMKz5Zhsu2qMAPwHi9R6VrRKrdiIus2QlM1UN4RgncnofYbCZP0LaMSAhG
rVFlMf8W/MFaZxyOrf1OVIYuntr4dDwsXdgASNnAFqeG6EHllqK6h5liotll6bdntGpd+fwwpC+U
utbsYxOzZEMnV2kHUKLZ0T1WsiPOMECDqzhLZEI1hNBOAk/1GggMDTpaYe4epFg/V6BrGHexVRQF
z9DAZBjMiJC2nGpH6tFWLnQid1LrZDlQ6KWYipOT1ZdoypgkZHd6uuqdRBd29jlrv2Ebx5DtvB+s
8sUmzbuGfW6b9Ssky6ZJhxgjnnDkW/Ta5Y4LTPnw1ckjYr+cYuHfO+W4av1S8eOo3+PcM82juJ/U
922ML47T3u0vgOvLXgnQHsiPATY6ZLhODL6A4w49N6uKf4mkmq9npMn5AA2I4eLkZRMt23pMSZV1
LHcZNxafVg+7aXdeKt3lMo1W18k3v9cnuGCvVYu/yLaIAaBT0rMtm8MAZoW8D2IYVVqp3VAXtXwz
TvzXdqlR+akl7pyHn3Ef16tV5M10zFPIOfcRMrcOtEY/7Lyc11IJ6TM18nU1CFPyMWj5g0AUmzAK
ZeKQJi/FiwzBHmUjfYUVjsBqhkpbyGq3YJbRfhdQWWuerMTO9LO4EA1VAhBW8vVjiTiIiymaGW+Q
h/1RhPzwggsvD4uPa1koPqcaba3TBWZsmFVYNGoNup9SYo0e17SYBS3GQkk3TEW1Tu03NqARmvnO
TFL3I1RgoJW7VCkhCOME92pEPN6lH8nAMOX8sP38+/SIGmHdi9HhzjqE5elr4buReFH8aN+jdKBU
sJBn+9V4ls57vUnHrLlwTgMRY3ltnTatjdImB74/oqKMGaNFpMBZVX8kfRjTdT9V0croQw8C+Kaf
QFLlcvzaWlmrmMOztphhnY2rWZZ52BxR9I8J/KfzF+qQWU0q9aSJQs7P8IBIZCF5b/wssJfVyHdH
uMpSZaVxkbS2IBo3su982pNj31toOwpt3wBBGRaq/YBU7Ly9mSAfLWpaszMGzJfyDs8WBFG+ivg/
bHYOUpBtD+BVtVNXAS65tQaMTtehalfzHc/gmnuq/jZLGV8L0x090+uwBW6l5+G3S/x+wtJzvWGz
yBxDJtTNpOyaUzO8TxpsZIDyU5p0f633HPJTixMUU/8z1d0NySG8/rTJiflcPdAoA9YUP3qTk8t4
HUPvzQ53+O45OGNLQmNsGBQ10AwcFGOQ0go4CeekFK5LcwSWC/qEp9J/FNPK0Gz012/k1+7H3cmU
F3UcKXTri1TJqF7zv//8Tys7+Br5jAcOBn3eEoqRw39mSOHIVdO2tvF8QgkB+S5YTJK93oELQpoW
YwkIqyeJdN1+yzy6+KlTNDWX2JhCFjOoCzXQkIecCzwV5mqzh9CzlOnkj6em1Ja5K3UEb2cJrvMH
4cqBNUnX5PyRki5f2+tETOr0gwef1Iwof7Xl0T1IH65cgrxJkdYZEcUE6LDSh3k0TtVcrwRzsjRl
fpyPoifwAMwjwPf506VC9RcGFNYXTGuz+10xal5MdhxjxZGHWWPZ5FPtXrmkfZIsZoXEVlk3lw/6
X0940Ted4XkK3wLVoDbtM1TrmA1HALqJMWxBQ4Jads32kisZCshkGsZASKe4Gvnl8NfSKHmG07CN
25QUexC6hBn0lntJcSA1iDs2asKcsihr0dAqxxXz4eSsRw9BPgVx3Y8I7ig0vyi7u0wnSPLHUot0
rdRAIeOf8wUiadU5ZJhfJvsSE/mF42JQTdsCuN9Zru+JPsiIWZCaasBEwsTFLqG8ltOfmRkKIV0c
MhQzs0VHki68Ug6Ix0jN3RmHs4kP18IfWl/j1sUJLuh/A9RwMEI3tMI4t0FOkxXMaPr/NZRJQ86C
8iB+NhIFoW1NJZoaKOukEo9ZPtkStfKY41JC+Yy7YRWvBrZSeKA1bgU++qeZdriVDI3+K1r0lFiM
0QyQdafRqGnnGefVO3zQayM1Mjj8+m8xraxFL01usfTFqtv0I2ZrBhjToJ3DIRrFFy5u7AUg9no2
VtIQd6iboGJvASb44r5pLXeyO2kFPkBjmbx0MImsFDn3JJL6nPi3I6DglgpCYUW3o7QHtq5GYpoh
milp0ZD+iubnxTF3WRA9XQk+U9pWpt/tA1QlbjuWrdTLeJodVYuKvcmHDR5cfbLz6eLd5Kc8g5B0
LfUksJ7IPrWlxbZeVJQZy7T/jaK4r8+dmiZh3c1d7QWbP/NDPfo3K1UywcvwCKt2FPu1doHE3t3z
fnKFJMezfq+kEPsH9DPwZDg2iUhtwjQAe+6phP30QTKpWVlrSRLRvzVDr9nMN+qfHvwFdHwUqCra
sU0jeIPxtjKqL/x54pjx8XsUczUNTduEFvn2Qk62oKEXXpXYWBYXdWUc8KOAeyh2Ya8fAOwESxWJ
U9vRlFMjjbmN803ywPKxdnAPvYQpnE56H/NSBTa0BN0IQ0GvkyrcavgCYZUu0c7CvTAgQZe2f+cu
UrCMyq86n89aSdYoFjwPyK2uiR63MlRiosvwRmdFitqI2ab1fgnqHGttAv1grh56HtgkFB996WxM
qqNEZ36jeciCiW4JG3YH1UTIntbd2PvZ+EOiNjZIVur7vv3im3jMVeIhlVljvi4I+fqBol7YRS6b
XMBAI6hKBWA9rlfSHTWeRufbCJkQPlSAGOAXNBMiYMmiIiYaMqqOjECwXBxEMzpyEhhGlpCiMuXt
to+C6RAigNtY6X4Eeykm35pU8O5ZcuVK0RZPK5VSAaBsZKC7FKze5KstMyc6vIyLkoqAI16eJT1i
f8GIPvU+3Lm0aoIp8N9pY/pzWMcaPVrHXGv6pqCX74IOVpwWbqV9uEdc0vF9Pyzlq/Y+FGeJBhoU
X7xXDO8bswcGVx6DL7H8cKN1KF9+18E1GEgyDEvUZdwmeHE35Y4dUrlq/prbUktmJT8JqwSYs4DT
V1aiV+6x5kZsH/IB2WV9D1wYvYwnD+AD7Aa7c3LggOv8E2WVpKojeWkE7pJEjB4sJxbQsey71Zsn
GD28XLR5F89jz3OhRH9Ap+bX8GSlbaul1sWlYdJV9KK8bKKC6bZBAdcl7mM6lFxbAVz8c2E/a1d8
X5E7SpLtgAt2mpj0432ywKe1eeZG6FOsQak02Xfzk17wqZF0vb6LL0/ISac2P0zvYU7X94tBT9i/
Cqd9dMbxhhD6GCydMD3qCGez0oBZptgX3mc6mi2JRkda97yWZDhEFwXtED4kBp75GR+8omPxhiP3
2yTbPVZ0+P4lR7CuHIxE89afZQO6+1rUA/pATzr37uzoolxqpIB3AL2Rqyk6C6VSQ6NyRBpUqRW7
klZOgkTaCKiV2+DvWN0TuSgNSfQxTeAIJ3ErYuLRQIK5b20sPH1ju9ciFlG66nok/8S614G2SKAI
+BMTQvhzpKgNodalKC5gTUZK7aAg1JeDbOI22N2KZYYAt12VdXbAUSxNU3MudkKr7nTDvu/oAHeC
sXXjJBXBLtBPdqgxdCGDF6eSIDMbTFSXjPjmvWZUYxIlmGXNtXqSakp3JuB+dBjnHS/fqKEJXoah
A3BTEYbk30HWV8PBhIgogCpJQ1A+jN0WIsroQqCY8KeZvVl1OCs+pBB+/LuEQ7IvEdTFned2QEZS
m+gr8POUO726RH+eWyZmS9uBWru+j5oW1gpKG9SouFbMVOvnrnKblHBpdiqKzE6aLXfBN2jZfPS8
xdatwb+oM6BHiMT5W4MCm4zuaU2Wo2aVsOFccEXNmd5PBlXbV5dvNOTPxn11Ntnnz2WNF8qZUc9c
FEWLdvtoh8Z+M91SFU8/c8NWWuhEwlVD/q+qRep10R6/ByeuPTG3l6PnfOc/AtX/P/c8NhJsqCf1
4kiBgl8gguo3yvWdGWNcGlbADih38rrmdKk2Ox2tnBK+AUbHyJjK2WUVhTRi8E4D2CBtJL9BYt+a
7PW0qg8GILLmQ45aud/ExqyTC72rLD8qJ1mnDUl4XDlxbraAF08un1bGxJQ38IUrJ1U99IwetLpf
NH3SGQK9KQlIuxCqc21gfMqYW8HZpFTXtIljDd3P589Qic3Kss5KZCgwgjOjHHAPFdwUz62YAtCa
JeCP+woiEEF2Y367xJ1akrdwLkYUux3NuxLYa/YKjVyf+otb7gjD9fZmALAi34FXb6UU94kKoVSO
waxtavoAu3bZEDHPGmfbQaMcdPfVODYiJCoZqBsf7FbgjmlzNHcCcdTatb2MQ6hzt6pBddquYEdo
wHXfeRQ0h5FrPuQJb2GNGAO97jbd4/Hmc/fRaYnegHCfsjrk1A+mpI3hxrt1XjILLCZKgim51Koq
E3UA2n5Uo7/VTtIpIMTjT6po4iBAxnyKHpmLwB36z730QjIV3AY9cnm9IL6Pyw7sqJ38xjpnWKh2
xMskQ/dD8kSU1xnVbB9QLTl3FGba+GKE2pi373bb4o1tgbQqd7K69ltAZJ5PGHhl0IrDpRU3fcdd
dM9AGWSfiId1yuuX1upYmK/Toft/8fY0z/RMJvsasIBLBP0rvrPNAwxyMkV6uu20CdytfL4oxbXu
bcESd/7uBStjGR4Rw5PebfiegCpDctBHGdsdwNVNh3GEhhP+iIssM7Lw45HUmGOx8HX4+hrkpNLJ
hYY02QgE+Gyheemu1uw7lQ+eZIQyUip0vMe66vIEqFL2OIYsZz79evN5pu981r55Pw33OTFsbA8V
qdQg0vrtd3SCgaorXWomQbTSCaxmkRPnagC47RIBMfLvZ0ZpUmNXKnvIU1CY/RzaYabTDhP1PZGn
mWblin5M5kXStVKw2HpItoxzMv8RpYEX6oc1TbvC7tTmajuPVGarJc53GIRL4rZWcDQTqoaqSiHE
aagI+WdKzh5XMLUukIAJ1d2SgfiCUH0EVghlYCtlZuQDdexyriP6dltW4iZH94s+1hsRIUzGhSlO
P/9aeNYjhBp9pSjEQ48b+4IGD3c7N0mjI/tRBYwStxLRxJcxW+Z6rlLsrp3ysnIdfIBb1k/NWYKP
ZQ6roDsBYVSFdfciwM6S0jxkoF8baRMbLU2qv/KDOIUbtpyu/FjqI1WsRgI+MNorOjpBNb2tyDtb
tG3cRj09LAjI+y72kHKGGvToYlMrNzUHCsZd3Yzao7jJDifybchlNivQnssuFiIRkG+qRUHqCDsO
+8pYWm47K6sdN294CYwrI0NcKymDhprSKI9cWtemf247yyOJZfewRz66Cs/WqomOy+JF1sQ1VksC
ySdSefVOmZaESjj4yiHR4Xrti+JH1Mwvgx6TNh6DCXUOIEO1mguz6XLpBjoIFJslVfQSa3blvtXs
OtJSmrTN/f2qIFNh1EM9R55CnOnhSeGK0TJOorwzHFUNqWaPm8mkaz4Gll8dz2j18X4SWxDFjOZk
TIr1Nq8JrpRfBrvLq7xeb3brzFoU1gIMY7yc2163bZe9uOwn4gwlzDraRN63khfNqy8/6CrXVVxW
tUi4CgjwiKgPDKb6smrIMC3yBJXHq79sdv5ubKV3UaO5K6b9AoCWO/vWkN0p6AArDcuHM/x1n/Mt
AjdKgyaM88RQXYi/5/tB2Qa1IcRYTwGw5526LefLrQkMdPo9wZf19qSh3FFvfKzF4cCZEJt1/WeJ
JwC9OaZ2AlfwagaJpv9fRwLvreb6Jh4ZIJTT3Iuq2Yqk32iRJCEnCqpsXRIT9m22+ThBiwHNlyrW
uxdjBFQAE0TgC4tBBdnrXlGTZJSvXH9P9uqHmOIaIPQ6kmYztkYT0rg4gMnkINAaMe6hTP/rB+FM
cz6cKxJv00D/rnK2wpgct5x5dlCaTk0fzIDQasdHoUF2k/rA9CuqB9RoH4tHmPG11/DveDaDPvef
uWqpYUeSfLZa86cQOnuFwiqn7QhLrKzXUKbaghMuhVDJfXywaZggHGDy4XDRzj/PQz+1un7yHgBK
Dw1c/KimZiAc0Zvpi6jGnM1pI+Ss/Zjw8fknAYbUjsS5IxRbNvHSsLfs8LjxNwK8VBrmWxtpI4jE
2D2X3wpT1i4IXpgG5Xnmb1+1s9sCZEH47AFf0njoPmSqaK7SOYUoxf2fSaeTynZ8COYQuOoeWdwN
HMqYO1mgnTQsH8J0QBFpjRYclxFNWXZikWpXcqKyMTR9TihjicryJIddLzr6/degkgtGAd4xxJk8
QGw50RpJWWU3KvR3J8l7yuvbutmJbONBDZOFuA6Qs0t2VJcDXaZk9nyfR1tl3dluQnKQZnQo2vwv
8XpN4LTb5r1M0zEydaEFUhPoIm5XDLuBmwSMj3BgICEmIXhQnackA9nskt01NF2DBkestMkiGk12
ypLR5NkE3eOx037N8ZS+wd4Z6Ii08OLkVSpw8eePu7tIbEjXWGJQmpGfaIsyQD2Vm5v6gGcveXCl
pZ9QNHVEwBJZ7t5bT3vHhlAY64zjbUPa7fXhMsFefPHUxiG2dld+WLFQWUgqB3rL9Ej/W7XARNuc
/HcB7O53fr77RPoC56vgcOWwa3wcFuQTqe/t8jNPEPKI10IboPFuccSBQEXd8U0b+BVxapjipoZH
CfMghkpAYSHKyXpcjSXwN2aQWJtO1pSlZ85QUN9hu/j8YrbHoGpq+/x2h25Pw8pgTzAMwSs1J2Wh
R0BkL1FqgKAszgf2egeP9ab0Hu3oxzC4+jbPBhZz8RbJaZhxMMgAqRFm4oBLsnoX0NRab/4vxHIW
Hrhj2TmYlUVTJ61YecD61ir1wUP4r4I4Pz3iAg62aaktzKsjOsKCp+3zKRHYTxkhNIQOo7PGr4nX
DhYeKYWzTKA2RgN4GP6jRyH1tHPRxyQ7a0j3VRircqq6+UcH+RV+6T41LOHLwsPTle1gA+ANXYGB
1j7g63/Ql7bqRqeGL3rizgxNXT1XFdzdM4/4SI6M/YVYOfq1xxYPVHQ2/1Ag+OPdOD9GcqH7XxYl
+obtudmfUPFgvfIqbO/TYMFF7ZL7mthntrzP5gw7AalR/0dKM/Lg8oNPOzbNg8fj16ipZopCklx/
mDq3KXNiA40RLCSGNNDz1zHFHCS9UYrT260sPIiF1ajYFq6i0Qjk9N0dNx57IeQF1PPjFB5Urx+L
R9KLk5mw7kCVz6uan4Lb3Y1OQ7q/zRbaNrmNcmiAzuf3/QiL9QI7eK19JYVih+xXrLSyjqq+pq/i
6Mi1RvD3kQX6rSFoob7quVZs9mFGelNTf1gFXve+AR2VXXPxIWwT08cIYv6Lpc0ZwGu3gLnZpcsF
9wH+aXbzLGhQdyyzgD4Cy3n3vEBeDxKdoK39abn8P7CAjFb9RZhXY7fsKoBe7G9NPGLqjM8ObqX2
ToAxu9IGYHiNjWTGyDJ6XPiroInqbB3q4gMNKouM3ChKUbM6M76ZDmodRET+ffbw1blPfaJ96OQF
ETEdRNh4GbnJj2y4r/byuIVLUIZke6ItzeUs1aUC6ml7iqCvVysP1HurfhIyKUGHlFZDyQ8RMBho
hoF1iQhD9y8C8V761EcFCZoT2dCk0LFjV4c2MZ++deDtvB7xBO6jND74o4xRGMi2QMJAFy6zcVq+
tJdA5fXVCT9SuYpUZx+VEruc5mjRBgTmoaWguD/8BzQcgNxS0v81IapAEv3VxggC4rvArcx5P+jM
MQ0SEvuaYhkDWnQM1HsNQ1C/s4+3QGaUUGZz+hBVEfk9WeV8KAOhyJyBe6/kFHDc04mdUYPD6ZV0
4i9NzeQMc6QvPzbIFuj+GKXMGeQZI95jUrZsdRbQRY9AEzjeMx0AH6DOWtVVRYh+DOXpJs/p4I6L
CVpnTFUCHaCiAE6R01gQ5r4s8aCwLcV/kvRDckNANc4sQrpKP9xz8ERDG3eMDrHkiXNAPV+QZWig
0BFg3oL7UXpHZwi8QOv/LCAsctwycaOsKTR4BYe3tMq5Ssc3AX/CdiQtKjcAJSlIaNvisopIFpUe
XTWlUSn5G6iodxpNyKVacMQ+MgEkE3hBoFKrEPn5opP7rJD8w14FCjkdcTJ2Wexd1/QyW4qJ1EFs
mT6swumGvuXHhdljp8LPVwT0KUrTLjWhm3W5rHl5ybKvMWg/8i9O/34sn4CRmJI+Wv7fLkACWBU7
DJs40gETbo9BvNBicmgWsjfKzqijkvIY/bDnxQaPHguKDJLfvs0botkHPX2C3/R015oja945xn18
e6rnc9Ja7ajeyTAItZPOEFIOvyBX/C/RPt35SlzSoZIe9NVZVqv5h+yJFw52b4x3XwWTpUvkcg6A
N4DJ2ZioPid/ulrDvA06qPtLxGblGVmgKN5kTvHRTyZgdM3Q0Dhh20IIKUSG69yB/0k3sCiFWF6c
7xGlqUnqab9Dzsvrw1tjKh1hyoHsYa2mGh3UqsGqtreG1qG2mtJeZ4b2V+orKaX9NA33/0FuiuL1
Ut8QF/4t76zF6h4MpSU7019iRp7lnr6D/kxU+Fz2q1riLS5IoCHXUiqb663kQL1CzMnqvU7f43RS
SwLYr8OM4MTROPrIzLHQjKiM19mHvzubGTBYrxT2sS0D4k26C1zXTidn2K8NZ+LRRg8765CB/fjd
Sef+nz3CzQkK3wMP0hHy6HfhYH9hWlTgJdSlTvsORJEarMHjv2DqTyjHwkYull+e64cTzSHsr3/7
81wQompBYtwV1hmPeRrIc+5uC/01Jy4il5fjdlfMYXTjIz9RfeDby2KxzHKED0FvoWbr63ngKqcR
8wNDYtVZajHKUmZTPPYlSnRfduRSbDWxKoMxqGD7Q+9MCG9lGq9FcgIXr5qZUcIN1fHIyEW8hE5d
fJt/Da3MVD5AyQyU/H749Tw6XGrVSih+ShOF/K1wMAn+Y5Klrl36UQIu5jkma4bVNKzYwzYUvwnf
xyeeiA1K0t1oA4zUKZGfU63PU14gpXbrz1xYV0FPqPPuHSg/JXsh3n5eErwvxudBmno5QYFlvXlX
Cwy3FFogEv9o2Csk+9+4zkF34I8L+7kIHezLf/viW5En+Ql11WndsMt9DDFDg6yeqlkemceef5QY
CtebrFiILXXBsjL6MiKX3la8moeivaqwXL843h/N+lp0BMqanlAYYN7kgrlttrtCxzRZV8coXrG6
Ih3HObwqCjAcDga/4lR1V6XmqVejFaGyYvWh+arfxM5UH+zvdSi9o/nz2OC+NFqkuVCiPfhAvy02
J3ezANQIlq5YthLzM/0Kb78cVb3qG4NtOVQQC92wcExRc9co23YUD/41VY3zWSuCm3TX94SxL52X
lZ8Xj5e0dOI+kXFwmPBmTCXp1PEF0k6bhxlCxWUk6VKmlrCflTzDolFzuJMFQ5ruhZAzXCz8iQiF
lANLl7X4LS8RHcDDq+x4ucZhvj7EGCFgLNxaPQnGGqAUpb0ULRtAvFOs+68pA0ClMrNo0NFsrctk
dOWyvo77GNVjA380VAgdZ5599Ik5HgOlbiuhuvCb4ZpYBoWKHCS1Thyer0uNyXaTvS2W0q9GcB6H
SCWPQupPog4q4oRYhYtTCCFuD2cOlc5MMhdyQWnCc36C/39AOU1E2bJVn4YGuwu/MJHn+I/pNXEC
7FWwjXVfgYn8v2S13phqOPDWrIgu1esEf4Vkz6ryFK1mVQA6eERPACgvg6VGCgiH4zdFm8QD006I
av1QjB5XZu99SUGj82G8/wfpKNJYUG/uhRuKURsRDtUdY0i3gY8h9W3mE+lWhb74SEX7IoKs5Yn2
2QWLdDmlcWWm1nFsrVX72EaxXn8M4L9luZR5IBjecnCMk1v9GM9xcv5bIlNFi49/AVg0uOfbm9YD
vMVh1vmQlDRaoCxQqubd8u6TuSPDBz0B50sHuTWnjwIA+GH0I4zuzKitNyTpMxcLkhtcFnXYdGLB
t97qV35CKPzR8MP20FZIW1bTxyAw4iSa3PlclKGqspeB34V7qtN1hOEizWnffu5fUQD1v5hVJNTU
feBOYrGkVm0EPD74lIjR+5kY23DR0sYqDV+hOaICddrfubExTEQsN9kzKDwzcDlt8yi/zt6DwmkT
IZQYpdzTgZS3VDCNnzpiMH0grGq9JLnXeG2DIP2rjmVXwj/NBQqA3e02nOJT6Vl9VRBgwTyyn5xJ
f7tbR3Epn9Lyf5um/CmFHv5qodc9ZwKFCvYeFNKhfcsHI4YEgqDUBDyxwCk7ZvtXKryb5mYYM3E+
tp5CcNUUZuyzujk9JHupvgxsBpKkaQSxSqvVVAFbgb+o9hYj63/tKgo3suGi7bNIlT4RwToVYcK+
lgpAhIB9mnBYU433L0x1payOp7K4qjVbfjID5AWwUig25UiRZgPB9w44IFvoOt7/blunGNSotLdA
BvBxJj5Iwfr7YL9oXFRAso353Ld7zvKSvabx/ddWUidLWWiCoMXS4LX3rJmTc3sKEHxk4yt4ro5f
T9r1/KmiLBK4bE7APGaRObl6V5S9jkU3vwBdU2O0ryy5CjRdLDoy6lt5xa2nxyttpnULs9gBAN5X
N9DuXV6E9gTDvIyRsB4fahpNNGkVmxiRGwjme9QRhnBYXQLPGOns+jBHYKVPvq74RJMq09iStR+A
Xpv6f5BhFiz2OqEbpO++U9KKt64Sng+/VHP92vGAhkMIu40D+V6qslFpgwZ+fc1w3a88j5U4Ka7G
Xt+pyqpS8PVauMc49d4bhotT7gZs8z2yBQREvMhRSYT/2LZxpJ2b54cHlgFE9Zz6x4lXZQdFSKKF
C6KValc5L0btDkyPKZsGjLZhhNEJm2MzhGZxjUQZYASv93jfTi7wveagV+0eu6DJThEpicvoekiY
7hX51Z240BDIATWbcG5fpXa30LDTlYleFl+39ltLuJBvTRBFTpoPANoc2dZdDJd3h3UZSFcUf4ft
d1woj2BC/OwkI6lzKH1GqwAFqABms6si53UCUNEYynfuagf3qwgdJVE/0FGUNagL/oFYPdGuWNiD
9Bqhwxl0XshVoWjSypRALYoMeRMts4th+/UQj2cMvFNLfi5/hJp55cJfhTu1sFy1Hvi9V+4yjoDB
SdAIVyYEWjAWEIhWdEoGiSlmRZ0EbxQhqpHBo5yC6C1BYIgE3VX8MpHmUesR0eGaKfvdnhmAyQiB
+C4nu38a+65h0xtMBJHDuwfFuy8rix64vZPMMO3hlw+8Yetvg1aBNqHyfxxA0nXFRCUHzN/Jfm0D
ZA0x14stpnJsVwdxTF3slje6OGGGTPIVWP/cPg5GE4VsB00wmwoeJOja/7aVhlTDQcbeNHpo+CFX
1/bXDbrOpH2Sq/kBeyxQt4R3T+FmuIgnAWQh+SpKi/TQOMJJW8E3PrNu2kkDuc7xWNySnFP4MK+4
UIpwJBp3jtoote42dKKXpuGA/2C0UI2vfZbjA7QpMDhjjjwp6kZfoeU6msNcxwghUZmKiGR1yaB1
YsYZhm7XExp0PH6HThzZnsd/Y3Wn5YwDEp+ncCRALnMUh3Ehpy02jypiLxGLnxsDpmQJLy1DVdfT
vGMiYGV6JSenf5zi8Bb8aIe6NV3iICH7hz/ihuGZTgc2dQ2xOKW6mwlGYLJnjk3GwEwhD0dKBRhG
VfsnX61fJo1m1lsCc+PEMXazkrCGb5bf5hzQwP/gfwefcnhu3U3pcOFFw56J1li+3sxBQVSL+Yn4
VZKB9obsJYonXf2qaK/fgyLn1QHD6754BuyOqwYbWwVoe9cYhLLI+H2WaZe/EXiIgQGZzH4wB1Dw
wVPaDWfLx6hGz9UwK8YF2gkpg+NEHMdcd9C3x5HfWTDkCTLQx2FuoreVbrmaYriIycLmv9Xc/p+o
7f3f4CaifEcBAbuT/H7hmTx5BzRulUfUIvmALKIcAyAmb2WBYcCuKM4JtyPTBpF1HCKd6hMrrCmr
gsyx+z1J2aFNGGGByqgvlKrOJNhtNQqvSjqdwU/0HhAfQTzrgxsn6BxVVhhiL6AiIJwrGvo82Hwc
4e2/HrM/Cn2uefWyfh7eIo70wIPLne/ZxTeuJ9aB2auisfP24+jSumGTdcU8GwkTCZ7aN9uoxyIm
xnyj6J5eFV3kSlLieGBfdtBW4wod64SrmBcY9fdU3zcMfx13A3Hl4zRtSLZq2l89m4dIZlHHZkWV
cjbr/XHIJE53iRvo3e7jFmtlIHUva7bwIElcmkelhYZrkAe60+Ri7852qb7UPeh6LFr0ckAlfZgW
y9/LedXpkNPUFhZrtYxJhlI79wfLYciW087oQs7IMuFMblCbQSrCLQfl0/VqNBARn4c9YDHpgiga
PmvdMEV00dUuQSmPxOPKC6XpQ/GQWBBGyhS05J14GlrWUtr8+2BFTtXlRuarj1CGPA9KZx1C8eYI
Oky0252uQKRSCbElU33iMkw54w3dArxr/PKu0sLQXUroYHIFvbWJDivRo9s+CyN0P/YWFzYW5o0s
CTbYWNCk4LgI2FHOJt796r6X9+9Xo8IQJr3jpgVNnSb6DByRkMaeKXk0i+La2o049pQqfl9BUfD8
ZA75NgdQ6RrQEhbBdNSaw6dTTqzJUP9ooi2eKRmLLAw4qvF0Tm7eMT8tOBpFdFctqcaBmXnj5V8d
oPkGDfF5B+8OEhc9HRmju1BU7LWGuWlf0djn33PAnTKhAuPpwauilozLdNCKLVnmx9SIW0c/Hotx
HmKOePzLfQHHJCUikUZaq/ozM5wGJjJNUUCdEEwA0MpAGuKw3EsXAp9jEeLoqQImJT5VPNSVkN3e
y1KibfeNiA0r3Uuzs7ry/JjEkpWhRsdIiPL4fFfLEEsIcyhcL3PW46DxKPNxed8iNmG1U24eL89m
kLTVh50cs7bDOTx5SX1+HjsLAxqgdsEUWKCQCO+a1ZcWXeRfI8IEJ2ku6XyNZEB5avqQzQFWGYip
aKel61FPgqOgmCTEz1IyQ1NiZ4htFQv5G384igI7iuKRns9gCK8033pq7GKFuWDzF3Dcw+ZmoEVR
9fvcAOFJrx79TiM9+hoVhl1jFAy7JeIGtgLyPPwMGBP/XJ7HkCXR+8Wcfy4OXYoT6ETKRF3OG+Lo
YFK75Tezwq7u2wjiiv+R8R0E8aqFXHkf59EjKhj+qqBe7dGe7TbAxPr6qK4X1Vez3aT/GvgsfCaw
ArucKlWMvR0UoamgcjBbuUfxpCHHr1u5NcY+Wjy0Nw+bHbI3WPPYIzYxvtdoAp2tjmPu+gmh4Hv/
1qf27hVzkD2ziaj9RkyfPsk54vnTWPvB5v3RrGYcri6rUazzsqLGwV+Q7b3T8Ctr4JV0nIyNTO9P
8CtZ28fhFxbaEq4VebNigrt6AmRiS/IdxdvqxideUP0qMD9rWk1leE9N5aV3ogpRPwEmOj47uwE2
RRWf4aNZLDV7Bwi+v7PopckgS+5hjb8ir+rQTuXLIN/0EVuo0tSvmLGH4ARdpWelTEvOvVnongvu
3krx7REX9L3PMoO2mRa3uPFZpMtiPbxoi2YOE8DFJjAL7vG+0ixZPD6RN6ey286eLryksikI8B85
ZF7dmmmKndheU8mcn3AFXFwtvsF7iRRWzMfCOUM3NQXkiemdVD1zp37EKcr0kL/mkJG+ZBrt6s0Q
qzw+HIeUMxmK5dI+DixSSMcGZB0dZkcn5OUT2jbk90941JWtU0LmfjtK3VkG1sQU1cAwAlCQCSqH
NsPlndWtgUTNrasPffsI2Z2qrumNODeFo6izkBuzsTk8xJOpe2yzwnCG7HgdHgfwc7eI7Nf/iWlU
ENJhvdDtsu3syEabXk7nLPBQbxASe2y3olOJe8T4bw5/bBtOZblV5yKb6CxctdtR1eNVpcpADfs3
VPnuZUG6xxJ3/3EpC13+/Q1IO0rq0MNFAwSoQowPOfvJdjJsoRzLWNMNgWPjOyNlTZOP8KCxc3T3
G8wvLv4vTmCfEzGkTkUCRWoptkJmYay3nkl5fTGk40mRikA2l2WRnYUXBLu7s2fn9J16AUxMQQ64
JqVXgwtcpBzFlTmk4zj5N9Z1heTJTZCWFKnhQpQVETBnNQbLrC+KNiYRWx3N/mN5DqiwVJ9wgn7G
EA0cA09Gw2u/h/NAgVpo5d6qguQslZUNPUQIuz4TRvgCDi/Zyi0+a7Ze5x8ooleShMyjYTaztxAF
/jpjqwCrKj33JSdL4vuuneEE8O0EiMrXWiXQtQBHXyxAwbzOA7n3yateBcrcIIVokC7WLHQPAD6x
sT5Cs1q13kXw9JLMrpYfCCyI3KiCfZfON+EK/0kdlHHnzjD60bdD1+in762NvQaN4YORZ2OFhYDQ
odtSWo+1RSSBvmq4/G95IpLe9rXBRjw/nPHaWGW68Svr9xRyiHWNhN1xAZphwp5VBgk07LfO0X92
rOCMOy0NmvTBrnyaMGkuY4lOAcjF7VNzLMz7OwlOWcNTZPNtIYmTEeiW2bc6WIeP1zyNx/k2161F
/nWnSUgZVDLP1zsWHaa+NGlAClBmcmvS+lrZ3IK5LW1tFnSz+b1nOUUJbwrJyE2ub/JhVwT4mF7O
9WDfh0AkWopHQMCZI3sAb7Kvyd7RU41ELBT9LDf4rl5+cpVw03l2f6q1Qqsd41h9eLUEu84gTa4G
iMFH9xWfabcdBUsOwd4f2Fpf7rJGydKJk7wTV7vunmr5xvFbM4bOnUhjDSq3j565WMd7HjaYvgUn
x0UEZr7M1pRhNbkXptdmwPGDeMJb0115mcsl3OnHiSZ+NRvZIGnO7u7zdcE2WvtMttmfaoqRQxN9
LjruOmcy4uBfmYyvQc1VBpbWMU42AE1JkDowTcy3gKNUOVjCJe+e9eeZoD9z7EANcs8ZdFZQuEKO
EV5xVQbUb1hF5b1RiYGn+iju8B+xA3loslfte5vN5kbv7u53MDCh6nQUAe/8kWGcKy7cKWApEdea
5Q99Tvfe4Z9wpu4vsLGmO4+wx7KOLw3LT+yPNoT4sWeHIEvZOmwL/HCIqppWVa0yi1bnVzPkuoBi
/KeXYMzwi1GI7Og808rPrOIkr6VTBShb5YHUWLYMauT2ADZnC0pLFhP1J33/GW6m02tQlpL6gtOm
uNYVI9yc6GPVbipaZPNjEHh/S3iJsng81ZnlHu+3y48TjndB6Bps/uI0F7SkdDibpCTVvZGrX5sA
6GALBLxrE9pDn0lWgTejM53RXQsHNb/jcL/FkUwCKSrdsjkA7xxPl+CjHM4iFWjG8dIjG5Hrft10
KwiXXM6qM8wKXsh553RhTcJkcDaA68ePsClVkNfXfnp1insd9ivYoIJY7XMsmPS9Ga1KzlW3giV/
ze5S5GEbzsNEIBN15iDJAhpQf3loZTgJRKJoCM7xdqGxMMfOnDYN4SixEBNh2A4440PX9e9E/hTX
oFgslg4wovLAh4cHasspd6scC8+FR4ERs5FNdZZLZnfW0trf/tvc/AhurSQ33+srTiWDQaGF/+CT
FVLuS2y7gwErPcepRFaXy90NL5ltjC6nC0O0jydz9B3SMNvi1Rp+rfsZWthvVlytjQNAY8kueL2H
oLO9zcoNJHSz+7M16UYGwQpehkVJWJi1M0nyCVcXamZ90BHL0a+07AlarzHYImFpqwMubHAZNlka
LyDfkHdzWCond1MPPROFCVaF9WdQnILak6Zin0ZvM0lRiLc7kCDY7Um7adxYTwqx/ncmRWSFJ+Ae
AF5uG/mthv8J207mPL06xZq+eGB3eBYTI4ByzulIObHr4dXHkMDjZGIM0tfYytmPnGJNTpIvoD+Q
ex2SJmswYgonOwOXGK/UhjOzs/+FQ/OiR0/neCDoXdJofMMrpV9tl8ha/T5nNxVJEhBbpXDAyQow
UKVCWDzI8E8ilnrDtFEN6rNB6j0RLe17vmcVVhLs/j4CSuXSoeIMpm4t5UPFBSOpk9VH1Ataruwf
Idf5kFDewpJ2LwtiNOyIOkwg0I5g7MmZR9sq0wrHd1++0ITvumkH2FPGup94TcfleFPK4q47nVBi
dEKU1dLZ3AmblK8Rfa5lSDePdhLaB6SlAilA1M71FUVshb9EJzGqRMTgLGRiBhD+cHSFx9jaRxxE
30nFLUDImePpKVjQol8dEY8QLuWTGGTdMEa31v0yHJqQwOuTczvkvZrFlMT2vbgEnYgQPTrZjlck
5t92DVaUa98r9pBH3mGH0tpho687Kq7rEW3gNOOaOvPq52Jfd/rHbUa+g0lz2QclQDDPUCfxSblc
Q8fFd/k02bIZjjyFb09KBVIODzUFVwFPMTFFNUroLbLe8S+aWI/HfKfReZ6/P16BCrynXwgHTXmc
hNd5Q8wE5jJKStXS5lhXAflPU6hGgg4RO9fJ6e7yTQM3Lqb8wTa7dNyMpKK/Ljyk++EBX8NYZJDc
VcbYqIIs9SXp8waw7YcM7U7THpjh0e4+j5RObuScnIy7AwK5zlo/utP68cuQEfG2UFGe8OcKf7lN
1fiOHog/OxExepO2LSJI2fC1p24uXtl1a4Ly+iulN9d/VfFMbKriFeRL2DmUkg6qKg1o07iIIjNs
H97e6zWowzKS25JN83gZUZcVtlg0pH8rn7RZ92lc7O752lHkF7oUoirWQ2twlfFoNdi2M3nvXd3B
GrkSBL/dY3W7mHq1+lzGFlQMtluPmoOUPYEmfOVjXRmSneY5qFvmsRfkDD4eq+nQrhwnCY1R03O2
Xu8lnp+x5qgiNi2wDVuezmCI+iJ+NTgcUVLrnjNz9IQ4GIRhMKxEtCjRgPNVBWtezIKX/6aaOrc3
XxtL9neQoQSzN3FFQvwG42TjMPt8Zfh474sL99JIuCGTFZnM2QFt6CqzncegJ4Ej7K24IC29jmwo
CgsU7NvZwcmrRHVYp5kS0fCLyHAzY9M9cBgNCYHI5817IURpQnoqAiU8Fsg1m/U80oStUfFDrf1e
xocAmKYhVDTkkXJH+mO3nSeWf3QBqpZ/w1oesfq72KhVc/NeBBBlpf4dTLWFFDIO0VtQu3tD3WJ7
Bz57Mwe5EnfNYuLiWxpusvFqsToKvPR8Vr6OJHY3M0iPbTB4sA1Famuk7vpdRhgDQRjKoBvsTmfA
oXMN+ljSDycF30RRBEkMnCjbN7SdecJ6XVQmoa0er+bW4E+hv23O23Lu9HxIPwNNOYW32j6LPTbT
YWWOntnYlNub0iDw7Eysxly+rQQ+GDDMghBi6HBzUy1ImXux0apo3rbnXeHsyuCLOR0rfWixG7KU
zWkWk05F/W3hcqtv1hPlrfijrDaIwultqEOds3nY8ic68a2X0ctAlc5GgCtykoyETjazOMJtcr7W
TnETC2rYc3Wp/lBC2tyaUky0DcIxxssmxX3gvajNuFjvb7nzXXjwF9O4iyZoV0f9B4aoQpgX51gs
LXzISVpPutA48t+QglONxmzPwtjNsFu5F8IO6XWC4RkiKfCtwd+WX9F192xwpi2t7MCVUDZZmzg1
9ZFOw7/ouvheahzYv6hhGfNVcFBtVoPsuvTlylw2uXqsObQfAfx+GC6jODVZm/XY4LYlQbx1MevE
Gt3Kmd5YNU9eb1OYfKF0fbxRN0EHjr0IbTMjUNJYGq/wxlwmFxxjayLhJedyoWQhOyPk8NDyUuo+
UwL0usfLvNE7lwXZxMTSIwFq2Im0zungAMTiFSeGypzGKeANL/Y5OPDJ/Wt3nX3cYaSoP7XUGi+z
5hpFM95vglLEjfNXckXjJgnvgZ7Vaz1JxfkpJ6YV1aUhUGaZ7cRktzmNzN0pXBdTpwJBPyp5k/Qh
oeXJXXvkOcEx0lS83DkX4OQHUDsfZ/IzSFCvGW3rwQ2qy2/vwVqcj8iGyv1GdJIjAnGTMSt+u7om
aqMO5uHHDDCBZFSaMyxItA5rMoGi+FW8NA+FCsVo5dALTFnit8oEBhxdB+xnfciuiX1o9zIBgccX
vhfBleh+pJ0kvtQCPW0MxGHLmwgmxJ0XpKbH1XyHTycUgBNzTQWVqUePjWVEmZ36G5gqX2bJcOM/
LMy5J186fhDCAWyjpKzhHhivuC09lmj1NHfw0Ptns9IxhhqoIEgDwAvzDSdY65SiOx4ju3/EwX/X
P1uEk7ia5XjYh8FMqYBLbwcDZ2mCZzPu88T2oimHVB3h492kKYJRLiHWWvB/XXUGrGilroUFkOt5
VbHGoLjFm3LsmAa6vczATOzE1wZ/ZQdVw5BGPchlCLrv/u5NgDsgF9bhVLZj6AbVi7ck5DzaDXtu
AllHxebmHWtEareHLuuao2NErb1ZbaHkf2ncsSq5cUR4oJCn5FYpSKkgEbG7Aj2gSUkfapMdpiwt
sz/fJXV/DoC9lm0eN3DbmFZyR1cnwueFMr7dMLLbAHN+9KXVNkOiWLiC/JMHlpSVT2ryBx3QoIBH
NZJLpBowNiSGhh++6AEYaDTcx105DBRhV9w07y4yL5fbg3w5NKbcYwqhkU20KrgQja8g9jWp6ThI
ZaSTvIyQnjk8tZZCl3mkuFZ5GVleK2BYAP86XTJn+LG4StGX+ul03vhnf4HejmT53VnS6u/TjcSo
IWJp/+XLopkOp0hphyoHjZzeQTK2mti253KrK4jaeMMaRCfjit2n01VfX00NXLwnnKDuQZhgXmwY
OzXw4EtO0Ucyz0sf80Z53CvFqJlLIizRHgo8UW0CIThAcxuwFJq+pIglRPk4YiuIFQMnhURoHlwh
g9QRR4wq5q1k5Crrwp6creD+BCZ69A2CxTGtkQXuWjnDYDKEUJbcuOlerP/UCmaxi8ZGYGe01egX
OB7KK3Xv1qedl07wimXZaQHg7lHa0dIOMbLb7NzeLCb7yuxImJRe0dQLrsEPH69E1YnDQX+9S3/X
ZwssutNgUkx1UmCBFxCEk7C1SesOIVN2E9wbbE8coSjnGYX5c5LKnbq387tzft3ShAMnneb3Aryo
qElANu9BJF3HrsXx0xpUbFQZs0ARC1IQ8xSQeMVoi6ZbMRdX+Bf9n2b+cmh00kwztEyP7KYkMshe
gRJMvB51ZwPGM2g9h1mObVmCsce0kmi+era5g3XGp4ZPVXYNyuDph2upNaQSI3Nf9LfjwT96ArED
+cJRZypTrTzsw5Y9XAxSGljfX9oqzduGowipxNJxTqi1LRvORoq9FMaSPLMfRRJPD8OxomKTZG0L
3gxV/ywMU02nMSiYcvkKWtwhoyOdk1EtZTuPI54NIUO+FOM2Pr2S2vCP7GTxvGaUdRPqyPOBgAo4
Gv7HZITpHSl100iAOgOvc+uGppD5BAhQ3y8MkJe7eEkgHYMFjyNehJOyGdysxLISSi1/CBl1cox6
cbpX88kBp6MJdicUwc1euZ7V+y+feLupuiRusC1ffcURCcoeKnPElX6uulGI9wG260HVtnH0K3JO
us8yjIE9+KvTCH4B7Nx7KMHLOqeq1BBC058HrTtCGGUYJU/jh6fMSd2vRR/NR6ZFurpTR+BpyGTo
8NzlfKGmrgeWkCUx7DRwm2f1Z8eWIARvtNeTUwl53+G6hsH9HaCuQwmXIOqtHJ29FKMQHteRMAZB
NVt8pMJIFy12aiQCrjpNr2A3tg21PCRqdXpxaOQMyFnBbFIF5b7UOzJgsaf6N7TZTiqbXb2PaDJm
/KWAEOqLBiYFsqloqDTWtAeaepzDkmCbiUj8aqAB3W7SsgdrHCo8TVnxgWLeSm4y4fBiW9pW9YAB
JREjoBBu+YuzjUKiX8emA2E68/cjpPEXfOvu0RbjRYMbc0sPasA+NZKNxqGu6aqEhI3LZHomauyn
ymmWVLGXxjlheI3RDTrmbEoWe6V/+2Ub9AOgB4aVWxyVlPpqn6yrYpKKxEgC1ztjJdv07VBjehPC
8P+NepzhwzrwtEafQIVcgJc9HkzOxtWpgVAtMF/4Ncgtu7owiXG42EFWDvjFXXlP9/x2WiGVWLK6
tdtxb/3Y+Y0z3QbGSuE8kB47Vj2AG6iDZQD1VtmPsLMDELXLxruQKWREZxEjGXK7pKJdurqIuZS4
Ie2uk2PctfNEMfaEr8vAJjQbGODYZkWJZ+I07peCcORxRYURj+bh26PnXBdUHew7NU07jWK7IMWB
omm2ulFClluxNkfyzaeE019G1LelC+tSy6Cjd1MMD18laqev2nbXPsJ93i0BPRyQVRH+lHvtN9NC
+UxNW8Frf9EWCf2IfswL/0ytzNiV1ddogpMalBsV0pjjr8FKqL7gnX3xAFuA64u7eE7WYwtXRM9W
19RVym8oIq701bR6fa75+OAIxERbB/nbZzacovHppuzwjTH+vflAO4vZE3DE0AVPHvRPjmMuRJUz
8L8PRFMB92VUW++cij4RlSdGGwpWL7cjCS4ospkRfU1+/C53OvDc9BNnB3cCsKbq8OEBxt9C5l03
fkyxlanydpaT1wKWjsEqJkst6+XhMboONThEgtUt9FvXr90cmHeIVqqvcNpwD3aoiGFDtFH04lkl
9acN+rH8AzJoT4SH/6KMSrB6kDcj7gUc8W4jtfHYqiL7dqXYb+2aA1JlSGJBOd/JMWoO2xuwM1gm
L2uDEYIR6a3Cy15SA77njPxGO9Z361atvtv2dURh9uvlCAGB0/pSz2mSFdTNk1zkUZoRGYWb/Xpk
jkYeWPUizVTHVa1F2MKBxoeM40zFTeTx3SxjBglPVb+4QWgc7WAlOmZYGQlxatMlpRolCwibgKoi
WShPvx0/99QP6hiQ//C6WLU1SKq/gQ4/5M8zZEEStdknBphG30Qo3fxS/qhY61JZgmK+iowbpNFL
YmsFGzPkak7qtTWlNlK7rCOBEKiOW7dsCaeVfbocSWx5mnf+qxAhZkqoF7C740bvxtr2g1MTlR42
O1z9b331ve+Qmyqr4B5lyKWnTyZBwVwliac3s9ABcJkpr+usqkwnwyO0H1ljc3srDEKcbLI75azk
pYfk+OTOqbe656XbVsqpGI0goYDv2vOUfZ/0BE0hB9PZirQU5wS6fz3uwRXvfMK+Z9Xdlzp9jYOO
FOdhPpZiEG4cYmBNIhOkxuPBuuIjQ7N+t5fanpJAOV0B/qQ+/CZollwWA3XgO89P2L97x/DhqRHS
OVUiEOfGynoqVWh4XxERLHAaI8I/9phaEwQkyu//sw/I1LTO3PnWdOSVmHxTzlV/Oqnj4421XHdK
iXl5yHIVNiS10hSzyhoduDoJ4LJLB+LBQ4E+CUUqPKyunt8Ta0wSSxdE3tE+TvYyeLBR2OyFE3qT
NYUQBmcIH28ZPhR0KhJiyLi+EZ6ICa1eRKexN0QexoKJOfb6h+d1DHdhgbhAwEY413t3AL1y98w+
dJQo7oScUenl+ShbCMq1SW0NE4dwtOKh1Jh9YZy6ZM3EEPegf0DxSB65gSYkRqXmL5eqvRXqmTD+
BQ+aQpffidVGp8fbzxO2WRgJo1cr1VRN6C+g8yF6x8wUfcx9mf7O0UkUC+28XEi2ZBd29wbxZE68
MMMegrLFwnFJwqIMrk4h71nwj56B1qGXVbG6ilo3fXfoWQxU7cnL+JKxaiG12ntFzzdaJrrp9K/z
Pc2S/STGGM0YuL9WJXf2nUq1lr6HKK5HqaEXE/eiW/bj0SLyzkqSkvTFX+G0dHFgPnde5T8PouBJ
c/YgIKsiir1TeeTUWFbs0MA3tEEgvBNKud9p1LcKkUWbTXhJGB334gGP/mo4UuleEpEXq8Nmx7Kv
UopgP0IQDGdwbKiUTFknh93dZt+YB9taU9purwHHYBelwjpV3ZsdmL6Bc12xZvRr/sKd10NSCfN3
jDSDImJHW3ojwt3mAWd9fPSpkkjProSVgt7SSsbe1yFUMO5j2/6+BQi1dxuIvKAIgkL08jAjO1BM
Y7Vxda+csAa8nL/qZE8pnAsF9ZYHbkhCx15ZzLepuGw04X9WN/1a6tc7QTwXXt2+P1XoTG3InCBc
9tXvf11X1HmOniGNa77EV0EY+HAbq4PGunlSEqWimTickvkqgKvrISngcrKIItPFpydrIgnGqVAK
dJf4N+KSwnbaMyPxN58VGs0Z2QBSF2fYdnoIurTRHRZFAeW9YFgd9LCM6GNq6qUU08A2uAGyM6WI
+sbp2n5zIJ89VCGsehe4x9uHCVp5kaTrp0GhTI1Won5Q1ZsB5GEJAhUsIdoc9UjXaj6WJ8hxs8E9
fpUTZNkBjrEANUl8vbdxU3kL/1833lMVfiWH/+rc8fsJ8GJ2qdVcB4F47PM0rbqrm9/uwAhzYFrY
9C8xE1WvqGyXxqwPNiWVQvgzrLfUap3KIbH2Jqzobn36sYSGYiaG1+k7rkXINVZWPJXpbNKHoqVa
P1xRnPAvssPFbHnauY2RisdDKlaZbzT4x0qAcvIE8f/DmcPtM1Ex9kBMothAI5MSxuFMaFUYlH4K
L1QPkH0wb8oWTqBO0VbsWs7KdopFb1S2AHPw48SeP3aTV3jJKiStrD5VTE5keDr21yll62oAzZNI
aHlVeFAL3ZEqp0LktyUsSyEW17qTgCI8k8h1nHiDretStP0NSAfHO0MuYqG3j1W/9wEuTiQBtCck
1ALhM/5DAggUW8q4lcNA56w1ZS0uABqDRU2euX8UGweuDoD9v7pTbu04kpiD5OOjQhyv9Lcf7rQG
jC1ditfVgRKE8JfsZ7fE37142F+JMXBDNnf5ET9DncovTlgl4muEusIOz8QIbAZ+ma916LPEkWv1
eXe+bE7adCC5//o38rHXWE0mgNTC+pk8Zf62B0wc2xMjJPJQJCrpjuqzgt0q+HtsfSQAPri218sU
dQZAdvSfi3MUmlee++mF8TULMLb+/2jnvMIoUszNlMernIUnmtlQntMhnGu9tXZBWEPlC2JSWAQX
Gd/yZfWBUMV53/T38t/PF8zZt2lI1UzvjUGfO7xdMEXZSRLi0k+JEtbe3nlJroJivNiTbDnP+vb1
Kc4VAbx3LW14bvK9xAT94of+kO+BTQXXsNvC792AFyqwjHRtcBRwNMaVGJgVRJIjbMmJ4gEQ4TWi
Al8S3ym66LvJYduDdntN9dyp2TwhxdyQgnYGhSK5yfb++CHqROYcfpLCHoLVwI/+T7s+F2XvIsHB
lhazJe9uz1AP1DhXY4JwS+NSU/VP3kIok/p8KfYvr9bmBsI4f6G9TIVa2xdG+50t1PzthqRvJ9R8
I8c4wtPmJIFBhpRfstjx2RhjfNr2wVy3tMZBR4kW8Th5m1Vke5pvmsmM60bRUIDlhszif8GQbISF
qDDFx6GwWTwruV/t6/pfnmXPhRgmMX23k4qkipmLXNX7WQmszgn9e/WuXgQEH02qwnK7wXturt9w
6475C0iDOPbG73pTdJhtxth70+LuwPH68uIappVYCtE43FYxanS9khlN0pztNCINeWYN4U+tT6un
f0ZNFZYAaqDrS7ai6oOG1pJmwSAyiCuI6823U67YvevXCw+56ctnkJxfiBfROeOD7PEyc6qpLXZg
QZHjl3aXVKIogVnID40xvDsqJQbG500lxmXu90Kykug7fICHrcdtbWxle+D3194fb1wJd7dbv3ek
71Ez9tiiN+jFSvCU/2lSyQ2Vkh4XFAxMKUKX/mz1tfis7195IVJhGfan+u87bg+AbK1D56AdUFHF
NulClO3RiPWzZuVx4WVpJgTCWoiM+QGmEU975YUKStPl1b4upNHk2OKU59/ySpFVX1pqJzXClYqo
Mr7X8Y28n02+UgS6Nsf42SZgK5OV8wJ2OIg4zsw427GCjPXws+c+CAFqX0FhbtkbEWolmfCtf2mx
s4w4msRWKH6uvp75/sxJRY2AVYW4p6/+nelr10dHGUkwagjJwci2UqBPXbhHx0Ah5HIS0Ds3blXr
kFANLfd6rF0C7r3D/Lmjyb42QLkjIDiryNV5BcqTRHmvw4Bfm8zTPni+06nYsUDeBaej8O4FNBSf
Is/NGdb07oQtfKg3WDDJcv/FYZC9go+2quIL1C+CpRj3IepON6uahR82p1q4BwwEDeI+bM3WDqA6
Uc63jvJUTJFWWR09+XVbDUoExZjwAG1r1QXIycBz3UAl5kCpziKmEhYiso2H58IUjFp1o6Wu3SPn
LgU8v2NpPl3X3aEnRNtu4OmsckmB4S9RrStO2fh3J7McczJmiR54g/AKnGF9B/v9NSmAoAExUmLt
H3R0P7GgkA6JgFCLGM7pZMmRZ62VzkfdWPZedSWccekI6H92EHgrXsVNKZhDsg/AWTBdBWgMrgcB
64A1/R6iEBpDPVsY0+7/Sztg8aC/+o/THOuyw7ZkOtFIU9YfooAImZZInRC8COORaJ6zE0U0tHna
kIme0zOqIOxEEsf7jIJkbitlH2zmkrDUQsUbVpKKJnFxye5QbAraMN7vJYtqj3jojDm0INwQSIFS
AA9y6Cccq3RchMpFNDkdSDovmgjjGrXBgt3rhZSPC+wx1keXeAvTSBwCinL5uD2D/4lBa7XXzxWk
SQf/3YYasT1MFrG5gc4DphRoqXw3eafWP/UtDVEnqKjhpykU5+S3Yl7TpTxRzgDpF7hi5lHoU5ed
ejn6f1a8MW0NIaGpiIpiJlc86TybUZK5S4A7J99p7egNNf8d/zolnBh5mZFdjYlNXbhgOO9h9Gbi
B13p9KxC3L4T5ofJOlQLx0/oYimoFDG1oJ2LtxPKi2IyFRyxvCeKahxXFspusRU5zM4rl3eAE6x/
qNOhr/MByAcsn1ANXx/E6/A3gkh/3dEb7RiZ0enI6zeF3qkqKuLylGOhhy9IGPJNVOX2w3sMptgc
Z0dnV7z+m3JcVql0ZT4I8BrpN4QhyHjDKGN0W675CncYK6kXNqC0dw/1fXzpiAUBy90nAGDdoGue
u+vFUyFGamWxCJxYNgzBA1sDQHd0/Px3p0LmI9Dbd9ZX2p2IYIzC/RcwR5Ey6ouXo7/6yAEUtiJ+
QD5jT1Fq6dqL1N81cs6Nk6yXGaHzctfOisHoE63CTRhBi/YYChdaTZs7Re++OxMrc7zQgvXlu7/F
QXfdJ7xRrix8TxTUJL+IB+lAjRJ7hwCyHOC9jJWkody0Y5xhNzMlLSLjvU4kphGQtmqMqmQOqZBU
ZMlGhavt3+EL7JXZGxj0whD/FuZmElkhnP/9ZfToOkjUAPrwK3I2rS38BJCm8LdEHw8M8plny1fX
pGEdeR6/PGiZ62XMyfK09CcppcdhpOzdy6fjaDqaQ3KrXd7nrakUhoLZAtnJrxG85rq7UzmAuuNE
fKNeWSoHLKeWj4JRAdaplomFeUvIGfL+MYc05Z5QNwOsW6+xHGjraFqFlJDQxcqgpK6NfT6r7Z9g
9qf5FfRFFMWRkYs/o++Fpkx9UZCSvGai2XPP3HJzaqrtG8kKs+EUBr4NJeo4Rmu4PSDMSXrpLsgq
15GGfnPlM9sVVTEfYVjJVfHcaAB5o41xj+YIlcj08Un7KfudN4z2e62K4SmGk3jPdCsskGXD5imA
VS2N2VjUPD5xEHpBdkLmjjJF/4++fo8VOZSdYOC1Mvut3B1x+qU6rfKVXJA5c5i/epDvqyHKQub9
gGxY6dQzaH/Mzc7Ot5mIqRz/GIWlLKr7Wl7KxpIKBUj5HKbRseVcEUOYEPc65D7JusvBFDZOHfYU
a2YaE/jtdy+YZNHfnxJ1ldmh/n0oeEDyO5IfnnhpniI6gvAsHznOQay6AdxdgCyeC3hn2DX8nw/S
MUNgqFGmFdbNmk8Sk1IQSkV/N1LeX9mS0HArIXMNEcBfFlO7CNHc7C+vmDrTNxAmchh1pJoUsUOE
cB6ifhIjMFvM8O7uWB+prPDh5DA0p4CTFwBs2jzEf9OzMXAtMzc82m+tkQ/zltZQPJd19YVC2LQ2
UzVS/hNfaxtxwLuXCf3tfX43h08kU7gXfyPBRj1LygRg1Ph66F/Ak5ms2YHgH6zq7r7yOKVq1evj
rmW0gIMsLZM+m/REbmpwulRZ3nt37hi4v7lbcb2J/HJuiIq5/J5jMSwse0eSU7+nKi0ocesgpEpa
snWWIyLdPjDl6EV5SXVQqs6eX2SyzaVKL10iIHk4l+tzQ4UhSo1a2A+5wXosgZtENV8TNTd7f6hM
kuVGcSYJAvh16CBv+/eqrfB/wRxGXb52kMc2tQCUTCx0yJmLMj29WuXiQ7osuVO5e4/2PRr8KlYH
TwVStM5lyFfBbhNxzKWKV4Hrsfu+VAc0LXIIlE/DIowoJ2xBCE/8u1z6CeFFh+nkPhvkBklglTiE
EQp6JVtX0klZ3NUY1/4oeaQDh+4+MymTltWV3FOzUITwqNmsx1OZeg92Yvj53NtbNZrHKwt+VMyU
wlbsDlivUXhXLOIurWTtt9WSJUzbthhXVBa8TfLImIUyGtLMAY/q16KK4s1+Ums4e0yo0Q4bJ/LG
37acpn/+nzEnqWqwg7TkJVipb1fmS1JiNbPWZl6clucpmIN7mMUCWzxExSUvz5C0mKQl4Kw1XxBo
dmrwHmkfz1o4juheJ/2d8awK/lTNeHFu10yyjeeJ8KrQgGD3xYEGRpqJmV5Wckzjt0hKGZA7LK8w
0texEXhQdxUcAzwlvJ4Dyz0Nbi2tAFjE1lHRlr8m+zrXrlvaej2zp3vVEJC+yGNgiEbVBxNen5xF
jwNKgT60aIms+83LtSFEGGnQ4tqmCvp3z0MEog2AyH/MmLfQUj/Y3qx1Xtthu6dh/oOP0jk99eRO
vEjgyGxsc3zmNSZ4epQJB6uHk3Rnpicv2VYcAKCMNro7zBQRVL7CcOhKk1lr3TwgPWm3gZWqAwLC
UvfeNLgZp6hfitG9k/ov1SJv83swE+TDTy5d6NSXwd4ZRPoFUv1jpG83SSPltLHqe5REv6M86dOZ
r6zEO8BWtdBlUdRVdyuKSGc8wmv/v6tAFQ/RIaCY13NDpQB33vITQ6ticC3goKggQUzBD+0y6aX7
owtfdsTNNvPdj28HWOfZjGizdHkDJymwo3Mzr/QFuvaUeRU5vHjlwHz/FhPNF4qAF/s6/SamZ580
X3FqEN4YypdVWujLP82n+7Yr4887vpWmOaH/H1wWoTAg3RXFuu/yVECXrdj8vovx/PNhrzRgMyxQ
iF7jlQ7WVp5knV6SCuSZeNLKSldbxjbRC9jFu1xrwsD9iMZ72nZC72NNR7R9bKLrX0w8RJkfzqju
pmc9bATl6PZV7omjZUYC8kQ2gEJ07/IQRoo7RKo3cL+dI99PQdEtoM0NBODCy9svinupJv6RFV3w
sSgIfqqCS5iJTSil/aaGWaUDmvWbY9bBK1PHB8MYnWL36zy8aGQKpD/2Ky4fRcTtsbciBb7lzBkP
qtorzZTtmNnT1NBn/TEbVDii1svmGc4woTlan5sRMt9oIAcgLay/hyEbaekfOdjaSScLslCtaW71
TeS1yr3wCaH5UwL3Oi36O4ZO05NoTI3Eb4Yxf7wbmcNmru/8fmOajpKYQ0IDsx0/v0L7E2WVvoaf
X5LnEFt9jhFSn1JzXOMGvsDNr9SiYQG2d4NgZaGbB/BZaaOAeGFcxM0u3fQSBp5Ipo0/gCky9myV
2pTuVW7P0K469AlxS/gS/nzrWPXARiHNasSRwbMm9yCMzVGHSKBCA9jk6KUOJf9vz0e3vpS/fEKT
2RRkr+1Q9wE31K8L5jvlHHZa6Sh7fdGhKWtk9P9M/YEQ2Q94cZExbB7b4DXeo+YueLpO8A9t8V0H
RofZWGOrf1a5XCsnof8zqccYL3tEmlGZccHcw33uoSMswXE08QJKjGq0ggs8aTMbjbkh/heVCPZp
R0fQwv8DywDLD9mbQCLStWvv4yvLz5mgz0yD/K74as7En8P0Pw30y4A7QCJHwEuU/QS92qtRflcf
MAe8r9IqU/JwUk4IZtjDsbyAQ4oWXeZPeT9cT/fpDZ87dTAnc2MDXbyHUOPQrZ/LomDNTbmGdaTj
MSHt2amx2zVG/aWU90FZiTAeoYa9gAtbV3XraGlsYzBrfA6w8FVwMyil4TKMHFSjLfkiI8ffclU6
4aRcAOabbrn30Xv1y5yzINaMyzpeAr0A1Jd7snryeZwieC4Z9toomZOL4N9hI+0DECGTgnGKeQ24
KoAzFVy2aeX9WG+dEyAm7FukDW03l793dI/RJiZMLa2N56exWehxQ7nWhLyXmVoFDqKutdMDte+y
xGtcdoF8hXorLLyJ3k4/ovTPb9s8lzuGs+BQek5QXacvL/dWIEh7U8dajK4hfXHcUEe6EMfTtUJ4
oBdDRlxmSZ4kAUfM01ky+vaLxMe7ad8WnS5TFTpvL1uPV4w/a9YEUdH0eTlymIcFLs0N5QUJEvbw
H9Jf82gwhiTHjHeXA4ePlpLoQp/McxooYH0vc6o9RIudinHiuBNwJvVTfkIf8xvhTYziv7PHQfjA
kXTDm6SXUfSz3yc6qkulrOkZECf2MEsVbLNTeibljlIg6IVHs9Q19XRik+QrjBTWa+6hZTQ7sPKZ
yRXftf0XCVKDhtYvlM//Gjvi/SOLbh7Zf/JM/BvUaJbCrjXcMv1jfqeLJYWHFXHC6VjeeNGV+3pc
TYLIPiuk0JOp6ldZBOPBivFI7gENwIXi70mV3hT+I9a93lAqYkm3Z90NFSfJZgqxEOfJRnjOklpR
naK9sdL7iYM3d6Udu17rYVF3Y72bS/CNHQG50WtKxojGxHEzk51//YJZ0PDU6CcndV/5kIZEYEta
9yZueT3PpemjfN98sSLSbfbQf47B1kczyNMh4lxNPOAcOCGTtf49/Me3MTsfwu7BkcKi6g8PbV2u
MoEfRjmNtXCphTlSoSiYjE4AKKAFFF99qlE7bLxNtZpQorPJob4WtxvLzrU32yq7xGN1qgG6SKmy
l0GldV5iwUed+5Vox9mI5Ol3/Hk/fiWa1ojI+3D/E4yT2QA7uHBO+Mb1VCJHTyPwc460EYIbwJY6
2MikbKnCppAirn5gyFejWfwsu/LskM7cF8uMu9DaQIiZ4fb0bCje3oXaf732LVw10tqaBgzYNngp
KAO9z5uiViBG5KX2wE9HmtisdcZzFH0fsCDiySA/LJlUZzfwo73e1s0nZzBMokymu1o9lyMEMOhr
CtFjndIcf0esC7pXW4KEaINqZSxlmC2Sfvwin+zonRzKvqzcdES1y+WF3kY+ZvTTqbQO+zNa9GKy
s7q7UzvzQKZkR75uHZJMwE28wKAam/t1yOXhqRJZm5mLamQCV+bAI6G8LLg6Q3xRJxiGLBs2g6ic
hoy8v8r5T0SvgX8FTQXO/gq6aZUvhylaqH92Lcz+wwDOjfhl6aGMq9G+FgX3uF52kCfO1AeFKkuJ
dzM9ISO6IpYEsqzSn/ImK8bXS+hCOtNi6lFOQOIetH/GrPVSNKUlfbptmidk1L4wCH1cULQYZWoX
IqfF2AaNxreook96AYkuh34T4+s9QkgFmmtLcuoh8aeuXa9i/wHZhDAmwZHOCkr8O5Z9xazGf6Dp
t6+3n2irbY2KSV4VOTQgw1vzcfcUGFe+E7lpCWQ2CsRV/6iGqyjm+sKY1TTqCnRUcalH+K0GLO+8
klu4EmjGjBi3xaxcLTZjhCGK6/akIwzsniH5xKfLfo7tHnxIisLOs7iqzlDwpHDe7yQCNBiIQztR
W45jiwzAl7fj1cjdi9RLIXEVdoabH2tlVKmxAA5HYS14G54GgCn1pEfrtOVAlmMx6rnPqiw0FfSo
c4Gux9VXPo/HF1IEWR6ty1GwSqpv3E4QwbdhJMZFVgG6sv6NziLWyYIRwntimi4smifipO70+0lM
r3eWgnUfYLtpUT9RSbk3kZg+aD70ZRxJr01NteJLPKRGwPQQiUSeF95S5ih5RP2LOe+6PTA374Q+
MDWE99dZ64+u7KxiwlZAKYRk8HRv0ZkYWeyLmOlhMe3iZ3NGH9gLkIabF+D4phkHsCInb1encnwd
r4hIgRkLgntullKRmq1RA7OchVCR8MlG7G60jceIRA/XX4rA6yeLLFoNCW+ZOji3P2SWbFnUHtgd
+Jc9lK/7V3Mu/gKmMqoEFm16O3PAuMzMc9u+dRnrqZUqs2ogAGsjxBkwwk/ztaC9qj1VQ87dBQBK
I4qVwlLI1er9TP6qenByakwVc1RPz5TLot0FGP4b4bXl/BPzDiKSUwmzjpaU9kC6jsEVLovUT3zN
Q9hnEUWBkouwkJHk3oGW9dhJASt0vShQSiYX/3i7DlKqKehHUf4nlR/XjHmuxyJV/CthETCFXWWK
ooyV6f1bVwJeVWjfKMaQBPC6FOPEiXE9/+WZiPEkGF56DYZ3M8phU5RljEXvEn8MYyQXRuE+VT6G
Ja7G7NkhL4NYzLCIkieEc56chnRHz+3ljIOehcdX8frcZbDo4N3U9HQAx0QXMKnRTnv/ef9E8xHC
IBc7UTv1bP8V2vIJe5SDkufS7STMgVTpJP9DrYxSjAw5F4dwMTLgxUQKnuE0xGfVLgjssQTJ1mG9
spVs2y32Hh7j1yXYNgrG9tlBXtKTjxEVo34M+BqypB7dcmc7hK6KKcNrYDa4qUwV97ARxHemUiqA
f9Y4/WsCh/Q+M8SbDllPK3gmht/20bbVs0JXMkeR4wqG49GhD42/VK1CB3cbC4TO7ZPVq+dKVSaV
gIazvfYW4ez+qsMJ2aIl4g4D6Qeqktb2lP3hok0szVFYGTij1IwbCrjyPVPbHUTXN/y1bypoPscJ
Xk7olQDL5dfAfpWfK/eBwJUyFYdQHv6i4q9mqmlXLYbVffXXdKuDEBhlY757IToZpZ6KBgHHlRKE
BUzd8JGXRHiuXBIed0Ihof/P3qchsqyZsDyF92om/DrcMNJB6gpzM7DKni7EYk1Ujvp7KXacMYPn
bfTTfjUZDz6MjM2LpaKGuPQaYT0j2MF+q8a2+FSDWc0pUqBRDfkawG9dnY9KOUzypLzx+lDq8jI6
2T/L6o/D4UjFRimsT4u7Pp3gcq+JJozr2CagOYh428C8hNJ6curzECHvN7tfXkaGOQ0oWYUUAflN
Am1qqKKW2KaJ9Bq2JeNlcux0jnwTk3Z3GaxnM6XZQB14x5+HY5wtW+rq2J4PloJdTRAp3/ReaWgX
LFhetBPk8pijoEn+jrFerqoaExW3u0LLbVPxF5TCliGjYHGYtad/sxhFnBINNJoeLTBbDa3vq2/6
mN5zus4KcAtA0Sybejt9a53mHC8aMh1BFDYWXYSU15Gs6slNZyXLEzxDuzZu6gPAuovsgnPzUb1U
05+aaxwU97wvAM+Av5aQmTWDMXqJaSpQIL3tZ620SFrvrL3a+y8mEsHYXamgvG8084iXX4mOfF2F
IO+A3TdkQcgkoH38yqu2Gxt/MM0F5/efnsZklF8zHbNAU1LQCaqETqh8l2FB7yV0TViBGqmrRyXG
S4Mnrmz/zG98MINDOnNfKKOjTuD/w/RaHl1aux4UJg8YJT1YFQuF9svUhFbGBDTdh0xHrsvefjUc
Ibr0dKd9VY53jCMnPR9TdtOaM0INLxb5kO7fIcWFnmpwOBOmC7jLljBb0nhyfeqb8oHkCLxunk8z
/MtWjM1ZXhrc0NHyJKTvqORicRXqtP2MY+lkVR4eBhp+A+vp/ffhZXxH6H0EQCHwbM5A5iSdE0ic
3qFs1Pqod2s8pc85JddwUHJcCMGhArJQ5q31afvAXNBuglz8pagcmA+jkAVGeahxqEau/NokP2r5
jFeYI1DQvCfzm2qU/DkjWrXdfJeYgwwBI1WCozJeyZFBQN4OpIWU/eK9KNvv/6IPRT+OEmx/EXB0
fUzBVuRgMQCG1Od5doLj9fs2zxPJgJo+izFFrLk6CO3WilxZujm7fV4mN4Y0miF9U1PKwJ8Z5TAj
9Ash9fCZE6VY910yj1RTjBpdUpbkwKvNWBPg+ENtP7/q7ItcKmUUoV7MJMUe9QxKEend+s2x7YFu
JDmh7KLvEZ8dty7TBDqyNdBaH83RCQZgwPai5ePbypu895ZLBCNFNWRLAxeV9PTEdG2I5LNHzPKA
QuOQ6Jv1C+oOFOQGqQ0yOCP0YuuRCAvDX9e1PGmCA1y5TtSgmDk/evEPR+8aN1o5mZ8TzBY+AzN5
tiyhEdnjzqH5/2zAq4bLXy/xFZcmKVUoHCDHDNFckJlGgTVONA2j3hO4aBqHQ6CV68TU/fsN+Esl
FAkEEtjZSK0spIwzHgVyunBG4dKcrCKjeZ1sIvA3Hu0qqzqVy5cdBasy1bBERgUqRb8fCVm9keLz
1NKIQVe1MpAg8rOMfTx7Ex1WRoL9A8DKBPisUjC7tov8a6wG54cQmvfbY2VFYxWNxUv7hOgVUpL6
WWZ14qs7HwYrZ7zSJwA/UAEwvZItsoBB0QD+7HI8V8p8ZwBQW7aVNM9+MKn17imDa79zRj+cDO9x
/kGNCjcHhaaMbg15kgjNyF2n+up8pn559qX8zQDskamVjb5Zh8zNFTGvGpMJwU0qCfYP48lTyoZH
MaxZm9wOefMhYs+dVTIAC7QAonNle3O4YtHGy4VSZe66VJW0qi9zayojUioOYMvmrqWwtdV6tpOY
vMgn5VF8DluMWJoiYPROZ94X8kfg+kz7OH/SzATcQcg7KmDWS2xxpaktxqPWhm9ybdjDfQuMei8b
3Vb/JaESEML0/lRU2C1l2sC6+twQJttyrR9reUO6iaz6prHYRQ3pvpPXS5k23YNSomzUntXeFWWv
hl6w/51NDoKVsBDz+b6BSgw756gbQXwM0V7NwqlwdQJUDVt4BBj2/u3SblH8tsvFzvgXBJJlFV//
D+xD+0bgKwCnpOb8+D6CPf32x/r+qTP0c8Quh/zH+h+AN5uL/q9yo+dnTxTQw0xoIWfCdOF7whbF
7wCbKBINtDCmz4aaYegxf0CqahlCHkv4AGMk9Opl0H3RthLIbim880PE2cvJm2s7OreTwfRAt9Nn
UuuSdw56mEz/DxsDsrknuEAyE1XeqyyFZFLueuw6dFgz/dHvB4uGod0FTix2SqrsMvl93YfIuhSN
LL8QjrimEauaTuGRDM6iEc3Q3baDNdyK3sSICn577KXmI6t3GBmuF5468BaUtbhYSTtayk4T/KEt
DR643GKnYDX6aGkLjJRMFSLJlgIy5rgCbh14ag48qj2uqmZ+6e3UC+Wyvf/2XxEpMiuDHRxwVPyT
Nm2MAI94HMZaEVHE29F01wNQr/6npb/QyjayDYUDV5IC5fxn4J1VH0PQY3kyN/GABonjvA/sI8RW
fhOUQJUaC8BL8rZ+dfX2iR0us9zQerjX5MqMtgPEVba1oLRcDuE+e/IDqjH8ALnpS5UHKQdtqini
uiiPfG84kDSKw0xID3zfGGGV4EyX6pPQ98lmTTqSlr9k3hzsgVTMEqJzNrxPRsrN6SBnJL7Xo9aX
mAV0qUXUbQF1SosQg/JTrgSLBDdjWJhAYw+5z9/4cExjrVcseJCUMMHeZwciGGbYiwPlaSXnMXNt
rRa9l7J6Zb0yRiEQy0rssFJYdUQrp3DC+ad9AAxtdJMn+DnvFxAIFaAJaZtK4iu+/IvNmnf2oKah
cIvJsK3aPUmQYGL3qap4347vaP7/WC90dfJacsRoXHwFOyF62ln5TCy964ZUXgd13QSnbFeb7x8O
gb7BAzR7LAXREP4eTmNGcdBh1SOwnPjXqd2oeruIo3oR9oEAFvWZ1OGw6yP/GpUBgNIqSTD+vGuQ
Ds5z010QNK+ehD3BAsox7kiUzETCi3Nr6RW0TdnD+nZ7yw5puxcBlPcCyI+iTy99RbYQxB5D10qu
6dT168Zye3QUVr14Ug5wP9xcQhb6+1MbCVy/Sa494rlzKwbxEhxpWF9e75t2USoWuIBQu49c8I8e
VzfueznJeOoHTItLOaeHsCpOO10yGIVwgnPQCT3Dk3TViyWjqsmR56YYAQxdis0WAoZir9e5Mlx5
A1QMzwfJ/DXqFLoPBmHO/fOIXX9xGICTwNablkpuLW6fPsaUW2DcOfy7YvULQaaMXfbZD09QH7cM
n41mg/Mxvm935mC0jkEvInHuO9qe7p2YqU6gA9urTrEyY2gVViUIYB6aCEOJhko3+cUbBR1KUOLR
yJgOgBua/k5TmPJd60MQZ3bMmSK/EGqZhNxDwjD4GCMW3+w6NXoxsImT+CXee0a7X6/Bq6IvOsyw
Ptb8m3ueGEK3xES1rln0to/kvQkUcCthnekxb1CwzjJtlXjDwCV8G9J4oVoiy50WcFcW87MpKzNy
kPuEM3rp3uXOIT8KpZSXjo1V6EN1wk4ZEpDiVCyAZPzh7mU7a5WOHxTMM5SzZ9zn/RKPJg//Wh4I
Vxcv6jTPi4eOVsel0dRMD+1GRtRG1ilh9ZSBkBeltDgT5TEAufJPKaVc5LQztiJcmpvHaPrahwyF
bNAGZQrZ1LWthX0/IcpRIyLc/cZ6uqpCYmsveffHiTTYZR6lROO7i32zKxy4hjIRWHIGzMKMT0fx
6GnVy9845n1VslRL4hd1KPPhbGfoOUNgRWaB0SdTlCu3oOyo3eglhGGsmeZzFO0G1T3jbVf4gHoZ
Di3Pgbb2FGPCjyIA9ElUxdqkcgSjggwJHj+4ZN6EIuOy22VCHaMMm1k7SP9OfOi6AjEOY9A/724M
MfzBbzqwSW2+Q74eBBCqy8LZ42qse+fnBLchZg/yfYOu65rxCXd31iKiKdI2fWwzrb/VKZkO4Yv6
/dFw4w/ewivLKtOejMz6TeEN7Tmjem7hSxwUDqSYs02C6vsSrtHYuhggZuOoYT8LYbljwlkNVMfM
6H5XWx1Jnl23oygzg8FSjnE+B+hLTc5eFbAhqNmQLjdFQ2pelIePBaqETTl4LpS1qUb8hYFBIpDb
8cRZwU50i35REU0SeYhXsnBgHYKKHudi9TAwEzoTN7VAUfZOs56dF36vILy+MIMi50ld48RKpS4c
1s2dTOZrxJB7iEBwFrUkeBf2l7lUYnrM+LPrGDvbgLso5P/6qNGH1qcuoJKUpAKHFZMKH1nrv0E9
Es98Bwxq9J4CdQlFCf1qA/OXFz0QUE9k5wpEHOjgGe4da+BQdt0rU120OIA+VjRjT4mQtnnbZ2c7
AN/7A+xlQStw89ExYfQOXAtjmSa9P2nIAV2bnrdEjLaYNe45GatxxElUWS4qH8mC7A0hi6uMQYgC
bHirh0Dic7g3Y6A2u7FzSyucU6UGmZcvmb9MzJwhKSAHN58gHRqQQzDJt1AdHlHeFZVy1kdOmtqO
2FWTkIx7qgDStooE8I/Qq5+2M6i+92L8iPkF9BPY9SQQ7hftZ3vrwlH480DDFI0Fu067GYVYw5/4
kNvhiZWcKP3F6d5OJojwaddyD+sjVtgQDoqEnv4OD7XVkLiNGRaoVlsMvAmQojgRIp1Y0Pwbb0QL
14PuP3n2ZlH3bTZ7dAxD9l9MFgWbW6v4BNMgQmwQwt4SrrK4Ko5dyln3dklwIVIQjAiaoPMGBgfg
uEcKMsMe2oLdRTU7d1yq85SHpDtZ3MFvOObvsJbjiFjCzBxnNtu5d6T36ZAvHUktV4oHKKVmloM5
cZTI9jEQKYZf/UVq3Cf/Tvc5GdTMrObNNo3c+Igdw1MmuPLfQHWUAvBp+b/ccspUdXeORKt/iW2X
jodDbMW3AMku9tZ7HOdaV41oXvN8+AfM9iG7JjKvUGBP4I3B9U3d9aXk3/hi86Jbsu3EhYqejoAY
LO+HN3n+11LkFF1XLbsY1k481Vjz0HwUiTBQAwhNw9x7T25xwSKHXnwOh6dxlizInC3OoHemA6Ck
kzWjp7CneFkJajre3FBLHgpWActqOVw/cgUNHWrbfoxQMOU0CXG0uOONQObgdOddXHH+M4Dwg6rA
NRJn7ow0FAyHbQOga8Wner+K2f6stulGN1cqhEEz25+7KQy/33wX9Vbe8MK4z3ENGNj8Jofcxzk3
cWEr2FeLVmSLVvfUvE+h2OV2hqGoY6h68fk5xu0J5D4MbflR1FlL71YNr/MUzd4/F97ov7ceSZSf
0X7kKjEWW37ReSJv9fj5dbTNsAqTTj+zeSXQ6DhGXz4vmOVRTZ82+lmX7bfnhpUVyVVjSNnPWTIQ
lzQjV7hePflu/9N4YIEJqjvtbMKBgINi4AjBAw6f+rVrXebWdETt8xIY/sD/rkX+0jdxnwTVVCPW
/FfRN7CIkIPNRqSPcPROACwME7qJHOisE/is150SyGh4Z0vEqYoDF2KzheIYM85s/VHGjbR4BXs0
PDdn+DjsU46AhPcMDE6pq+8lmNEarvlM5+zV5gO731ukHl6IPqzY4kosMj5Mtp3oO0h9ewXgmxvs
elf2aemK6hgVobEev+7EWlGtVsRzp1WPb8oOS5GfZY7rAZ84Hw94A87uQ/TT6oCrADRC8b+QYr0U
M3NzL95SlsXOXX3MxL7er7/jytv+AFad+vE1kNBCKxIvGHpntHE7B4Da7ikaqjhgwxwIkRUL+0wa
wEHePgmkWc++bPQUO4cVUZsxx4Vo2a2OSa/6IfdpMr/C2GTxUCa7ocQiDUnDQXEEEiNkFdQxuIgM
PuqWimr8REFukEdbgZzGodLjE2xfRjRjb6V5Ru5aKD+vnN+4txQhjxPsLVjW2Z5MbI1O5yklMdDa
nF22L3CJ+HNpzmrN/ezxiiioA0aCHjoT6xzTicj9ku1nPCE0K5tvYuvlCA2RmL8Oe5Vd6uaqCY9P
JF1xoMiH4ydM2ASehjDUq0OGPHrWs39xDTzEi9asmq1FaSYcKo3bP8/+viTrwCHbO3W8/im6cM/6
yFp2uF9d4inid8Cq+Kp8RQW+loNtDDvB6yJtt91cGRLEehzfjxr8IOF8Zd6G49nI1y52OUXybUWT
iygFUPYSGAG7x6Ct7F0IdQtddK4TgHDDk4CpFeEjmbZJjcYgnoCKk48nCyklyc0Vr/s2Z0GGy5Ai
uS8HXDlO97DXSAFsNcoF1yaHiqhuRcw3/c5xerK1EvjrtuT6LWY4C7KTZO2JJ9iC8O0DqQ16TRT6
CrVGMM4Mdi+UiXGxTOqp0ryTh4bQmYili7IU1rrpj7NhsRe5z9fd3lb0aiTM2qb70D/TqXMl4x9B
lbWYtScvAbrARM9FD7Ztntp+DexVfucjW/9qgzPXSuO8XgwwWqmnJoTyWng0jJL92kKJyiO8+1AF
AJftc2lO17EifGLbKO+j5Nb0vinhIm0y/S4ldZ6jvpynjdJHwCYel6Gonx45nXvZasntwM5PhZa0
cg5d3GsqBreGoPayEQdhTBLxlXNF8HIWHnbdD1gA0T4CpLFWQ594WznPkyyoZ1F3pNeATevDU0Fh
2GOaVARMFy7XTDfMI+ISJvlbKZzjpi/VXkcwfiqTjjfMV4aDqDMrnyYfJ7F7DGcuN4fSZ+gLrBbB
uPSK1UeK7XZ0ydBe4e3m5WO2sbSQyY9IV2Vz32/x7wGs0UhrK50/pK64kdqi/892J2TA8qQPFgXE
6k4o94thBDgORa9wbr3Ejr9BCljGg+4UA2xZAO2eTd5YR62W7UFlskB6bV/1kX2lEQ9ggCgcLH18
ktOBwwjLu1KvAQIe4OzF+Monw8S4fJAvoPtBVKZO39IBY8vAiIyLfd6tgyrYptAcZTh3w/OEwaw7
dH7+QaP1nFwXzYCVO94wrumozZ7tyep7U5cF9Acf9TxXkOHavplxwkQEbU4u7kZEopaTYfvnUPDz
TJAHJoF0H9O8xfaSYN6h34SeNf84b0Z06F7J9I9b8dxXBXD9Q7B5moQiJ6pCyUJeGikM6vfaPbPl
xkgCa497uNnPH+WYlui1Eqj8hD2h4qO7Azi+yOCoUZ7v/N+k581cGUeHDTrmvSkpVQNadgV8nih2
fArQph0SVxjjZ7Z/VRgXGxQZnquJFriHgufBsBdG0Aa1GYgeD43BN5kozsj/zv04fMYrRK0wJMza
jdGJgZbEMHTDV4jH/lLQm9y0VkTBFVE6WD1KVMQzN1qLM0IkOZSBlPflQ1BPuYo9evBccVmJFe4Y
eK16prriJIWUHYNcjyoX/CFF1thDfQkRGG5fs6SE8wIphsVIoQQpWYHGE8unKMgqJNiT0N1OAG97
kl0YVLecvVhh9LReDU1Sf5koivZ657m4he1h9pIfVc0EPV/VSYjC9uOrIqr+FLDCE6//ZWWk8UCm
p/D9lmyL2G6oTsG9KTe3OnhV9iOE3by4TnmBUzxEsdicCPoW3jBS0qReR0Pz+ksdIUrLlcVxD90M
W14M2kPezOgJYqBFCcKop05tcv4XGyOJOOsxct5xSIWVqJz4+k9p6fghnxzcBkBghFajf13wNamB
wM/iBb7iRpdgtORTpnF5u9SvmEXr3SUD06TYAGFJ8BomcjV1dimxh+zhdxq2Nr3wawT+VLplur++
Fij09wcSxy5xN/12HFlaNuTAiis8qvOINh4TWD/e5/7ZA7fntWYIhJvwR4+CH+GF1q7lKWLrc84q
r4DaLMmdheCkTb2wbYT5G8Pb5E6YEMRgSwSA4c2yCSUqNPe153WUOKWfYygx4zB8gm7fAOAsO111
kOvpBWlG26hoP1hnyXqaNdi5bx5sTbGtOZSwa4SwM+v1sAlOEhGPrk60N3q7dsYztcObnefIG2FQ
wliyO3cpeqht+1nSNJemg+rwkqYlGeg8p3nj8PXDXLe0DU8OokF3GYRXKAE0Ren58JTkfmMrMGOd
nAw9twLkqsCF3qv7IitnfQFPpqhSewQxkiCiGPVFQUWpVRZoMwOyChLDV3DpJ7Rc4g0AnobOTLqG
z1hmxI63nYUGfWE9YI7OK4y6gdkkPora3uQHQpOH0JGr+7R8QbuDqnuiBctUK13p3ET6/6cMgmB6
vhly31PfzcQOb1JsCyxS73DTG/E6gp9xR6/Y2MKGlzADIcexkz4el6/VVhfSbYO2ruVnwYY+67zL
0aPuaWXMZMx900npqdhBJlyGAE5TOg3vmrTOW2oVH2y8iURSOln5nx3eJV4Qh4yM2glNfdKuoyjW
71HnVUILKRsHgcbkzHl3Tsl63wSR6YFbtIhN9reldbwSdZk/UPC7F04hx0WuMuf5kw7mRIjNfTe9
nunUKMEyz8ul73M9Ut/Otlfxvquijw2VdWhdXbE1CwaIbNaDvJincoErMQNoYeusguZyM6kMRw6U
4OMiL3C0IUNegClWoPi1x+RO0uZKoAkDMJvm7jvLPDig8ek0lX3nMKB3es4gGw93K4pqquAdBPRs
HTEefO/Nfy0hVHHhwuGs2yyOQXgs0V1LEqsUgmmYH4egXtiFfe3ZV35BqxdIuCGk0YwH2hNAilVx
Y98cpue07IgHICX2nzq415R3A36kykLgP9jH/hAVfgMlBbrqja8zd+mwyG+RL5whLat9XzT5UR2H
E0SGrKSvg8EZrBf3x4TU3PciB8qy5atop6PPH4CggSEgpSciS3/RtwiPWkBF9eae3r1WPP2DG0Xk
WcZAgH21X2VCdHH6OUUa3oO1wVwbN4rzF4wXN6zxVtwnSmaCmwCizc2MZXK5WPgJ5/TYsF50xI8k
Jez+nj4aphKfn2knOwLcGK0UUaWaQ97LDE9jK1qdUwyt/8uOzBlR7TkXrG0rIGMVBu+b50DxQRP2
EUImzFOiRGuhr7jvNf9lL2hMOWdlAxltjsi3hBRiAUjsFEJceX+/nISzMneBpm+Bo3K8wPsFntRS
KpLIbeE/mZc6RtO/4Eu126mzPGM3FiuA5DJHPbtof5EYFs8cMtkS1tISu1xKhL1Lyuzc0I5pd6GH
ErWEXwjHZtoQdLJJK7kCpbIWUIAzb8F1BbBCX6nW9Zw14TOSSFTD3NpcGkhJuzd9dG+4wpFHR3cc
cOKL/Lcfd8aLryNE3fKbbiDeKDwB7WQizZOR9sYwCo71M3xpK0UWhLHoEchjdahM9xh5ctD+5sad
UMsUfDrhTWIIvb17blh4cjvrssRS21laKeGYghvJRpEJRW+VJ8ld4PB/+sVGsncbNl0cmFGsMYT+
EKJt4KMqETi+I2/2nBuKAe/vsDzBdqyctHD7LEU1TDcEIGlY52OKi0JqLzzfZenMiNPTZgoaf6NK
jFU4/1F5McgzVaXury1X6pPc7kFk5JT0f8XjrgTGHFQ103uw9jYKHCBF+HgHb3mLKbb8KgM3gVx+
bHxpd09Nc5bAjs8yo76sV2trzcmgw87R50+9fldZENyir9wDwF3Oti5mmVH1B30ms9TLO5MUJP3b
IYksXJBfA4157eol/QMSEp5wkIbbykXoILb/L8qPmMJXsx/OPC5bTlnlp3xmDyMqHNk+QgvJA0wH
YaXKwWBOSb7WXAYWUkdWbh4X/tbbQ7CbhGoShiaONieqzZ1S3riSLYMkhJQSss/2ZGcY+NsIeXWW
F6OPWjcQ0o+PIA0lOperQotpxFfOyj5Fy+YrXo6wEAhwGkQMkDNYcVGbFm4BEZ1YlwrCeLt3hn8C
fmJcmHSZ9V1Meu0tVNirPokp740VcAPzau6143CeIY7zs9W9l5HT5SjRqXecFKyzlvEE6q+C4AZR
gOUk/NVUXqEtYUg1jY+tdkwZqwjCNWy3SDVghBrohtFGZvz/LJAKPaSOwQ5zveWuM5QfxaqjtL5n
ym3nGQAsU4cZxJNyp1UngGbVHFtN3zOb5ATPZHRdoUq50vezSQiUPo3yxUxOsynaRZzFbld5L6eW
ioayNyZnXfK4BGtz4pOaoryjq0p54SWjywzbrgNXZ21RSAGPKG+rrhmeJG7E+NBzGPgO8TYOmZ7n
DV03g4sA3UaSx0YtUfopy5eskioj6agVGzEeVleljGlGNwuNGu+kHDlW0xtOVhRa/ostMghVQLa6
ZBWceScR1T16Boru7iBnmU6ZS7/gz44Lc4WSLk8Ca2KHISusgQZTvljKYoE3Jg207tRTOlq3D54I
+I+1TvhzMeSBKWC1XyaJjeaDMIB4S0UkFM5bwCqPd0rMnNoBH26uBHdGp0mojWJ5qHs6tqQSNHx3
L+x0gdE1GSBHQE7iwF082fosLARVGpPRrg0GLqKcoNk9DJFpGqR1iu0/M6qH8LFxHSMouwRGEgTv
dyiSdVl1gbSXmfetzOe1/JLD/8xYrMRKEWd0iRDTaDuLN8mv7F4cmRua4PKxJdW8o/QCFOn8zYKz
OqByJg4KXeDYQGoe5Gy03ugRlpmqTw/KwOmpLEbkyQa1iHBhBA34qDqsZkCKlGfzzVq30dmttMrp
PXr14IHQzwhd2X+nirJTX8VZeF8SoYe1fdLtwHB3p+RFmDOWkbLBY0mL1gjrtyEexyst7Aa7hnUI
1FkuYfcRiWjAd5LDn072aHE1WY6Kos5uUHsne8rH2mRPyMqiUOreXm4Q9uhLKahxlUgBlJVa7Nlz
AATvYqv+FxX4T8RQr9Rskqxh9wd/OXPzXMTHYviMH3hkj9jEC7dLbXBzxTV4UGQ6ZGALbT2BISgE
9g+eJt+5I5e2vwSY+oNrQD5XVcIL+grxm8zFBa8jOFYZ4mWc/1U9yLfqc6K5b4AG4Ph6petbd0qi
itikvCq1feBx6bR+fndg5IOa/6xQmxB6zmgu5I3+eRGkuh8pIz/0BrPJcvONfW0PjUHsDttfL/+F
uRGD12LIhOc/GRnbgBoUDnuhmh7nL92aQbyUr8+zBX9/Yi8y1dUvUbo/gB9WvaotnTBGA1iNnZK/
IlCSUZQu3g8qeYaF790Er3uLIAB3HG0LrhNbF00ZnebGIfihY1Y65w6oc1qcwp+DwjzvSbMJDkjV
tjS4s5dJZHNxjaAZUoQAJeWzoAYnYp1uamyqJm/B14KpLUx49iXmOepRd9EhDMiAru4XkiceaXDy
TN40IquJwAubPOKPcKqHvLDfXQ+yTzYvM5VDU2qOK6i9vxgc+Rfka2uYpxI81+R+GmfU9CQxhdsp
JDm+1JpSCF/XkfisL89bqLZMPIcmG4yesg3czLD/+D8RlCDJBI1TO7NnkL3bXWMXd1Qz+4dVW3TV
jsM+SE0Y6rUaTajdCMLjJB8f9qwshtMgbLTFhQmnDPcsXEc69AYhrytPWNk2GP5bmrNk/XDjL/ZL
Jm+NUbxOLjPcDUOdAcJDHcLsRWYUdLuOaaUwmyKRamgtDqOaq571/Cf4ptAfGvv+U1QIPY7Wg4Bj
QCxPYSFMFyd2Gt6VS5PDxFFn8dS6h9d9OQPCFfhoUgzqRoFGRzETmT2xrW6ge4FEyr+BaLWN4mwi
EjICFE36zuB1bh938oZf5PM+igAw1vEXF8Wq/ziS0uDgzgjyUVuo1RX2M45aEAMsH4sIpanL7pi9
KZ7SEA3A4HDXaETdk+oXuG1kJhlwoor3JbZ+MNl9VFhy0EG5mPCRp2nnETArssmhBWyFn4Mg2LTo
rPauKIsYWSHb6AuvmSGk3nU/wLdsulXK6e5fKrGnOEj306ftKqXdOb+I82HGIODco/tbcZv89pWb
W/ISyeVtjayZL1HTKLm3BfUQJ/6OjYYnrNN1qVBRHbGJ6atzBC0+N1k1EHnfalxegS2FHEoKCJUP
31yRuJD62ISySzZHBDOS6ifewf1F9lIQppYu3CZR1nDolqdk1rEenPcXrOatXbeZtbKmS7PnSM3z
sNXGMEzNCJTlY5QhPY5sVnTcwoaRp8Yk6YSgXf3D4dWXcPzRWxrJ47WPqIfw+mA+EPhkniZ7s7U9
z3u9i4TjMK6LzVUCmKUz2Gqv4zwO9i5Kvvs9K9AdfiF9cL8qXI8zDjVJRfB1iuAAsZkv0YNeYjYh
mXmFuGKDF1GfhfH5ra7m0LAq0T3eHdNvYncGbz8CSGk3ySYOyoeu2IDpQa2fWhONowRi3HIU6kSF
O18xqXXE5ni0/UOkq5x3X6pgtHid2iinioY8hiTzpxDHmpKmXtPtO24a1rUjTqbJCoOoycHaXVE+
y0G5OiGuIZQEq1EhUTn0MnX10kah5VLwsqAkQ+nlO+znw+qk3vHKh9Uy2SXMAjKWfgY3yNJJnnXS
87DKK5KqtOVXgU7J904MTxf5mtTY+64Z5Top5DPhXPWqeYMPUElNnP2s1IWtB7a7XPgMsOqzhMMS
LlYQKBk5TWzNr2jHnQzY5OCxBQSZsiC9IGGxbUZgqmG1PBHeYBlLkOYdQlJdkfD8ic5JPyKOO1i0
VsqByJ2gVM6YOQNGtn6wAUgQwmW5bwaxv42s0qHNoNK8085zmhnDQRRzdgliYynKsfsJcz+XS4LH
zmiPwLV5+46wT2BTHINRh+zxkQE7xJ+O4uIDTtwxpBHNjFz4Msxkizp8hHxnTdYApiJrkmady9W/
L8PTGBLpu9uXLjUo+XKjK4d86rKf2KtR3nZbuxoRYJQTX1eMWz9WYkmJ8tyrbG6GO1Xcf2gUwht2
GYryKUEAIoem3MQMBh8P15DmWFvnsrK+WO0hSeWMfTkRUos6V3KsMqeKO6SN6gObkufealzN0hXe
DkCiTSzQMhgdugbHF8JHCR2/C7XhNiNA8FtbG9BqP/FG61I5//KiRtf3Pgk5mFpua1sl/eetVf+H
pPAMxPIqTwNOieU45rZz+hz+7loeMK7IDaUIyQKMpZAS2e+H5vsPvlzoa2QKYbgyxnMeMIByesa+
EnsnEQlQXhrqPYwMle4NR9B7XXYDWOQMFdoegqQcfAG7dCWYWXrNObkZj6iJ3YsRu+Y/kRAZJug3
NySoxZcugNF91ntgkejeH5GebDYb7YS+hT0xreeLuZTzk5269DxIm4CR8KGK2I3vJcFKfE6QctZL
wsSiSjyxIfXHnqdfNZwBSUg+kLgtE66FIH3av/YuUeQPpwTIzJgGUDXcvwugMXbMVUwovblqyXWv
ouZUvdRYgBywQ91sOCILT767jgSlHmRGGlcNjgenIQrlvlSDZ9NA8R+gIXIn8fLGTcLg3pO7CI6e
6lGzOuqczh5HphcxdKPGrEkrC1KZK0zFOKqXprWYMK1Z5DHBfnQQsagYKHvFeJQU0UlSdkvRYEYN
B24XeS/8cCNAVrn2+ISBeXmZfjK0krgd+IQBxQWAEgKvRvmmjlOklOUiv8N6ZwdhAiymkAh105BI
t4yLbl1FKm58RJ0YClOP4ZaNd/18pDkpPf67RunE70FEahAbmzgqHP+PKvdkBWg/1oGRDswIQimE
h1smQNm6NPZ3F78D+1+V1CMlbtiyCtWrPnZ7Uw3gYdmLAO5//MC2yhJJPK28xDPak3HJpe8g3MOZ
b3gjVC4C77fE+eOA90WruCFhkkZaWOlG+ufF/RnwAWkC0WgB65ZEOulnVdBFugHnLL7c1vHk6yzt
p+Pgdvdzq/juqxWb4PnqtVIF622SPv1ptRMVGX99sHKsNXvj/WXXTRAWk2AOZC1S/ZLySULjUUTk
pq1c9G22vjpmLLgmR3C3DykV8NvieGeqjrvPxHldDmVfeiOD1bqRquCb/P3W3EtaGPfjIr9F7/ep
JQzvV9PTprYw3X8JgImQPEzv1BvD2bv1rIpjrhl/JJgh63SSfqSN++ieCvbK1R/QuFrshUQulCXh
dty37KoSguUMiSzoaLMf6fC9++zUlbED6qu2I+KBAkaRyz/ijfDtvprd2lbAUhVminxjxrExUKPT
3U6QSEiHgd6J+Bg6evXA1oVxvKBcjyXsaW4zs1bkjSTj1drO1XyZ6YJ6yAzZRywdtd+jkre3KVWW
EwGgBl2HZI6SIGBN0uMXqhjXBstdOn9KF6BEE9lM7vs81nx0HIlqZx6AMOu5+TiCYh8LFuvj+jVd
lqKXMSOt59QOG5FW3wDoggtrksyPhxMOfZe7P3gbt8ZqCeEu645fEXJtshPk2HYo7LjtPfeTyDTa
fwJkDcH9VpDRmHCRQTK2i9n51VE0n9MQZFLFfypZCry5MrPkH35f1n8n+rj5KdORQa3DtW8niWPR
GfRi0blK0DdN7kE2EajnWTv5P7oM8vwkJofc9Kw980Myv6G8/P7VxeBue7vqUwEhZJl4f7mInbQ/
WgH9Aie6aHRSNeBj0Kl+MmpLUtnaUQ/7WnGthoKzfXVzYFJpX3Xdwlj4MpdKnIeEIDcn/7Dj/AjX
Yh1OyjBJOeSvR60rXkkOKygAB2LsodB2VtyPHkD8WSDOnzfm71WMmzS6kgL9tabJhZ4OLnop7uIr
a+mCncZGFH9DNT/Z5bNEKjSbKcvohhaMnDKYeJqP7Wx55HA2FUa2ETL9zDVK0TnYP4806x+fLc81
zmrkwAZEUiwinZ5lmhWU8hIUdN9dd1LLjEFd9DruHM/ixBPKP6Prrpj/EcdoKZEkgqsLa0uReTO6
l8bYMhkYJ7g+aZBkwa5RNVCZfIOSe+TOJjXifjt/SXCg+CVnSWXYi77NnjgBritw3+XiqhpSiFnF
EbXtZXTTK7PJhv8zYfUT3IDYXsbekgjtcMksSnBEVYmTOwDaLTzD9Jy1gAblWExb21hKwddOPgNr
DZrzZ3rchyg1+w7/7JJUlPdisX7xdRz/w1BLbQnIZhxO35tRISJ2o2ohh4nioZgHSEPmPjnEcsV9
HV7C7lhTP7lXXCxDtNXJpK/KdeXgV2NkKvLConNgGIqejJFm6GyXX5HtlRcqQ85EZkmEFfrbE+/1
nfmHTpxbDUvoXoleGOf6Bzzd01K44FQF1xdD5Gsby2NX4+0ZGNqU5PjZgeZv8/NhUzQ1qA7qx604
hu8R6NdeUsdlE7Z7qYNzxA8xfTrul3j7FU0zJIdkXHXM1/PF+e0YQnE5NX+cPhiIdFXCEvaWh4BB
zxtvwZD4mSVZER/FugOTCuRrlMEhSEvNde+35SVIKyfadXnUXoeE+epOek5fGIyFWxjyptF0VA/E
B0i6gSfUtnInDvdRdqgNGKj0Cf0eJezRlOePrgUH8JKtYIZQ73N+ELAk8hUJNj/pfVUeMNf5WC5d
+1/O0T+dcrIUmToWMV087Nxuw+vvs0FCsdd7G6DBTjhVwx5+02OMYNc2fIEQKQft2dIDWxtgajOZ
nqWy6lBXMXCBPlM/p5dTXlr36VVm0UOLdCltqqskeMm2oME0/DHiuyShkBArx+Jk93ahtKRGfDuZ
hpZXk9Gf7l3KfGF/WYv7eg81ah1kYrdLKsJHX0NUDf8I3AvMVibsyiFnoKz3iiXm0hoZWcWibmfQ
twYvirq3KoPzQfyGnII76wvlzjtDl77wUqdXdQiurcMO5+2bmwirqG8lt1dfWhHl/cviOXd2yqIP
9cxc6TGBSswrJ1N9h2alJi1bWrTpbEJsxVaU15EuE4KRF9KF0lXhJ9PbmLgQ2Rt56IfosGxVGlmP
ZGpvCQ5XnCEyjjHGQQc4mtoRK7b7AqvKKXCreIKAx8tuh2oXo9SwTkzyGgzaBFdrmuEYnJ9/H5vf
0wZMkiqtmubRYPzIPIrs27vVdYWjlULcXovRfsy+IxtKC4Te+LJsTc0p096vfg/eVdV3YAgU99yg
KyELLl9qu9Jq4hvfDmo3rZI88E2EXKxyFf0fKQ7g2omC4qg/s+tpIn7533aoQw1PUhTVjPnZoU3v
uxnNqX4IVWlw0EHlw2K4RtU/4Lgg8kgB1cczOZL5q+qf74jcSlejnE+0u3Bf26GoB3gPcQKkRtCy
sPpsw88yTD13J8PCeKWB1ehF/Akdd/KCWaq/DEpHQ+Ey/fWQW40yOLY5/jgozRAnzNmK6L/JO9MX
II5Mfo2Q7y+1aFb7i5GESXwvhfVSx7n442owrOwM2FhXty+smCnPuAeR4jLFsMTJ4M9589u9/d1w
oVuTmBQWyWU41MnvGN4Z19z+KCI6m/a/PTFzCdgB5Xbi6IwpmuGGPt7qts5vqAtVsATRDJIxLxMK
vfjCMJDSVCrG6akA3hgK8O8cVVGQfY5mr2zGdpPNOYnwqX5pA7TgPTJvhJyVFo6wvqg2jMuWazFi
69q2Ez7lzl9f9iNzdyWmWzNXG4Nxx1AQIqbvqCgrVAuA3EwQT1YIP5CcatQS/wwV+XOV0dU+BYCE
UeKthqqdsuQ4xC7YikKyJCWQiqB+yXHvkT5DYo5h2KuqEW/t1yetPGl2Lh21qf57PLx1E6df5sCo
e7wWf71C9LZCij7Ek/CZXAooIql9ulpTXYBRqxOpvKcvQtznYlIjH0fLmXSBC3kB6hopKoGIES4H
/kj4IntFAQITZ6cm9Yh7LXzhKGLdETA1p4JwqVilk8asAIvMWXtPtAqK0GRvhmkz9cQ8gRRaJ8WH
IkTnXoiEubGpz6FXRFjtwFJZ5rbRVCQQzZA4+dvWokplYrrJCoUE4vrYeKf84t831PrvN2Y+w0C0
VFV+/AtZWdPMsYAKRTpGivQCyFphCE6kUDWMboFNxq3T4MiSS3AN7LiZF8N7yrC6EBvtNRvWXT5h
TlUNao7a7JcCau3PyFodrfUqgoRndVHEDW1cxlJNWx1NZScLHUkc256rmLhx04PZRnaURfPXvlJM
TsfYFp1aMYbHskepVsXPYhUR2jHT911M3UeU6vtsu2edkdMnWNQ/eVMdha34HzaxtRH7JkxB+H72
OzW3raRdVHvPWR7L/GtsJHN3gJ83IH0tE9/aaNZYokxhwDNi3455ts86tGIdjFBP3BI5T83qyd10
W4dr2ZFfOPWq8Yd0FkVNj59pqdfN5LNxdadPn9NGR6DpENg+wxfL3Xz3OTu0OOCrhZv2lpZ34oW7
WX4olaEmYBgCaPsJmJVYaLJoUsnxjR66dBymF9x7qDpHCQ2wF9kgFrdOsr0r1aBr8kuS2M/yYqbZ
5irhaKZWkmLh3ScwK1xL52EW4l5MeDflw2yHaxbbw9bc0R03rNELKJ3yJAFDvo0hE5ggto/K3dwO
+efjyo5OC9s9LxKRR4mXBeGBtd818YdDHOQk7L5TuDihZb9bVreuZh4rzerICqTXxs4kxydkZq4P
SBiO46b3cgnanb1vetIyhepYt0SUkLQFnJY4y6NmDsxyVd5aFAsyG+5gg3wqTuNQQePs/cn2kyuK
efs1ypDG+1mZY3hVMq0UkHxvqPJyauBVYc7rYoAll17yqM6Q0QP7wNdpmylbSkYZmfKp6i+5QyB3
G/ROIihFEWppFYuJCrSqutI+EYvfBRaHkNhCX9hNgDqj8+NSdiAHaV1EFPowso4nRuMR3dcD6zaS
4/rtqa4KO50xyJPUKpdwMxbgD1qM3GWjjGN3mhaHajz6nfadWPaM94tjC7pnnQLp/BfZzd8o1n0C
jYzXyfQVDrTXP1mw3XnQVnD7AKEfVjU9XI98GE+KQVF3Ld4/+xBwodMzqRTQDC/yZifWOqhRjSZt
+dDQmNJEULz3HTLmy5DYYPsyx/8cioi57be7k70eCrYLuV8lXJ16c/da+wag8XXd0G43odnXb/Z/
IS438tOTbB9TlddAQTdMjyHDYmoBnas70h4GjEsEwXAV214KPVhkZXQzRPf1onVsRsC3beDcUP3S
Pv0t2q6WQmkg8Xd7Euohn/Zm7lKPzj61vZJhfaIWvpDvjJxg1gH4nYQxephZXEZI+v/bMnl4nd63
NZRi+u9TzCnrZhyseNbDgEVgnljqARl9fCxaUUJPOmPlApDSLYbEO+vJtchujXSABNcso720fe48
XOJFHX75qNO4fyxlGlcFyYhgVWMRGUJHixBXkGrWiD2C8N9e+v/r8pzaS8KVgR9rBe2N8vIHay1F
4ne4CKdQKi9+YsoBgJeOXOXcp0q5V6vbgPyZr4bBgeajY47DeVW4iJarcWiqtC04+orRd10H9HbR
ChRyaCQE2BLPcsb+3HDXJggP+OTvkuMmfFFhdz0O4j7axXIH2hcfxiWrxsuw4HPObnffuEt036p1
GBtvh0c7QT8+xIiAoITcnoJnmY/J9j+0NVzIG1b0zSNWRczyyXP5A+43hoUI0Cs6so/5qy2X3a1g
Tlj4vDLrymV0KXnF1Fu2H+Tmi9PPkyU0wr0+Ni022Wis+NUWvlIkiXWvLeXDH0Ay2VKUqQhDQygD
KYOWuYWtrj6kMQHnX0iWEWOXIm16+5SxJO98QvGuuFvvlqJYaeVcCqCyI+FmPjfLYyr/zSyJEk90
X7pVY04kznlD8A7/NvJLgKxewzpjbIywGFwqhgBVkLkSS87cKWKvyk3RhP1zxq0iovPqyc4eO7Xz
WJsDBKNTi2zYjOHzjzvY2cm/EwIFLEhNAHZTwLPO50tQjWjSmYhvclL7/M4Jcz25h1JCbvPNmFf/
HlaqRo0GXrcF4K4u5E21Df4npoPjqtOCzvvs4GlDP95DYbQ+6OnxKY3N2P137e6uY5rnPTZQzlXs
8rAZM1qmc3h6V8DrMYQxxjfKvkq93we3Y46c9NLPrQygs8xuCbN4Y/Q0vhImlYSXS/i5o9XM/tTD
BhVuIzyW4hbyIWuLIEFGUrij9AL+FJfYt+12voZS3VjqbwaL53FQg07JD7eY/WzBzNIHVz7n2GyE
W/CHkNWZXm0GfOz14jv7rhh50TGq5qtX2wnAWb2ZxKIlVIDAeLWYEH8JLbOHezzobnJ3lWzBl+tG
WG25yH2n2wd9S2uM/CwPoCgaRpcPLIAb/ditDcS9pWeMgutAapSt5vEeFKU8WIaylB2LBjNi9GJ6
rEloN+rUYcfgDox7j/zlb6FvzAlvERv5MGWVQb+544xKyzcSLKSvr0wrt3mSlrMB1toKzadXwECM
oAE8WZ/KlW1gYp5Aw7qxqxmcD1C9B+eWlocuBvkH8jVDchMW5PgSDwuI8aQEQOlWimqLUkqWIPX9
WfW0Osqs8Ya2gkhXMGNDa9Vvz8opkgKmqikrxCuCPd3ccQ4CWsG242WyUQSbpPKlazxJaAQHU0w7
f8y1PfhAVAHEIK6i3scOPpDrN8d90g0eYI6TIOA0Lc9cEU8IUibfdvggUuSFdvsSPSesiHHgk3QF
j82xbk2iSf4WciOKUEygOwXGN7j8Ls1e1hg9/d8XBvXcEDkVYuCMwVGZNZouyr6DSEoOys7UduWb
5ot8+u5EBqT9ZmfbJ/BjZP0xU1QB6ZF7ZR5mhbkzgueb7L0QInzzG4zxMb85xR75IuYzG/XUBhwM
Bw4BnxtQ3zOd32dAvi1tYC8O0L4e3WHlSH84vpTLtNZ9SHgjddBqvrjq3r4H107hsN6PvYu0Lw/g
j8h21CRSGlZHS2v/cOT7WgIdkPzys1ulX/PSX8gkzMl6QOdT7z8ssoEfhU7lo6E93n33k4xCwDFE
B22Oxwt8R1crLGL5NkTc9dfkK6v8FBsdcDnzMETgOBfjcqSzLw7fENIdI84V5yLxe3ET9t2heSj8
oP0LutSKmYdexbygLL/jwfjqhu4SuPlbQs4WlOTgYDTVgfk8k5fUf0BevORjU/mSdLrnVgPzJ0Fc
gUdwECJUr21MnjB13DiKRMlKoUTwCcbYsK6xtqwgELGs3GDP6866S0QuqEwEvwSJp2xNV8022Ezj
XFc31fA9vgKEyGO4PjStvZtUVFSDS3IqOlE0k4cqAVb4+yqN4mzMdpmStGdVRb1Qyt/RstCE7AQS
5YsO6JrDL1zLBfl5m9aiV5SIyt3v7aJL50KvQkWg/HA90+iR/WNEb4XSiAa2B2Rn3LDFyYtQXNCY
Mh2H6CqvWFibVuiR0RPcepTJt7Pn7RrMkma77cpaxVBgZwBTFQCt7mPQtskm0XS3D9tZ2KMGvE3Z
7xjwqaRa4REe0SWy6Hlw+7qsOLOzj4xjRIyzGveHeuIIgpLX/4esD1Yae7fLeHyuUdE3ucVk2UIU
1/vXXbHfZSZ8p3SvtttGj6pmHU4dWkTfc9Au5Rj/Wlx+ya+vk2Uqf2iSIsYK6Oe9g66PSBi5Xirl
dUkki9bzmJ6rmD8zttbIMVsq6tA3+tQRcdiAYH8GfVTe19VHTKu3a4qXruzZs2UWUh7RHHsKBnNZ
SDp3VN3SrJgY/oxo7lkkUsp2dV+d3+4a1nZF/tvHfhB6LICRHt6M52xNvzT3pKsUMH3MUPL7YZcd
OfzJD/mz6WD3l9HBvXB2glFwn/aTjnCDLcNficCyhldLzAb+fw3fLy00toxrkfckibM+EGoqMWWh
AvwUpkJ/M5Vz3tWDmi5RTulCtXHa5l//2T/TjgDhc7jvD/HGViYVPiuSXnAcNsZxfRrPBcTGc03J
mzF8qETD4+elIedkMXLsS4w7rIUt67N+KcbuDcqP78awKllqvi/bEEJownwTQnn2mvdlNoRGIH1N
xejEari5GNIhfQd/MkQEY5s1mFj3xANshfpwMegp3aZph2CQgD+X4NYYfS/zd4nluwgTj+Fxh4zv
94yp40M3ffR1LI/qqjhwjDC2Na0+ShRR1FGNSIPOaW/2lEf2uwrGypLZMrnO2DkQtGs/FMeYzx6t
pZCVU7Jz+pqB3IBD7/AXyslfo2zzy6tDff0f1aKuIRbrCMQPCZFcuPr6mNo0C0R1UNqgJuiNo49m
PFWkjMplAxGWd8gjUWLpvv0T2zOhsERDpt/avv48c0vPxFDLUA1mH5x/GTjieU1JZZ6HPFabWOmc
qPcEMlN42ZqABdlmaKLErGB3BOkOb6XtBPTmNpd2pb2S+eJt8h1pxgAbbbTx3JnkAqqzdkBHEp0L
ZXaCDEzrJozAWHKl4Z1sT3pxAZwWPRr/ouv3zfMZEhPKnwd40aCXsdZu/U7Y8i0CyFNZziRYmjaT
trxjFyjyGCfZV3NId4byphCHLPD0+mz+lWPKFdm6+7mqk6WG08kc1+D8w6dNd+fGWN/2SOK9fhXE
wOc/jlQzNgD4wFr2TZjWhjutnHQUWOk9kj/KPnjpQJgg8FnLlqksZagG1uhUe2U2R4CUq2Ftb2ZB
TDE27AaoDYfuZ0393Ch3Wa3i/Kz7xvLv9oXbDBSX2sJV21wG2I06tQ5gPOMaCP2A9P25+HvTJ0FC
BDg5YDZpqKk+sLHzJt5fXpPOaxyi/qrcjmNHmM23ZA1ukxemQVf7Q98tjVnWX91YzJ/UnEVapYx6
UH5KE9Mvcz/YdYvGTitlc/ZeGAWt6ITcvDdGnzerJ6j9P1aWjsTlHWIWL7O73BHGlpMvQMGPQOMH
H/+sPQttkdef2NSQnz9P6GrqrpDw0rhKrELMShk9Zo7ItneD7QXFFQcCpy0cymaMhCoEev3avWq5
Ykh0a0zXdy2LScFnsJ7NIKaZ2kOsdGPvYwiToDxtJHI+zST3tNvbxZo4cRNodAxsMAlhnUDfoZXw
1U+xzpNYUOK9/quXXiw3yMcUiSClqvXdaSSjAaJ7wkuQRLkwOHZpblGxZNyNMFKFP8PtglpqqmWX
+bAv39ht4Ist1NyW8KYER/3Q2maQxoyEKW6mMR39jBUbaMLf1ZZaB8liwQXvtsckNp9MjJpMWNjr
Yl7wpEtxJ85TZ+pMD+6Vk13ZkQB2FXA6zloMehfYRePtRZU75ITVTj5SRfqwYCUoQQLztP0u09cj
BDvHs0xXTb71AF84SM05jYdXyJNd6NbfSOUzFLS4B4aVGtX6FoVUtLsVfboC8LoEOrIOJOXInTAv
vEq1WsXcVVyGH9g4DBZkY05vsEOjXCfOM6VpSZaY1AoCqHO93wnycXtjr/hkW8vc+JxsB42XCHjF
nF/Yy3B3VVuOgrrNUng69ouz8oXiHcHoqAwJFzVDSTzESsNcLL8+vobOgLByeHo0/cYLtOs5UaRz
cxZ0tzgRsxkvhfFifsx1WJSE7h9MTVlgY4h26qJDBmX2joTe276Mw1OEdTmlQJvXTnzRbeV2W2+E
oleXVKemP4Ig7/yNrDslTK3l7/oVJ2xmIrZuy3SX+N16qJnDH5zttJ0jURWd6uKI89Dg6beyd2v2
6xAzZxY9WU1bM5QVMTV26OhIHjH4Uq3tpjk2jKxjD8l4sEYAeeWk55GuFKVyurDUSrjTFJAuXhQa
QNbyWe7tWTYS42NjNcTTLVQlt2D2dqt9RoUbEMRYZebmKP+UvinU3kKm+U9n2hCTMDH+3wonoyyA
ThvEiMu3rQuCYW+8hZPt4pbI1dQ1lEGmEYZYxKpx93izagnCYZ/830PYBWse+YermPTmvIiAQMlv
+L2UEFnBxpAkVv00gkFiaFvJaM0fBnQi1J3O5lPcmOV77YAlXbuoJXLqXloIE10N1LiYfi4PTRF0
h2rImy0HQFJ/qhoH8UV2p/5SBT3yQtEL6jMlm46htiHadL5AiNK3Tfgbn57leBm/X7jW0BznZEvg
hlbhrEp9AADDoafZqmFAi3Ka/zMssxrsFZcJgo8bNmAV90AZGKB/40VCkg9VDNTRXT+JpeNlwWFU
w2Xhy99bU3va1dGQhO+kp/TqtBpALBVPRPQPBjK+U8AZmDzSnPTsqi1UlUbBFirZXoivREHEycbs
8VisIy/dQpX1yzb716YrmhxJTjofVC0mwfLBVSqQGiuQz6dmMCWApliO3JnpJ8BTPuYfjkgiXGIx
fgDRIgZQXBtp0y52D2IXp5wXhKmUWzEKN9QxvqB6fYsm/mieaVqBaSnptO2sENCS1lUoQDLkW2Xk
mo74qcmQGqRvGAzJnBMU8wAK1kWUvI0A/Danh98ULaVW2O/P4thSNuVuLt+GVMZExqoHoB5ImdOB
xIlRz/Zpc2d3T7WmLfTWIa733GPEitX7VmIagHBj7tuwQIvinr2wq1shcwvR1V5CwIacsiY90B42
om5GWBhay8o7PaQAeVj8UNbjmmtZ6oc0G6ZbAZPa1DWRsoNwScxD3vP8lYOec5vMHBqW7f1zy0Rm
Ko3MsBArC2uyBqoQiivFEDjTHE3nA7sgQlXaboLm2ij2q+TY1uYWKj4hjphAZJBzBKV6jAWGQvzO
J3vXpAXrsZiv6dQ0DLbB6MpCDfHGfOtJQTj3vfmJzgBJ76nepsucLlpWCQVyuCym4AtOCm9xY5IE
CbkdKOvDJ0ZnJ79EZ5AMLgscNEBFzHi0Xh3Q1tnyHmO7zC7l7hVI7zt4c5qFQ3m6Lt9SqGMwP8YJ
AOijX60wrUHbD76dQVE39io9jiFAvvmKxEUQMXPgamxbcq8EwNPY8BgKLXVmxQWNV14DSE/GeHFk
sF107O8SUerK2L//ELJYrhhMs/qLfuWbvtMwd2lUCwk2yHdN9mD/Y8wb1eywo4eLGwlpLUvmS/rX
G5f1C/HfoFd65TLCEs/ftLj/n4nJQH947bE7IWaAYULT+bsDiqN77740TAHiYSrUYBq1lWaI40VT
ijqp1cFbt5T4MzQ0l0p3Wi4DfHCYahGWlGtTbQN1epmM3sA0RobsrHsuLxSnsWtSssTtC2Qw6xGb
jfwqXa26V9zTrGiawMW4mfkQo62dVlRCnytt7FwXJXWErRckiulG+aNVuViieM5r4LP01mN8M6e+
bUAQZ1E+dructZgkDCn8nI0f+JCTkKRsvPrxOIiKgMj5Hq/pLZCFC9XA9zupoPDfZ7fLFYMSmLSH
R8JI6fbAWq05R+TfT3shkthCqCkIZyFo0Qp5b0K56xYeWTR+ZnHpFL/cygMBdr2hOBJqSCLCJHye
CD/xa9SW5hZFzlkqzwii6WD/omWl6g6kX360kZD/lmH6g3LRBlV5wu+ZA+EbW6fhfEaVKgLalFNN
To51GOiLukTEPQQ5MN0lyfvoV86xsEEnx8xVGE/J1DbAiAj0Ryj40I6F8HiSuN/aozlbPXCnFbQG
8Skcr2CQDqhE7JUY7+rVPHELfD5k9K8UPHmxhQj28lWZT2amkC2YL+otlf/w/zPmI387WbUn2+Af
zhKSX2gcej+HxrQLfdgYGZ89jHHC+abKz9Qryi4RHLY91MhE9KLH4jHc94agPsRAU6VscxSnR3kg
8CXfzFBCm0Pw+ByiUoTsMY3oLjSoyOInY6Q15n72wviJM+z4aqd5dHTHQcETHU+jCsPbRGbG+aZW
UiA1kG/k77hy8QbpUMW3BjVMVm7+yjFAi9wt28l//sEdowqCPK0Uceq+kGJewp/uhdP0YV47AEX4
JJHM1W9rIk9JRU1dIau38UBm4zMXXAKFjw9LMJ0wUempGTZVzZIAPliT5YJD+5BpxnBxH+9qmTEl
5D/Hg8Eiqj1XoZvGphPt9cH+sU87XkaRBTKjDsBrkN4E6W7x/x1VhRiWCEAqqfNPHciloTGMgaGK
B5IWIri/rSACgRxsIBmqG/z9QTuKGuKeXWReom4kid6/V6Db2wWaPM1kKds1THZXX8CMDCp+4Ax1
cTqQ7r6gzRFUtxyclQlCqW6eDJINa4JAhzBQOCwzwugNl6Ejkn1XWYyBnyT6qwXmtVlV+NdgJpkO
8XNiPp/bBrOjmrefexQmQn42ui7Z6J9ehS+VrOOzsvAfloLam4P1vTC3wNfAqjbh2UY99SRuhxMo
gjFVnYh/7YyabW12Uqvp3SA10deHCj0Vfa+C6angVY6Pp0fXuXnK9MJdKr3hPe0M1fzzhugl4fhU
xa55AxuQyJkH5r9z7k9Jn5caB4TDtF23G46DfYUvADRMpUhR9sZ9+e9KK3rg6JSdGKvPAUNKrqv/
9BWkDllnvr09Kn3fXvu4cWcQbnuSCTG80uxkBQUXJKqaF2HeAMudd8rV1mXrdxcf7I2+Q1Vj9lXa
yxMQit1bQHFDRYir1CcW3kjifBcbjYDnY0OPDc2jAX9cHDM7FJ1LTK3QfisAfd9/ddWvS/wdjTpT
bxfnzXfe5wfzJBkj1urBmTmpCniY6AQmzS8CQSfWBB3lgR0ff+V+h1Yj3bcvxBKUxY/UH2Acbxmx
bgnrkxZ6EPGyJhGiMzD5h7TiB1Q0LAMz8/ebKoNUZt7ghQ2J7b6fR6M5qHbx/XCwI6oH/eAkMvDw
c/cjYrDhIZ9BX2dmq/zSKnJwGDnxNNBENqzOua3HXsOfwsK2hC/av4Sjgc85r+GOwe1y2G8ABRXb
cz2+yNb3ZY0pzDz7XRC9EdbgqGo148BFhDScyptSukYu1mVr/oRBaR9UgnxCJESZQmLj29WLcf7g
xhX7e7oNFRmFaMLkhWH4uoy54eXVhvTM5PjvShhC5RhWineVDAxs6HOxQ7d+wurz4u8E9Q+Z+iA9
qRC5oFO3j2nYHNQtfrNZJFCajtDejfjwtk1NSrHmYs40XJuxP2tGAhdBDW3W5wQ5iMAjiTzqqYlz
0Ozic0Q9YdAhb8x3zsjsCzHiCp1v3iVQbwh002DnxUaAzQt3cIgHKx3ZupjUpbDH0RQ1+uy39UEm
oCI93Ep89jMpgNjXc0NIh0d1at2hzLHFAJ0AtMazeprFCxFVfIckShkVPqOxlPQgerBMCfBttajh
uXrxglxmlpzIbVvfEeFOk2VNgF2fBqO5qLgisHVU2zAjZLZCige/vZzr+IIQXvbwGVQXdGn64HKQ
eDohhcOfNh8iJaZOimydnHMEXnCZgUzmo1f3KhrqLoH+8+/y7Zd8INLKgj48q5/3PlFM3xP6iLDS
CcyDJRwNOqEp5yMT0i4dYmVXbJeQh729dGDDOOGrI2hIB3doEi6XKFOj1PiDpQxzUYHbpynIYImu
vtGT/X9gvLA2/6x2jvFKQL42nvfNFc7aNeqC2XcB+JWWOeyMCLT7HxHvEf2X42KWE6ytu6XANVyZ
QrrgAcYw8zP9xR+hmvY6+EHthSSmVlJbMSJUqT8BpQ55oJEAH6Bp/nkc53pbdD96r7mKqycnFnSx
kJUIr1BHu/8NyU14NpU3vIYIeUtW9HS5uzkbf60/Ri2zSTCX46F0nX5+UfuZmQt3/4krIPiIgasm
z5w2vKkIkepwjWlxPNqTPpkcaygtNDU2ThieOO2yQsbMHAFt6XIR6fGkMxUdiFHFhoQf+XMZYjzj
l17E9DPDIoiNYzIT6mymDg83w7n/bGrABjN0fnSq2OSc9c4bzqylCiZrNdXiAtcbhN0hgdVsvItL
YedDGGK1MIivjbABJt0ZOIStG14U7ujlAmGv5cPuQZAPLk2VTnybWQu4VD7C2+jZ+79fSMoF9vFi
i5IXoQOdIPa/4U/NdogO5jOmPMUu4OuF87HFgyX5YCaZzOBO/2MDax1LJbB/IDH63MNRNoE33yIE
qbMAQDTSnSO/IVaMzimtqtbmp73zX3Xu+muQC4FlcpSq7rN5RVy9AeYHVPiIJ0Nibv+MscgtWovJ
c57NARLcubgRk41tU79y8eLV0bSFhssqrnS/KjsDnr52mo3SY7A73xynpIgcEfL4lF04bpb8DrqW
WuWVnzaxbOnSYQQ6Scfn2vg9osdpHlp5mGlv6b8yE9XoHLA29uVSXu9opec9ZAQ69K2R5Aoiek6g
82VKkig0URd4qLh0tt+GOCofjsMu92JS2vj8DehukBObV/7b8oUX35GaRv4uiEGGsrwOQ89APmi5
QTcScRdYIl4drHjLz0HyuPSAO5/6r3DyYXdV47WU8Hx3iDt2R4efux2EsfKRhdzENDH4pD4Toatl
Lslgmxd6EW5ur9zhRALFdEQ8QUoa0Lq5dF/0Z35pfD50zbJxdIkupInw9Wssj7//8p4NIpUtDVNK
QXjwJbwvPhRC8GKFI4Wr/ZGsA0AUfrhy8K2BdMkgvfRAKSJ9lRFGHMBmXg2kdi2d3U9sJOPxZdtG
D3OZX5zHqvDqdJSTeeYmLfslBO2s6zHrSsHe64UU8Qb0yoxNpZ8VX4sCFdEygY3D6FCpG6/R3bsP
gY56ygz6GAubbQrTn1kZWuXFCVwu0xxQcFxHxGil8YMH4bjQbbfoR17R94W0mXh1zYzYXnVSIY4y
l5ZzXEsrP6KkIZYkY9evHHSzpSn5aMZGYGTctWE+Oc/ajSgzd0ZFq53SZiszvkf/aP7SVrsJG+a5
FdKjQPXt4ydfmSYA44jL408xSEsNmqkLMR2ZzeSD35Wc3KvqadCkrFRy5KoGMORKe9TiK3xODwsi
nRMQp6RRyc1/XXsS4Dqq7hGtM/g4ePY69bCdhfHJ3rr+qObruWrFRh5DqnkHeunKGHwRgtSSaf2/
s5RhxXrwKOhYLWBs6wpwxKB7ycawjtJYxeUXMx87XfrQQPB8IK6aqjJFmR5pYASKt3AmA2wsv3f3
NIne9K5/Y2XRuzs8jtF1o/em2iq3O9ILYDIsy0dHU1V1NoMimr/mLkbo4B3TfTMUl0Lxt7cage3Y
vAvfFxoYf4J9Al/zHdDfTbm/hFbNx8aiDghrkU0mZejZXGayF0fBCSHcCIGTjDeRC1UTXrPJmMO2
WaSlCKvMfmGvxu8bllecrYIuPIf392f0AoUSwTzB2Hkt04iP5oWIF0gkTT/DTJJxZPRSrlcYEG+v
2eOvjigNctgXj1dnt7qbfNcZLK5diAiNrZofa5Nfgc+r8ZzUnObruNDF5vU24LlbnYwmBFR3AH3S
oIpic7ibQL+nYzXqvtu6a3wANK++UPCMW+m+vCTgfrsLZ7l1wyXqv95oiDXF/gL157U7dExH56A3
vZHyJL5fMslD8nMmR5jVAeqvWZwdLXRbCkO2Re9/qU/A0uCShcxYcBejbwLHZsCdgCu+na7p4cJa
YiysMc8LjgbigGUKyP/CEFdoi6IQf7xiF/NgrFyVwNrqzkORyCe9FGmwnJ+FzhMKq3LxCnJf517f
oGmdHFbiDQX26m5RX+b9XB53Fn/gc3EQAiG8pnGsQgO63NVC7lam3hznarTb5w+9umnbgG0ruNIS
+pgTur2mWPME/lyslCsIwUXWLcZ1d7w9E4QGqfwOFicTEIovFld8zM2axHcnEdS1vimaaciiZv4n
bsrsGcWzIkhkiGZsl40xeQNy2RaNN0y4dJuH4ePaYGd/9PJw7TPLdzz75WeztP+j4BjbwGTJrzSj
bvYHJ/eHc4kW7MI0c821bnHdpekK7XjXKhxmbK7kTbJDMgK579G6ri9klj3A61kL697oun9DeeNI
EkQ/VYFA79pQop0MSSxM0/W40h2fThyF1q+XxN0yXCtkWqNMhW35A/BModNV6UrhUzHbMF52qeSV
7B0hxSwkuNaAYYfSo8j7qKTCs2Di3UfzhaxWKaG+6Exwa67GvGIzhLLiQ0JZCDy478Lc3lDBLGkW
TY6LtKEn15Nk5PyLAr+q+ViMln3HUrlHebpfz7ISOsjoZf1U3EXMKtv3K5rnw/fjN5VuXuYA8KmK
PBmfobLhCZm80R/23KF1UkxQjSo17qKQmOz8+BPt8FAoOAqtC4NJP98k8kK5r2xmh2yYhAqD7hNN
4mtFd6M1pgo3dM+exdTyPTeEZ4ReUEuTEzGqJh+2MYzNp4O1oU5r6Y1V26wOSkS7rRpoMdE1yQA6
R9ZXeU4yFAg27/QEi1hecYToPz6CCQXl9Xgd2bZJt3OBDRbUrBUdP/u7axEY9aQvXM+V6r7xoOlS
YelgbF/o4QmNnQvtSTvhjjtkWG5nkUg3FlLbxnaY096mESemeNC60apZQ/c0uyNU4Ygc4qeKyc/6
kcK3NsUci9c4YzPhUuEj5Io/MeeAg4MRboQbKmJGaEyEf/m3oko2cHk/elYwsXIGIlFeO1WqnUtF
hzk8nv4v38YiG8ph8eWFimO57x6YjJNf0AHUPQqwBnK6Uil1xzJV/Zj0VlWfl4jwpofJMzZZymHR
GSp2sDsiPwCWvpYX7DAZbPnsF+h1WpUcwvMzNBQmpOg7j1Vik9W+WQaxGVDsRuyF9kRqmIdIfWrg
fXjqEg4MORFNN8pN0IDZOTusEcYVosGqNRkzKuDMCIA9rowbafhcEheBPtHW7awzzyeg73QHq+Ow
PO67Uno2/nvIClVhp5cT0e4KVpSJfrkeeKK7DzQU9ICbHlLWrV2sYubsszLoDmoonhSTDo142vqI
/Bw6rLwgETiFYPQEsz4uriw2CcW11a5Y1Z9L1fl7RCMralxnU2J72pAgl6aNjxJBX07kTeh24tG/
oV8lCl6FxOIxpwtD+3Floyz5/CH47ciHikGAnU385bOPRZ2VPVonFF3woSbGJ6BJD4XCYzUamutP
esIo7L9w3qfRAA5r8kwuofYTJDesymLMBcRwIxXimY8sVorewOjX1fIP6ME7xqorkGB3cFNXEW0H
t++/mmPYwuxUHY5TurjR7CMmvp0OQibyVpwYgiJR3jQZzcohC98CQjKl0LysU2mp26nNGZJEEa3x
hqQYB0w2qLMuW53zeDw9/GzmcMmlzD2T8NGEWdy+Qd3kqwh7UUuXe0tFSRmZR8GxR48/qJFrSbEs
SOOfWUpuqvspcI0WdxIna7wQY/LgvGlzHVYYECmDk1D2vmgPmjHaXHs/weWS648O14NPTdqSO3un
b3xN8kkUtpGCFvloo9j2GAHY6hqNqMaX743YABYt/G6p3v5iFcV4S5dd48pnwQ0zX2bLo1ms1cDD
aT6aAEQVBuRM4mMJK0T1StpSgaS3KUwESG4VyYZepFJwV6VwnOZozTtJyh8UkoEcpGWyhvsoOblD
C4g9nLW7nRktP9jcnkjjKRjXmhlqg6r+iy76SFYa/M7V+lI9FXZjo3pBVmZdgTMvnyElaJA7d0Mz
JMYvwngR1S4OCvXjzZAn0Zuaw2dgYQVuQoXF+kyT19SrUgLCbcXjd9aA3k87eBRwrW66uuuiZrdi
XH5rQ7X+UoNp4pTUYlE1dXEoXaShafOXze1nu2FOEx4XFJySRmPZkRQT8GGwH9JYxp0Eym35tuRa
xeAVpWc9YQrbhUd0ixv/Qwt5U/XgEJfPlV+qgJTKw4bhaH4pHO9tAhC/1xyQiEa1xF+CGxycq/Bi
yHZxCrF4Z9yH9zrKCpKOsov/BblVejvzNmlApfdQYamwZYYRPaGIm8r8vStCkIJ5WdBNkUtyiJZw
ldg2lasGJB0XBk7KTSj0Cue1h6cYpjkm2uKgpdSTct9aIwN/LufHQlegZFHdgoYroM2foKIHnUyV
mPjC3TyVNWEIa6kHSlugmLK8edeQkDQpaddKEdCtbmfBMuugl0iDxBJsHXKT4fdRdo72FMqy/8zS
tEOBc6kArlkkOg9xFFHptdydi/XZ1xG+bZkDMlQYOn3g8+eES5+T1rnORk1kWL3J0QhJG2MDHxjv
vFBYzNJLTuPoCBiTPD5Dmowq9HhIter3eqlk2QUrfAjzfEXUDTtUH/wVOCr2nltJqdVY7vBp+I2H
julgq+LQhJUkvoFipOB4HslXKLk+5cKBtHpCuV4vCsDFVY2m67URBDNkETHRRDKAFMdq8zX6Ks1D
w/xFZ9vU4V11Tt+z54wz7zvsYX43UZsWRpDyRwN9WH6sv3EYdxCGV+Qt6tutfO0TjaEcrSc1aqmq
OCJ7TY7j3exW6BjZ5qp20y2AFs+A4ft4XqsrJQWP5yyhvDKQkIjxZy8KuP6p51MIVKPt6eXN3iKS
RwTHKGe3n1AZ1c5LzVIuVFNqhyyoCebPa2TdwpzpjN35xVlB7EcA0wwfyaGURinOkihCpmDJ5Qr7
F6D+2tEYfV5Wwf1vpmo1fSabljpOjBnM3t2DKQ3YqfziQhlX+s/eFCaU0nseK2xcJ9DPcCllbrRM
hToVtk0An0OAdzeKnqSaJB1K/sRBmlcsNrFFJ3gyT++ltm5AWoDDse37BLaYIikenj2X897o9E53
Nm8tmfCYMwjN1iVUNsBBempDia7cllnDyemfgWJXTKShDLR+4s431EHRuPaPEEAA/AjyP6KLWHIW
mxrIiT4Dqsc3VApl6x8fp+UFX6BUl9a2dZmvQOD5Nl7PUHe1zivfBe+LkYWlNf2NpjosLSdN9dWt
x+oficSR3H49aGvGdcIAjrZp30Z/UXo/o0BcJDmwraQChXRv0BDioQMf8M2cXGjpOsogSesZehqE
tJ/Lc+G+8ypKa5Wealc6bEqRN42Ebz6E1S4DLP4YuPy+pU9Qua4T2HxCVN6ReBTHhzNnb4aQ+Xwq
TqkzsetHkliFS7L34MZbSD2mcdQq3v2qU+JYaq7G1e4YmohNc1jOpOeiCfVWQ3CtiJyy2uc6PWd5
mvSkJ4zUNRNrktfPcV4sL63do58Fo2HvMleN1ikvuaf7kCzqy1NXuoU5KVZFHSdZlslqdct2mDB1
ItshXXLDj+HI1XbRIMu12Qx6MJdWubLTAqIpw1Ue7LnSAT58h8ZcAWMBDdZgKgj+0HFoyk4HM6U4
KWuA98BSRAiofOVLxiuMyF2aDtJlvbLSozvDV0nS8tB5lvg4crtsdz3H0R0x3MFDTwjApcq2gVjU
BLTagdqCjbHLDsZGR3ArhdQvbOX8GTkWTF6hod2atIZMMVSK49znm6kL92KNrLWd8mr00YB1JSvB
ctmC96Yh/tgnoD92Uq9z6EP9Bm6quidNfXL87ZfaolInsxbpTHARljNlUlSjLFY1Y38wIK6PJeKY
IOaZ1KD+fvn8q88F2BRpOk7Hn3yv+uv+0HBUHQiEGvwz8qNYm4LaktneNy1WSgH64DmFPLY3/PCI
SBfHEOqxMQMl6Ka1Cyvnf72shItXc2I/aAR3U0mVL0XR9Rtqtc7pxsDyYNoeHKRYpBLRrbtQEn/N
ihi8qrqlYvFJeTIkVlwqgK7vCt/rdgjpwwqZPXYmkZn5eDrN5fTMJkVliHlM3TFa3j6o2u7XTTnl
MXEGbxT5/WmFnSRFVkX7d74PsmoYH/cdEFOXgOtaJ/s1svCsxpf0M376SlvSbiOcfGTPvR2QKwVf
+O9OO1002aB7Xsi8jZGii1J6DclYQb0wB6UjiXwWnYDc1OfjXjSUf5biyxZuuh9YgGTHVmvN1PAZ
teiRa1qC+ZYt6xtN49h8dUYSgS+cINbKTBhHalidbad+k5hUZ80qsOJStWh9BDDdNiX0cSqN/09C
N9poHlzn6CpiKKp4EWvQWXrMJEf8wbOUSipbisNZClbtpXJdu396A6yjzcDZ8Sj1n1B5KOQKLzlF
QgTvp0+DhBA++xuDlMJwtWzKyIQabJdlswm2uYUCfXMAwa/NSjoqtKux1l2huRMtdpdFGBw/UWpN
zbIYOe7i/2dGpd0pIu8ZQz4kGZ2tCsVBFR/cY093Bg2Z7c90JPZkOOP2PLucE6/xJaGYGZU45ubU
ZAoOPXZ8oX57dAWs5qzvvCYYCf2Bx7g93iUiX1EeCEYpsn5Kyo8Jt+qto920iwwnZ8ZroFwFTVor
v+DguQNA+6vKAI8pXUsK5B+pab4fKEboWa9yc2TYNkJEyB/1aB3PUUE/M6CEI5huc2lRCfGchlg6
p2uBNITYXcprOw1dK4ORZWqIZPHsMuYKqskMFEJa8NyRr8cagH1/B4NdGWFkLYUS1LM4AReurPXB
O2ifIF9udclCmy4pf/TFATuddgrfFM3qcVKswem6g9iwqpnTNqkN3Uy5fvFjrLp11n07jS179xl0
dfGQepODfBS3RCLLWV21rBLH/tTKFjOXrZhmOqVm0Q2uPDpUXgyRs+/TeX+CddVNW9Eoub2yfWMq
uV3sPXo3U3D/Hu7abMepMKzJpQnI0IDQrLb33r21oGXDM5hA+JArIO+iWMF0rfhEwlHszFq0COzA
nmUkn1oWdWNgknQY/9QI/rvLX10nK77lIOihYieWASlXkx/VXVeLuHIT7NGi/q09hN8nnikKn3NV
AMwS1dtJgVL0p9S5PTJLeM3TGOAYiawIS12zjhWVLdUSYRFJBl63LHmmWlXwMG9PqJnqZlr4iNBj
DNSVt3VvEyr1QKAxcShKNfsg1HS29dLlbwzBRwEYelyCT5x1c8QYgiEGvi54Rhxnfz8BwuqAgPdE
7BAWL0/mnN+AJDvB/ZXwz+hn3ZpgltisKPj25YTwtRLvsQND+ebuJLXjobQuhK8WUQ2+rg5bnhkl
ybh4WIKjWa/RhRez+pidIyGs2v3BKLcZSups96HTP9hrIcus75kDwc4of1fcS4SjcySM8bqwxI8p
goEmTJgZqMrP6wUHfN4Tnt6syefCdxYTJNImyR5pXJaqQLxRodu7fsXCKHC9ngT4kgWoBxtaHDkV
5PnPRQXFPMKOQ0Y1/zvpAZmWRp6nWKoSS8WV48Phdigb/hdtsN3XtHwFx68PPEZeFL9zE/oSlNcu
PTvifw733G7ymlwuSKi2nNoITa9nVbp3M1HkEP/k5EWyk8PhgWLUsz3ScG3lQplrWlXd0u8xkHop
nvISpFgOYaPAV7KhU8MYXevpW0ObM/60Zr626xuwc/hEStruaL7urVH0wfEQI03iTxy+C8+N+IgK
zElQ03fFb61NuzZnf6Ty2K+xfa2z1+ItFVIFPdkH4Nbn+Gp04p7furTy4QRPx11fBrvNF/nuUEpW
dZZc58U3k+wClfRFS+gzuPUCmOkUqYIuIQrO/AzCBVhHfWVIs9hGlkYgfw/NsRnKiDXR5EdfmBUv
LB3/xuj5Z745fJ+Jun4isCwEEl+xL5OuibBZWzhoDfjyfY5wvAb70wmWOrNe2OW/w57Nj7yfyrA1
1QydmwY4nF1tvA1e0NfRI/klt1U1uaaN1u+DdLofKLVEBvYHWvmpxezOeBT4UDB937qiwNVh6/EK
2fTw8MBm86Eu8mW0cN83MDWS1F14japckypaPL3rZq2ILpkCb8Bl9qqprbWWSHxIVTKMbS3H4Wog
3E95QEzYnXZPmM+nK49CzFPZsqE3HKi1uNNaZzgLK7E4MY3L3PEGHEeBbJENLoeuzEfTe+XWZswH
wYSod1xG0tAVPR3TNKbxnxwLPi9IQ/YJ/SQCD5JuD6unjwMgfmvhoZQukISvXs4XC5UIaLP/9MMb
tsnsvjUU3ksbwV9vOk//Wkff+HMfj4k75UeEoz7Yk3IRl/sdDrcn3hrbqkj/7ojl+zQlDm97Q6DC
hEmKI97E0cobbmfE31dde1+YZT8SxzrPTt6u49jSFebJruNmyiFqTX1At+xU5XyGGh1PVWZYumhy
hlDZunX8UUFjIPmup0iQPV2iqnV+FbTaNnEHC0i+hjPrdIZrUySY+hfhxUpviTG4NBLDmAKXopTf
XIIiEio86jvsVUntJoeevmuzBjjh00f7ppxUKfaSTDONAD+LuW6G12M297tVyGdIvSWe1EoHeDgu
S19IqRy2uEbqD7oq/rYSJs70EVO/bsB2zCtVEYPPEZ8gVlvkFzbRf0ezZZGb1EMsTKYSlmAJgIuH
4ZwhseLFD+G7P9fbNWjXF0ejbzNlJyGq3qu1TC0cdWd01i6c//5WLTE0V9qCiP95mkzyAR2M0vIJ
KgfwXdOmKl9/ee7wjG5b+SrgBT/NyOw0+eGGjDLoPTca3iicJPNnvUtv77S/nv5B92Cog0yH6XYj
vIEyGgx90Hg4CSlElwGvKQyiFVk380k03W+67QpmuucNgB/HsW7n3hMpvxRbVeHcHpWMSJZxfzOl
dDAJodbTk42+wumqsj/WefArM+R/rxdVvOPcFjBuuiW7hmRmeTLo5ZvYseeUByjs8lGSFAzmrz7c
nAtc1QqgEU+zMqW94RLOnUyt91uAhZPDQ9I5lQlQaiQxW956h3iOLasjexXbQfpDwhcCTooB1gNM
AyTLbWGv5UlEH5JWStQrIYxvXvh79LXS1PBTKG+GLniltdNVa52FhVc74uXhS+tf2pSsKTgyVknS
S0U/dj85lX6ZrqT6y2oQ/TY/b8cNIWpf521xHqqRCWjEMQTHmEeUvxqK55N9QN+68CZNARazxixV
bDofxrtlrrMJS/Gaf7JzprjYlm6bW2F1vPOnl62lwoUGHSVqpciw71p0WnZ59t4n3pA13YgCnFJc
NIU90HVvdFqVVKzx/p8nELql592DUwZMp9hoDyf91yY80uFRKoYUSyuzOhxYs76ueImEvPir1oEn
2/L+GmV84ozOmXlfRZZO/rVCSQ1OugLywn6KLvHJobL7EWG8swbF0TfZbzZil6KETrdZIXsw/LhD
bdb45pTrk7CHt2pFMD/cVFfcLXULF7mZAwTlkLeOF1V0qiJ4wo0YSlB7S4u3uH7JR/aWGyciH4QZ
NLw+T6lG9LqHwOWrrJtChC2s0aD3T5GC52IkMNvf+xyp3+QYZg7/cFbxWhKFQYYE5HsIVSw6Lszb
3RypGbDvY9s2xXv1iCoUUo+Jrhtmv92QGZtZWwrhuvEXOVo7Z+A1uT1Ybvpm/5c+m2LXqTpbur5P
Dn+c7bjlSRc9pzNeKQViC3FThFy2OM65Xu05Ae9IgeV3A2U5dswvxYX52b0VYAxz/T3WPJ5E6Zsk
Ba07FDmsi+Zh1fvUK+30m9c6nRkMsRJJ4xVphoviKfys/b31kjuoOTlAQxw9RR+FLr+vSNn2dWAz
vsORi1mcLukWB+U8CKCVrf6iwSNscX+INWDzZCTk0V2iL3Z2nZc02wEumbG/kGAJMoVeWrZAERKb
1BeN1tnwpV0Llz+0b53Ob5Yz6DBGXXVokNCvtwafVgdZ1zHGUO2nYPJKKR6zF7jvou1vUEC5PFmB
vilD6fJj3XV4eVraRXgOqRczh2Df9yfwewbZ4+LCFkLVnHPZS5ZDI24diLFoN392rlKqKR0SSHfs
LSL4OfMbWureXT1rkHcZJ8/D2yWtAUvysQYq8uK8FUs+i9S0JvmWXmaeXveiazxuggJ17pze1Ua6
P05dgTCwd7o95xHQZiZs591z4FWKHcua08BkuR4c7Gf2yVjF8SWzp5js8sLk+vG8YiWTR/j/D8K7
RX5AQQdmpT3ekAE8eoRSRueg5+SMdNEywHVd1CD4KBpMjCCXih0gCnrhDE/DHJOX0k64ERVg3W3E
RyauoyE3wOZNkagThu2y0AfXmGvBv/XmKbPqLH62tXsUw4wzmeJmnKbEfIXRJdVsNrJHKUJZmtdz
k54GyzERlsDnQ3pYHMiv3P83L8p3HDpQPjr40Ucs22iuEk4Wg2/2fB/HoNMPef3R0xcdAu4caZI8
8ebowOlpTQt/tOIvaAxo3wTXw73FVjFBCMhWKKgcGN3/PVMqDI+E7t+nGic4HjffOOs6qePOUivS
jNYmgzqjP/odMo8fcW6Op4bTQ+/dasxPsJZz7fmeUVw1+7nEPL+32tfjSC9G58jObcyFZJf+qy9a
lmi0CDsXRUwVXc8ADInotW5HCQqMCi9qmwqfmuRL8P73QcvWjC6beeu7MWKWGUlsAwK6F9bq/Vsf
5hYnbpnoYDckJnjWOBPRLKEwslv/TwwvjTh9Zkfpa7pmt4uh1/C5h9hE72VyjVGDY5wa5duSv9cJ
naoRwrtGrKS6UgTr73awnoGGm370HopHO44LZi1xbsy+E7paAzB73P2JTz5OzNZS+wrizbE5Upvn
J4cRLBUPQi67HSSfdOuuZOC0GYXxGeTEBjRhoRRgSGQcYQc9RHGNA20FcMJ/sRYxs5Me6QiLmmZN
gc5AGGDXxjKjx3DU8pC8Q90ErZsPNYP6cK9lWWxLhP4L7JWdpo+vWWluIuC+DA8e5vdzuc5p9X67
1wkcfWguU5fIaULO1M8EpVr3SNa1uG78bjKn0VDwk34hr1utGq1i7fzNhzxqxfALA8Px/8f026Cp
zEOKRJxL+YVWT8XhZUXKwqSnFa9h/+RnVfDRrI4xHVpBqT4FvHdBXpvI0KI581UNJ7/slfpXu1hl
J5E4njD8d9aDLvipQHnQQMd/0IMXCM3fwidJK3HzZuwse1lBb++pdzyIBTTOVccphxvZdceEDN54
Cd3FAMwGMnLKxM7PtD9ply+M0/aDUkYkoSnIf2YR9mezU2FuKxct5pQ0uGJrkzxARmK6ig23Afqr
FHCu4GUFHto1UiXfTlK5JbkrTP7NW6HmnWVzejQvIkldjG5ocQYIlr9917hWQAf0k0VyLIJlqyeq
dK8D3x+u074e2Sotk0Jof7kw0DDNORb+Po+pSFoJ3teY1UrnfP/b2pUvAilqk2Ou574dbxPy/0n/
cioOYNioEhNo/Zz0BtAT4Cx2TkePet+Ihpsq+AEKaD8FeFkUS47qgl+Mt7CoUsSqcSUK4eCZ/chf
wDcLMtmhL4XCztdnLHuHX/Ay3Pxi8uQ8uGuU0FVGBK81EmjA6w4BaQGSjWSS0/kHPdotScdYIzCF
ECOktNKpdDE/5tiiRF++iU4djUn8UwwCUCr4u6R4OriuVmqbkGQhlQRoqUht4dCD6POBSX3zvciE
Arg9G2bg/jpfYU0wxj6cwMukGwm0+79jex8MIrK+MFfgFQOpp31cj/Dy6B+SpB+xnfiQjaby2sDq
V/ZklgYZ4UevVLNGuiOAhCGlh1e2EB5mHGIluN2d2NYEU7Et1q/FR5kxB/0MDnuwjAvV/NBsO9Gx
CTaC0jD6nLr/1d2ubf+3pt4g0ExevV5til8pP2bzqsS06qGZRd1pyC7ursL2gig7cNRE3r2o4bPU
rM2r8EloN4Je8bGBWZ9mmoJTK15E8j6rKkiTnHFEt+y/kz2VBuUF5qMGJ0mjyn8LKICz0csl2C0W
026AmFoFJPZHoc4USAN7uwFkuCpkE5aDDyo2A2X+yqh3jPOVBbpU/3o/qqIY38CxrbtqragxcXu9
t0mqw9rBHYe/jt05emsgPBNCETNQ5/47mJRS+LU9U1W8KnMsIpD1cZce4PoK8pXXc1hK08yLi4Uv
L6ezkqi8Rv8a3woEI7BqSFD4prDsmYAcauhig1muGGXbtyUxJ4oPXmA0euKa7tKYrQauxqt8kQ4V
f5rLCBU6gw7xTMHeJWc8Ns8MyQb+RzURj7Vv+ioZ/TQiojaSpaVFgPp1Jv8NIBKK46zZL8TG4E52
HAsfN4FsqGUwz4qhxUf4+BgwmcauiFIlFpYdH72nbagq4cpTsctILnAv14/bvlwT/6rqBy0weKMU
OxKwLMephjw+gyYQF7FouQCsFueE90qR2iYnCJ5ZI6/sp+RUy5zA7z5kXuVgr+s7XfutpNEMeVJ/
1nfFRmuk+nvbph30fykq9xpV7yE3BIH4nFP9r5fp/kpcWGHVtOjToGNF0WISGzNqz6Z8rDSD+Dcg
YASRzJX8Ge3p1t8hED7Qg3folhAdWe9hweS0i65kAxq0QG1te1Aj/KA1VedwVsXZGTLczPrTn/3e
u0sjvmdHyT/N7E+TR8Jfk84kMV8D0uy4L3rw8G1gGD7SWI81OkfKKJTrYlNWI8TGwPzt4Sf80IBF
Ucs+ROLGM4H8fBLPB3SjmU5RCC1Kq5AvjmoMKSEGGhTCuLXnCkTZ9iwpCW7LVBWZzJtWqQpU6/ea
poeWW/H50wdpmNLtamLC3VT8kzN4DpAlfdutmGBQID5IbnEZhcYkXy2d9iBcYl5AM3Gj33z1b6xC
D1A0B/G2q8ljEc16tvUpqHDSS2fwxFDGER67We9Kgxeg1TPPUytGdimlbybNLr7e8hKB/pNIkFbX
079mdWX/OjtiBhjU0OGxGtwOGDLtHuKUzW71vVQqDJMBH5fhYfc1jviCU5IBGGfup6c1FVl8H8wl
n9Ybmlyw2ttBnivAle4kXkhK8KOX+GGvfP9RRpGUr7eHtr1ZQUXBlrcTjh26iaVxp3gcfR6zw1lD
Z88UkQ+Zb1roEi6vVeKbqb5hLsugj4WkIEtOBf0DAjfdIzvVGZioXC5hdXadw3NO+a+T3pXPbJpu
/34xEaj7FagjuFgSsSNUUzCqi60jaIpv5KF2VR7aiFLnZ5dEZkenFfN2IjjOFgAASFJBzNvTW8Tl
Vymiy25Wh/lhVhN/lkFJAsqrsQLRXedKmtrUzel1G/S1+p6BOMpCWq7M3P1zD4bVN4KphCPmBC4Y
yzPQ3WZS9EOtqjGCQh9Ruz9yncqvjxNi3rFEvez7PQomI+Lm3otQeb46aoqYhZz1nLAYMGBVkvsR
Xh8WI42r+Fw8tvEx3y3rcLb41g2H0h+ZmJvA4e/38PwYXL75zzwDkvQTrzeWDA11HroZMsfBY0QT
r5eht3L5h+sByFGE9io4crCk7u2BgGX32QcTEARGi1bnkTaAaHdQFqnx5PFFmFcncatHNGB9GbAY
IZvOtwbo6YyusUWOT9LsNGP0T3TZIRlr4+VzqIgU/3eQzQbh/Mr3GfowrEAY6IR3HRQ031uKhoAh
HeUrNx5rBvzv/ESFefFDqFcfTMpU83DtLAnfgFsTIQ+AsLs09Q83zFkisZ3mGI9/TO3TEMOMGa6r
B4UhDVRhZzgocwMxkNWWHaMvNUhNHWN5i9zbgWh6prtDG9Fu0S6wrHq1Ooc1yN5ZCfIEkXucLX7/
tWxFi5cANAwYjXHHJ1FanLweyFQ+3PLBY7I5aUNwp/cpjpJwasmlkkq/eklLGnCC03VnK986+N2r
ZvPdKhQZ28KtfVUNJs/D3X6sxFG/s7/x5d0E+L1LewlpW+XFhHti6+niOggojz4kKzo1SToceOEj
mkSWhdpBVd8E2KWMRfg51dSCnww470Gf6kvSS0vz6DG4JfW0qWaPlHuCnRMAkqn48Xa0WAEHNtrY
Cb0FV6q8VvzKBpfCK+5Swg+ionKcuB88NjlRWjFX8GAt9cL/1Gbu9lFklk8dptXrX28OdNilLlgt
b0/x0Z6CScTPSeYAWmrKIvXjpcSUo+s1ZuvfO7UoeszcQgr2JbDaYpmm1JjRKPtVOjv5y/PCifEw
jwZ/Qg95ufjxgmVc6rc0eoG4TvDeFPbz+QBERHVU+huYwYgo7f8dDre9F2ATro/TTD/pkz7sH7B4
xbIr9PtG8WufLgqNZvnEGqfiDFihxFyTGL374eQF0GCKJGIf7pWfB4AQTInqFnhSRWuLJpobd6ul
tB9lSeh6WNNAL3zYy6HDciP4YKBXldpaKtZhivm1KRXG3nAyzkkWJEsmnMBZixjxhk+MUpNqHI8q
LPh5sx7QgmG+6XTdTLgIRN2iPXCm7GQ3fz6EWregzeaBL8q0oaLKROosWBf0DYfpAAqcNYNZK+ZO
i4H7SFtQZG7xhA6C8PLidBTGA43XtLHAMWZOolumjRGC80A6WFKgj/a5gEuKSleON41t0iMxSGzk
+vsKFAfx8esZ+lHqzwim+Wt81ga6SIdTVmu7C/K1Vo3XIO+XVzILqwLA/wVRDlyg3UhtcCZSY151
uf7xmkt9D6Sj3AWBVvBNYdHq/iMye4NnWS8/GgJ63YcHQjvM+4OoRR7vPvIQjUChxz15GTjPhvFZ
mzI3i9xSOvNNXLJBj5/iz8c5AC4d/qaddQsib5KXm/4rMdqLyC9tIHmnPYYw64U0jgqkXADhxn9N
5WD5D6tzjI9KVbx1QhuQ99IRyXCVfbGcNxQGbHu3vOKoDcSVCcBwsS4lI8yRr6Gl7As7VqZdwAo1
SAblaodB5X4t6kez7mXRVFHONwafaDUJ+SZSiQfM7wS0gbQLsOypJ8333XYM5tSvWCoBu63sy8O2
9uHay6dNvqIM5qFHKo2lfpSBsdUGIrm1RSp3s13sj3rsoSSwv1sPetucrxQr2jwg3O6y2mSzO2j5
yoNoKatVWTzdD6iq3KWpX9oug7REZFZf/4iYNYjTh1s2RxcDOJ+hjBgsvcSMUITxXhdOE74P8XMi
9mjsleQ38BseYTMLXI5drzMVW5uBTsazVj1Hm3NCefl47Cn1Wml3FgAaPz2gwxOS6fk43j1kFcsP
I70ACdjLycVV15lwefWTGNwMuktNjdBkEEN4sxuNb62wMdbua9PCpsw6s8IfeMxrVrHmzvr/dIyQ
jHsMgG3X65lj4y7Nmb19et6NCM1k5MC/e8YgoBDFHj+NW5Gq+yBKy/dVElyxUwC7a65YcHaPcz5w
69NVee1iwe3z0eC6c/XEwZ/yjTVatKk+ElhdKRvspP0j/O5rOJSw8nOJMyzmOF7kNuIvICDf7bSm
CiFvcFS68CNInR9yOShZlEHbJTS8WmkK5pktZU7UZ5GV6yUMpzGhxjxs3Bet1EqmfWk/bam+jcyS
1xyYSau9j9sS+nPCBb7AOHxP+XWBDcwmeVYH7xd/ywpBDpI+jICxwwoE8N4icAneWbMlj5oy0rhj
sMUWRsOrHUIFwkyGmUgb1AAeloPJOU1vGcP13WadFFu+o2QvFO4l3xgO7liYqeB+0lzFEoPypEUM
FbxiBCNEJ5X3uH3qFBTcEWZy4FgD8+Tnxf07WyVxYVdXPoYiIrtl2JbJLiB0gV9Ry33ytcvVDi/P
uttfOYvTHI7rWkpRTBiCI64FCkEkS9HZbh1u80W4q+aC8AfySPSi/AgRFk3t+acw+mc/XiqwzW5P
nVBrtJGaLCTwgIVsC+0vS39mmO3VETrktiFt+2FoVr3MUlDmreWxd5sHVwKNw0Xoh/xnLmBGjS37
GR58+AwpYuU2NVGxciomSRQVNjy5DVPRc6ZBt6lfkxQfDdo8uYfUOnvcC1WFbaGV3LQoEdQHBJP6
oFNtBNFLhxkf9T87yJsExGb5WYU9b0CmyJsydbk0QVepc2zTOdSMeDlXg3RAOg4wIshAWLR9Y0a1
gmyRcAqfjE64XvZ2sAW2si+wmjGVTewHW1AHOUxSQ/p/rb/phuduoFM+Qf1gj/FvhtisLPvfUKco
QLlVusgJi/P2slBgNubb4iaKq/Au6MQINNZ58O5Rc9y2bJ1yhraAwnm0CeB6gNIKqf8SqMwBGazH
Cj92yWcronHoYvBj+CpqwES1dzI+sLlAWgeH7VysAuLwryta0MpPiorD9wqqAl2h1EJE4PYteXFR
tF4oF/mepj/hU7fjadbZ9pbYBXY6P8ydXjZ0epbySF/wMOUpi4SgCNTUGH+XSBqS27RbD92uJkgr
b32bvPLgmJqmxhI/B/GGhJI4yDqsIjGxZn7hiD2OE8Bx8cOOpp0dQkrm02PbTmGNdbZFBZFRva4r
34QdeC+uw6hygCFDBRLIk2MGeO80D1J3rpT82iOm8SVWbWSd5msrC0hO83kIAmKsCHdBYQitaPIn
Uu+8C1GraNulhOoBfm7UoH9aZP+Wqe1aaXVVjV/Y5atYFpsP+9a4gqQKG0KDGz2fa6lkXxU59iRh
8rBILBi07xpyIrqhi6hOk9YGHtU2zp1WRb89iVZC1DPhLDf7QGPNU/MhPYWcAKJgbvdxjvQNcZf6
mGSsGgVIvETwG3/vTMfNRTm07uRuHukJMC0/XxnavIdUSVQ4fUqtOfgXtlXaXA4suRc3JDpmyAQh
1psTc7EF+xFLGRz+vm0rhu6scJXMztchE8TiPiHEH7KO59VpP2jxryibDlJln/QifzsimFo6/+EJ
Hw3Cx1r/E4L9jkxVQ5zulHTE78457NHgVEHpQgfrcnUCg+BPCILmsNA+0sL2UTVBzahwy0P3QXms
0Whj5CJmJdanz8pEHuivbKsKg6jOJmk6UaXXcypH5o8aVbUYkD4K/y6WaN8ZqhRfmA305Fdb5f7H
nla4H8ZNwVGIbIcoMI9shL6moO6nSNTLx/RzoV1SV/cBHMEoHfqrnM9dYLASh/kHJ7uKsn5544GS
FHn23sTNq/bxSgbDZTeG0qk9I2Pup+/XMqiq3EJ4dfW666dbz+jF4LurDrXfNkbp0xq1nHqE9B/R
+dJGWJmVblzIxuF4FKZKvIsn3vJ0GZK78n2Zl8CvWmRsIgi+hDhUVvJLKoN4CqxV/ucW7u+PU1t3
vSC2NGRJiEykYsGUhttXJls4wOeT/pKxw37ueam08BfYfDroMm0u40bqmVfkTbtVBjCXls+TG8en
El92hRhHKBK19sC+1pf1JMUV9YlenNYAv29WGtMEPNQKrd7WNgHBYK7Sly0EppD5uJR3PlkTvz9m
cYqI/c0U143wesO5Ogb26/c/Bv2qOGhWWOlTn5kLSyiDRS67cOlNTz4QOAbabv4EWrUlT7Jp5UXS
2Y5Dea0Nv4x+72xKsZQcNQnv09KU4gqxAWw4e+H14dFyv0/znydDtXrIj/Rb9pcVZSjxH/SegG7I
R7Dlg/jWheNK7ssporpauunxZeX0Nar9xQ5yZa0dgIcbkz4cXUWOB47Jove+yUjMCI89Byl0h86x
jLTX6j3qQmQ+ZPwAY1SX5uzLgIuL19tVbJ3brc2+SLymVaBgsyJQaa+okvtoq015cn7S93jSy2Gp
8Wj51ksr4xpD89OfL87hjY0/fV8QuNca2QhndFv3AUGlknzKvAYMyRehJUW9FMJvGxslU0kNfOs4
tj/1ykIcLDdrs3JAcCslGnvnXP+jVV5c3IzCh+t32GkzaorwtujFChQtS9c2gsgSgf0HczClVLlc
J6SvnM+EKdtYqkTlv7eKNQy/sctiMLynRJUM9I+7zGG6CKPaBdq6HdQ7BoUHXVf3SgECtFM+WrWG
+PBv+1GSRTwJgLjbn1KDLwrmM7NUX8V0rGBB93B82RqflC+3PGSq1DoLjoUGBinO/WjiZ5EQIJEX
FUAbaEo8m6uxwnAZX4khbZlz3KM7kdumayJByEIyyssxJ0YCL8fzkLLFBD1+Z6FPVXpfkL36nn69
2ZRldgTMlpEoFL00Xz1aLwzNWUt/BmaUSpzvzsxi9qQ4SAt8+d2VsX3uQLCHXQSiiwBEYKD557mT
/01akSlCeD7SXuUo3a5AWJK0VD8+WQKIlJnsvdwMWNgkXMiUIpmhX5pciixTXKTueNpdtlcUloXJ
3H4vXWU44DOwE4+iBYzgzcE8T37B3y0nhowTUUf6Z1qt/9PCsH0iv2M+9VQ2NzzJ1KU3HW7kj53J
4ByA+s0Cyndu/+42rVzmRmPL++oNHfmj+//ajZyiPHbd/WFgPDoVSBMiq15OA99ampCRnf4MuERe
cylz2F9ygOt4hurJPF6VMK5l8pn5e3zTmRLAFMQ1KloC9eH73Mpx89Trv6F6IVLuw4EnFYP8nzgh
B7Q7RX7wVwIFXhR4PU2piGxvjPwtWKoGNM7hqufa2HEHAmUvN8ABcX+pM789luvuylCLXqN6KC/i
yKMYvq+LHEQ76tNyPR+qFuVr989uqa8mVMfP5PVmcQodH5DghNcRidmvee+AyWMuk7XkBrLDnxs8
bGGAkri6hsiaG6RAps3vQ32Ej7YImn7fZaXYoqiDmitYDYafB56bqbW7M+G8CsZVFtFNazbkKMVD
TLp/r72qT2qvyJ4mmbJtAYPmtAajAwBv30op3hLg66A8aGljK6TGskixEKLq0RiC7F4zdxnZQ2Kf
OfbHcf5Z6pbQfUNl/KwbD97NIzhoUTfWXBSdJtNtYwiBwtov42Kv0ockHh5IZvmKCYIlflUjSt3F
L/Lcyf3hvCEY6e8AgOYfsZ7dKNGZ6u3+rsnJttbZfR6ivTClxK+30iDu+jSRXESWoSPE7UffiGFl
gWUhzOaGH/11ygv7ZAVh6pVLco005+ZJc1vAJMGIANPv2KUHPAkW2QdFLOoF8S1k3qM39NR2yC3/
pyMVNbrCNONLNKUhMeew7Za/PQE3VKS7ZKX4DC0v9d3rrixqHCXl8Oy11st2t2A9/xpw5XErOFEA
6O/Abpgf0v0pgfWVIOXiE0UiJ0mygPmDv3s0yuZeWea6w7JXrGwUy1u86kelJ6h/Uki1G8dV+h17
LCdOR2f5yZRlyd9CNEJZZzwezNAnZGpA2dGPbrGhnxlOUzviGKd02vvfE9ypWYunjaq6Qi4Ik+h0
FRIctdNihwcTZSeEx4LUiVRB55dPwZzxL79PU+uphyGoI5c2n0ECh3yW0tfFM2Fba0LQv2TWjZyO
IRymkWrve4q+4pH3oU8BAdzebjLiz31mKp+xVAT0DOM7bTWaEYyOPs3uQ8RZPmnRgnQTFw/KuEjy
sSoHFlCuvQ88IZ/q2Csth51TCRaSzrzo8Oy1gvPOhbROLqrO3jYoAraf52sh452JNMBAPvk6Ka6m
rPfBydOs3asnKT9MPFfEfpRpCz0/eZtTC0vbBNAE9maweNlLXngoBrYtkuaUGrClqGfdKozttXbe
NEkX7+an6si5W2N5krZuDEcurjPu2+J0U2vseSbzYaj5ixkD2UNwgjKTOAbWOjEvazOppoN2HT1f
pHasJPTQBqH+mdi/WluYJ38hYR9S7/ZBclsSE0J3NpOyHJ+cLM05FxcWq8eW5y0zXXN3vLEPv3fF
WcXL7IA4jskUOrqL71j3ufH+YOV1MjLCFvEeMq1uJw38VLx/RX/LMbYW+6AHYuIJ3/NnYXVfFQsS
HbjoZ0FmngEIRakbWa+jjVTQylaFM7Yr5TH/8KKpBpY5JgsG1318NYU+3Rvr7a7BpVFVLymjg28T
lq7bkdAHGPUgXt4SYdVp1z9RHI55Le+cPUW47FTnGO7CtkTt8k7B3XFnwyKg3IjYB9gfva9JuPGV
+ucqH2tHFDUm3M5ttvJ4TFRQWoJE9eQRhNcx2jQr42em3kF5nusHYVn9BxpYkz07WeGk216KDtEq
LDdUtnMGHAYIrCGQhsBylAGBZjQJvhIykm8QHzzBBHquq/Ivgak4jvtg3I3UYh+uDd3/KbeosJQY
y3tPVkmZwfXPlRnUMYLRIbwUgzK7pMdnloF+NI8i1BKLHRE3xgqBMsPh8TonZGGi0HUnuDIjsAaL
zPF0sVhgwZ+BGdqggJP+kTUqCapIX/5PSmc9dQjTqMLMinEH2nTulFlKO/rH/bVsfnB0p31VG7rE
yG7kPZS4zSWNu8auJ422hj22pmKuLHRIailqQT8d1fDoxKShTa2NXgmRgBCj43rB1+5GXVKpRLQ8
nVaWo2FzAQ7h8OIBinmL7LxNMz//PTO60zL4/WGFaM+QRF/pcS3SUhwm3ARkOcChK0qfRvA5NZgh
VbVAswkS/U0cpGmcMwlbhHbyh0n+dzvPl9LduP6H73iw86qrEiKmZ8HeUd49U+i+XQ+WvHxsvQdT
SRzHb2JvM5SYWGAVoHqI4D+x8FxGPt5AaVKyeNmJY+iRhlJSfEU/7aw0HGMV4qU4djGTQpWaWW+m
MryHnWZNaC/UkZ/6FOdHP33/05G/cHC7dSnACwV6mQ1TAys7XeNrdKc4N6iSmTEKDKyZonEyBkK7
xJbcrUGFeTLly2fb7jCiTvU/9nT4RthMVmdEWfbLLJfBhp+PaKXx0BL5U59IJ+44vt6rrbJZxhyM
MTxk3iJG6uj6AMP3Nugf7sLuAvvxw9P4U23DbOybdJFrn4nai7HS7SFodTUtzHQ3pW0o54SAyuk5
YPgDS5VUAP5bjD0alzNZ45FFnPtaPI5ft+ZJoEAiIb4GaFsJ8glEjgqYEjoBkCxD7XWSKTTFozHi
zoN3QtMDK2WW/zxnT94mq+fKtqgcrzpcg7eesm66yLE1cYZHivGJoBgwFATIljGP9bkJywHAOuy0
NcBeIo9yHDA1HhhoAAy6n5YCSP17dDcEga8kb0ofBS3nfciv568IJKEEic9FgpPqp2DQPNr5gj8o
oge41RMGpRO0OcOeguLvMZCVXzPH7+topC/Cukw8h945VNqRGC34M+3OrNNFP7jaH+uhZInBVPWj
wURwjMzwQS8BXIc3qxmwRDzyqC+4vSXKCMNreaGvqDWoihcb8naoQTgzl0M2PM1EjVgZvPmz8LIB
J7LqUTt3CigJDh054Sbv9jlG9Cp7/gNbjc3HXiEoETfRD7iK5S5tdQTAkQpW6DqwrQ2k4gyO5+l4
mTadlHlKkXEM94IsAiinB2VXMmpHj57idXUFdXkpWwhEruUqTBm7SluQHIhQbChX+jdAEgH+3+eL
jSXv/PEpkAZrpfAojOy0YaA3SHjMDUadSAj58IvxQiPW/r/AbO2ysGrEb2lmT7Qz3oDIqqKjzMmW
8iOJwlH7cjLPryFdOfI7x/vUWVEJqiYPZK3QlfyGkL9HqDTRRJFktxlBUnbdSUq9mOjvWHidaSeb
kUfz+HeMMJllbK2Ac/4LmidqcVeG4B9HEqjsqCFltEOp7Z8ErhZSxThJFJv10M6Pqp3DzurxCMQ1
usIf1X0kGhQHeRYvau+xTKTKmiA0k9sb3Ckvpo7ERLrDFptEi2YGjnO22wGerk9xjBLg9+AbXSIw
TuLxoGCWROi6QTGgdm6di/ei39wSje9dQ/+QXrkmx//gzvOoBsEt9mNj4N+63mwgH3eMirdcqHAM
+Mw2aYjpL7E5Mruz/+ku6OxYE43UJOeWVhyKLHtCj85scvdDXp/o1IA1jX6nUijiVpmzIeGEISPu
jD1KgFDEfMhveBeOjt/5YOYj3ADH1fXXdZj8b3i3vy1aQJ1MEjd7okAo1FTo+VRPPzV3x0KPziRW
mERNpQp16ytUlaME192+vieGn4qEEl4lhNrZ1KhYssHQLFlGDnPBrcs/IWIHSxwl9OG/OBZcqO/c
Qjff97VhdMcfBqxE2zJw9quGejgKOlEPxOHc/+dGSHjievzwJrHKDkoPhSBA0P0z2w6rv+mNp8jz
WrFrNhbj7hW3oy4FxTe7JS36Rl8YCaqyeD/LZrgNsYo/ODPBIbE4wPmcdJc3mbA5/t6A8JN8l4ai
A8aV2EcWW3XnPj2rDndwv/LxyjxX2r1AIpSOuCQq7+NbD9lHl9B+79meFubvKDMm6LmBXnvcEv6R
lmwZTveJ0z/U3g3kGexLGxVccRApIEf1b2KAQGITKLZXrg5gwOBrpzQhcA5AhFRV2CY2DhrY0lS8
Wap4i9ZBMqcZBH4y1IpXKBXb/yZ0bqQXIVb1v7rLQp5Fg1OhbQemvxXIrpbHx7UUOl7xGj7gDIgH
KXetbEvexSd4FNi7SgrRhu7jnvZBMguTeWj8BxLS9ION1zRwRUNEzruEGMyGaotJy8wXG3r9dQLb
vl0/MWGDMnvBR+mLQpchEbWdMd4GbDNisshS0tSlnbUC2OgHFNWKeHI1G89UYimnJZXyriUEOJKs
oh2ESvpu9EP47LvpmoZETx8CdrDYxSbXQzbYAUG/d8Rtv7CG7n5pxfH7jDGbqBpDzbY3V7Z+JvCo
7O2ynhPbf1SjxtS+vW8kgNG9BvWGDgzFQ6uUcax14JnfeGO+YSSEe87MYi4qJWn74/gMHD6a67kx
iFzdptudjOyDOF8CUY8zRDiTex3/VgonOH0Ty4AaN6A/ynmEtsT0c124zHI/hmY8Kv07tBQ69skK
B05oT/IqriH1t1/KZ0MAx3aeAkkgXsRCgL1fsyERcyjlTr2luW87fKMzTSMwMb6fbNntqo6OC/R6
APNPTGm9c3gqD+puzHR+5OGACiAezz0bmRYeH7ssI+qZji74WouL0tow1U9B1xJeF3zboN9U8SEp
Z1MT2pqQZ1dHoD5kwS7/y/epEbj7Ky40XQk3nqmPL6TB+nQgr72rMHWdAxlatokjJQG97/aqq0Ys
njKrtaNHzy2BszOvo1M2I+dR/PXvGRbOVn7JDUyjzdh8o7DzHfgqdYqabPNI07qq3mJJxn7nzIcc
SeaovUFBMlLNzfbtgU6WLKO/32NDh5sohzDPaJ2ziL1phNCRo+MXWath4mQ2Gbdj8poaTtTEmQ+4
GSehRd+10tYYrjqvNdie1dFRph1ybaZcnGNB4zq1vM7PddbVwo2tABZjdoMpspz9pVtKlHWGPZ0K
nHDKF4EzIf1wKXUH6Kc+9IGk0iMa8N3aHwg9mcmGue6A/U6xaXK1jK2RxD9me9eJUJxe/aTrJafq
jNx9ycuUxTVwSuB0SSk0MVDayLJXMMDURpP4QewgSz9i26laiHurvSXh3ucT6D/pyFF2/cW0riPm
dqE0yDdx5RjhiSH9HAn6kvhJF36ogfhTzmqX89lx4DpVZa9ixXZyuZlrA1lcbnygKfgy7NiWiBf7
VKQGfaqwoXJtj8qrsZyxTf4GV7AruJ8uZJsmJEdBb0qBVyJvqxyhRiLZLNes4+uhGLWRiAD2htsG
S54lJFqz2pbYTDa8uHmTPLHNro67r9REfvyuiHQh6MMwtNRnVQSQchWqLN5BFmIfgazjn5roPwUk
J3IvnsDsrXvugagn8rBqeAD6yJ0p6pm+LDgPpij5zuJ0IHVdtBUWcdWXWSkDST/BJpSrqJev8ldJ
3FjMDPgiuoVt8siUJi0Fzr4qYt3wC0SlrRsFVBXwZ+Vvo0iVM3Gfkz7f7Wlw+ziGaKTqP8FUdiyw
jpvf7eAMUiiiehSMlREvxSqv+J9TJ5yQOfrkpeUEJefs7LHKQTdZm/jswY8ayAml6/b2XqwPsUue
hnDhM24yzmLkjLpwjfwv6rTsFXINMxek2KKsF/49gswI4nzVn+Xrz8gqUl8X0gc3yxQS0P83B2ur
3pT4+P9mmnvJ4zvqZ762QfInfDegc/HfF7RNHFOpm952Nfm7+u73v0a5FsGNgywo5h7Gw3S+B3UY
fFTelRoNumCfc5tJAEcu9adPoPsXxbOAAXsVBzEdytR1wGLxmkGrj6gpC7+atrFTYnNBKXTxbuqj
OX+O2r4ny0GL0PEOhC+WEJzDQbZAVeWr1ZV1qWXIcaCyI6eUAOgHoWKUvRZkKXNZc/x/25ZDPKOj
/lvp3OPmbyeiKd6Qn4FKT5upM6tekkrUbOVlthI0nCFeLPQgswQK/4j5+TtM1AJviX66p2DstEKx
3+GAeJqzjXu74bPOLH/2wBG5aiarvU+nLcjNUsTzHBtTSdRg4Avzr1jLFM1OZnVqkCFbuBrOhRoN
Tmu4fNciG2s5PqrCAWUrMTUOaZTJFCDzSUgFpah8c+YNgeDZUKSRD9HyS3pOfDAGo6hWYoAUtZbV
1FxXtaH/L6afpHPda92vHF0BEFwrfwJ27QlBy7m+zXIsbHd/JF/JIEPmeqSNeq1MB9oRgnMQf9Jv
FGrDynl7YRZarQKK+03qhSlo8mUoCT+Txwhbd1bRUc8mJMGFw2Um01cYtBLHTIT0TXH5Z3dvzk7x
oU/ChfXfyO+yfMwJ6iHQ/SKv1B703uiAmyqu5wC9E2o078BbEjO1fIMqmcrWASFHj37Qb2Hhva5D
recivOQqdwiJUleEuExkzL9/JVfrDQs7QZTvLsOrEKXPztcquImSLm2Aw6JLa/X6qJWXn5FmXoti
cUG6nULdbO2y80QZXcjSZvU0093JGFV/DLSKj/ePV1MCgi+HNR8NMWP6xJto/SK1dxOcXXHJOWOk
7f+Hg2HEEzkt6xN2cz8PsoqwwgYL3JB7NSwmS559zYbsgM8+XOhtRADLSFfWXXrQI0648YaASaEf
l8pjISHXlVrap+P+bOmHTLfAUUw/Zr1NeUTNtH4ZcH7cGPgfnwZ0TsvPxIgHXLptD1d1Sg+WzusC
+zakP5WlQ3b6l0TFS7EW5SPIzJNG+iA0g2/1BlvNLtMI4q3O+iU5eadmyKKKQurkj/N/H9FItV09
4WMt9Qq/MqaX31y1tqFkKJivK5F88Fc6dgbr8PlrQGJsBe4T9HbpY56pbDvvTgitWF0G0Pg1hTbl
ySk32RsSyrvQreSpWsMXv34Hk8eiKhgUJPNx5+MlD56vIncZzIByX4bInAMiVreQOneuq3beL1XE
4zKBAQD3GtDi+mPA6yW1jND6DkEyO3csy9oQfLx7qyJnOXJmiRnSPX/v9DXgAdw9taVg/bHXqAZd
1l4ep90c+VxzBsVw7p0+OhzV6z0dr/ZIa3P0w12BL8ikMEPgl+scwLU4udpN2/9jxr6qyz6FZM/r
IM1QQrIQp7ffCdfn0pBcNduZ2Fxh3B6jYjq0ybrtUh6/4KECx0teZO+kxVHWePpx5KboWeN9o4mH
9q3KZNbu/JpNqrbBJYz4aahmEK2CfGY5/XDrIUJ1XD9J48e4VhGKa2mGgwW9HEx4sAlflCFDfnZG
2CcP0bBkLyJUri8veGOBFe8kTCE3xLJ5b8uAzmHFfxVlNS+3D58d7Jyg85bUAcCgAa3kZIZ6tp1T
5gFseqHWkcdPcc20yxTCrnoTlSpP9+y/cjWlkktUXS83IkbdYJI7axENRL3xuHw6IxE9Ym2sqDEz
+nFGwtkOKuvnM5k8y4CdtiUu1/WsaZ+CXYwlrQ3orRdNXYmC41rGxHvd0xc5eutwl0e33iwpVk11
DsCYJGTZqV8q/gnD1YQTvGoNQbh8tntuLa74T7T8KqYxfpVYayW38iBzAwZ9Qd1MWWcfosMy0DtU
i38BDy5FW/KAPm98SeyALXhR1G49DUPe9q4X14MSsnwpebFCj8J6ogKCMfi0rORoaKorIpwhSdw2
qaGNHkbEWnDSmJJMdght22z634oiV31nH7aVmqaYO4I2VeyGL846vqIS0NMDgOxE8Fvmk0m1Hq9f
6ViSlBFVuAnueHxwg+eFllGHjaAgSZWOiDF7eYCPaZCbIqcKsV/enlKk8JlybuJb0x10ABgqBLXQ
agqwW+sUfUFngEDjVxvrDGMNqUEIekzcATHNyS92BSHR3LunIB6OeoUeynWd++CfvIlKkq/R0/3a
gNFt6AQSior72sFdnDgD8gy9M2+XHjaQR7WNDolWorkk/r79VGs96iHnfH+BO0pZFY4mPWQUYJGT
jT7VVZg5HInJ/j9Qn7tjQ9UPs5z5h1GJoUPlLuibcsQ3S8OXvgbkSStXz7clS6yMIk+9oXoWO0AU
IjNhGM/wADXZe5UUy/OAa9MYxvCOSehZoAo7FYMPImsfM6B61AR0Bqb8mqqNOKXRU+zlqp/Nd82x
b0qG4pRDUckYUVNVxoHleRyPP+k8kQjVQ4WQcCfFgo0v+YbRgoUusvMEA8/8r8phQphxg4tghY2s
5SJGURv7L8GtNDj1XMOYFvQJzUQoIb8IN3psfJFPSD/tEY/qI1bSkhgeo8zPQ87gr9yOkFaYXfLo
qjWN/C+5ZDJEh71GXGHA9vuvsAGvfq69Nsw8uW+6q/rAGOZlpO7BEys0QCJSD7vWXEENvQcvskB3
iGSg0akqhFlt2IkfyEA0ZiMHqVHLE/W85g9mX68HXsP6alu8WIzN/hEWgc8TAueWumJMNB5L4ngk
hv/DTr/Uyqt8cb7H0/C1DIiCLdpjKV+Bn2B7+jKPjwOnUzIisehfqM60fDMbKHSKdGq7WoV3tK1M
kRcmgvYeHlBZy2cnQKW2mT5TA6x2lvtTQK7RVLGFjpaOYVrLLij/IMkhq6u4wx6Wq/LilhcwyE3G
Skce9ZbtGHkMAsNie727KtbS81m5pInT9NMyjMaZfe6OxzYnxI5qG+Y21DzFh+4TNMiapnv/lLzn
Ti8vttq3CMQ+k2DsfRsVy7OR74K52KYoVra4QwAVy/QYDF7H6yjWJZg77JRp9tKOURV7ZqjlqXT9
UV6WCN4LaMV4el6Z0Yjb3ozgGG+Bj3QglwECkoBnEPZGxlMYexj+0jO/sWI8YykzoorzOEV+io4S
MvL9fHE6+NwFSVOF4HYb/931pSthAJpoCHP6rUIQHi2OIsAOIX+HRhUnMoJ76J51oZmed2Ljq8F3
XYPJOGB6FDLxqDV/biaGNRyuHWUaS0F/SV0QaBH8rWprOayB+JXfg6OqmZ3hsGDrutRNY3IsjngJ
q80xQn0nAELg8nyHE3CrEXxpV/rf/mXOKPuZK23dMurFyk5uykmhf3Yy4o0RebeWZRe4YrfNUijU
+a8Nt/LBmfXMnwn9ZMAXEu696C09+9ZD7BjQrmmEbYgFLRRcIY0gEHhdqbgL1Unh0HDpHSUx1dNx
kSV8htbxJ50GfojfVVDMNmoa/ffgeHtFHPeA1I8XyweDl909q20+qhD4pdsHYk1LyEmp53WKPTBe
uTkn0BaLEsbm69vf/XXTlyMSAxVCIEG1A/hkPny7I+oZmjxcQhKYdLXTQ/pBmJLehvEYyavWvfi1
sTqgT6S5ghD3gzfmJxdv6Vn1k9+4zfJYjwxE6385M4GqseNz1gD5qPNDWxD6ekZ0LmiP6z8zpemY
jtD3W8bewpMwiXdAJhtNdPWThrPydSwC9fw5hHlG2yuKhC5X1DwxAgUYXQllP25N4bNoR1fu+p4K
wfrgQC1QQ6VXDZIYoYSjOe/AfBHJ4Vlp9QDo07inpxh3aFYyYni959Pvwh0MOqqd4ZsLMBfl27Ot
BjZSkIZq8jJXz89dM7YASe95NYPa9cGmigbCFg7Yz+5jCpKuAONrEYvs3KvKQ3EjUbb16VtBdh0p
BKhxbTxYZ3G0JsJ8RXgcECpfX9ABKUnhn2S61kHkk6F7jOKBD5OATiLjgzvGjEr1AUXNBW+x/A94
IL5jW6rlHC7k9uLRwRQ3HJuYXTnpgW0GWK3gDlMrsmD1+IY24wf5G/ZdZ9P8syKKLk7234TiEGxR
iNUlyF9kyfV/wIZb+NIvc9BEs+ROcSCHWW2HuRwdGeikndCBjzNKovA12Jw9yA8WiTs9npfiCKon
w0zw8O79vc3ezDs///rK+JFOWg9Tdq9jVeZB9dCpCvhKWKLjGv6yb1rDFjK9O7XjP8qHap4D6M6L
Kg9LJPpuq+KNO9rk4RR6fPoGxBrXgA6ybnv/7tOj0lgAkQZK3rK2T4HKh60eptsKmqSQjBAHCLi+
bFNRb5xMxfq/DGVjrfWxU6rdHXol+BBaVDrsIXnLeN7pzFbgJAxgdzL9CBlKZKZc87gFRwa8cB9X
+wGKIYBU4RmAqvlBhyIADYksGqQ5I+jXPIO5GhDToa2tAVbmX2a6b8piThx4xsJT8/C2KGPyHBud
pzr3RS+VN305wYgFMKUKoXb5NWaL/7O2tY6XqjmSISxcm6hXMLiXSBwImlCddJiHcA/xnls85icz
rBXSnQrGh2TJaICtNRYjgLHc+avMVjkH5P0cEPozSsk80FG+50GlwU337aMNLqNVV8Z0+3YG3z1o
wCJCYaiM5Gy4e1P5mfFS8NwYr5MMrXuHCJuZTFJK6pEAqgeiq/+IgD/OvP6ExfEK+Aq7oFnj65BQ
Xbi9MYN5aZ6CO8L7GaCvDM8NoKUY8P7YKUy8/2CONMS5Ywj4M6oXXff0a2WLZxxtYVcBujeKBegH
p5KetIA1Z9Ibrl5fWGYGopeBY4g9YWOJD6Li8ww2+lej8AbQd3Vkd/VNlNYei7jCOBocS70mbYu5
83N4DCivNEvq6360Tj9DpmanIDW89Rpdxm8uGhEHrpkGnCAmwYde/sy6QSF1A7EWXrsfz9ViiVJQ
6/URgUTahK42XZz7ojkzOswpbpF99r90QdKzr3JiViapZtc8LZtsKXeRyeJFl/Vq7XJOtuN/b/9L
73vHBLdtb41l5DW+gU0o2wdOxFgdPBZaaI9EntDDonfWJ+x3OdUXGWe7KjdRusW+ehKjEocW7Mg1
ZcVXX/Sak9SXXULvWBUJ2dx/iLccyTPGBUUk24EKapOvaI9MQ18IKRFri0g08wX2emHks4DGgVaH
HwpY3MLkgs8Wuj8xzuIpyvBRWivPEzL/i2TljjHg/mv5HnzMhCtDTO1VAGdJ7S8Dwx2NiqsbwlAX
ZfLDOLZT8YLKoU4i/+aEgBzeKk9GPps9UtiyENXdbwtsFnEgS9+YTXbMhTRMmQyfodJ/tdeNvNEU
R6yNS8IPTmMRHcmfutzxGCMeUpprkHWL0gjRLC9li7K1wM4jp0jL3u/Yhug4VrGYrEsDSUs/Z49M
xbWGlnSF9IviIA+8vOCTnhQ1hAYbsfOYoSNGsnVtpt0k1c0jW5FAgZ75JMEXpreiUbWhpwBHG3bO
WoYVrX1Lr6spd+7EdsByPsktAv6qrpfuFE1HSLnV0gP9IdS3dEsxdmLh4MKu8IT0LWHa764h6aWE
IOjOnbMD5vZ9gA0Blug/ExcDZyNMgUSS93d2Vox9b5RS6KogthbMHIGvb+Pw409Eyc7gjcgwBbhz
NxiuedW9KebQuYbxCJypklEcOV3z8pK1AuRnV6o135HvqP4qT0dPoBMRSzsFm7vl19G8152MyBSp
iIQSlz+iFEZFs+BCTWXoxffa7HpSVDeDpB57b93f76GgjrBaU0/QKbsWrU8Kre/q7H1Cr/22MwYn
mJpfynJ1+/aYwfHGampQLrgXmYJz+U3B3zTDQ9l4bF1BE1tFw/ZDlByJXSoBKWiVgo45MpSzEu/B
JOzwPY+L3axiiZL75wiFQ7hRct4h3goNsq6qaadmQu31nNP1C1KtjkSMMKGPvXPHl8Ph/aehbsrT
pG5h6vzFhm7cDSn9XXm+laD7UAAxyZBrdpT+uzB7oIZYM4HIFFhIzpec9MmPZiIwv1YYoYXtrnmw
mPnVA2KIDc9oAOmOIZS+3G7XVlOPe9z++UZVbGV1i7Y6mHDcgnP3AJqsZVhD/tA8kYgmPbYFliK5
uZt7DAAQf7lP3X7UDM+TcIxmJrWLmZOGSdFB/irdNMDsj0MsJHYCM9L0mxYH+DWD/SVIncbB5yUi
09FTPKG5n8XXA6m1DQ3nKLFsWORd5ftIw/ULTpuJo8qXRZ0fn/wXgASGbuD5DUGrMG0JVz0Nh3x0
3nJAiT1TWqRlMeT4xxi8EUWiWPe6R7qYPhXUDgq4ndoiNZnL5g2yjv1wAoydDbJE6ES+2hyN+e6K
eU9Nz07rQCbhSlnhRhxzZEhwD20tG3q0GWMGeoayaRNZjJDVoFVLevKZEDjqwQm72tCvtTrbJUhc
MZGLKNwRgHr5AL/qJBgzhMJS6pWKx254wGh7iSoYzt5bL9eBPk6AE6hYeofIfxVF6xYLmeakNLCD
6Xnsv9YWaX9PRdLCjiob+OUBAWVpouzBh/RhBfKlzOYS563BNG8SI1+ZRNEQUbLklYqJhGTlF8z8
DOlka9Oq93/kj6U3Hg80qxUyV0aFkOLkViMfIVHPeBSinDiy1rBxOOva4DleEnxAaOfFDHlg8hh6
eRnmH2hNetWitwzEteHQJww0X0vt/PpHIv8z2SHg9i613/igSje0PztNZoD9/4bRJuQd2Bwe1TDP
AJE3Ech4OoBsU0NIU/3hvSma7nFbhzPUyCYLWwa1pWVVN6pcVf8F1N88Y99kcqRcskPqM1IqiKxy
agNa4+0RYFQ/qFestHV9osQDu1mW+TJ1WkU2T+FiKyU+juUxdeG9T3zx+RMc176sh5rYAImWC0+a
Gf/u1ukybUKpX4sQI53swHKcwdOybWZSWG+OFEXl+pQOzBLgAlLPvZYjwJm7fh6P5q6xwcC3OHwc
gClzO1o/BtrqO6J3EBqv9ma6ihkfibHpq04dqwPp9CBtv86brkRbATOeSJXfNbGM0mMwLnP9+toF
Wkv1wPzjP0I68Lw5hkC7mThjhKWnNdz1RxvXn11LLkF/BYhZMMSug6XoBJvz6g4o0lxvFmtzBMh+
FKHv9jiABFkZflnY/Ye3C3YbXnOlREwFsWImlGOnOsq9FKtXo2XoB/IeggRDYr5777kyD3CKF5u+
R/ABCmLILkO5qFnR7hTlVeCOqePH/cqZw12tx0nkxpHV870A1LprTDm8KfjLj09LK6bI+6QYStpZ
59LtTqW3sbMcdLt1siKJsoUXcA5rPbuIwgszW/HwTmzzVuBSV8xCFcMxAIxjdiP0UvB8CNS72JDa
2K55ESZVvY+EJ2p7f5TIUG/jQ4ohCwdF0h+1TJotmEpVdYSOrYR9yzeYYVbecuT19/gIpSQaFH/Y
/UAINeGiUvdKEtiquREvDrSRkX5FsUfu95ClgWohNOM02VROCNb8qBReGzJW2DV97o7l3zWcpKe6
2ZFCchOPI/vhJGHuItBYcy+90kLyKZ1GyF6/VsF8OL8bjOH1df9MSX289jLo0VdXNQ3HX0QrKIuP
9+sAtPoVSvvdcuSwtKdnV9TaVUnJFGSNhiDAFLHHdyl2RicgZ8GhDAyaSazGzJwGzTZnXL+0zx6u
tN9Y96SLRF1nE5ZpcxzaGD6HGDi2XHE52BI3T2Ugc8BAwwpf4irDvwWCWG9Gwg+egI8l/NeAgXM7
CQKi/ceKUFKJhEu0yhBy3LoXAEx8ECTIm1hyl+zfxShCtBjdW/zfwmdvIt8obZA4CE4cTg0EChO5
Xle5n91938XQe1/LpT9zu9nbIqYgMFhfYeQU6+k4UAw5EPjxoNSrlmPm6xZjHNicHY+DHe8rOlOn
cZFufZM4wrKxLB/Ed9Al1tpgP9+xYNmaHF+s3mvuRaKbQuCszVLpyOGGdHmTqdHv5dQIz97LF5kp
VYmnHtThfB2UmMuVECBn3ZCuA/BkOjm+iv8KUoTNztMtkBJn9T1ubEOlR75OjCjqjiGy1RuQJjOB
lzmZucuMuIbsexQrg4ecrYmeNRFd/B/b2XSkdZL96XpzLnB2OulGAYz1W5suiZXoxMIvWvCoYRkk
FbovYE1y9RD33W4gX4p09QtfAVg8Ejqq75Go3pDGL3AKhOZG42pCSzjS5WxCOATe55SHK5C7q0mr
pjIGP/Spo21mwTBRWLrBlGIn0H9SnJm6fvs4vU2eUboswGpHq9hOWV5kcONO5szgZlQVFwtJVNBX
TZTwuiybBC0zvKNMHmwWYnjmOlWYxssInWk7IfLlOfqakLzxrUpwMgHwDp4nvQo5BnpJv+XcluAA
/Zw0GUxxv6Nim+g8ifIFmV94PiQ8Ymys6y8iWAnjrmrqiKnyK0oVW/eL3UllUpNNJMKL2pXnXXZD
fxsA5D5Nird4V4nhDtwf1tV0UMdeMiUgRNbpG5HvzO0eGUmudgt/NnZ0LHT8aML38enLA9zticnj
tmkmpyYfBQ1Cs6trJya0H0HD8+Ja3norKrEA32VCaumgnSreuph4W1wzeekCRHCzPKHSQPJzRGPX
rOXnx/neVIO1QhHmyxke0TyGHGpPiTr+LDUUjtdHAiFivJB5mkp5pKeYsOioV8GinCOIeUiFHQOL
7Tfsc44SCPJT858stKZak5+GcBIP1oMJRRG/OqrX18R+fq8u6gk4YvbyCoRTS8jttAxmHLFOaghd
ywOO8wjn7mvite1xVXSSVe2zPSIFdZOnOjLCXuWUb+/lRdiQFewVzZlVgfzR8/yFm1B7wKtEJcbj
800z6QJmTA++ZsCDFUIXfuV+c5d5irRrfUqfwrOaozTktOx4Fr2IVzq4u31QGVZQky3Mpl8t058b
KUCBM0sYROZwL7pY2tHp4rB0pwpz/LWZRMC1Ztz1haz/WYikd147AvZHfvu5Y9EdGR4GiLxveqLB
T4JqHLgDBLvjfTkqykDUyOj2S3cYqG6IBwUzStwB4ponvMF/fvfmL+mJ7ikJJlIvubtuD/U1Y5WL
UE1x1qB9Zlgc0djdeLKcr5cYUfT4jKBrk7fCtgFdH7Vos4cRHqUjLACIPwf32W4W3RtyQP/a+60y
0ENwtszIFDJyH2twFzkquwQWhjhfDxhxRqbYdPS6ShOVVp///jtKmSizKMu8yKbss+3bj/M4uma+
aQjE9vTJxB9SKcZcNvgHHuxla6bejs4KGyFwIq4yRBlmlRVaJbIRuj5xwbST3WfsLfJ6GCyNnaRn
2bBQWPrTpJcxBjHJ4w4OTnImXGmqMUxWnDUns4JCE34kIMvbQFAou8NeS6nu1IVhtDFTtKJHiua5
0G5dvfaVvwmnMZBOlm7SHisORKqigmXKbpppRUe4BXkIzpZVNLLNYaWKugHUVQFbZdyHRsoSQUOJ
2XGnmUj69BBOHsOtkzQ3rv2wVdEIZfFb1TE9gMoM421LcI83/ZyzME237VIx6b1LSrnqvSoEcCEw
1L4vrZI0eGybx0PbuPfk525cBrIMI5ppe0c/g5kiFjxYGP4Feymf3Mi3VreuYYHPqdenbWARbJQH
LnV9thTce7VZUXEnouRTXnun/AlDljbZADZ7z37e82hLX5zcWwgdfH9EPq6WRSZXLJrsB/0ZG72g
TP0ovIG5zooagC4pYqnmAjSHfzfU7LrNyoRzrv093Jt2zywjDH7r/cZL8foHMlA+B8fheSFLJC8A
K+bA1DN108eCQ8DtMpgr3HuiDn4dayLIxUoNXfAZ9rSqRP1RHgMjKws9Zgte3tU863thQsX5yj1/
/zhpgoJk2Iytf2PX3thHrjzRXk/mwnjq0ROppqJ165kOL9JTCPqP6S1D6lKUZAh3g5B+gTmMcHJh
XfvWQ+AwdNuIFloIuRT51dkMnpTmkWkKlqxc85gNomMhB4YktM6yQBEKA026Q6RspMGZCmyJYWAS
nER7RYTS4XrJIHWPKnYSiAnUl1rUfTE6tctRIOGG7+haZ3fyCXVqiWSBjCDGKBWzSzoj3gZAOQPg
+HblWwYq1xQImJmPou5hUiO738E7AZZmpVLJhhba1bqoYaj1WKWVL5OgmbzulbINXhfevCzf/Gjp
U+ug6VZGHfMajEgGUFlzgCEbvCu+LYAy+I+dCgAv6mpyNS2XnaIzlFADSBWicrriXShfGLpsCdHV
z4IC6g20ZyBcbF8yqCLYTAyKP7rRup9TVFHGxLHzmLrRVhVtthUN0ZxWFa5DUBUCpAqG4M0yPDJ8
RQouRUJd91CFp/SSYN7ERcB31Y7tO60N4AUxUTX41WGvwd99ZySS7pwvx+01rdffW8cHEuYyy4YQ
QTNT1pO1xTSEZcWSMMK6FTwDdOj+q1Io2jEi1NhCDB3yGRprekMtNQQAnYtnAtlp1nmwxyFvSSE2
7zbCvyKPn7IvOKC+N1wla5DgRjx6p77c8kkHawgNlufKUWWw8sDIZj2KEkL56BToRo0mU3f/E6hX
K/zX6ShOyWFrtlY2RPNROYWoSep0rElWNslx+ZHDDTeJ0qMplDb0oSYoDxik2yCzxm30nY9rbuww
Yi9pfYguufLIfXW+BMxU7COM48ANrK22zB1ED8/ADvJu1zNYojgsGMpsh52qAOOSKA4cjUfsYRyw
cOQuaxOXB2+7MOiqR+LYRnuu/7WneKaOdcMhY8ox/fPcVIkqf/09Gg812nbkWv+1YtSd9ldOeijx
EBG+6Fq+WlfpkUWRFieASOc6fpbdkpZGEChnJASt/QMKTxI5sZnujnGZHFFa1vsga1/vHsgOHFLw
+OhacQsXzjJn/1jUEQSxpnGLWpyTk4GTaVwhXkuktK6qDkszq9RZTdMV+m3zfqJvkfcGQXnD6irv
WdJDAWSoPpFqKt5K6bdILvV0xkKswtej9VQyq/NkGCbDuqO2K90pospbyvgLPhz9HyfR0dh4KooZ
38fd62UKwG14SzCDW5yZCxMy/sRGm0OQEvTPmpaotGdTnmTMLNKyb2G6j2lD+5P9A59I+1D4zFCJ
MC4WnFWgGBRuqDtdhozP0r9wK5W0HTV8hyTGBwA3yYXqBfojsNInUR66LrcsmtzWxpzOKmiLa2uM
/9gXMcwsMDyPvXWPa7cwsqBEo86IWrzu+Yhn9W06Q7L4SWCvsBzMAflmDDyV+6WKOtuckD1cwcsz
e77ksQaLSvGUo2du/pyX+iVKGYYq2VpomOXx/9RNcC9HKV6ZudtD+VUb82fcg36HxNE3OcDnoYHa
FQwR8Razc1VPzWsIpG/uv7kEuN4f9A+H9pwFuWMXl/7QIlITzGOGHotFDj3is7h+cWoFShH5H6am
OBVYP0zE4Ix1D0oNev3Dyg00NkzTy33OYmPvWF0Zqi15nykF2v3RFw63zzfRrKJ5QE+1Tc83r9ZZ
+W6Ft+3B/htE/XUrErwoZFpxE2MnvbEPYspek+QWtxOBMJvnemcAoOcrtQEV0PqBP3zS7JvEbA4A
sUoN51JgYit8hewv7s4a7s1mq6S5l0oYOADM79yG/GRWjONWO/jxs4sZ/t+Tq9oIak+9Egwirj6d
OJ6/o9P/CnmVxu7vMWV6nepBq8ss+UV4nLpJTsmn0WRftI8Aufvg+HCP5pDYB1+jP97lBzBF74PU
geOyVot6us5Bk6f/3Hk6gpMu5QiclD8NCaeNrXbVm1KmchkGxZ9eyvqmT3sjlpv695xuJNlNNMBU
uHJv7W47ug7f3fxMYP9VCYd4H9LuEiR5DfJQNwsP/Hw9scUDqJ0L53RmgU5YfbhBr8IHRWQl3pNf
xUu6+aVzTKFtWPJ+kZ/ZoHMr6QJHOBgxFlS3+I01XGEQeP5xnuqIqku4eZfbNSz/EkggdIjr2962
r/6jVdgkQvbbna0wuONhFuf726qpSmBu2MtrgiH9t6+SQ8xtQMGXxu1hmc+qMn+rNfSsSrJ1NOqR
ZY2D5a3b7aK8lHnU3c+vQIK9bOhpAaO4F0LNsl4pMIXK6xyO5q0WN4SlFNYna6PApEX7eO0emyHW
+AxKVUgPjKAn3BfnRLfLuguE2pGCYiyffYrDYoFEmXXvz8lwY4qCqIJbfqkZ4fp7EfEul9Nh99rj
0sGeEhWVZ6s98zKP1hn68oRB+t66Z2pUBTH7ANnuDL27v4YlqaiN6EAUsznTQi1oLDs7K98nxhPC
Io+Q17xjlj1lSRoVeCK33u6Xmn1LiS+iBq7ePsQvtLb/56eCsJInFOi/QG+ByvkYSYqP6Xqu7bdA
DWUQf2Td1Y+49Uv7BTVZEM0YaeuIXgJ4TIeMr24RSwB2Y8RzbPSKTRyetZXkdM4i40mEhXCYXbfC
zsSqwbI2zb47pEWOcAtL3ooGqP+BMJfi5hOzLlp+gliDf4LUjucYF0KsiXZ4vQgn/54msM0sXh5k
O9S3+Va6nmdRm68RQYsW2ouwlgu1h3cJ8xDjlxevK0y4qhPgFC0DM9C7p9XRFBaCDdu2vkCt8xFa
cL3+5Y/qQLY/R6xKfhR8/yXnreaEiK3hvtvY0soI4k8gSIvpjlc0AT15DioxOh/3h3VJLYcUnwsz
Y9g7OEUxb72ppvzxCR45oOqGsS/ruGDijLwzM4gp7UR80uCUkg/ELgVP9fP8Kzffjup/KRCDHj0e
tLIWo1utZ2TS0/QNQCbg8zEE01sTgXRh0nw4UuXtisbJvWkeRidJJybiG7p/WS6KiXaNH5nAUkZT
LVXyJK0/4jnkuJhImPqRsPFgSLBrwf5Pksd6av3LE64HrBp0F5QKv+QY81ENPw5y4WYLtuWeXu7S
7RpA0Fgu3BmI4ZLSLsyhlk9/S0bZl9HTwx+3VpBRWJROOwmFY096Gd3fEqHHes6fAcRJ4iqcomkB
/VzzbUdnzN0eNsN1CSxxt2w3QjmbFQJChNXVfA56Ssxgd5cKSOKcs8/W7Ctji9MPJjtlAxAoSP+g
rdLREVZa6Llg7HH9UZqWShmKSQV3EF5fQX+DO8ocjYSFsLbBUs7AG0yrPcaAPtmTxA0vt5+3JqQU
UnOZAue6oO7Znb8l00RWaCiol3nVY7YD0AIU6tg69J2cHKqhMWN/V1z+mZSNBXImc0jVF37tcdBh
0MEl2FQqs8SXjBrAZP2d2PlrJ7vNVO4Y91y3/oB3a5MOFVraDmWxwfws8mK399+8hcKSnrFssvKW
/1CvgF2aXbv2tOKX48jTWfXVlnk7LyFV2EZ2AcaGYgI7kxecP8Fx69DIi7N/N425PR3MmugSxZsh
Mx8NzPOY4V+yAG44mxcb8/cYUj2KilYNWVSQKfjxyIiGUa8BcvrGk/mfzV2j8A3iC+/xBG7wA3/A
S060v8086gtWlO+v/TCrNCOVxo9rBEHBMu2XhPknt2jSNWg9I6iE2a2x2ehpkulN1QM/MKE+VyAV
Ozqx+9+HsVsiz7AJcHKdBaKSE+RTJNOrM3HD4JoNqww3oeGFuajblIU78nUCrqMHfUpkeXDiHwwd
NW41tM5nPEibToiF1b6NobjkBNk1IlNMwduf7bf18MNM8vmE7rCQDBiqxID45SXwqgpV6pMEYAMs
7H9KKZvThMEWBJqra39eOAhN1ldt7OPMctNtbyi2PzGbu07sX24MknjDlLWajJ6yTUtbrJTdV4dy
2/E8Q7nIWQHAEh/pKe0E3eUNrjw40ZOUc2TUM4At3zbzkppK46nhN5tZIWxgb7pdBTRu72QPS6RA
m3AMI2sK0EHeD4uo4tXVJwFmsbbpsiTwJfmIKkMiVY8LO2MVVlC1ZjLa9VPU5EQaReTZkdKviRek
clrrrKpfO97QNPvdqQgvJYZRPuFgIQILsWnc8Y55YKz44r0e4sAgTbBb5jwGb1Qa0KYc3YHP4m9f
HCHbuyV9v3P1S4BAe8B7Ce+8IhmYJSydnTh/LGGFQdWBN3S0D+YWjNNG+D9eVlvXd4tEA/a7AMsz
GwbW2N7nqF0R3TMwpAPtJ/rBIcnm33t0DvGCJ2JqF6G2vbN5VnIRunorBtnw0axohiO3niDft07Q
zPvJCxDvmr/ZPqSB8XUroQD8fcOIQ8bc9ZXOcTMyn4Pai54ifJdJNJW/IHt9qkwE2VxMxBusiXuE
fZh6Y3LTTZrSXfEsw+R6UFQc15RIXa/4yPl1tPIKvTuk37Rkpv8nBcq2bQNhH/85hsZc9WItB1iZ
nCErcYtSEB7hFR2CONHLNLsiSsIs3fZJeyiynD0wDmfllnOzM5Ebh3SsT0KzC+8Xu+Qcf8y3P/j3
g+YriqWXF9LJEdt4QKyYbH5rdd4/PK7MWHD6zcuw3qhjumI1Qq+bhGGZsW76QqPXlxRSSsCfozmJ
A1oKhV7DtFI0tZcR/ZI9u9SNjKFAOPIgPCKuejymAq0rcxnHNo08Qdk4OvCXafTzYO1Nv56GuxDs
0RpAHxR/v5rJiXeXlrg6oU6Dg8k8ptKJS54p4K7fts0qlCCuZpk6XwUqkI4qg5wiZTS7nWkeDA2n
MlDNpez230ICzo2clnAP1koeIPW5NTazOfhl0Yy4lb9gNPyeikQwRAxpbXCYViJypNnuxO4ZCRRC
dunlpJw4xTxwaODJW+L6Fmpwo1cBu1AMEPxNMFY7EdPmGf7aQcbgf1nWH8i36/JbkdLb51vqcQ74
8JMowlU//+cspZ7HqfGfkQWTszMUWQhWLFTpOE7KqB4FhY2pTD0xVFIs8T9zW0U8S+SYsQfF2/6d
sAl0OPMxojUOwSXAeUH5kP1G8zCai31mDBGaRXetG6AlYAH5TKWWvgon6v+Cc+RCGBXUE5VUDUXo
lhiovC1O6caU2/YpQkP9HM9+ftSeihc9w1/AkVZ33DETuMtjW7NbXyrJcBPFz0Oy3X2+1/JyxlWw
gYJsuyUJQFU0o+eawrqrVBBlwmXJbLmWnUmooyj1pDypAeZCZ88VyIHoOXM/w2om9mOXJNiEPLRu
/CLU8gEkFvwLOobFfm3GqW9JNGizC7rCGiaQIEBF0A+Vi/EZFOEv3FgLlqzQoWa+N9C7VOIDAtax
67aWqk4uDVnX2V+WKuXV2oS4F7KWsWihevMlolMzxbhLXji/8XzTi624P+qJjMxQC+CQMvn9C4+Q
2egF72JFQHgQewVmOHtGn0bD42we/kNGZhTY7gHAzep5vQGndzW5STVwoq5al2OW4FJ85debeY5S
ouTeUv7mY2PQuqYd2xZ2wuaRhdLqZ7xXEBKcg4P4RiCPYAqVvAhpoPC06iDp7PwSzvSN+qKOyWlR
9dUwHZ03IYWLvNhnSEo977xTQd0fU+gB/SCIZa0d1tkdGUQCnMHTUL2xLGH4PIbkqKS88kRcW7qZ
B/VUkNqopdb3TuZ6SV5hszCeFLwmYBrU+pYxtuwIeEVOIXt1PhqNnFD+RMw1vTmbeSnb3sGX/go6
qxywx/Mi+7fvgFefVXFd7t4+QytLu2edjYxgyHTA0Fuloqqbfx+P9aLlONrmh5eptCkR3CKsJ4f1
gXkmw5O9AL4tkxcKqUtKkz5vm+9WUYPsC95khE/KHFov/dtCl44EMHMe69OjxCeMtovs3Sh2ZiWN
uHUhpw3ZxDATdIRg+THBQZuLFSzzS6munNGmBJ2fOJeB7nYhpzKEYoXrVDO1FGr/98RSapW43N/W
3jj0USLzW0skDKZt9PpUn6yy7JgmklxIH219/vMpa6HqjQZrSYJab5gBswkHXdzhFAJRCCxWSadI
9QmxRkt3gtg2c4xhCwfp4nj/RzSybL1z4CaD96OB6HmV/FE3GnrUdR+8hWPCeCinndbcB9XfrCFn
XEW+M3KOZIcyQm6HXq+jyZ1xNM34oJAynCIyH/ZB0SV3UySucRXCX6hCCOeRx3Asw7k3/1+mCXYD
N3n11myUH5R3OPuViWGJGY9JrexI/AyDrNT3uB6BmSn9qU36fMjjNcdgNiwB55DD616dDOHgR8AE
P/NzjaSw5jBq2/TD/VSMDD0B6SpB+AP8kpJ4vAcjW6yv7w25zPZpKI42u7R2evkorzOJe7M0DHhu
VEFTW2XFoQyGw4lSPOa5fygGIfgsdtKPCqiRyJN2iFRsxPzhJ8W4miSDIQ1xWkliD3Sb5+x+GQt/
dOLSvFbYYbukiwnz4xP2wHORvwxYW5m7Yp+6dJloVSl1hjKe5CaJBqRDa4Mf9ePvSwVzf7ZRoyoO
BgUxFCIxVomuWNrePxwcJEz7z0uEGMASxfc5jBioxChIDFbv0Z7gPOctLbmQAu2YaAuUlMc/rvaV
G37Rm+5jMtIdpf7HAMC+KnL0oYN7vXASSBCBPQjzBwBo8YBmXhvezDjjWc/l7LEetn+kbgmN4iTj
VYp/4YFmd8/A8SdFL7Fpp/Om/LmqY2dEX0AnAKkWHsMpM1UE0gwzPs+4XJpwqeEjsEu3ryY7I3TH
MjdLkOTsB3qts6nMvmsP917VWDlnfGFu5jhcRyAhJH/JV7R+TPx35+9WIuHTg3jj++4fX4px/7JF
Lx5PjLKFQKqb3nyaWmntShpIlHxd3XxHMeQwfLGuVqF8f+jhiJktRuWEtoev1ANYkwnl/wk9WDCc
eu5QkZqi2KbBtajJx4PYQ7tlPTzp2vYpDEoUbo1Az4bWw9O9A84UZk/jiURac0Vt6wNX3JMs5tpm
a66UKDUKVz4ymb3xSxDFkxGXhCR10MU2M54Ljr1amB9VIS6uOrOBxcplhLqVfvJDYNjzfvJQ5vXy
1NM++ZLSlJWPCMwoYIPR7baRhD3nyvi7QFYxOBBU8cwl3sqCr5PyQIww3QxqelYmhElsNBgoz+Ix
Cpqvr49ZmhWmooTuZFEfmIfdZ84MshiDbnw+NRfKuCdyyGgBBGT6UHYLXzxl969LQ8M9BV4nbnAe
/qO0FVVvNfEcRzW10/eJzOk/qCNOFQVmR2bjj528R9u7ZRNJiNL477b60lLpNCCvPISx+J4DfBZm
HzCaU5dB8x5Q5nvpPBQaoOBvQnt2HbSaHFCu6t3cgJSRmsxBsDooXnthpcmAAWvXvQZaesJuxUmN
BXIrGeMgJv/vnzI/u3W2msIG1MdihcTfNK5Hha06fnPrk2/qT+HrRl59eHHJzqfCRJK0MPivwilL
NsunS+QDluhy10kU4/RLyz3l8GJW3PZOYT8Z0DrwkhowxGLL+0yZIV/ZPSYMeC74knB19Neldsdf
G/K9qIRIcIx/xzMQRxPGx3GwmfBLhnF2yYb2QN3JU2Gm36lnjXUY69kpHH4at5gsJX1nwja+iZvQ
gpYbRCM03FO63Wt0YkVZhcAVX13Hr+r6R8TemjHOA84AKtONP0mkvrAmryB+TF/HLkhxat5wMGkg
215euc+6fFnrjIssVe6sLLtI54vbyRjWjyX6UPVrz/lCElZDGnhQiaYcVs1RWrVgBZYVacBakG8j
KDqxk1Pk71ISmyYixU0IBQhefn7uPTDbwBO3XvIkKd4x2n5nzyrGUBr5yC7GV7RVlZWw7s+qiSUa
tlWS+q8UxOkGRuPxvydLehTwM4YXdQ9Mml/Eki61x/cNa4UvDu5dAC4W2dmAnKlzqMMKbRgyukB7
C7GjIks/VhLF9jz0+oZfZJgh/36on25bGHbx6yCGle8o+pCeQOJ3ZNptE3hAraRbCzXZ6vroyDHj
yTljaYlzfyLSsmUY7FXjXNfoKEoyisklTZF4K/U6sgLWvqQIjkFSLA9tYuwo9i1MOG1XOQ1mkmqI
jF5jFGliT35uV5vzSlHMWRj8yVBve7K43VPUk8/PWAzIl4WkbO0RCDb5BjxBtZfVVvx7fTcrWBga
VAmy3/WApibcQELh2uO2Xn3HJ7TwCoW4517lNt9uU/2FLQ87bRFMxNMTqcu55qYCoHf07on3fPfv
oCMKMbkBVj4P9SAj4WDFjfE0YBR4V5kJmvb1ZVgQCIKWMnqMIIF1UlKUmcqUB0Yp8J2SIxmieiI4
DEsknLcset3ZIpdAB//vEjsXaDV4CVDngGaEXPL2EPp8L6KPVWR075/OWKLj4jXPYmjJFVVNQKSZ
2R4f4jXT5c6FGQ6kwapeDYtLnPVTbAJJGmufN0wEdNoNESl20xJexU2cYL5I+mBUMpDm6gULMz7Y
W2yi/OJBmIrsBrSps92V1SZiIRGLPeqZ3J1d0TCqr8RgLBQvkdpvT2zPQ78qPa0gy6oNkxIPxU5Q
wctduJL2FLGf6RWwOC8WaMewkMuJ5ic6cPzxIbVD+u6W8q0tCrho7sRAUJd19Kspz+ePTuvovxTj
/xIgwpYfvbQ8cPJV1zziJP39ZxFsnBIodnWF+eJ7dZh0YmAtAzRECZXFwwMNx6tmZfHnrfO2E10z
k5H6gragxHszDt53bFLoAza2UFn4cUSSm6gUrZ8m9Tp6I1IxUzjJK/K93c1n/yKfVzRkMVwOUSIB
GNHw5M9RB+bhvy69F3mf35qk6QPzyyOLxOIVreQltUY3ZQiEVbRFkB0Wjfd4m9l++OjZ07KLOGRz
EBqGGTCjJZYK4IVFbKGHV10Nn1fXfOvDWFVeCjPUMONZp5wCb1HFa2BJ2Y8o34S+pe0iST6qLYj+
RrWGWwdJ+PADW6OAdokWFRD8w4k73vuyoZ1yAhI4z1C9uaYUBwSC7lUXsYMVRgC8R7TTET5GVwrL
ODLDtLchRehGUU5Ba4/TG9rR1zrQ7ZqlN92h5DdwMU8L6fz8KhB2z28QB1snFqjfpPgYnoEs8U6d
G98KX0DaMNYK/8gYIZ6q3ri2DbKFgJILjB/TNi6J6lV9J/m+5aaRjSrNWv1YcexnLc2so5hfQrCg
a6Rf82ulJDD/zUcPFgw2yOrFlak6/XjCnBIHs6yP4EQ2qWmFuLPqfR13x/9ypHeEmo/dN3gsN7lC
Uzssm2ls3wqAtzXPbYcAJvgN+Fpm9e6mAFVLJTH5K3R8l9J48F2EMDubSpRC1/mc0HDVDKu6w1jW
RYM2DFHRnRqNx8wLVMs1VUflyV/p5WcTrOK9GZglR5gpth9vA7ysfYjFZaaZuXzc6/BHYqbc1mi/
Cyp3tDL/sWShdICSjbh+j3Zvw7/eJFUnGJCE7HD5RLz+Ya/Y6SxqbjEuvknAjs1xqkLEKPUuDsnJ
KRL8+Wof6boYqQShpw0XU2G3f4bT/nyt+mGM2oNzdaNFyhhmUZB95m4gU5OKRh5ANeVzpXPwL9EI
1XiLCHYkbBMo84YuIYedxPGM/EwuAkun1BOERq4SG2TnvSHE1aF+v69wPNrddQG5wGJQSQDhfThY
SzkN5LYuMxGQE31AXntf0aeyrZhKAQZ33rJxsYERvgG5G3iviU2fin8cDTkcRFgXdRdY1/arSwAB
fkU+gBsBRHDGdzBsQz8PGzxZuVZmEyxLMl9b51bf6QbKXUEoH2k/erxTAhKOuzKY5Xc+Rq+rc47l
3/hzgAoshXhQ0ZN9pXC9loUqrpnnQBJzNrOyhb4/yfi2w71fYHieeYPtW7zo/kzH2gKWNNHRUWiA
p02cDPz8+qfvR3a7pauORjtaQCfAub6FsjuAk8WuaeBBoYimJ4G4siMBK/to6i+z8z3G9A3zEuHz
COoCDZb/auI71mw6KubxzMB8Ki0GYN7B98cEG0s+xEfDtPB/0BktdTdSoQYzkwnrKLS3aRilp88+
A/RMfmoW+UYw+8ouWHoDxMTpWNACknISAQwsPk6/pOGv2cBP3/iESDWYGfMArrt5mEE1UEyzNZdM
dCX+cp2AYaocKZdwNwNuceWbyNGoc1OEZQTR72hcWnikXHPcLEYLbUlVTClqMwkfxFJ9BWTI/Lc8
211wDbRQN09Y2VxiN0CajbfiVVRYSmBw+1Nuv7DTuiDPdN0rkr9P2HVOAlzG5Er/Lbelyzti88kj
0QNrwoQV9xSoPM736yt70HFub4hGxBx3K0u4q8bg5gIdO4tekp7romzoVwQM4etMDuPRrHko+JWy
2+jFvwonAolb2HGVZCuSCtXUw9Ob+H3D33tCJ7GoO7E7ytXYTABNLYlHOPEYmk78QQ+ME2Z0rAZu
qdvO1vtRUQyFMcxEyz0+12f+CtC8fVaQ5smNKaLTrj+8ixATicz7T9eLGuQ/aK5VDTo78XFqndwJ
1iWPWlvqVXghkOWaOk4Q3KKo/cyjiNd7IFywdwVh2v0sd3Nackm6+UqC+lkfRDdW0hUKgLR20ajC
b8wTFpUvKrLMFMV79BptxhFDD924+erPrkfRW3B/G2SyUoHR3oovhGCBiJXP4EHxGn4/hOoMhNOh
xkssrngIMPOJwBYVw2pieAv6S7wYn7EgvbpoAg75qb8fDGzKn4YF+utUE/63RVWf7HjaFXCgtwtq
0c1k2T/DWbVpFGIt5PZzJgc4O2Tz/p+SCbpZQtfCML5PmtVW4echTQ9/I2xVyhnQNGEZe1GWYGqr
6PPHzjJqd9gbc8pXIJnaXaCzi8qFXtCstjbnp9y1BEyblxxXEtIcSXRh7pG+aJQXgO+G6pH3jZBx
vEqBprhvdZT9fpmKmMnBwxDZqHocPFscQ/NRNNoGKfZNHztkm0f5+qdSMbjc1v7bjvEcU0jMYaQs
Q90WvxRFa+b+dm1ekbBhsae8CQ+DhjSzwy/EY/T4w41damHCNhKW6pZVNrkvqTMbm7tx0u+tODAc
8Ad5ne63yJ8RBvvcb5U8x1Ymvs+76+CgvgpCshfxQkwKiRuvKxMEBPHMspxrQL3IHZqVUg5s+f0q
4YGYb2f3H9RwwkrFb5cxj6qowYWXdah+HNAFFY3ZYO+Vbd8A96oA1Foc41Ea0uELReiCgpxqcvye
2WYWo7IQ1s44c+IdtyzdkUO1XdD7aoKGD8iMuW2jaljvD4ypZItEkR3FXmGQzVA1NjwX9VRP+i3n
S7kS6BF9N63QxVML81syK6pUuRv/OVepSP/k8CTAMqFwAxAJO4N49QLJqayVOtJ5E8jJbBbLOVGm
aJu+j3ywi1NJT41Njh3AbfOwp/FWmOpizqT16WYHyQuTetiu8kC/TPQYDt99/Mr98UZENjLvkiK6
mwsNGuL7PKsRCbndJcSTHBl7tDg0B/mwq/sZeLG66EQApXwfQYH3BjlXW1tEy/trX2PsGTtJpzCw
fYg0zF9ZvV6qDJBbiYJD3jK1EgEzwhu7d7USP2SoTB/PrbkIeeKgTPOjHu7NHBZuaenq03UhnkTO
RB/kr75/cO2UEkXfwA9rx0wPfwwnOZJwx9rUC+qL8ShsIGDfKIo8SbT7EbfJyPmHCBZlWi8wViTR
afuOoP6IzdJGf3mbNUmcLWLbU5jOA5Ac4TZKRmYIOPo/1CJptxjDUaRwX/Jyvf4//BD2MhSabUQw
xvHKOuTQGgRYeMDx5TKxQZVT/0vvs8BmL+H+PM8vT5n0RD2NCFQccJCreGBw+6nCiR0VstioLPcy
Gi0KjY/mNTSJ/TMW/Q/txteMrRpKaLX1/BVghq6b9Mbhd1kC436Dlf6m7wawpdhmIKgpjg5kNQck
0986SmjFxygLRe26l2HnA1ha9JtR530z4q4WrCzIlm0FOVmlW0/plxpMdFui1MjtxZ9uOOI1Uipt
avBW153tFhWfnPguprDfALuJKd554OloXiGBnnPKwt84Nm+lHP/GjkvB9mh1GTfgeqrtr72YKRVZ
4nsaxyc+pIFR7JJp1XWn2vLQM9A3AFfpVQB8+/1Z/iiDW8WRk9nnj6x1zdDJYyTxuQMpZYlDLp+L
afL9nkK2qCaY1EfXw9Vv09jiOBgcjhW7z41qQWE1S1caR0+9fe9lDE+gTgnobvSyw4o5ievlDKyN
NyLhOx3r7WYOF/5mjerAwFRevP/2S3Ej+1CBR+2/wpa/gqV4LS7uLnBwVVma60gNgaEWJeD4/U9n
mLmxikyIsMU1RXX9ga4kayGUR0Rl+9saRTXlUy3vyszbbcpvfppzf1fh49EF/XyhFYzhYgWYGcBg
a2YtkmWwbLdDum0DzLbeYuAZH3fcrbjh53+4fvTWoA91ZOBCXeo1NnJVqJS3kExWzXN84Lyg5AXZ
fLwEZ3+T1NnVU1qV5mvS6agS4cVWiZxMhNfA9zzpQ1JN6soBEsrFxR0canBpoTuEeccz1TyRVVmc
xeOTDNpWA6UB0Rsa68qKQtlP43fiToSVkW1AmGPXrovaMRP/NrEq0WjsB+6prvynEPJiLySOWN9c
GU8xUR19eprmiT5P99LMse7Xko34aBEEeQ4RB5fvq2+gaFKZ5YQPpazJwkI2KE+t9qaf8pjPXh4C
UV7Xpcd6EZ21zGXm8sakbLHpTO4ry7FHF/AqHbucwQ/0TnFL4ySZ4Bsd1lvmNWm8ZUcZV2nZTBFn
EnofkJa2ONWCPrdAfvGqN9FNHDs450DvmZ/gH6tcLKGepweRFwPt4F1QU5yp1p0+yED2N5XVAK+0
egD3urSSpB7N/BZxSdn57e6DBny/rmHzTCmk0vOceQ68EGuG0Jyq0qD6EJia6wcw8K53HW4TESzA
D34o8TS/lf3A//q1qoaRq8d6A8C9eZaVs7CjKxJ6FPp889zlfgsTYUXh1YsbsukiX2NODmt7YWqv
QP5sBfvUk+rKHeS9lpQ/YdZ+WMG3iuaeuUIUteemrsEpczMchum/yHJgfiBx8eQbLOhNjILtTuxL
DF7gE//UquXocjH8olOYV7u0Fuw8zteSpkVWd8AVh4LrBWn1iN03cd+8fJKPi8J77AiLsRIBFFjO
ctp1BEbzm2lzJz8/ttrsH5siUJDcF2eXAoYdgoPyDyB6i6A60HZJ2yjQy75TUGVOAF5u7G7T7/Vv
2ouAOEUzD/MG5NoLXjMCBjgOUpjOgulx4WkFIfrHDSGfwv7ODk5kEZsCp+Yroav+1ZmLq8PpFvSv
dzsuR+N6kVTSSv4yE8Tm+/VhOIiWrCvsdSeFr3salFEccuv3buYXmxoP3uSGLPamUxQqQdtTd57S
yBufPuZGAjFhSjTZlXdSUz9z0wb8aErUnrojqHGexRulKrMgWVQs9S/snMVigjNHeaUpEnOEW0jb
SgdjfSwbbw6i/6SQ0goKG/fWlMcj+87fOWhwDQINbdkcydf+kB1jPf4No3gm+FdBM36OX2YnBPPX
oL2G1gbM5ujfnzxwX4CcXTwiNUUdr2Kt6XAS4teQgmD1/Ytb0A/WFynUXljf5M3yCAX5HjoY0cRg
Q7lpu+BLQ4z2JvHhIqPLj43MwIC1vkPxN9sV9yQaKj5wG6tNQcBGww8pPTYyBirX0G0vQa41ZtoO
DD+3uoFrD6aTg5qHNQb+YFSf7glEMi8jWL69LXnHlQi6scKJ6u5uQdsadQ33bC8HrbG+UrcSpLdw
+Mpv0uxKah8gONlDFEdL2eaontRLl306yYOcViMd7ZXLx+ceg/G45dcikagfn6cqscmEF68BK+VJ
DyLUCW7gNrbd7UZTKykUR5O+/VYs3loVkyOSZdGk/H9PqP5pWnyaxwLvRmTe55Ewu6D4MlVg8+uy
sFNaYCSubQ4Po1rs4mo/IskLE3U934fGbpbVkR34VLvlc2B6s72mjvELXhli+FD060o8HyJIHX1A
kZDNjNc8pan3fIOWnBO9Lu/Qflq0/5lmLEM5LEzgJE0jnPBoED0IxHZe6iG60o296AFttwrRFE1I
KdG8svfF1CRjknVD8ZbyaL8XGC0s/llFRt5wN/ostow/2hTSN/3eRZ3mNOOBc/Yb8jvqma1tZS+p
XbQMl/Fp82zOK46uXsp48IrQO4Lidu5svmqweItBEQXvUdWkVBoU5AzRoD021qIes5O3rvNv/kVr
W1YGg5THohQWtUFgP54Qmiwe6a2urqeXVBmYS8iaDh6jxwsVkjR7Dl4jdk5D/UwcmojDenfxJMJn
D7HFqmqb4gm4mDrHrUoJIn/pMoeI+pdk0jo14wIiiOFeTavME0GPgovxf7MFvXya5JH2Cy2D5PXI
aIThacjwXF+K8/NkxHqldrucCiK7+2DQ57+uSu27Fkp2KAEPtf69KKjR7GUJDvb9Aho76LCPORBM
WY0SdD0+Q7aknVmykijzVPQhNAVwrjZrwNWVGaKduE+Vv+ParKY+RJy8WzdDOf58QPwI47Hhv4o9
MMLhpG4RCAUJ8Lcckq3kN55z6/gxpLbZt/CPJ+/cL+nYhTf1ITjJ4hoI+DVXTBj8G4BAVvdCpUA7
PJQyaMvxcE8yfnnb71cDaJMiSZ1akW7wQy+l78hVS+jxdir5fPliTMwaXOGz2xHr9dS7sPjAG/JS
ug5CQWEMN9MidryweWmQqmhhh1xyZDDXc85GS2uNjiXVPNm++X29yoIDu+esrto0ubEYTXvkqerg
VBObHeJTE7OL1V0vybWnQRap7z9J3CbOpKpFLfd4csaBHQvbledXEX/oO2NRDFPH81b+TY67UIRK
gLTxQeSi1IzNcqMfbMUg9BQHN/HXvMD97TYt+HheTd54vBv6GV8vnAcYkfW0mVmgta1QkXQdqP5r
5PJEb4/x9LEP7GNPUjfJoQeJhbJ6CCoZ/qwr5F8j1wTSWntjfBGpGS2tF8LxqT58jhTbsMmiMY/J
8sstqrrRsHiIp7W9Sr4pBt1IwzOzaS1iuhnOVN9HNX3ojxs6bXF18Qi9WAwp1oeWdXu/qqzeYf2Z
gUD8cLGNdrYwVGeNoOViVHWJ7Fo5vFVOCUUfxEjB9LxIIgCHJTBH4xaVUkNZuv8swsc0QR9CG4aG
quJxfc6//HsCB5EFHk6JVEruiL1FREWBlX+d+CKJe+FILpKDKU8YAuq4SbvlbfEFfqMOzHtyxxAX
NC2AVL6VKv4QHI10OJUJup9p8HZypaQdc0Twu05Jk7ufpKnunYaEhl3KiXkTi64I6THB8mJjAdUo
/O2AzAoGIRJhzFLuYlT8M8+UoSb4cqt8VxNVauVdtoTHdKNp3UW2NjgyF1/QpOBn5aEfhKxboHKK
aI/i87SUhtrKNX9siOVcGfnYJaNtmynrKqpnY+de0Q7PzJyLycL7R1Gk+SY/RX2drn+9ffnu6myB
n0wkNz8SRbXdSIcP7zuMyPZ3j/WJ2y79IVflqLa9vVEYulvWYH8K6FHM6abcUrXZhdtrZNti4lkU
2TtsudRo2rLyAnnk0rXtyIpHGi7qCNfz6q/z1NKQkMrLLM/SEk/zppZ9jNfBUHS5ERKP2JFBsrE+
WQM8+ACItIUUilpL3L2gWVPzrQslzYFyLF8KdOHu2ytx+zhsDydGNU4JbAJh9E7TVOnGTZ88yq2j
zG/AgJ0sB13uD7XQ3JZEnIE6NMU9i77TWKZEhgBo4t0Qg46HmEvjusx9J5HixYVBKWxYIhCc3lW/
MLfgZexVkf4Os3HepKZP8FrNLKg4mbD/gH0Nfudt7SKZxLaWg8cBTvqC7OHZZqTx+tlTSE+zq9ro
JCvxu6q4bjZnRxXlBMpooTcJMNAXiQiq2hxDDjuwPqJ08xcfBJCekdKjTGPfyDwZXPlW2EgBW7Ro
hG5qQeBKFFtHuJrc+64MFesGJvxF+6STcr7c9lrTfP8jjC0gZEy8dRZPL5QR8lFITAeKNgUrXfT7
zky5MlsdVzzX5prqwPhJF194QZnqIyF+nuyANmDJZHrhRLXckg2o1/LVNLv0CZ/loMSlqF48Xr8S
CaBhpHuixrXD3EWr5nlfTWCTXXPE5uPHZ0yydLRs069l/gL/eLygG6UK0GTqhbhP7MVJyGLGlcVk
k3qUdoeQqN6Il0+FkKYrEgFQgYzcwItAt0SRECk2YwyW6QHswMe5hm4b8wXEf0qP24EN+bcZuSZ4
a6OFMQva/Wt9wum0wv0IJGwuBcvIIaq3QwOVPZNFoPw+x78R2/ZmGev00reVoh/ZgR1wIaO9c7xX
q9gjuQx+ojoyiCsLBIeIiTkwuWeRiMpDJLCEXftpy/yPnNAcaDHtR+Q1VDn/RM2nxP8q60Eqz3Wh
ZkyZGV8V3lL2+/8rLyektiGqwSKq3cWDTKEg6RVV2LwAYngi0GPhcI8Bz/ZLlt2W+zEaQfBOPC7o
fuKDkP04C1xwOzaNNm+stfGfnhlk7PgVggYnQlhzNB1/inpf4ZRaK1vECWsAfJqeQiUVOyFkG6u1
u6dVglPT8MW0jR7w0YLF2n4x93bavppIgnE8a5TSrUs6Q/pZO9QZBZ4GHVN8257R1f0VNBN+k9Rf
EJqXMcqqSJ2CI7l8I54lryO8z+KuObABx0kl4dQMVBfeFqBp6lHpUdbJl+z2sMhp1eo1kwbqzuAh
jc/MiTwGvlwO8foBX79P/uGYcGCRPd7tnYu7gqmnz1eTW4C1jOuH5gx/MOghLKRM9UkgVptPz5Mk
i8T7CQNZcSNw24C+duXFR0e4R+nXvHtQxduPRK+w2O00rnWbiyfnOhh7RDXAVnPAUSjV+Oj6EQtl
bizJJMXxumVl3+l6AEh4NIXHXnlc4WMZT4LH6vZnC9r9n+VV+juGXbHZeNSx325eEdNtDodiAWg0
w5gYth2IbZqNQBfCpBrzXkEGdYsSVStYBGn73Bkgb0uPsaM15hoh319PyAb6g9EhFREMC7VMptLG
wMB9dUzufu6VDPNrSQqZgvt0tq5kks4iA8iymaBkEph0uG+cXCOCZ0meMfT0LLb1xL+ttzx/4Y9K
NibYd2n6U+5HMwpYYGdueGZnKCaCkxzCyNQXLIArI0v4GfzdReKXiOn02B5SE9VytH9M3w1M9VK3
LT+3FS+QnLBDlxsowOJ+Zk3LP6wRSvF4EhaJhd4J517zOAxpZjSP0SPgfo41Wl+wOz0JgaQ9orby
9qASqyfo/2oFSWeUbjXA9ZIarCoNBBqZzWUvgCayywcnJ/ejfvot9AJocfps+I4yTBfWP+WLazSO
P1KBYsSKJ0MsFgS/zXU1nHWGc4DQdFphI/fH/c+RYTi6ZHXEDhXhDm77lioJkh0lATI5wkvYjeq8
cZjYsbCigZwszsg2wxRNDmPU+jOqiGwU1WwQ45f9P95lpoFuRdk628QFDfaYky/Jv7avl/I16k+I
V07lyy8v6qhfC9UkL/R9MftYkGUe7aNGoszrMIBuh0OEGxPneTYiOzMSp8JKTnNVNhfSR84L8TYU
oK8dWETaVHSXRaFcotuN5zuLqUD9WegrCMIfYzClZP/sW5DYgR6On6NdsFYYpqoolpiTSuDoRTym
k8OL7h01yJWyhnzlFMzQwCuIDbAqaDFvKumG3kaMAMcU9+romGDkB0+sl+UULn0uB+yWrBrRNgHP
ASLy7MZK7nbei3AQGgyj0h3GtBkGgPweQp9WmNfvP3TkRH/sW4MgfgTQweff/vnsed2oHQ+seZPR
GvUiHrQSv4wHQ1tW19E14jpww7cKLFVzPL2BtXn1OxUaRY2Z/PkabntSVkTl3tvin+PT8+f6pXcr
qSaqNOSodegcg3CcsyMDAGasz6h3rZ5dl4ZX+I7fcAdL/WrHKmd4QXkYOPtMPNiZYjfiqHNTeVxf
kiniXVag9NxATWSnJIK5ymaozk4owSNzf8xjqJQLO0+A8bdTpAChsGoQspe28HnKG5zMZQHHoGRW
joVgKNfHIJd3YBJuPNOUOT7Yv9l43T8ScWyln6GswC9XjjvO53XcdV1jzDbNB0rm9w7CkpZHdTt4
rW/i6KNTbUnmGk3IWjAq1tYT8KpVJ45JyTKrZhhLpClGa+Kc4XM9ji+dMdwacri4xda76iOxgTS/
MrF3WLjX+jry8f1dUfN2zTYNMhpLxYbubhJcJdZhywU1VyiGyeD12fYz5ENTxBHh2gllUszmrTI4
99fsQT7Nd3K48AD1MvGEhM23oTnGAk9UgbAOg6SVECtGE9ZQKI3MhdsWhBwh3I5wGu+so9ukuEuJ
Ui+KQX/IaA6ePOeBPQQwXgVFtp8j31pLyneq7DcDNj8qM2ddFQLKxn08qPJWkloULIL1CpjfI1dT
+MWK3PgTmSD30LlaFwCINq/W5jAYQPIemyuaALl14o0UF+xLOL3ogEIzevXcZTp5NuoZ3bxKx7cn
6MAxShcYVMSsZScIrFOul4gjBRyEElz2CiEkvm7ydtOdIaFucDI7mkQtwC9dkE7yGGQX+etGO8Wb
1cqYhc1CEf8tERKqAcI+ZYzjB2eTK2SEV48oZEcoE4phDwyJty0ny5JsEvqqGKyFqCujOmjWl2DJ
lIbyD4f+13Y9fhBnxfPm5cHbkSE2OsdXntGEJO+3X/dwPkkqzanIg3MbxUos9z5iy13uxmjAsQgZ
Gz5Ymd4dp22Cl2Mu8qQdbTBHsyShQXwB+KevGoFNgJVZ3nrXKXilzHA0qHha0HyYEzb2a2hqsB1M
PUzIdqB0/dPQDnwKXqdmxdpULZqSpK73AQE6Fd/UQC9Rc1fV4XY2IVJGSR9B6ZurNcJjSAzIggH9
rwPUfRxoHqbI4XxO3JkTk4HB7sVVTNclgTpRHbgxTofMlHeA54Y7LM6pAHZZmSIptvh8mqihqT19
J1s+5198lNCSOxG2KTALizrdDaNfrqgYPlBlo+cPyS4Zvi/0g3n9zLkpzkJpKz02BjR/z5D2fI2g
GGFPsSit+aOyDwXsFwH2E7kVbbhitv0YhZh8W5ph09vE75BKyH5/wIkxY+lDz7uZySFMKlyrejNu
p1EPgyXivPglEtbmIFckSIDy0Ui7I3ehK9w4/gzDEN4q8rAY6yqDZI9xWsZOnlAzXX2vuxIxmt8R
rhs8ARjmU9kTa4tnHcmhTlYYXxKJ/uk6LMbhaePtKYSL1rQ0DCfVleQ6QVhSl0vLN1m3BtaLUfmx
2Mi+By9Ogbz39EQ2lSVOKcW71BytvF6vFnKpUzQNF2T94z5As51vdP8gbYNB1ghwGSlo42yHw/OT
LDVWxwQpwcVVqV26eoZga97H/u8StJfPE9qmBWtYIMYu4VScWlCwhxg5X9VUM0HigRmh0vMOF8mj
Okc5ipOxstZ8FS82HOCgXXTXFb3tw0KDoTAWjQzE1tdGYmCtsYHe0d/pVUy4sr5srV3rnb1MznD4
klln56tsBMA7ta1AbnTD6zfbRFd7NA/vGVwc1iNdhbdeKbO9RoXJu5BXxyESgNiEY5uBUs3ALIV4
gSm8aUaBw28WVbOJ3V5ZuUnWb3ST4HI0lhBD8Ylqo5VAdNofd3AyCQcC8po5OHaacO856WKM/VcM
xkR0gbuI8LX0kRvJ9KVC/QNAaWZLrGOvLjbUomYJrk1qlEJCr7pEFoZ+/AHUJy1NLP23gvVTyuqm
WXBI0gFSb9ic/9GjH/+ICtDN21qWt29dR7qKnq6040/1mxHja+fqQrBZ0x4FumTvDOEprqNWup24
ytHiWv0qD25kMV3BZ62bDCdoTUCj8mVOVr24QhXo3HWyAe5RHKFFfIJ8CvNXejcILOk/Y0L+wqP9
g4DtgfXxcFnmkNYfyvJYlyDm3EzkSY1ctQFYvyINytaC3INWOYUMfmarmX2ZmYURMNVq9jFDP9nq
D7E7UYohSyYq4Nk971UIsJnEZ+ByfeNfpwCbVxj73U6VHRuz0jFczXpmfxKpQ1KTWj75ymE1jRIJ
di+UXrc94x2tDgK41moqqKqtnXtcQKDQsHVI3FY7zSBpV6BepN0CKzoRkojo2PG2itHZ63vYjI6L
q9yjHjzOgfX0z3RwY4XUeq8uMebI2DfPy+W1yrRlA18/CPRexKhIYBaZtBpqOhp/ZxAjjsrZOy0L
IRyHOgTc1OOez3AzVSBMPsCrmYybu4F4bW+aYE7H3Sm/T5UwddQyghdOaTrYM17KhxarEwyuER+L
H/eSGPhCx7g6gSjyPetfi31iP1ecYYQwTy3BbznRrd1Xpc5JVWxzUeLHQE9kN4P5M4kE+Y0HP8hj
YS4Jv752X41ANgPTgbBkqfIz24MizuxDRrVFKyWhNjH3hkrERMRZbUz2YyEL+YRfjDdy24B7a5IL
tM19DOp9XfHTSIOy9DkYB9uoyF9wBXEg8PL8HzSFUrUTUo7tWLdFZQ2y1DI8XArLIxnD3Pchr6tV
qxFkl4/QjzPhhYlMAnloDwhZ7L7qhnE6GHF6iM1qH982OkF2ki2zG+dkfyaBMgEFDA8yuuJvroKV
+7bXM6mBSxu/qICUmY37WzF1B1kZF0a56crG2t2y4J1y6XMo1f/wlTmkcU2/1BtYed22I8VMMiI5
RA9l6mUp7BATzf+b87fgV8lBUXgAUgIyH4UJAZ02XFTA208Yevmxa3SqlGS5SOW6xiET66nRPpUW
MHnbDNjXYPJkUrcQ/Xt+2m9mHUSXes4yDzmtBJUsnj4/Hbw51Zch/SR+ExTOWX3mOxhl2QrzQX7j
mySIApi7iD/6fqQsWBqI7Z2dL/gJchdGTF9QubL8k2fBW/FngZt+OOrr7ljuQH9IWKVieDG5tRuQ
0TIpXtMDyPQm9k51a+68Js6HyVBmZUH4A1OPaV4+GEqYK2dI3FhVXGNPMPfoYf3h+ZxPEucvYfU5
FFwlUdu++KVVPqLeMiirMhHcDKjt6dSLHGmaNCnoepno0Gq0wQePIddLpQJoywqXd4oxj+xFL4xg
TCmxpDRt6csmcPULBh7kfoyHXxu9aMw1sqhAJYptnmr2AyqyD3ByjmofTY/qr4rE8aN82au2BH+b
e6LlJiJiWOW/RFlQ3qiM/ynzEdDTxHpieVl++lEd05uExdVJvs1gPt/qvvMHnRq9BkLAo8uDfS7k
D1sXeYJ7toiGkaIP1X7NUUeG4Jquq0olwBvn0SsyYkKG1b90KeJF07BxRP7+Y8VasOOVnGyVXheu
WAZkQJWhEfJAXUMl0999UN+IRAs5keZZDyZkFn6aADkcbedm2qA59cl5PM1HGqPxVTiSwXcmXM3P
ZK8YgadqYK0tPhV5sbIlRva4b65QEcDSXXcEhrmkN3ZqSm6S2Vi6KMWplIV418A5ilN8sgqihzWb
zEjIbYaqw9JkXRnDv49g4RinKFxX87la4zspLn9c+Vh7gSC5m99YLXpgDUQ50FrkTd38WQoLYRwN
YTmgzNYVzjhPBQOrKcYDqeT5GHY3LZjO2+LxKCnQM/YMOyu4gsKyfsvY6yUyKOaCR0X0aUWsn9ov
ecqBFzPxq1BkLuGtY/MA+qS3TGzPEoHcZ1FR3L0It9nq/Gd+0kvff94s1C98S/4zrggUzte13lP/
qAVWQZ1n6N3nje1Y8j9MLqgZWP/xafFiBSSWHeXkgZIzD3oOvUd+BUTOSOtu0vUzY/t2ZAbzlatq
mZupi3L9HTvtJQ1TQspXQRLg43PZW/GMa35mJRCLqDOB8TMpWqrdch8XgwZNcDsoAeZoJVmV1PHt
CiYkT5PzK2ULMqgxYsityXFLfu7Lgfp98qem81r3p6fH27cDMn8pBF4DXRRmH73mxue5SyWSz7L0
bkJqcviixiBiHUY8UnrYDz9L0lvNSZOm8I1ku+D3L0hGVuTWZGEN+0r9FYM9vZNzJgintaU8VG7D
2mBDV/xRPLZZzkrl94GZMhQUcyAz1aOuIrBdh07BlZ+SGxQyyu2SIzLhWiQSO0Ts1rs8p97/AMwn
Ltvd4XCwCbGxrHFk6XPAoKCmhxns3BGgwXp7CFkOEvnvHkGM29x+yyrXf9GRiJ4UIaRDTFfj9oa+
kLt9+BdUfbsNY2Bl7s2N7c9IgekYhvJhkS0tw2u2beUBJmvmf27INe3wdVUBtt5AFP+gpPb28fAg
iJ+v5ZOSkg7A3OXYljamUJYqONjC8Y0bN8r/K+bcN1a5l5sbOABJ5D+3ApQWlU5CglnhpxBOV5ZX
39bNd2RNclhatBOLBoPLM48tIW3tA8rLkspchT/C+G5pNDIZErkoUBMb9X7l8/JH2N0e8hmeMgK/
LTJTgmLCI6YVWkc2vd27r0H5HGUS4ICY7310c8O/GVFpmtKRjFxFea4b2me1i4/beSsnK2UfoxJL
aJg6X/z4AKIZD5vVpBJM0duOnmOdhA9I4d4KqYjyirR1/hs8nhcb8nmNjYWNIQm3J2IBmVdhDfiG
gnFGXCSmS1rNUmNn14g8vW4M3tjQclE2+tB8j/FJkh9Q7R+J5DwnoP4p8gGtJnjcfK8ntFMiESx8
dgAjX/Xe+15j1cDBtlRVhhKltPEpVU8dDLkAVs0kIReX9nuGpBU3AidrC6acdzM6sD3OU8PJlFhM
ndH7L1/0NLy9IkaSd1Uv+c11MAMR7gp5VEGB0CBDKXGzIavg6uY8YNJY0Thvy00pLRI1L76V6b7Y
yASsZWsj4JclJoCtn3+jnuRYSaMWB7N4UYbCwj+Lcj9uIuFc+tuN+329Nndor+SmFIUQa3ZuB/K/
9Zyhi60FeU8e2xFx1xwGsOoRIEyJw8IgxdXue+AZgw/nDVuzO+Q8hu28eG6q3Sb+uuK1StyknHUq
Fc6TyFyt9wU0kZea5mu91D3+kk/5Y9OIu3WeOag3eBsDL3BaGbAPLkOSL+wsP4XzgbscZhI3GKtB
P/iYJ+y75xJGHmpu5kQDuysyyTRHe1BbtcPZI3ZE8NIFdwaU+FnnfLrCv2grKvrt7OB9myFnZmFg
E6ebcH8GUbkqbvJWaLsScK6rQcS+32FeE9Ec8kjOH56YKJuHVR7fwGJc3wJEXZ7k7ouxDp62RpB6
zZCGFMuh9vP/F+pRaPmvvgnCU+XxYiwj098Xu5R1GZ1RJsiWjD4j4k1AruQ1lsYsaIO4BpMcVeiQ
5uST7iCfjxJ56R7Uc/C5qzmN86o2Edl7G5l2rel7r9H4QYRNNwY/bnNu8LsaiZ2M7xj7uiKsWEb+
65D/FPgNEnW66rp3sSAgBargeX0d2O/+HYuCf0+D50mQPPf6Ghq/IwCf6aPu5XRB40ZExhDF/WRT
7mVgZU/9H7SL7Uo2R7yZ1g7VnsyJpAyc3KttOeGM1tm/LPwEVjPcnh0ulRG8AbrbfFNC4ITWqnk4
gN1GAsX00t9k2PeasuDyMkVNZSAUgz6cRtBPWCGNcgdYGsxhP1bUt7tVBzt+8aO1M00OzRVvb3Vi
2CVTLii1i97S7Wnv1j1pebCLX1LeXS8JeMKtuDiIS3L8NQDmw13YbBGgpTatQFmH3nOp5/Bf/kGX
uAwb0kLMRo3x/Mi0y1dqpwUB0sK7LOblkjjbkNCZzn0BzPTqA4h4rzWA8QZiqW6hMblswN1H4Ljf
OVFt0HBH7sYfnAdNw3RRYD/2QgeQPRhHNXhXZgvpIQlw6kjeaZkx99E8qJdBn9iyMp0Z7/T+vAWY
bZYFKhYL5zJNJFYHwjaS+ImY5tH2QoBlfZRBSRQtnKj3RsV9JZr9qKhRDRH469OMo/AgWRlmu2M3
7Jps9jhf1MOBh8fV1erJQ95k66HDx4xG25O1FVf2oGXI8RwhDPFmd5/Ed1feUfKdZK8c5Ru/yXIP
2NHVst+bdsv/vObTnWxmhgl11T4BWJHdoTLo3o2C8BYFW/BsltXE4R1EcpDmUCGl9lhtZBZGN/uw
YYfe4/Lra7E8xp9389FkFb86LEkpdJAN8hmkZS5pIc1wpu5fWfT5F9Q1axWlmnhPUVryofKdQGA2
1GWoo4T+Ojw7joFBPFwVTFI5YKH+rC0URKHmQblufODZiTAYjj/h7v0+UmFGEDRWwv1f/wFWB+05
ab4r7TBpGiwdYnkHGFfudUcTrGaXP+IfobnlkqN6ljE6S0AkQ+9lI0gu0dzCimnx3FcDom23bqCf
vmcQyUn48d0XYHQfjjqFzXd6WxrZE36H16ZsGmPhwgSdb3KlO13kbQ/+QG+8eZEoJidNja9bsX7F
L9k7RPj3gUy4aswvySffq5mZi6agyZIRcqWZa/s1wXwfPjGyEDlQGVknJYsc1MGx7Qq0nK2TpqQr
jhVqFnN/eSSv+lwcvD70Yvq0UlCMeQPnwAi/EHchm0vYGwCHhSrj5gnHQhZuru7gh0kMLLqo4+V1
NEyzXy6UakQgft+I4gaxTQQPkbLLSWCESsDNfZk6IQ8gTiDptKCKwlFUM3Us1knlJs+hsu9dyvMB
Vw2ltZVZGT8WNSa6xZ2eW1t5dm00zO7frbToHwnou2gQuYHR/vMpiNsc4X+ojAq75/cITM5mEC/B
P/KDvzNzu4O/GG0cMGzKPitr11lIFPEV7iB0UoCB8BPJ2pL+mWaKjN4Sms3i0hmjmvXJonVPYW/W
MncBNbEtktYKeSAtbIvX5gkwTd2OKUvVfegXw0nxxWP8P4HiNXLYKomzUIBo72gJi/z+3LBh+ZOb
mmCcY+tRE0Dkrkc4MADhB/wRqM7Oo2wMW38R473vM4pQa/akhuZnbhNl+FlpJ8OiDiosX6nDYIML
uXZBOyA5DDK2ZZcZhGQnk0It9iCtRYnp5TMxLy0syTEW4wfpDFKRZ7IOtS24l0Nr0w/RkKubklZp
mu7/kV5wbgR291p1In/U/4b8d4cdcu9ZWmuyBrzg7qyQsGG2WVzmpN5xdXZFkyzi+yx6Wfui2tS4
Se7eF85jZw9WVszuQD1nbXYCs57Lqi3L8VMAtKB1rgBOoeWhY6ishXilE73MpTlVWAen2WKZxUUm
IE18yXGwDLWBRd24+aQgQlT8bzNtJRLL0MvG7JXJ6xLdZl0Efj6ijI9FDXj+c68YTzX9HJUfXohw
NyRvWEtiMkUCWz0XVxFTerpIIU1ZPdOx5zJkkQ+lEr8sGgr2JUgVlTi++iL+0HYJYM9RbwidMNlh
eMk32ifIfXwHfimUJK43ExeCCiUXsHlU7EzwfYVai2i+697BBoH6EoCJWCavYqmcs5E6+GhbuAd0
ZG21ecwCJ3NORdrWVOW8WRG6OxKLSIlmFWTkohWDPEFp2jZ9RuiFzabCPLP203PLgma0fIDoW2LU
D7z6ZpTEhk1LagydZOKFHFGR9Rl5FNCx6L1CrazkcyrOfGRqoFnTfbvRFt/pIfEQcRBt4AUT1m3h
MWRAnJpc7iIjzWQpqjs9S80eGLJ94+f4giZt9nF5ZfIdX69/PAWzyYTMquDSspxdhngaKhQx8HwM
ulFN4qWbnHtzi2fGT77GYTX20CyN9bVLMsgj9NXoW8VukpojDSaSbGtfLzFIyrJvI6V8FAFW1VgK
iUzHpsYl64tvdjvoZzfpsQaKnpaPJ+f3dixZd+mzlvGgNRCj1NiZ5kfzp3gRO7w6GvyefUGCDj6l
MxyptpwXPFS35BQCF3iGQZQuQoFhz2tP14khmyegJPx3/nzAjLYuBU6RwriA/HcZvlUQxkZHHKEx
BCdwRoUwAF6nuZ5P7rInoLPjWG1hAB5I268OEJ050idPwHwFamR/Q31EodnufwjL+mDZJNB4ronH
wfvHXgdLHLf2Qc4Lh6ab6uTYYrekFYB7fzAwdoOh3Bok58V+stJl7VP7kpdW8yr332eugKVayfhC
T3KviSiv7OmtELxlHfMNPSIjNFE7XA8TmA0/K0hV5sYjE7cjE+exoQl8wMjON253r8te/VFMxtf/
Dx9O5XNkqT9uC5+l/2Q/OCEKvYIECoWzKjMPuL27itBBmxcxtj1DR9fNYF02bF0HUQIkVojMVW32
0uynCihPDBvRgHkTSqtE2+HYxs/kony9bxQQY4FsYp/rTC8LMBXD6cL3Q9kOVd2fCCAAtqvKGAHy
T5dYIeXV0IS9w2bRzEJDF7t2Rl0ztludi93aCIG5Xq9BgWpsf66pwQ373i6Os/fmbC2mFzMOKTVs
JN4hR6ny2XvXKIn8vPN5+bFQ7gsVeChcVWn/J8BesyJKuGtnWjtxWSs74/XCTY4WwX4/xE2HZ9as
o+68MOZvZDmeLxToBr8CYdDVrheKrKxXjHKXluY1LtlCSHhM9hJmeEHtxXwWTP7/7H6rJlHqP8Pg
4IQuiK7qCvwkStwjkw+RZBIb7vOZTvGdS6yF1rg3fFYE8VvY+urbsKvwjMaQWAXZNEvSJ01ZF7sB
AObqlQRh6fWJkeqM8C84lL6Y9upLHCst7ga371+2wxTL9jHWZTIil6Bhm2ez5ufgSM+tofFGrtde
AcSIAz1nyHXYJ5bmt8Uimt9gXXvipmJr5vxYir6arU4I7Ns0+zOQOacCZcAwz6YNaPQGp5SMMsgu
Vn5AnZtQ5fqgJDeH5xu9g6lzlNwd8DEYu6iTBh0684Brmt4U3FznadJ5sh4afHPBf0VLfH7568b4
bWeTYMMfNZHo1VVzDC1YBXPy/temHx7ePeMhpEh7vgyzmuZFvvgxln+BDJJX/7EmbkcWXi0TIGH9
vC4Iy+w8ELUaOm2Fbaj5xezeKmkOMeyRUCUSXFPX5WILHTfWottzgQcDIr19HahSjLwdPN5IF+oZ
KmcMvVko37nddd/eDRjePXxr0VZ25QxRuCfNkcqWmNO7AlCgXjr1nuLzZYSp9ULplF0kyxGXFagI
6GrVBt+RTPA0AYLypBlzbOoivCpbzI16bBDQFz6ZV0F8GZq5zECXhEpeTSpVG0fjsQerkxxg7ywr
AJYPvdZyjkRp+bSFBoxmJ+p69XG5YoBYrDPOsqbB1ydsWhY9YgnTBtozSq7fo+gHIVKrfNk4KCcw
LJuZ82tNFKaFgkvYH9Una3lb28EK+v11PXNWz7EliL81gDh1lrCUke0qSRB4d61DNFQa1phQ0FfT
GmL1UZZojERQrKzaj36qDS+0KPOxnOIVewJtHSTeljZNr5skOnTynwdv2xQT41dLq5gxwHL9+90R
9jyGFlgjKKi88y6LwS1+7sGjNxec+G1dUnKpqYw5ONikNgZVX+WnYVVerDp0kabGTwu81jUkuqtR
N0X3fKc/wAtC1DRk4jESstnlCSjdFbNKjxxMX6RYY+/M9T6kSPpWA31N+z8vF+Cwj+2ukj3wQYEo
wzhf/hzqbAhBcrXBvECrTHKETpiqW960FnExI7Ddp9w+EeKPVS92b8nSIWF7LEhPLCf/mXsjK/HV
uHuLKM1ELYrJg/DM5FwQskJ/bDw+mL/qHRpHm2J5SPGQ1/kdI+FtkPMCxWyF0J7pXpw1Zgp9/vnR
v7VScrfGJkRTxKEz4EQy9zU86+cLoyi2PBUEWw2d7GkM5VQ/RgLqlyXF0NyiZbEBX92OQK+OdoEW
n/z8iZ4DLt3JZBPxrM+GqDqd2W2oYIZzoP77G+zYDPi51s7OucC9E3fOVhYfWsy9bLXs+LJoWHqJ
++2mQcTABkD+dcKSRyfYBdlcnUWw5JpRxx+QjEx7yvpFJHromZAbrUBZMMLonPL+4/NnZfnQMQNm
WeV4/Mxy2MrepnH3E6aSu0AWzdrXL1eEvtFVphQRcsKrbn+rXcTVPK6eXQvDGZvzJTd5J6vC1aH1
bDK+qEVUsdX2a7GWpmltY78t4ObeCiyLUt1aNEq5kbbiI7KphOU+fbIW82YpwLlQo5GO9bzxcUsd
AzlMA0jtMIYtKmF/tsAWvc9PdeFIdthQYte2d3eMGSSgf5Hbt2ifOHfyM5NggROG5YrH9nFivEQl
nbYmoJIkN3B/H2mBeFrhBFlL4SUgm+Z817ce/SOSyZ2zGiCDwpoHH6skZgV6eHJa00FosjAQ0wy1
15aORtM0hBQXdwkokQfWZEQ9L367x+3jBJIU2Dth3bP6fkdufVZ5byuBM/IypaecjeYkzEMbfbDX
3cKyUG/0YLWKOAkZ8d99LGtrDudm3J9Rnt56NOXUcJgj5WazfoFG14GypHMcBbDwC+U0am9/8xig
k05QYAoSs56v9nBSruepJ52ADrPZtwxoe+pYfq6noTpoj1qEKb5WzvXUFzzEqlERmCQB8FdJ2C5l
OIGBjwgaMYNmEvm1HSda+TsZ/uNie3vYFDQa1dSSrftafBQ2+Dc5HtS1juidAJCgriddio+U+UyI
/nzPbp74qxNAEICNs3rK2DBaGYeN1mZoAajcCiMC/sfWXqpNyrsIrZi/TfcURXgPoWv9ms3IuWWB
SDXss3khOSeZ/xlqnLLNNW1JsPKmYB0W/GMED9mqGWpginNWkrufGzR8RHip6M8uokkM82j/EyvQ
1I4qvKNl0nl6bTWM05CRbaxnI+/rHmEcpxNzd8ATGDKaIZ0a9XPjABQPgv5VFabLlM4dQ1g4hhw1
DtqBxdk8pON/gsb3+1IFcSQhGdoJ0Nn4TTEj2eCrUQEIQvh/HyodAd2QahPr5uGmQHPXLkW5OtLD
5ll/9tiK3c0l0b6Yl40+x92V1EVblUB2vjEzFPci+bZh2TVhejMo5EYbkB4SrFnxRs4wrcfMDJjQ
uvxuOoWB/xELq4ffBjjNqSGypJKvDO096GTgZnnuj8mpyUeQE7azoIhI6IJN9gORaP5lk9DEg2je
sGlgJmP+VQei2eYrvRnnJYDB091+mTZk7y/ruSZeZKFjb1q68eWe3XtWWohHoByXiBzpRQm1MN3k
2XfoJ1sdc5owglerU14rQNf+iDTkEqBQGvc7LURM/OcJkfy3eOQEd9nzI3Rj0EOd3ilTzJOXCA+u
E265ksq08o/0mnVf3VRWTH2EOssPwVbjqrH12852G2psRITuONjR0Asx0zcmt4Ux9+9PibRb/JN6
9EDkTF0EOFqqwVZSv+TRry8HKsXhEV5Drn0axPb+84NSvM5fTMio9Rm43ENfLS0lpSWrw+EE+tMc
r5k9NKBLmaiGf6yw+6Y+Rq5aYgLtyXjgx9RrEWT0PRC6Tbq5qKxr7RnuzTcNBKqEdhB0fMm3NAm3
JmidxuzzWvXA1vp5ZH1APjXW+n2HQtn1YGVBCH6A8pappoRyOkAhAHcYptw/EtFm0ZM87wnHSBX/
EbNDnzmVWSSoBuvN5KbvXd3u2MsbLwj1cFm2mVVX5UBF3dzU5eI3XGPylQb8OXvPM2BZyFqtxRPt
GeInrRn7orPJgRIMhUiJqrgY6vU5j5o44goB/dfGUxIuo4SvHjMkrGCjXI9ro1JmfaiAWx67jDZg
BeWySWPKSCcMfLd5w4xtkAv2kIBocAljVPDxfzRpOsXQkDqq0jhxbF4RVh74MG4zFexDofNhhqlW
oA1HYWLPoVpLPLoOx71AWMZJcV5rhjZh4SZg0GoedS+VViGxLFWNPJ0dWz8WDsfS7yNJeoO9hP+u
fepW/wsQU35WnK0ZwmkaL0uZvuuV7wHUByeYl6Z47+5BuKuOPTgP7tAj/m+L/nKAzJ++ZJynjsvp
o0r/hKOqQQ6jEcXTAzQXUqa6VZZy32iesW53AmZp6etL/z90I6I+91xGcz2JVC4hsQI/Z7maVfwK
G8/N8OYx44LElJasQQYv9h0Q1ShdIUObwZ7oDfdWzmml8AumJfPvxiL8Rtaakwiz7sPOYP1kV0YR
grhGpriN5uSCqKtV+h2C+ZBdBgKMlK7DrqftG6bFxJvrmVtoLc0wHaoa1Vf+SUhcwbPwEchUtXRA
vF2b40s+AzvLn5DnG7jsAir4miqEOXmRg2o80/BGaUqfa2mdzfOioXm1apLSQ3R1qs+jQKRieEd6
xEoeFt6oppEYcyuLk2+Wfq4ZtTf6YVsyVaHBitfN59hxNaSyeZ1HT6FsBdeDhPnCEoWXhcSMbh3t
gdgT/BJdP262T4T6R9aXlcIpPaCJdtMQZZ2vcKhjSvlfiEDwR+/aGNMOlP3DOT2gI1D9F+uB1LKg
livzL2iohmhwpCtBIfxwBvJQ8y8VOA/UtpKPV9TIAd7oKyK9h1kmqJJbq6VnK2s3okxt1dSuI+X/
mZR69cfYkopmdxwGSOv9FMaya/Z6xJTD3azIwcmnfQS1oC4BA7cb+XDGuCo+PvQx5u4LV4aW/d8q
j4OnEpjEw65FhZTtmChr5d/4CekupCL/0X3gegBbCth78e96N0DF9wST8WgquJNdYpAO4zKwlTmu
l9+w55d2BQcK1FhqnVYuoao1V5PE2KVqLkJWZH0boMUoue/Kbj4BpyL4elWNgF9sO2qAZ9iSwFvU
cu9DA2IiwzwqesTtYAnjDoaZom2LtTp9XBkbfizoLIhXkgY1ZsTM6uNA6u6ALrpQDI9FxPWrngGf
TycqS+PKO/WgnIcC71PEWmu4lhwrXCF2MUih8jG8BMZu0oeDo3NKGqR6lyQ+2GP5qVzOgKX0W0pP
ftsmbSujoe4P6r7TdwKCCJbGuMGhHv6hWUiB7mEn6qdl1zOPDiTqDSrLwU/8vsFGwkNsduP8Ak8L
GqGx6qV5drrFg+NKq0rWAtT3KwNl11ReYLRa496yRoVglKGJlmEESUOzkcVT1hofLj/VMHbJ9gDU
jT9bmreOHNNP4Jk+Z++Sq/EdLeHu8E6Gm1MDtxDiyWVaqJq6Bm+GRC7cUsmKggJb8xzpxFHA2xwJ
Ln2hi17D27vMKQCa9SH+55yJrKVRfQ8++p2Od/zsyJiW9U9guLVr9m/0/rde7QGkv6oN9CPf3gAE
h2QHhktC8ysA+gIiEMh7aUN+/fm4lwAkR01s2ezc0CyHJCVZDKaT09RbLeJlPK0QlGyKQ8tcpR1O
v070QZBW9DMvdsHeIOJ9BAAN0nYM8brQJD5iVbcGi1E/QgGlLyiDrHeA/Umn1oRhKfFe4Ng5uzMZ
fT4DO3TA5HETERuwcprbF4zTD5iBu3y6v0IoWIjXR+4CdhziZSBuMSod9xfqyh91WzCk5+DxWPYB
SL5w7GxhZLygvRt1jbB11Xb5vT8hObu3IgRt/ExO0dDJp4mC66neZsWpOp/DthsAIycxlejV4YEZ
0MbLVK8XhUEaEul7B+w/Y4kvUiYV4To7PXzNRrOuXtZt2U6exvMlt4epJzcanEAsIOKlQVtswHnh
9BtYwOtbrXRUXyLJHiQApSzeabF0J4OUy89sVuHNPMafskhE14JxFEuRg8/PbQ2HPI1etJcwPh7a
MzXAxsiawtVJRfXmiUlMBDQ/UbE1agK57JlADDh6FvmusHqkfMZlB/fw4g7jYSHkGNjcsqMhPNJL
ogZuhsuiqLVV4Ws/LKfAg1b+HUt+YtnM1+mjzYNzypSJ9yyxsp9beD48U+JUCQ+LhNvrpQpQ6FzY
OSGoZn42j/QInHjz0b/5s9XtgcWdhglgmgh9Le0I5yRG6p47hc3i/qcb1TmG+EEVLsN5+KHAXPJB
goPpzij7txc0i3iG6IsGRgHe1pn0g4t6iITY0KmpZ9xla7FRjhfe9fXD+L+hzESIXLVtYLld2W7b
n+D7UBom24A9JXfY0uef+W5BXnMFFPHOXuTsBi4U93gIwGK89BrWkjE5qeyc4Wx1eSQez1uKwDKI
n9dP50j5a86D0NvJMR+pmzqQIOeXEDpHU72T5yktpNR/PZDe7KEgVWTeAGTCB0glGKFdjxPJ0QLx
iXtBJuaEy1ONDnDZYOfbthDhc/C0hQkzpmsnJN+FadbkFg3PhEh9eJB2mA//Gai/JYYPwlk+G4Mv
jCVczxQQ1RSXGl0bu98S/ZtagsZnXoGcUhlqqQVA9GfWFHKmQkdIwBb+eruVhZIU4uZzWWCGLOtK
A4LETrLQSA/mOSoQxUb5jxQTPbFWKKS8Cvz4lmLODCffTlFc5LfqNuG8Crl7eAQD9Dx4HJ6LksRG
QxQ74Lv76USN+k+HDSjMDvf+Qjgy6iEr7E7AOFvjpzdNly2ThbTE9QbqVBpioxTl4v4yOtZTlVDt
sq91bXASFrtjHAxC/oJUGwbvIuwXE5jbEiija07hx+GOKYEiQoUBaL8u3EHW8GR673mIYJHe0/G5
gDKKb5MSkVOn2J8R6hcP6Sd57IBh+Vla20EX9uR6AYwXCi9fBR6ucrhG5Cr1X+QxsmZB8+QfHzbH
7xCZU6d1OV7ehjMctChrHUs4gdviDWEzWLqI+6AATZCjJfYC9mu9S7REgXC0HYTJwuZZoY6ccfMJ
jwcXAVTBcM55xlk/HqSK/sdET4fFYNCsnrIOShjyZPIdIfrfL8AawzJVEgAQNpTdRcosU5hALm6j
KpXVPcCeDJA28j8V/JyowRCsyZ348gvjP24MF7vh0Eqstm8tpEb03QUhM3ZPxRlc9WXFadTLCnjy
rX6oX+ExpPyZO+a4A2GgK8IuZQBTpHGrNMexI1AHECMxLbO6KZI9WX/VaI58cFRO4BA44vfAPiwu
XjDuywXq+8MtjzfjkC4HsuR846Oa7sbztqoOULakmz7BOoeAb+WW9XavVrhaxRiMKJ9oBqz+GTGK
gPJvA+pN8PEt7zU7GdDN177KPLt/Xx910ZIIr4cVOQjKxqQ5Aywok4iC/YNR4GSfnNGnTA78trjv
WCxaZvdWN+svOF7CLlJpEF0j+EVI4gnhtzz3m5VxgqDtz2yPHDhWbuXO7UPBRloXeIXK4xsaTbjV
2eqrVvfaUC7X7jrwcjDfxfG/iXbmSESMyo1uIt+Qd6MQUXJUloAM/doNwcR9WJqjvrrccuWT0Gr3
Dm0kAm861RUDk/ytDM5cpC9bGJ0cvsFPuPSeKupXkAhUeoQhFK7pTGI00duR2NQ6uRbQMtIIR5lG
60LZnXrkrGn/E2I7AwGTwrxXrLh+uWX2PVllepbfgg/fVkxrWp8hwavkx/V/O6kcBok3QCo8QTVB
OFkpzfRqETNJ9kC6EPROfyYkUnZDpTKNyGplAGxcc1rHxrVYpXcVT7VHy0K1Qh/unwR9JTTmezwi
xzFCJrnaf2w7WGZICsKnYyEq0PoQ5tNkNkMa+cqQoqepbWhlrOkD75bDyYTBO1yFvh65CNxZhQyj
FVRa1X09mOkglBrCXXvQS1VAWYPVdFAd6XX9cr8MTNcySNQU8Fhz47027ZXH2OJVqmpfwBF3+GC7
2f1jh0q1BVU5KZEvSJL5YcwdRRFNsfd1IXMr+S9HiAQrSHDzLR0glScAQj11Cs6KciGK8py+qFTH
p3Mxp+YBCHnHDgi63eIICEzFUtG6CWM/d5ee8ABT+mHdomGDEi8kHby+hllIc/EF11xs/QPlZhHZ
f/VOaYd4jHzKQeuBXrySlCLi1Qt6uDILwpiaXI5oz8LAZWM1vfZLwrtWh7KY2s6C9uCgsg1t4UFm
N7zZyj4d9xwa/a78QTzAJ/AfMmqPBQ6ecS9jofyyzdZAQUwlfRpWlOm2WRF8zL5+ec6L4+aq61+C
ojxPDtf4F2QyGhKTM26qaAIFV8lJbnBRPIx4kkolTdA3UcYcPnIMC0eldHtaCcQdsBnVSLqX+N/+
Sd2VBzBAHfI3XNT6zEBNJ80QcUlgIQ/kWKQ6Cet4n4aeqfqnhFERgQO+GwyH2xJXKr6gXpnvyHHT
IG//UEdX15VSSZepo4LZRDAKeQdmGKBUzwqeWrP8fKYZkKm1eu9FnpI8dJ24aUE1e1RLL0N0774L
cXs7HslSD8ri6hsIPYnJvvgdqS12veRscMP7HbxOjYWpQzMXW3fEwGim4jeCol+N7rM4m4gG8lhe
fovdu+feiQsx4v+vuWZCn9rHd0CGuJ9qz0U/TUyoi19go8Cmv1d+0Ryq9auBgZq45fn3QCw8nD2u
lVHBNTebDWHviqhJKLfdbpdhfGcekusMVDFRN/t+xayjwgWYq97aMf2UgcM8DOKBAzNdUOTKveDb
e6EBkfGpQGfqQjvymTboOPunGkQK9CzdYJcKvdVW4TDDSijxnf/MNgg55Vdw3IsIdA1PMt3DVrNX
iD3J+/kyw0RJC+0N8CdBgSHXZVYtpPsfFCOklYARh8JTTG2mt3d54ydwGHq+iP8U1XZMRqs//ykM
ZQMQODXp16hDVFvPa/8ig0rObLioeaYreGtVzVNhiD1AccPnPjjuGS2T/kRjYUafrXm8NvSryQr8
bNrYzeP6aPMhDdCnJ4hs7xs7Gj3mdXxGQKoUrye4Cf7CkkYzlG7SzJVErANp4lFr+v7QGxK0T9rk
1IUzhyhnfy+05gqgbh8czyzAqjyrC6cgkqv8oDiNWv9ej3QAttgJ7dz1OP/giIGWCVy/evR16/Up
2E/zufDpxAxRv5X60R/e/QYTB5M342uM0cZh2YOli/AJALjwG03h6dRcqeHv6xAculG9kmvID47B
JtkuYsM3qQ/+Qsb10YJOVnIGCsHrUk+StTwAMHt/L53ehap1U1vSKs4B9r8ph9p+VxZ5CJq8tKUj
4hkQObhxvjS7SMLSNpKmsjELu6jQrdL58xMhSaeINezwq3PYKIRgaDfKktCDWGXyOSWjuotMa90k
zU5vn3xD6UcID2YCFN/9l5e4kPjM9e/WjVzVBXqEbjszANKxcartAkOMzsizdHJIaFOaH0+TUhcu
DLtVihxQ2Cl5GvaZsfh2Ww5m23SW4crWw21/Fd8dnYBuJpVRJpbMgDHMRUwpQnKbZTrxxewuj9j0
XxDJrUS2gz6XT2g9J3CoKbdjsMqJ9lq8CotLsXq0ruciLOms96CwP79EC0ygPID+Wfz1JqeSoKe+
+ULthp+gc/XABGOjFdZ9u4b2mJ5Tc5RTIW9kwtaaSMy0BcH1e72NQK+5h+ZQjKldDyUAwxTir4xo
BCf+srSgnZnwJ+qI5XXJg2wHnET5Dd98Sw/mup9CFZOswoynPCjtV3budzTl9MH6aEl1eQc3kIKs
LjnCekEOjGMhJJo4Ua8Qv0Y/1C1wYk4qXjG7ftwi9xAqdjqKkIr/nQ3K+K0HNV8C45YgYjx0rGhT
ip5xxBj+PXdpAB9dd4xRsI2pmMPthImK5Nf6O9V9JkLs9X4dD+VdboegXhO8EeE9ZNw8h2I7aacM
2sGEWw5R+fcPvlraBb+sX5GTLgbMSBUBQ+hv7O0BUTuhxPU+2uGLQx2VQrl01fsNC5PhfGpFgog+
xgZ4yW3OGiB0zhR04m2Ng159b3qkfJvMcNTRAlx8jhizovmEsADGJ5PXVgtMWCeF3KjDZhRTW5es
G8aRNeHeuf9AhdQRlybRVXL6dp82yFHlFSxCMz4NDKVMPi19UVpgrxb1xvIKbCFPlkR4DvNuz4QG
XB48YYxkcm6x+syR5iWc6qkLpI+nBAHVIaW0A8BbrIpWCRD1XN5iMBPyap4J6dP3jFzgjR+LWUR+
2v6gJ2JCla14ZKhhrxHwH1ED1nplxSENHBnTa/rx0sT0Lm16rO/oDJlQoqIEF/OdM2V/mi2Jg0HQ
48s31GE34sL8LknJ7/Mw63+T8aAyYsXU/WF+CroK2hWV+S90cOX8e7+Hxq/GaQbDQkPHp2M4/UfR
fw0bCZ0eM18zYbjLOxg8kRQwr/nW82DSGwzUn4Qao6fa+DBl1If9+gTn8cPsL2ZiEyzj4+T4TcrI
qleB12y+YpozM1sQ5nYkR2Vp/4rMUKnpEGjkxFTkkmQIxl0TTUGrXKTkxIJErkQKe9QEWN+Dh+Tj
z0cfbY7JjV4GhP/j5GOVuQ8/nrcgYlxKMa/qIdOIiZeG9p1tqE2h/I7WWUGDBSw9zn6Wd/t2Ud6i
mccEYRXDhJdl6CDosmxSrboCMpdh8M0TsCmhQ6eydr2XH5YbMN3OMzWw7EOBIJ7jGFcuVw3ySgQy
QMKNV/PIU+AVFl+3TZCmspsYix2woywbZbTUnS6238Qy7yM9EADjiezudFb5/6fJ7di2tfRmqA19
JTzUI80j8+5q+TWj7cCzUHChp3zTu84nCkV109pNgx9CjARrN+KXohYhr2qwy/E3CV38WTPP8iCg
TXYaDBrfVjUC7pyoWEjLbUGqjMG6tuH1HTp0UW3B17u89OTzeqMiZZ2QSu3peYB0GFAZaQ+9U5OC
T891fUmbyXD3c07MszChTLPgGrEiTa4sE9mwQlnmoAyWNmmrwmdFe7Tn4zHaDwjAKFW14vuxBhyW
uKDsHn5zDaBtBPRjfANIWhOjyJDONU3uSP/zP0Y2AYgy//2hLcHlbhL/wqk8rF1fMCMdr7I4Jkwr
4qhb8Bbhe4jdaUo3hfVe/v0aKDw49JwFD6NL9aM9uOTESDEAinf1IxRy3skDHjoGPRZDbbJXqGQN
Thg6nFsp1wztFFmUVRXL1DsErFpn+cOfPP56MIuW/FvivkeeDj1ybgfS7fAB74wHbQHUdNrCAgLI
0RNlmoaVdWhkbSUv/w9L6OeeNX2166wcZV6nmNsYdnbZwdM7ZI/Eca12W8Pa77SWx2eNQvyC5Xrt
CUgydFAevjn8ky0IAD1ya/bqZrF+ANxt3SbZK2QwWXYQVZloZFbNC2a67HxMTTzTAl9yPjMiqhOz
dqBVflm9RKsIiu5AtEMpw3ctjahPmlASdaZM1bhLnsltMmR1wf0frb9rzNqnNqenlG0cLO9yyHFD
7JgIyFdj7KR0oDSqsTQ63bvcFvt1eUfS0pw4H9I7mgsdsEK+Vlo8Dr5HZpXz20bvZuyMM6TtGxOb
KI/9jjcgyM1M/fGlKcicC6vHpvcHOSs3VYuFbb3sXrmQgb0f2n0BQiHzhiiIbVuLJlpzBGj3Kj+m
yKwv+ElmCNqlpVqpP80xNJEPzYthocdv2ujQs3oJzaKw18x0zwtqyjLmAQI3Rjm+yrxANtY1dhKv
2w4EzsxVqfrXM+wf+3AXuRCSSfaumQlXdtRXTadXSyJFsAbzjSba2Jf/XAgnTaVxlCthYrJqw+Hk
AMsLSX7bYXyvOCb2zrfdALELysORzWQm46BqnOnWcA7TmzqCNtELHRC5H4gy2s8DveoBeE7o1Gyt
W6CrOflpcfdDfDJASdv0XeC5pOCfGGY3coUb5pGYnal6PXVC9xpPGDE9ygg+ltiv85jC96e2/OSC
0qHyN9i2VVBmngjMp+hj/QszmUMDMaU+dgrjPA+bg8aj766gKjRd0cRsuyzas/2VnsaG1UDnsQ2R
E34FjxXBeIiT8nnIZaJK2jpB9X12UMOUhddWQEJHiLWUxm+8IJOsxfYVxhbfbWBw80y94YSI3+jo
JknJt8ZU2jgfW/LF+5oX/9xE+BL2pVEkBwl2SLM/ypyQouRX9yDEzQEFLrtHhtEH/VUtxG292MlS
iSdLHowDjG4B1Dn5WneTLwgNM7kCN1cj0ZiFhxc0iaa7fe1xHN4GVd/wH3YFoIIf8Q6qRnhMAZKW
4AzgeqcsrU3SubKlYc4weeaWctdSSlhT72M48wfMv8l6+rZBB4R4pQzpRyIkkQQMEHtvSa+Nxz9N
aEYzYO0ephKP7PJQR/94JdOvxEHUwnQtdIdNIvUyyirBJX/za8wr1dt+AIag+iy4UNw9CpVZYyPX
pAHKCrXov1ZaobPk2gAP/hIwnYto/yhsyuEuyy5vLO+Qs0XVeQHbX34SKM4qOxN9T9PerwHtQKVe
+15OiFiSO43WYvumoq1w2Xy7EJUXKcnd/kTrG7yFn3vj/33dv64+nWMdJ6cdnwX7qN5Ie3HnT6n7
/3gbh1Vf1Ye6oJW6dywD3n78jljWedoKE67b/nxBeRv2elZ/WlTKuS43cwzjKsb5MA/phiT2uLHL
TqPXg/3zSnauvYNzN0wR/RjsbjeJHgc1U6ieQCT4gQXefvN5bw4A9Y7c0YODEKws/VUyBm1c6vE7
f9dQblGe4X0ZbPnDLtqLecgNsvN68QSGKHpTG5K5dYInAagStFrXcRJLDyLKH70Jaug9u6mbhThu
/SLGZ9OXyQk0ocpFeVDeG+siAPE7QyLFe7xvXeugCttT13tXzPQcxnIlGuPoXXqnlZnwemq65y+4
SOdrCY6Cula9DYm6DrLHHfdKNOB+TGlJlwBMIw/DuvjLFJJ/uHUlJATr0G7NEx482Zstot/9en1u
+6ubx+uTFYv0rrJ+LkrFd6tIAFi5TKfvFf9hekbjEJ07+fr+w+6RSwajoSPwozApBIjqzSyPLLFU
/3ov0ZmL9gQb+UQGIOO1OnTaf5ECZDCqbp7gFRe9tlMKAsodIdVuM6sygSeXRija1zYSB5Ediv6T
bXTUcfMYpCMZlHyay1zrcMpvSitIGRrGw8IVI8VacwdBwMaVwAcbYux4k2UZ9qY375tVLoSdpIyi
e4O0+pdHep0j7KaALq4bStGbIQSkEx+tqA6v+kJ9TQRY8LTp6x6q38GRXi+s5yNOoNhPMIC6RKz8
LvSEW/6sbRdmPkx4YSz/+oZMnkK6oEismJS0IY59Erbg8iyC2i/HgZPuBpS28FItZitG9q6i6x4X
820GzzlRahBOorsB/PyJ2vn1Dly1c/Cfhi2RF4h/qSSgwYdcaP23Hb7v4jkyl1Rd3Gt1RbD9Io1p
N+azdkJlIIK+HvvJYqIOWh2P0K4yeM6CJHSb99Y5aNTFR4clzVeke4EvCSMOBhpV/heva3BH0bym
Zm+7i9H1O2E6FziMqXuNLj01iYVw5WfPfuuUb/Anie+VLOnXxOIyMT9EJ6DIxo8Hp2O90upSW0zs
gbL74/1gb8KnV4faQeXSVCpAkUJE35pIWo3VYZpp7Dbunnlp3+KO4QUraPYvkzWx5xOwMIGoJiwf
eIXSkTnjz0tQq+g9RZuMgh9sZibfPDzLYYdNjMZ0e3LYrejiXAAfWk1dO1nIImh6+BwCXzTZSAdI
qMtiVPoZyT/0ySO8+oy0KN1G5BPFTY5QcLWLAcKhzQ92oAOMfcirsHkt/uxXQQjT0FRFSYvZmYlf
25f9/cqaNvdeNWfKwzMCfL43cOIkI60Z685wbgEMLXhGwTVSzN30snBphLLYpj1C6zJuGEXsjmxW
TQacC0sOaVYW9jeFFnZTDBXQYYPrZrn59eNGmgYKZ5jfoP2Vi5AEE9XudEmeAWtKKrECLWKfD8D2
Kgjav0PCIY07UwRovFW+YD6l25LbqB2geD71aT+wIp1h7jln/5YZub85fOusQrVIe0TJYAyg0PTv
SnLKVQx3UQU4Z5nkEkzWCNVsge4wohm/2nRxfqJG2JOP9HWnZeUye61m/bbZWuSkm/RDT37b5ihC
Y34nFs+KXG3r8EjLLWsx0pKZTE7U4m2bbG73joTYax/+q0woUQv0t7lMIoBT/B5SoMylJ0rdVwr2
KBCII6jVZx4avcysykTXczSdWc6HK/CIC4f6cADD3U8LXWnTGKlfaEwRGuNvjZ3zxGqtfEMhnQAM
VijMUaXx07gd0TpKzQ5OsyIIfVCI1IGfHTQS6zaVPHvWeNJDpdFXMowMptZLwv9qceHZADSQan1B
3ciO3sXF6nle4FHrk0Ig6d2J4aTt6VIlCQ1bVi4EllazBKtux2hRFTzO0v4lvF6ucNUSe0U1yqsO
zMjcOcZ1MWYtKK0pTZu7s7kP/baDR/yCpr1l2hDbPh4U5RfKOCd0GoyZcy6M/Fr3SguSTKpkvMNQ
B7e5fI0g628mBrxntCYmlY1XaNWzKLR147qJ4KoVuJqd5v8Q+WFH5uOof5EAWfpTlQKweC1NDIC1
i244GAS7rZU7G6LEE3gOg6OMs6eDcSqnQ/gqNqDOOwn3oPWrDRy6H/QUmFydRz18iZEajMfVoO5f
w5BzjoxGqWt+1cAxnY1FPRk3m+YSctXvQoXIStZcW+6riRAhfkBaYyD05gLVjCysAcu+SebS2rjS
denDo8HoPoP3vsTysT4vygRMiB1OJ9B/8B5c77jYq87egtv5Xq57k3g7IEez/xdgfVLAArEvdnr5
gWnmDA1gwZQXjslqWieys2WoGDxJJoEFdsrEDjSKvpBHuzBOOhyAfd8okvYVRCFBAHhT2jNQMpDA
m148dCucZJDO3NNJMfwd8/BArEsuEZmT/yDiQasetslgC4oQI46vzS39+CBNEvFad1noZYLE1+7g
54JwcrtnWj9ASem+bFNRqNjQLFHbxF72VXixASg2zPv5SzV9KvRz+rAs1+h/u0u24ZFBYj/Fw3Ad
+9w+y1PI9Rw/RFmYtNPmcbKRfU4jDAIXpkMKchMheMapJ3Jie8o+UPwUzxPSL8R3nNWCNW6j2tmB
S7JzfhI782ToRsM+50USIqjzi3Pqc1JToFiasBIYtoAuezByjA3Ks6A/qLTWb4XwnbR6SmFAFcuk
+sR2v+EF87QPUdgvL9SDR7uMrBrOgJZg7H8RglKSEuDM1PAhXSJ4vz4QHO8M8RrXE4Di0aJ1W3cF
7EOLlLEvDShCTs5IdYwoLqSktvXYmGgc8uI7P0zZieJsC2j7BHdtdXh6RvCTj5bpqDOa/H70EsiY
CwRhgIp7etZZ6TDrusJGsrjLPCu4qQfAWxoSL0UfBPmrMYg7Jc6qQ599M05P0PKGBRxO4KJLK77n
k4fQQWoGIRR6EN/k+gC4Ep6ySvJunLOhaV3+BcOVAdqS23HI+exWroR5c7Ok3bZ8VuNrk7AyY94z
L5EoEVa1sqrsMWw1/N2L5HaefjOfrlDrd3YY2AtePWKJpreiPUbVUAS/XoiMOdoqEoZ4lhAghG/E
J9dMDhKPP+3QSmi7aw5Lzh6kZb5d9vSJkRdLk8lOobqbdrjM+TpxvzxzT6CxDLEsuSg2rGS1J8RH
gArteJbny/ilG1WRytUwm2AT9AlIYGMDvfwFEyqMHWeh8mT3YvRtUUrD4ZFcbDIh1SIZGZoMoP8Z
xFagfPE80V8Tfoqs/o31BdrrLQVTLknZ6nNyhrmaoangkACmwqNCP/vJNn1lQdtbbLjhV7dQKh3x
+CxxoaHMFmC3lAGvtUUIJpOJee7sYSJcLS0i74ek36DTGKLw5pxsK2wbUpCQ4cQedTH4+cTOJTzG
pKubNqWn+KRkwq0ys/Mc6FHsKVq0kQ7p8M450nxB1esNmMy95mKeib1I7KBw+ycxM8q56aIH7OnF
d4WkQjz5ckR1E7K61VqmvFX9aen24zDCMuIHK6sipbWCZVGC0w068jEbRm2W+mwfovaZGGjVGi89
NrLdoO3usWfKy4C2phH6+6oq85kMsGs3U/otd1n2VTfxg/SaTSid9uKIvk89S9sYSRUcd5AW3qpe
5W3rtkd7AxC6ZPgM80oal0HrplCa1M3LYQt2TcG3aHvisNRkiWJFknBt1UFzUsqoOsdUV/MXxpeG
7Vd31oeg+ybZQei/gvi4g495rYNXrOg6EAKZi2M38zdf4ZPoTZTYV9++x3E/D4LpJTUPXo6x9ncG
0UMtP7964zbeK22KP6Rqi9nTX/MvNOpILaDC26sbGAoStMIaEniAolkb/yV3ct2zDRqwPCet3vU2
f+4c/l+qn8NH2wm/oxp6J72Zh1dYgFdKZk5ZZRf4OwIjd8y4TqcrK7OgTNvTVYqbDJTEcYEIHFcc
+lWxZg3fRxNZQIUJPH1T5vgjR7199AALIjzeBKzh5Iwa+0+fUb+0/0LqcqZbotn1BOH50KPBVJJp
0EytRVjSS/c6Nl2k6/BbVCZiqLCQ4NSiTmieVBr1gjjvxhfqDFWunY34NJCTIu1PGv8tb0+Xsg+O
HjP/mSElngLdCs5Yuup9lzawaTMmfxhPYej8gda1qVyjFCzIf76NUSnZkzNHEm0EYgUrvdVMU1FH
JftrY/rEBHN4uphzHBNJhbqcmHDKP/MQ+3b9qdCjLZvELZgdjznt7Mr1ebktmwGFtnT0BT7jixkw
YHsjjaAgBZZujIqvftHwYCtnON/+Mua4Y1IkFRpyTFtuFl4TfHppsv4xMWmmrGUzqWYPMpA4CazG
VaO1tW2n6oxXqTd6JxmDDknwUUd4gt8q56yMPKQYNcFBEN7euZkmoUumgTQMZVIpeXOVMZ68b9Et
arC9vpX4cvn1mEUmwYM4sNwFVCGWZDA4rMq4ePC4TC6aFOyYI5P+55zQdoWRy26ZyWT/XFPkg9VM
jU28zWgpgsw03LtzY0t6nxX9GB8qkcbHmAo69uJ1i/6jA8SsFLgJwYFIInCe8WyNfkG3pNzekIsL
f6e17cj3cE1MsoHjkkE7oXV7cCBwq7cxmREH+xoGCP4/P2heQAR8Hpk0pBG63cxdCLXCK36VmtZx
tYsqOr7qZj4b4rSuGoVwvHw184GH2VBlHdTTXeqeGtJ6eEXUW81VUH4cmJ9AerlMYN4Tepa9nbCc
l/2+YCUpHgFmA98i6fVQY1YTondCjlmymWgWGXUahjDcp0KGW3Z+JzsXGVp8mebQz1yqFDawKPre
daLpVFCQlDxen/tWW6hNQzQbWcGVqzzZ32B4Sb7VTWFL1GsG1yKTvlWCB7lZ3ILgqieGRpDAUlMo
tzZllFj2BGop9pY9uSJkaoIDbDBTCtnox2DWT3FpB3dfBxMnVrsvdVoL/5U7r0keU7ld3WscrxMz
x2iTv3OXCf6+OiWdF+ximDEMAnfra1F+kMt30wgNibnE9H4Lc3Mk0oep5P+J+JcNwNfOXGdzybrH
anbNWqq8dTDgZveRvTIqwG5LR+HOMdAiZ5GjZFZjq+6auzkloaN+XTp/VvUAf66QPJ5l4hFtizg5
GsdyRjGDl4URva3OHWFiRFQWrC3itHv6LoJ5VCF9t3EcTQpTqv/jgrNXZURr0pTwbEKneUFgJ6aR
K9oL6pokNKGuFGR3P0yt7Hz+nYbyR2m3k+W80K03hfx+4vz952Nui+8TFaKsnhpHvYCU4TPC9Kz0
v6Yo115bl35sroUQDgs2CIAmfvh6AHnS2Hh5CwY5pbUzmG4fcigpJoO+FqYz/qB4a4NR9r/LJCE1
tFmaDrWSwDFHqcZ7d0h6gCHMhUJwovfmR2A1/2kUUJNP4GAU/z9tMdEQ9bxNl9Qs5zpVB1SXBIee
TpDsv9PoKy9u7JIAK7QZ9GUAAiQXUDmUZJrrt2ImOuF6l+VCcaOUy6QqgaeKdzl/ITQ8hHgba2R6
BLpZ/ZuhJXlhVjYTQQnvtcCz2dCZ00LcS7Jz6v4ag89Dkof1+W5c14lzAjNscvrvsqJA42+StPCn
UtACDjJ38yQR1VGCBiLfsM3h9w6jlXPOf31ViXDtcD2LC2fLPuUzhBobLkAM/fivDfIss6FouQOF
eIhNmOrZGMXGnD3Tg6ow7BcF1E7BtG4Am5mF0rSwZyPHbUa/S81IwLp0VkCso8XpcIl8wUBBGwNA
OdfaZAsVWBDi650Ec0fU+5YBnDwOe33KwiBnXwxpzbmEAiqAdRWK8sDdzdbPlKbdPKh8Ykz94fvl
HeJ0NCqc44M/8fpiZGrTAjfIlPW3yw6m5gXW7kk531/eeWy6rJbaQtwrXnv6MxcGqcHomQKVCXlw
pU268QBIEAbIt+tLXQRYSaWU4jJqs6j8/FveHTR6j5tINfRz4sf3pgAIedU9IT92uo2lCLFVaw9h
re7nuxLG07HVadWvbM9qHKBXesUpKYttabG1k0OfstiEWeQOB3nlfxTUslLAq1cvSfBFENATAGn9
u8JY+EoH93JuISIw6M2CqOyWEK6biSQgXgMI/64VkXvddC1+Z1g8bf1kip8DY4xGORyZ9kb8tKyS
KweqkV2G06ySf/kQ9tPEc+96zzD7pW43OqbHz9+d4BcwjBZ3WaUGhIXA68agXcuQQozNADW8CQCH
Ljr+oHLn8Fivt8CkiwrXMGho90UfBqAC8oEYoHAxQlWjn1YDxuokdXSYJ9AtYGUYqymX1/mxkzSp
T1MWEdHBWUHMclhT+Illoc4GY+dLd8BGCuq7E+CtstRD8f+1UGw/KkS+QyJAArRA9r97vYRmsXXp
IBilfHMafIxi4v3QmCgfnQ+TgyBEr6oqyIMU7PU5q8P2IhzK8zx1S3TAniUBaxtq9oRRQcrvE8Wp
X3qt5uuqSIBvqTvhQtjhTDVN3GJpc+KpjJeUcUZ1r/P5GM9r1ZZEYFoxtp7Ya/9R/lWCHzQTM6g4
t6j2Y/t9L57P2+x4UP2V79AXirq4+ZsqEQU/QKV6ICVRDxfe3l5pSqTv1j64Q7PvFkF1qqhwRvdG
Tp3d1AAs4W9oqwyMlEE/LF5AkoxXtQ5qQfOtiS3hWRRCtnKO2Y/XPVRKJJpRH1OD2pGRtNFN/yU2
4rPuFkw6c9yqxyGFisSiTKb377ecuTyho93pLGRTnpGfZPHnuUICmTnJA9N+W02fiNAeplv/azl3
YLt7VEFmorvxxtLyOOUBCd1ZvKHnUc0i8zAFGTp5431omhcNr5PQDQ9Eb44ruxn2/eMSBcwubCJI
hEW41GCIw2SDRbKG3dKIU5IH8hYCwjWkdbEcqFi2HMjBkkp0IeX89AIvyqLKyAep1gj3QBucwQEn
fohQ+P7IAx5AOqauyFHzwbTF2jhsqCYQDPhOam5GAa6Ij8kCTXy1650ujbg+4pKfeQj2eE1w4gLQ
Ww0BHZ/JXsJUzQyzJTOOQiExr7gbzdO9IRU7AJgIkoVoFygl8JbEubEoR46C3UHZ2NX4grv0M+Fm
BVBHkwQt6dVuC471yQ8AIC8Gt/MRqd22XzNWjiDIvUGLooxw7WCRTnvvxlmABi7OB7Z5lzyda1JG
P5zVocqRsgJ95IkgA7PsuWk2yNmDxcCAbGgsPLNQmAO3cat4bZCV3zpr2LNkw9LHwL9sbuvWoS2T
98m5B37sdi45TtqYTsK72KY03j3YktDXcsfecLgpMWL0fR7DQuH/YxauA3O78tH4Lz6BbvmoAyNf
VzfKRHJiiCoSkZxnR8DcrKyMdmIhx+2kLKEqDlP4H0AINa/XLoWlyRfzeFnp2MMFXOa7V8pogOZk
rGIAb9U4lR/Ky3GNVHhVjpHCE8TOe6wfiC3YOF6ODoNGZVD4wK8XTKEWbWKLIPzOsAOwdNYDq2jd
yiPuXYHe2MrPAplzoQRD9HywBdC+iFzYkwmoIMl6GLAblKmKlNS3nHuzJzeHjEPl7RyCWE0O3OW+
mOUWlZk3O7aea1pgMx2+k+aMXUDoHX+x4vsj2XkOboinAlg/F4PhBGmel/xLrHfT5tHtB1aBL0YF
PDaqqRtRMhnidnXT4JINqBunTq3F1MTIK0S6c7EOVuX5n1lGq5XQRWLQK1W5YCXgrpUyyR9hLxp+
tydiQR2/kovOZtVungEONetJa/0gLgeGgp5jUbQqAgRytA7oZHpGR907FbQqmCBk11Ok11a+zHAF
LAZa8GEboXww7/lRiCmBjXj+p6Mel/lqQiFj15laIThnwDqt3qwwwgLOGCQgnlL4Sd7PIXcX1ZWL
6zj7i/tXOpMdX7iDofaPUAc0gusRbIC4iuwD34/paKkVEP1u27D4yNjeH5vGYZ70p9jowO+Sw1NX
ip+nloVLH9sF48iMMlHAukGKvoDcvRXfJsT5j+yts15LBBBG3WkZ+dwRQWidk9dnN3C02N0CXwG/
x4m3ckC7AjVSKPt2nGWT0I0RFBqWvfcrqVNVlUwkr0EGbmMvifGudNKLUQU2AJmXGldUgaagz483
Zy8AiZuMC9zMieChJLz/LdUo1/Q1X9wdADyL4cddcjQNooSUwEfwTDHwKszhjQxFPJAACEKH7XBV
0m2iVJltbsogqkzlz9BFQ6ou4EwhtC+2RsOgusai7O04K4YYF1ixzFfgIpeSpf+Tuti0BG71WF3X
fFydLivLSa+FxpsVRuW3ncDI807SQd+kfUhNb+Sf5PNNiHwS+/DdFYIv1nME61ueekkmJmxj9uVX
Pt5EM86VThM6eLJhIbKsL/lVOrGVyelyvGiVrVj8DniOt6E5lYi33hX993uVG9zm3As4vXlgolii
a2GzxzvKPFzuMmv+uF20b6ifF1fLIzEwDsz4PcqMjx+/rq/PWW3f4IlVnvaR7wTueRaIRwMO4c8J
6aJM97+pZH5HcEF30yeH9qwh/UA3SQ++Xgl1KOJQf7YWhTNZ80CnRUcOEoAo6/4u/isVdjs09JiB
FbA87493+91SwJOZ7A+hgV5uCRO1l8eKhgPXBu3qyRqAZbA8XkZn4V73HGkP3XPEWO9o4RKZ/onX
/+UmobZCfv3S5HN+CNDuoEMGN4MHv8MCsSddTFGk2QFhLrAKQpiDbP3ZDIQoo0fbGAzWwoTaeoEY
I6wWHEJBitxql9YyArR3sAj+n2WvltfMZWqdWIfoSad739aEjBr3weVR/36Fm8gBhUa7UPJ8q56i
NEqKcEceZMzFFSbue6ldGku44l2/PFymOx0Lu66y81Dbwu3DX+iHSO9ZMcEXYn8zd5LBLdEgJZ82
9PLtL5YVuYIytviSUVV0X4yefgizagZIQK8b7v6VsqinP1VpibdEDW/teY2FHCSN2w4wMXzHByw+
v1OYX6mbN/W6Iq5t+/pOtPlzEX3eysL2yBM/O9x/+y2fps7UzTvE/txOICv5GVMqX5fSjUarG9Vd
ZQOflNdib3JagH3wY9GNJ78TrsWp3uzuWidXpL4TmmVKDHLwXdOJV7gcGnuPwt5L8JcYs5x350j1
09euTdLjI7JxDePH9lddrzMW+c8Upy65FH5EpJvppYX6bGuroEVQuvlp3K+dgiSmfvjqlzv2zsSG
91lO4kDZK/BTR1JTVKzNuq1kV8XHrAwVzHAWf9yVkFXOdwzV3stUWjdHeqeWoWMRaM7rFAoaNdgt
LOCigQaOCYdQHVjjJ+gCWvi3+QqaZ/7X5nbGpuAkBWjZ1CH/HdCV9V8UOjHbolZ+yoih63k3/LNx
4ZvhZzbAqj7ZumMkIcefbUofAvaCjxhV4aiya5ZA5Gi4sKdFtgWvZJ3vhyGl4N2NEfewa9nngCMM
2lq+C1zTQOcNSD2LClGU/AEowyfveCByeSZF63AEjQyO04xfnLU3QsvA4h4X3B8L4gu35kEKyF+Q
X/Dj8uidx/yoU2JjUG3zLSgK/DB8T+j+LTqmo1BQOsIxNIV017+S6aDGLd4r9aGm//uHAfo5nK5f
wc+4YPub4MHR6op7mXsGyoPWyhVo4UnhgJhfs57+rHTVpDAjUgQZSFkCyRZjlLKfvrG4sTRPkgHc
rwEqRFeVbGPA6AhyS5yl0JtDQF7N1fchkWHl8brT5r5eSslAgJ3s5ovNodGTtQrtL621ad4Xhv3G
qAKUQHlmOYDHvSEjAkSj5JaoY0BBSanHVyNkpEGy5o1BjwxeA9VET1XbdoN29rJKg7D9uma7xjnO
Rx1VThXivmYEWiFon/bSjbgPJjQWmTKh8p8XDKBFq/rJvqBRpMpmunUNYeutJyzoSYU8K+okfieF
0SYs0+qFFGJDlVJvwe5wJxNhF09zndUlmX1YnEp1XZqxwDxpnweVBd4xTFflR+kY22mVdzqs8xMf
1NrWNbHPoCCjxl22d6hFyQgEzJN6pC7uu67ts6WpUc6xQp7+D77ThQWrVC0z7eqAqJFuvqWDHLIH
LdW8deUZIIk5kLHnuBlQFYw0f/qM9l1/N+/b0SQzNlyzmh9PFVWsA6Xfa4YzYJqolqOdxPvYLDiX
oTcdyMP6O33dxyWjFpSI5Xzeez5pGvcpPFq8YfruDjfE9JxVY6EjHdsWUzusSAT9khl/+CugpSSV
UP0qN2xYjdoPk1lJW3xSoCKgWOQ8m5DEWfTv5VV362FcTeg/cGo5yrDRtd1azuG68qCkMqq2DKSz
TIPxBpgpKs1eB0KEKmLjNb/M3F/UQ5WMX4yFbIYnarvJt7k74b3L1FXjU9zOnhdOC5XDzoUjp7VY
T0DwO7UJFqcBfXZ692M9ifwQvVMZbpLsKzrnAacrqLp0ESPWtZwcLDRmMeqnMPeXQM5r8UDa9VYS
igSk4Hc93/iSJxvy2yl4t50PeKiSXf15P8kxlTBtX802xx5IHLyvb8cgaZThL5sskRblaldpaQ4W
se94Z3TylpviztUqKtBdLuTy2yF3X6wvJcl+2f4Chm7xDk7TdBr3pVnsk0z65bAhy07pz5VtdQS8
vXMmTUZQWgiMCRsu8Sc3yT5B1Qc3BZRNz8+mbuAQwBKPllwWTssLcX1lf1Ha1oT8UklC/aykENI6
BpexLMqMxEK3oyMfPu6Gar84/FIgNp1RkZfKMUO70dTPIYZ2VegzSM386ZIEHBKrQeD3fovt7y/R
rG7UXeGOaFQFgVh0LCH5CFxQ5NGwUPh/1ra8aT3yjDSWXVny5YZnZaEmco+1HB0owqwUZ/vVQEqS
v5ZuEZnEOYYouqVmMfh2nXcFmY4R00RXmJ+Srj2cQAmrQJ4/1E58TjwP/Fg8A8KGtPBhhzlFqwxy
IF8lWMVBQupUHivmgwApeaj/wwg+T1+hjCOwsmqrNTJidq/0u12/VJwkSZ2bN33bVZth+C+DZsDY
VtVdT9WAuGbqgTcERCP7R7bqBWOuYt4GhSRnlA5YuGXw14wVwFSF55hlh5gANoBmPCTtMLiBYmMM
IB3D7jZSCb9RHpF0nZIxSLd9rv6CmWof7N2QYNPxRNRFObDe3ed6KAvSTWww5uRfBAiJEcPNpsXM
pV19D3CgHwsxi5FL5lu7rwzvpl1D4rQrSMcmdTP6LrzEjcgMCuTXGXMh6IlaJ1BKPUwpdqNgtiIT
95TKo0x1vuFKUhwApaMLTY5wqm7A87B3aEfrFa3yO2PYqcty29XqI6Whhd85qCpQbTLN4VcsN8JI
Wn7cE55mbKTbYBSSW9fi9lhAV8BxjkvPiCa+le5HPxAKRt9LqWkQay/m/mZxJDtO+I4Dc4T3qfVe
pt48vlF6xOFrMksBxrIurUumGdE1PL+Jf5oWzQixBzUnt8tYiKaiYcpKX6kiVtwAKAV5zQw0A40v
JHZczhDgFndLqmTioJF6NCYPf03LSRAjpPmG+Se1ic/Aib3avLrfoOAQxPO3KdC4SaIBAElIDeL9
tJBg8nJRSzQvz2EEU2bqXDauB/UI9le1WXE6qgyfVAefg0cgC4CCdWvNppXSVZdGHDR4Di9MzL2R
wUCPZDeNxPWMbefoLJYs2ZJajmU34Jeve9FjnMRXqVq2ADXZdrftDS4sriuxXs+qAHG1zT1rJ/4d
6WjkJwKbyjc8YySGAeTaAV0xqXz6AIMR3xJMyBheEp6ajZ5blJkHbiVkIcBSwrzfr1nZVrDq2/dg
qIbxB6XbIToOzC3KPQaYizUArl0iwnehJZIzXEus1essh70Qj3huFIC6tQ+1RFkXB+mo6I4e1R81
ZQtPDf+wQsklmoKYEF5NLK1j/yKWf2Xh1Yy7LlXHVbKJNXfcOXxGUXKc4jAp0Fk7HDzTjm8AsrYQ
aQNw8KlTX3LSX+sYmWDJz6vvLnyZgdfaRPOrbirxql6hV/KS6i3NySfjN+3TwmEzk5mtBbuhaQ9c
1wu36HERMSuZKkcxBbhxjBCBDqTPm802C3bzJ8G1qvkDYEq2eOAgSGM4r+PfURUD0SRFl7qjjQ4d
igHETUCpH5Oksw+G+WQUYjhd9d7D39Hvj2o8v2+X6E3ErMVtHhoOdW7VYS7puzMoC+7/yoB014vN
xfPS9/jZDsZS2Fkz7ArxOMOOD97EsnMjUu+tZTYv7xGXoZfJmK5Nu/RkarfPC21jVx5XiHNIPTfU
mspRFFZsyvSG/T3AjJBSI6mvAJipzs2FtWkgam1haX/Gm7d+7Cd4sMkNiuLwo3qmLUvR4nEwB/8f
2aLdxmi9SZhyfPDurDfMugzbYsu/jzAuCh16mZ51i0lFrNxOlLmJD8FxgIoZPWbkZxaB/nan08IN
iW1HJqhsCTX28j/c5yVYLsCWKTeLfHNZHQP/VxzU7zmNgHOAQQMcUuwJ1ljst2SHrvTZah+tLBcA
aiIy91XsEkdaq8C9QlaZEqQUy8PFfVvQLIQWTmbM2advfsqRf/mPeYHmFFedu0EppD9791CHZo0X
hhFVF+q4UyFlVTi8GPIp5u4QmUWQHB/gfUaaLUNik29k7hsw6pKplQS23VEBdW7FzOBXFhsp+Br8
OLJrnqUebTd2bY0nXqFtr5wa6lEeCTeT/XJu3vwMUOxJL4aVSVw/LBFW6k6uQozAfS5tdGd5K37V
jJRTNTuDIvjsobs2bRHefUYO8WRapw9KidElS2FiQEP8J85jeQqD6EnU/2ep7Guni4hETZCiZjrN
175tKT2IWKZdHwb8WL7DKQ7mOK2hZVkeYDQDgQvcg3t39H/pWSfpPJERYmm/VivJAHXMETHSCl40
QLfrg39+uxUEKy79rwQ7eXXVGgpORUfH6Z0G/LaRMFTuDyqMJKXI13Oyyiq09GPmESHmKhbylxOI
t81ge3L8NaqZ4WPCRccxZYv+x+9S2DeeQqPVse6hyVcLek0QCsAJXfsniAWBFl7so+O7zd1KLy1x
kpq2dtbrpowDIu3Hy3+g002jVRjnHE3qKHx4HVtxu+5+EteTy2PAroX4lgXTEjE+TPuUGnL5iFph
Gxxpa9on9aNipsu+lT0ocpeLZvhkNpR+1dMFpGqEjMfA4ri4veg3g0Cm9ekH5oJYXYnBROOH1YMi
lFxoA3kIYdt75hjuUnJ4sSQ8juycOmNHtk+1/9ADp4paBg27SiAP6c8LGsE7F92gjMl4U5Y/a/6y
CYjZnhuRSvttq2O4RldqM9YFbP/FCQ3lRqYSaPQRspu0bdC4gd4S7TW/yJQEqipjqtm7n72q/FMf
iS2fl5j6nrHQ5kDZpj3Awcsi4cR49b3qrvbABB/p+J71gfkKVq191B5+BhpHrqU0/ilqPKJKcWtU
i/0w6xil+RUXZR5LLBs0Mc1pzhue99apcGLWfn9Lj+8Z7YJODfRYKwOc0PoUJCot/3QuuO4TCay0
hYfGrYxVGErHfEbQAiuIgTeVNlyUlAFHvbiGIMeS/ynOr3RWCA37nsaA7sBf065QArvLvPVhvXDM
Yx8qGeKzuB9e/mnHL3NiUAS7J28MvwZ/U7u60Od48u/pgI3bAUZMx+M6p9hJKo/P1+eaPDBije6w
Ba3wf1FF7I3OqC3PZesBxQrufTb/bKHU1UY9oBDzTGLPdFv+CSlZ4mMXpG0/MCpgIMD8cXa++U/h
hTUvmWZkC9LnkET7puvSwv8SzfdW8mJhZV0a8Fg+CnzlcRuGfBlo9atKcWIv8RXlUSj8l+zer08o
y6NChRqLlDyARhVZXLaV0gtxzDIIwrcybC3cyQRxi1GzwZu5C3B8+7c6yUoOiY1egtEBJ4Qg3KAh
LO9ZgnKGj/8cXR6mbHKtiYF5wySrWIkdhjKzymuep9Q3E+1IkYbPqSj/EYGLkDec/vAAE3du292/
TemV8nQUsjzkl1cN4apSCPIPdMcsoQajnR629WCRjBJ4oT0uIZm6hkogczx+db7WeDKyp6/HZPQx
sCHyv4/+9BeGqgEVE3D8lVWNlRfta7cLVB+1hUUwpP0bGbiMHTGcBcdSMOzVKW5CMH//+9SlMJa+
/1on9z3WFZyakSUe1jo6edS0HErfu7yAYFDmK+vXmd2Z8goHVdPKaudcRlM9S7x0mZWsrNk4sUeF
BKQSNf+Xc1H6s/mQQO/H5Y8K+FljD0JFUwJLqKrn/3lBxH+hcLax/pUvh3XGSASz2ikqOolv9xfu
GMa1JcIB3jMTbCoEK4CnkdCpYKTFS3DvhN0v179I8xkFdaeyRiOuW33QDxuQP4x5VxyVCkGGvQF6
YOLBdvOaHbV1H8LbF66ElNDDmP6y1jyc8zoKSz7o0CASj4E2Me/AxkZJVTnkoiITv1zJIuldgrl9
kR+abQlN4Y83YSwqZqQEP4pZbilILbgu+GC4KFA7/ah2blaYQIHFm4BUsDA/pf5QBAGJUhORQN0n
Tttpp5omQoTKpCOMv9h2aIkQmwmsbNXbZAlxNr3IYiXlABG9MYS1fRL0ZCqwhsiEyianQOefen3i
uLqHRUfKNpW3XxFYF4FztaTkTKbFoP9BVACwaumtOW//lYZgZSSW3ABO/0OCjapqUrZKIjNARTCa
6zqGh1NL5xfOveDo5PKHY1/QOX0qiqKwbBu0LDLbUFvK29bFuVtXujqwjLur6NM7PMLD+qEtmjjo
M9eFd0CdfSzeDdaG7A/oUxhvTc0RMENPBd/kGgalMvX02B5TN95Ntlw+2lUVo/1pLx1ilxBvtuMS
VuX1Oilz6+YUVuDaedNK4E6n3QbnRN9fD9HB/+qSwdZirNAm9PudIxBLDpMDNZUQF/vKsrk19+2a
09ssROmj6jA+qr0Jobtclxm7L5j42lPpaqn32twBqR23epzD80MbpGT8C8Innwx4tjOh/K3g3M2Y
OmLVzwcNPjxSyYM+MTU+Dyiz1PyuYnOByDTg3Bjd/v8k/C9ctxmpQnTW1t8ibu7EIsdFjfJqZoTs
9K+mT7gucuhe6vWcmG5YOH48tsLk5pRrNZWVTYHhDs7q2cmbsM1QedRbm9ZwA8c9g7k3Ox6zSl/l
tbqTYcYsDLFhUZs6eHrCPF0rrhwDy+H7/JGsgWeJaJXEr4LZvuM7lY4hD6GAC22HGtBtSGiCewa9
O1Wq31t0lUvg5XgIyeL4Wg5C4AggBeFvvui0dyoomXPFKyEr+v/Q/252aiC7S3b5KjRDF9IyMRfh
muHxvx+QShCfLfGdvQvcyn05Twv5ucnDNNjBr87NSjKyO9IHcxflaoLIEgf0FIvzV+8FjXT4glax
Vzgxljldxn0ilSYGOY0h6CzlleWjEBh2WOkfY1TEKvKk62NoAueqJdqOJgZRmr8jKqE2SB69bWHN
ynK/84fmYfie9U57rFXMBWg6lZK23L/y7lZOzR6hj5wk/lJDCn2W+o3cl8XFwHXYEu7IOU7ZcKzH
LGzkqb88qwpiDjVbM4m/5KPCw2RRChWy4ZGuObXvCDRQV868sOFAS+XlI4HBYPoQTwcKKCzagnxN
ekjiwprBaTTIuv9P6Y+kzSDS9lxFaZOfPXLRQJdVFXFodQ+fzOZQztVtAso5ZGfutMxdLzVqbU3t
QEvJmLDqVfb8+Nf4y3zeNguuTzHio3RneVshTVolbZeUqj5josWncJLeE+ly9YW3qUBfH/ID/53C
OEie3yl97DtqIDwcEz1ge84Td3DwUECJz9dd51noCAzfxvt8yrsE2+n59VVg4B4/zp8icWWiAkIX
ZPCZx2fPgV0MPHpMu9Fa3ObKlmCCnCO7i8k7yIDv9jHkNJYfWpW7k1x0uqPCCgQw0R43SFM5yBkg
vCjk47UDfFRetLNVbRspoi1uL1hTJjAmE2XCAJbPsTlmkxByc7nrMb+AkxDQtruUmQcGmJ8SiEGo
4gkq0ex1/uP+IcXmoefBjsb2mjbKR9X1kUUEnH39Mmy4xkuRCUvQwgge6O7vVfA6Rjt1InZ8hYzn
pq80Svw1wpTW3oxL+E2q5gfSmhG5awlBpKFBH2zSRzqCRegth61uQoHSG/N/2M6sRLIjUOUYEphK
hwaqnJDuxqMSMc6GKAjau7sHk04Xzhb9ogx/Y62+l6fbTHvtU0EoNIHxvLVoBBh1W5gxxlcmopw9
k2EZZp8rar++35KMpIdoXcWHh7zn8uxjBqiUuhULqOUk40l4yKvVH3bp0tZNQpPSSR6dQdZxyAsE
8Kvda2WJ+sLyzDcZNRfjzmFbNuP+0BTrML04OJMvKnrSVhgvV4O440ttg6fFuKznNBVJK4LI2fuV
MmLWMOMJdCyjxmHZHgznsT9EZDf1mdUHeEpStEHBbaCjHrEV/Mzl6RGFEKEzi2ko6O7cIOKPHi4s
OvhtX1V8wqcyXxH54R0eViZwkGhR7WiHArE6DfMuvPZo2BQA3oTv4fAh+2O01D5YTkYpsZyMN5/T
ZLNvrRPYOWvU6/ouSHjX8RIMol0qs/G9T/IdU/BmWmpNNSJ25bxrf4FRtlie7VO/HSb+u4Z4wGtw
9maa+1GWnfsU8kNY7SN29AP6CmJIOcMRFisKYjbd7SJLgsXShRGUJCE7TlnHLdf14WwvP22OsKd1
aK2BHmVeIbEFcMPZanF6bi/Ud+OAONj3wM/BH8/5bK9wHNE/La4sLpwduvpHgR3gje3eKfS5oehO
lK2mn/x1IRHX5usDzsH5VeOSDlo/IMAwz7Kb3oYQenGH65+n4h/ungNK5q6pn1WNL6C6HrjZEtmZ
YeEvl8CVgkbZTxBmx7oZVR8hjMewy4yUB0aKPseb/9F/lEJC5eGQWsp7OMeH0TmXDj7Q/TRQCKSh
ufYr9wqlw9keWrQu9U/59D9+TJq9ep07FsgqYkJEFgrYbNdaLoRG/qAW2eQK853GC8+W0HUgQTLB
S4fqhi8zVhM838+MUxDsByfyEjM7/jLrFYhMuY7lol6GwNytBHePcG79OWtUARQ8gKldt2OXWEIO
a/EpkZ7H+ZxO9RBvrvJhbSyTIfpYYJ7pd4ySJpF1ZPh5dhxWTCXtezXhlYOT4JK1/tKGOGWFkXuQ
VAtJF3GdjImZzfa1+577sf5IMQKEI4QgSQDgOWNawDK+aihO18CkwOHOKuE9BPUKOQKF4ZlJJnUW
nTaWHIvxDG+DFoT2onEQt0vLNvFayx7RPHTkPTHLjW9LAbHhs8TQs6YkI2K1ZNRNc0XvV3suUIze
lTO/1WP8KVUDTq1Cr/GTJl4tDLqsdCzO+nfYucAaCKMhmAMIyTHJuXyRzwxupAryCDwqAEVpz0pn
m7pII8s1i1/h1MF/omDjCmy4pk22FbCx2fdNRePuKn1vZD6rxIxHNJKRYPSupQiJKgQYBbu2HTXs
FS4HyplylRNN6fImh/Oaz4ox+Kdo841yh9B/pYivx7buIfRLQliuAWAsIro9pDnhrkwvIWba7j6U
0ansJrlltVeCkLo6Z9hK1sJNG+XK20fB14WrOu8E797Y0JAg8rAH8UpSZPLsUIx8obPu2LttvMkq
Tk+NMRQz1yLZ0Qmdw7ChrU+IE5+AHxXopMmLzuaZigBly9DGZuDH65V6wvLD4VHAlEW8c7tgwWsQ
VuWd24mfraq7+aA7fftDY6BuYL7060nJrjDFjW/n/0AqRH9oxAwQw4x+6tS869asG+eChZuhlq8F
m+tZ8zk8kw3CFg0tKWo/nV9R+ZK3QrgahI+FOy5RvAoVOUXdFnUdT0WjbljWH9mBGeM6MDccv8q0
b9GHs8cbzR/CJm85+ISDC5baq+7VbJzzgk3/2+nBZTG5kKmV9snIpSEyn22pvrUFAo5hK21KFkuc
uuAA7zKxQlZWPbSOFi2x1ClpJiHGirIkXjFeQW8IRq/PbQJOF4PHXJgrc3mt5CK9IAO/2LSwhAbw
LtvHCMeVd3oH17gx+8IZfESxRu3A2g7fc+oejGnQWg+oNrzop2ANov1Ue2Q+oJfIssfjKmmt/Xfh
o2W3Oi55zz3sSXsR2cY8y/at8Wq+sRNis34vwLUgn9BsxJRrMQrCWej6Cbj7fMSNIabl6nFqGqdj
hBI0rQA8DYT8ZlCnOFUkWaVnR4db5g6wdDXRcpT2BMeOI5tVKXzkkeHQ8EslnZSbcUDzE5OeOljO
VJsIo0pxsZ4afpqzRHKuX2va3Q79tTSun//C7lXWeyLxKsaZtK+25SdAh8nDlSb1dnqRlKYyeHlh
ayTcgtrEogfSsTX3V0wOYcjE1SV1kPb+0Fi5k33pG+/rMnRG32B40K2zIrc4p8nqc53JHzFZcRgW
OHVPLus2hwdYp/1KoKGcoaqEg53NnyF17GFN+0j9hhmCeUtrGejnaZD6J36lYf5PFhQBGws/lVTW
UL9BfRETWtZc6PvWTZFDiNqod2qqwEZXMp9ufE4LUbFIRJtmlxu2ZpJexvXhrzOpB1uupZQaUq2g
9eaBhmwm9o0bvwTEYTfLhBOA5zFJGq8CWIq+7Wha60MstFJoMl+PR+icyJWDgWiMdru0ZSm84wT4
9X0V9hQH8w0MFMd8lQ1KF/i7a3s+xJhvK/wkRhnIYQh2ch/d1CltvcnSH8yCNNeah/U8dSpnPciP
dXgcU079Bij3HJTPp8IyNT3FMLxdA98+x8D9DZmnnd1SGCXxWhUhyIHEtqB/bby/mcQknno881bt
vnDLduFFVnToaMuxKjoMp8j/FtNMy6BdfXl/Vjg5LyPPg5DD2kET99s7srSrsb8eDoBOuTRintT/
UcyASSvqiPLtskdq9Vt531oq+mX+PFZCvoEijT785ayl2YB/37pom8E6ubn07mFGPD+4ZVZs0yfs
mOl1gEmhFZRdviltZBxTsVmWVdMQwd32EtHjIdjbhXmnhBl4KSej0W1LRAcz0ZNz5Mot9eGQcwoz
475yaYxu8KE8zQBC327Yk3wnT+6OeOFJF4N+cli4k89/kb4yxYfOgNGPh8epHardZ4mfAj65iilG
apYf/AgU54PYNWUBzkb4kOxZ+33OKl2IAtu2QpA8SDFaqNHAMM6cyV2vqr3xAjlYQ5/cVJPC8PLM
g0wUv/jLS8wGNfs4Fa9O+s6sRTkvLXxQkrzds6egMQPOK2aPqmXrDRpq82NzE8LbqFkyI0q9+Yet
qvV7/YEmYzpmKC3GK8CwhkSDNcLJQa52KbmdHoNhsTwyqwI96ZRvYis982V36YcXh1xBBZ2oDcR8
CiE7uXmfsIGMo9WFGEBofjLmnTK8D8wLwGtGnHc5a2jHJpcT9a4Kiaz+adz77/nF1OaiynaabJHD
xvGeE62fE4YnVitSIB09zB8o5uAcGM832YwRw/fodn4j7kEXmFnPQHTTLiVZuUftKngSZ3zcKCgt
jzofni+T6r/8LjXVGXkmLiGUswUw1c4q9LgEXVqvm4ZwyC+BhBn0Uj0iJ94JFqtzJQ8irwhjOHgH
qqC+59PiwQstkrM7UoWRvI1Ro1J8YIYSkTFqM89nsTfFsjMV9thHRvZvNsG8jxIAP8suQ68RrAil
0riVin14swJ6lxeFxq7b9yk3cc0/xPe4Khn4mxqcq0i3eNTra8FRvx8L9vk+V3n6CO1/ORaIJMpn
apsDvf5u/9uN1rY+a9t9BQjob/t7XdeZEOQHi8UK9QYlahlGPTMm62hwuENQBKiGjdNpI0pOjl70
OWI7EV7u6CV7nLffDG8EPanSmpovqhQpJPgSRxnPr2Zbda+ug238IwR8pxp448vnurZvLeJ6NHv6
6lkjTd62jgLG5gSJfLXF5b7AbfFVbbF3PZ0gYT9pouSjG6/ZYJlnb8A4r2K5RgEzl/MSVlYogP9d
SmbBflfRhLI+eaWXlTdZDvn1j09LzV/WvGOUuYXLbpmebdPD+rA1YiM/2ruffiVFTKRDPVUSa32b
7exb6pZV4wUtMleB9mKP1UHxI/wsaag/W6RXPp2qqUcu7szGAJPSeo5+lAee9tRphhssOMAIdSNR
T0pSOmYAU2FOY5kIPiqk4fyQJs0ZlMAD1TDQ+USosB4gd4QFPbGUWCSD9tFjpsMjcTgRfW0gbqUu
fOnPE1fdRDm+zwKYnTV7K/v1VGUCXBiI9gygZoIox8gYrRUey02tLe7hXKcOhVz8XQ5uOn6uwlIx
yXcCfAwC6v/lCNevIg0w4tJfroF7bPnUP5oo+vqEWfRJVxNOWbFzvy/IGXcgdezD1kjCAH6PTR1C
nwSx/5HzbtpUjppZsmOqVcY2yVGA+E1hwyCZ7Me3ej2TfKC9d6CCDXMRy7Ly6ZAumqy2rz9u9VXg
mYJiDUu+AJ+5wswm8ItPeypWW0XJdyFYyIBMwQ3A9L3wmh60s6srAWxTCFwPt/9+LhdfDkgD+roT
1VMGkZ9rr15Y3aXIyrcxertIU/upxuYxep5WVBXnuJ30mhREfpHkIqOEiwNqMEMZ0De8QHCVJ+DN
7iumyAn92xBB5Vhf6WIh0j5ACjpHq2dN19JlfzbTOsfwFrlEqoCtFxpaY97P/SLjri/V6R+TsXOH
bsQKKc2X/61Kr4L5ZvM5ADHh229+q5D6w72I8297xdqQykAe9gvMdmtFNt3bAehBdqt8KA97jQ0s
EQdAQvDljDLmLMayAYxFvzjcTLJPK44QMebkpspP9pX35MjR0Fmpxh2ttbXTBtTBGadQ7sPSWOBN
z/Jhor1AQ8beMvcoWJGAG+fGb6Q1s0pYGE7pP5S5pVcXLhqnR+MYvN4DNk8Zl1IKrshF2zgv2v+V
Hw0xBlrJpp5wkTAVFzmk3BHJsz48L6PN2EvkSHNn/V3IcRYhrF91PIB6DyBSR/KJk3TDcEl6TIU3
92dpv4/L8bi24H0SjFw8AuPb9So/IKOHPsoYWAAybs5M3MyBFCsT5Zo4P7/gG38Iaa0guzGUuDmk
Hk3U8/w/1hBgHvuMvRHZIJShGxJABcN1RzeUPnjXQ+MkiHi4e82Xz5PEA0PlNRZys4qW5tHNhkEx
f63XyIFbZuhorwukKxOm5ik4m+oEAnOTaEPJjEhohfPnYx5rzTB01QRt9zvGAbRXxMat9tm9eDnQ
wpXtN57x8MynpAN0LmlySvm78Wx+nGXSSvRimzBrGg9mNTnrXogOkkETQs8vg090Swn20iG37NlN
biMpwDB2XICF1PjpQ2FkGwuuO9M0NvjgR10hD6AoaffLqfuWbkyOvjEmJhV01JoYvLNjGxO9D57F
NwmI6FEbR/iGJAwhiVkqOiAJAAamg1cPvIf1mvUuYDt+An8GGySsfOC+maL7vpzDXjOOoeKgT0/W
t8fEmuE+khhtwxgQsaZnzYDSQ0UsrWPnuxEzhbnZg2qnHdtQbGw8bo3fCgQ1HTEdmBd7qvq5yYkC
XdvUjpNMn/typqFxrVvNrB9ZYGsgJfkyVB2wHMPECXbA5kR0+1BCB8nEgyn5XetCDwjzAKmohkt+
hnuOuNlJVd8wyRSSvZg2lllqaCvct2G3zdvqsDvyw9pex7HnWRImZx9XwPgt96112Aze8K7uE2z+
rUcYWJKw+3eZlOSYJnuKyS4hWBk5t/0JHN5ji1TiOvhbOS9KFESAiyEEabFLyg/DVwlcb0H+jvii
EjyiMHa3hMBeKF4FmHaiCwBhBMmwV0Mh2GGlfE/IezLWmm2ugBOA2GOLoVWe20K5668c1pcOkg7T
IA64jXiBD8iMKQAf8JIukzBwKCnVn2PYcqgFw/7IDePe8biEhSvOeG/UwqTEbEQM6CfIJg2r8p59
iKls/LDgJO92hqEKVHwBR9dw+AR/ncIAPZk34aYiB4sCxzJhAvFf3r91asclhy5zmNC4RRPQJOGl
OVlSo/9PfAkn/qiRmqqAJQxmxKi1tupKBgHBIbz4imlirxoaLWXQ4DvTvFt9KbARNh2RTazcFdXk
hf+p1VNG767kawwoHvWvv4zvBppe4UMHbslNJen45BdVCMDBtlljGYE+Wy+U4MSs5UZYCZRE6mkl
bvaOD0c3q+i4KB67PPWFbYlglPKs/BHfP2a8pszbloHtEkpPfsso8SYALaHP2NswVKM8knzxsRE8
6vqKhrWrWo+0FaXUaBB998B5pfGCn6B5/Xadp1f8SfCh4+2PkCILvamZk9kwSvdAVI6UcXiEtzJu
+q8mmsxb3UaaA7g47gCjT6fnmpZa6CSiIEy73TXreGQmhVM0b0ss6JBh60nYWkZMsPHEMvgIrn/d
M/jX58STo2x1dBIN8Fj/06zesot+k2kbHTYB9Wzjv4PhSKfLG4fjQVUO14XKWu2M7misT3EazzZc
UFejnzpE4PwapBw8WEpqAQp2e6F97kOVRgDoN1XjaxGSBayS9h2YHADV4ZwlJ6PMSWOvSVnmo6Ks
jf4Pc0guG37aC4aW+CAb8rjrxe9GCiElmplFmJuPkp0NRpQQEGaO0Qy2qzQgI41vxC96J3CF2wI8
VufLT4diW5SvcaqstTx4k/K5Qe/rNJ+HIcfIclQ7fqesu+4h8BvvBKzygW4qbjeDjSwaOCoMdmem
Ldp1RadQCRLaEA4L9v2kuZQmcwItoc+PQ6E5oRWycaGgAXgGOoim6r1IrSmCAzGbHctqX5dkwCW0
VgBJKI1nAdfQbAwg+0uVhMgIzYBIQ/B3c9Udu/qcGSAh2BnXfxvzp9U2FnNJCBx0/Dza3XjnvEnM
QEjzvtpqxjcGxkdBOt3/sRwxYGrKYiWJD9RDdedj7vc6uv3TlYW7a1NrWXfRLgEPO337gxGC1LdV
tNNi73smRvyRVwHQTavRTBIuYcZrPlrPPvEvPYvo9C4NLi0lUmQwSWo+gVkhrHAKuDBTT6pHwqcA
bKvlyhhaBLvF5xW4yWdH7nDif331mJxmpix4ZWhi6UK+q9mwCl+uO4Aniy6DRDrUYm9S2sbNBDS8
qmfqSyKF2w5egMtzaSSXam3TgMxzOPupo061LFcVkJiTCJHQjOebs8MqnWp/vbTkz75+NlhKUzdI
J6W/3BiCaSS9TwOK1mOh5hy6SQO5ci5XNJ2zlEnoVjusP3fp2+5y94m0ZQ+xOhFAP6Q0ndKc4UuS
bWK0LYd0vZPxUGsBZ7ZeDHTON9BbOMHEryH+DCecEIqfZq+zc5PNpF6g7a8k203mtQhzfXQRrFlZ
jut+4BrTU05ep/uMjqeGFc2WAPQx3iPhMQagwhUHeQqFS79RXAMAX0et1sU9uoFpGyPCb3xnD4fi
DXkEE3coh9nWYsnZfjrdKuNG5s37CDi56qp1uEGKZ1WbRSS6mAa8Pa8FOvk7mffS4wYMCCHVB2iH
ZPGRC2QfMH12Xv3tHQp3e1MwYTs2LzKdOa+1XMzCuiRf46h7YMVwtyHE/ayFEpDQChSUcWjD2YbP
dsue555dXlFdjQ3bySP9hNaVIa0avCA244n+YpOVLjhOIzmMRzsfcqTfYHOzxeWskSIdvtP5zGdj
XNzxjtjBDlVsSmZDLub9zJEEZq2J9/Vvddh24niyrSb8MxarNOZ07cfAhmRNGtJikWH5wsWg/cNv
BPGVxn6GpWHJRghkI4dtC/HNXGrkUEWBmBb1x+9TjYeDnHMj+dGuOn4LSAcfuR7ohIoiTo1m65pA
/NJR4r1Ah9y0UayoWybWGdWwF6XWlQVuTTVnr+WS3LWhuwp+hQ7IsnvS2mXvSD1rAX5/zxQ1WqJk
3nsrsHZpCWcjOdga250zJUrkHiu14ARrrfIuAAnUXE/6RBpkR8g3cAtrG8rc9gweClmY5LOyxJ3u
jViGxFnSZ37iWB2FIbyKxK+LUeq0SoBlvqzbORuaMH2AxrhpnJlqOcWrEwICV+Y5LarAQ1w6c9mr
twgBCzaEqWGitty0wDBYFmcsBIByNrBoU+Q2ZihImM37d3tae6PWYPzlQ0yTTIsdj784fHFe0Tgr
lg6iE+8/arLqQ0jE2VU1Uwoj85M8MSOIJJxZdApQQv5tRFzUWnfccg/Brsr7Rm/0gJtJCiLwbimW
JSO25cJeb/YNVquo62j4edQdKFnFRnPeubWGQ8mnNXVj/nTZkRI3Azjj+gREmtPBVEDyte+skB2j
EWX45n2A+Y+AU6fS97mTTGAGLZ4f9PiaHhwLVbf2wbOg6j65A2qsmqRLdHutxtDTmnjIRrgHGz5v
dPtRPAm0+UMn7QmmWcnh/8Tqovb8O4xGXAIXqEMgZ7unMvWEpIdbWSSu0dSDoG7158gquH9Yuxgh
E/MuC6PWZZyl/uHFinfk+Gr1o7V5l2KVqvLwdwq0DCicL1bAFcj0Gh16uPDomdMQpFCC2cpvEEcw
swCejCg65fVMXddzcT87reWbdNfdD3V25d29pwv8/JsMOHATWRXFKLS079IPzNCv3q8fAS6pb8pD
5gIsvP4RMV+jUZt9p3N20KUHMJc5Ah73M4ckELudRj/m/aey3hRtbH7Qbyxlz1YOP+SYE+FEVwR6
ml771TobhfFBflpTOSD9qke6hF0B0tw0FAtzSjjRua1ELI/fvwczQypW9zntGJTstMWtCECr2vuZ
sWwmYQqeV2VVCN5xKnQBUVR7eTPXRSDdQKIUPUXpMLBxGqbIUA9UeVbPGdXJB/yC5aWEvmrAZ6rY
X1ZPbjVyhvIHejxjLPPO8hJYtxMJlI3NO7bli7Txt304BmmzMbNUq6CsWfhBfqzINXr+Z7Dpux8y
FPSZzLc/fo7Fr1t9k78IAfHclQRTn4HBWpK/4gFoe9zH3kiiJMwe175jY6ECriCFPoUh2CzoSNq4
vResWAyhztKyy9sH7p3KZtOzbA/yg0y1o+iraywQndgaIr7DA0yNkAp7dY15jhe3t1dRHYdP2oXe
DLYEIloriXAd1EziKZL93cBIjNT77fZetMvyEs/wNEacLIjXfdhG4byN2YvHkLX107Aec7NOMdML
79ad8U8G37TGLkbgpBtmFxl91N24RJ6+QOpMZ81vYmVrHM6gvoXSyKYo2YEG2/oI9TJkGUQl35Hq
q0n33nUk97t14E51uSQ59bFXvKI3e2/Gt1eEtZjTkYmBccji94rBBecVEwPSOwv5NrXanOSIvDq5
b8NNLAzFk0Iizpayr3V/zkqzyCXLHbHZJ87MzcXPseuvdMJ4DdPNOsN6g33ZAnVJ7h/vrAM4oTgQ
a7/zr0DwPnUavSGZsO7UsK6iifL/AkptlbyAAzk5ZT6D7s6GO1+zsAB8It7Zifhj3T++qgYHIvSj
hxCU8TuJWZn/1JtaTBl1bZF1fEQFlMdfP0aBJyxJCbdo7vz25wYjs6x8anc/TYMxo7WnKacEfOyq
RDEmXjwMDY5oKpYhW/5qVpjv5taOYyc9lQEnsJIPCqCn9ramw+Xwllapca+OWm647o6K5P+XXJnI
DlChwubfVaa5Vv4b0LXgTYhZ2zDRupuj6ylnZub5QruX2ebQQ1fRO7coEs/FJkE+X0yX/fBYFTRN
RWNpEH5YK3VxdISlcZYXjGQbhqmYwy/tLHph/SFoGCvJpi43jgOlvtuPLEzvrTOsEPqTbRMv4Vjf
uqQ+hnyLGi6FzEU+komZj1bJbPabbTxYQa3kd1UItCP6o3O2UZJsx+uGlYio7X3eF5yVQxaMz2Pq
bD3WOBvevgklPLNOtlB5+AKjwjO2nECOkzHT3x0U9nvSt2nWeehsDEc6jJdceSJAi+0NfyIOnSTf
xrrXnlopBVoJPz8rtDr1OZxdY4GeuyO5AAg38+/BiLVqL13DPxxgHM9jRPJMVKS/r/yBjLDwX2gR
NTpyObgigupyRlUAnotuyKMGaQUvs0ykvBMMxlVPajG/cnmfVXjWxi4STVy18IVy+8ZFnmZyZARx
aR+WQfvmiqlrYmat00Wfm1V6qFl73trY1YflZ79QnWCn/WArkud8u0rdjr+SPDBkb1km8cK64aBl
1ctTOomzai3oza0Jl1n0+hZ+65LhHwXAP13Y+vabmtq6NVSJ5HX/L5rkPByADz7/FpU2XEIh9lnD
1DUXOuqPsrjnUIUMwFngsmVHPrcRn3Z1lcTgKEolrL1Iwe+cRptBDdHhwjYJkKdmAz5r+VWLijbw
ci6jCXvHVvaJM0rD05v5KWpm6bq1cmGiTU/Ul+pYP81+zjvdAKWmqfTHiY1UUPw5Wz0xUxA1kk1p
RhO/2PWhsPL6ywUbxYgxjOWkAwyAdniElnbS5Qvzq1aMflSj9LEGMz+WUi9TXJEf8siPY3pJrwpi
sOO585ZacXiVW2nk2CtwoCFRZzCQeZsg9lg8/FQt9LE1aXkI8fqE5daRpRNXtp+gXjEzCVsp7GOt
KUw/LMlotOMBQnk4JLqYnxXfJec0PvG+zqfWN10QPWrnaDaQu7zGWEblQBojywTycA6eyJWOhdnr
pAIu4Rr0R8LMz6W3UtO7QN1Rb+km43u4Hrgz0tZOnQUT7a5KdqbwGt7zNjkYHNMdi8lFXr4iiUxV
Yj/wbwnMAfWQdsV9xCfjcM7kkRxVSuWlnZTt+/rUC16lEr9hwLiuJMEirHzfJwQCDQvgYLEbUqmk
4txPeTVg9FpgEOY81AIO9vMi9Vu8OQYBiwkNAZLEBNcyDlGDcBUnaLsAneBCui2kGrzkfMfLJcH3
Br501heBSKieZUjp7nYTJRI0oC7vy7vuNkyOBpLVrJfp10K0KG6RdozNd7fE5LUlrvTQmo8+j3TE
dYgu3+ImCmi42bLd/Gcm6ZMO9lGTHYbk6ak0cxOV8x+G6mcXbwrsPjnYiLnV09PgcUuvwWaHdVpd
iY5UAIpTb94jEegDkQgZqD+ReLzNWLmCfsNf/iAuOKSbg/DnwnDkXXRbhZFVdi5iP4eWhHvJk86s
KfhAEK575UYpUnagyYB49C/OObqinrKtFJ7h5b54w665YWFu6HTUp7+ABDyAZ0V6yPh02lWfCbwG
8zwVpsGyGXOrTmNLkfL37ukszq1tckPKpS5TuHfB3TMHl9YdNld2Bkzj/KGzWhTZLk+XvhgOCuum
WR5ZbW+xG6in981QimIknX0MdXvSeTrbXDzXKSiGrxGOqKdUkd/rLkok/o7csxug42w8l5xGT3qo
NC7XGkzXHWMp3nw7YSuvUKngABy/Qcl4dWzt8woU4aodxiCCPMVoX2f44mc0IC3jpKJa26q9yHWu
YS0MHUfFuArZ3+8SL2tw66xQJsZe1fMDEs94+LpdHPLegLLMYE7ZtvMXltE36eEqXYy9W0SJ9anP
BW9n9zBNFsSunhzbN7xGIrSV8cv/6WvFTqaw70RwRNRvLHFQeoxU5bkLnaVtdar+lVaGgl/wREDe
aKambV0JKtpLTDTPC5okoOb3xBBszqrjY5z1kKXcS/3KxdQf1xv1+puZ2UIwnURUIcpN5vH7ZSYV
V90OPv4SHQ4DzkPlGrIPzQQPakcjreIIx70OqtgDUv4C0JaM5hz52CXFP/ETu21H6OcZGBAP3MIS
qWio4z2psFRk9vxAox5ccTaikCsiqlfrQXJXlDCuMXPPE29RW7Tg+WBe9Fo5klrndmxK4yVqhmkJ
uVvVYixhSmp27n6XsgU4E6mCywHJfVV2GAcDVuJcF547Nu3Iqh9stxanphql06GgJMAJiEZSsAql
GjDI19hx5thF6ehw54Zs6qYlQNeeUUCQSd5kKfJTU8Pa7Fe4bnQftyLeHjH++ryRhZgPiDVjIep9
vq27NGKfDLwgqFy2Wil9PWI3hI22wxHL0kZefZrwDNOC6onoUcOF0JkhvxdSZcy8GNALFmODQZ+c
4YOrFVUbf6nCX46nuFAmPq/Yrcyg30UF5hI8nv+umsV/x0d6r+J67hqKACWxWpaZTjfRCptyhXGQ
NslvcIiUUIoi9uoxBN8o7YfIsXzC4WxpGsRLRuwN64/KhYb8UETIk2nTp43KY83eiMJxbgR+Fn27
QmgGNoIlGo+zOkdmKcBtJj27YnYd8MIedA32TO3dh9rm1zTfrR1XeCnCMPM4ivxs5e/i/HCtZ5cV
kzHwUaALI1luvCbUNWY54e/uFopqg9pB1A8QwerRIi0MAld6QY2fGYWn/hzUcWj/AmYMjXyZrB/n
mTI9SgQcLzPi6P+bOX3zbACFB+2GDkGdohAPjELC4aL/vlGD1YgFRD5Y1L3IbZb38sipX3qAMmok
wnr/nUXSv9pM+iR+Mik2VQ0KrjpAN4l0sTkbfqIvrFP+CC77rMVtkDRAaCtvMzLrZp3n924J9Vyt
YJeDFAneAGhIQi3EC2MrYJdvEXxe55gYr9aQhtzmJeT0wXD1QlRoTlJGkrRtlJEpgTHJHNfe1BqP
ZmlKXJb5gj4o7nPwCDhsLJiM9QnAw3F29LiELx/e/ByeSeAATlNwO7grEAFlpOaVxiabr1vgi0z2
EFModNAWlEB33iOZYRHY+nyLICawNfp6udemyQG8NlgQPGSoBCa7dXmF6fUT6NYDhRMBfglBGQuv
D85JwCs7J+I4KCfQcbhS34KrnC9P7INXi7tQbU9v2TRiLcJGonrHfOoxUL5GFdbT2CAZv25qlR2X
gAt8g0jzS5KNWS6F28wdLlZhtCovxKEvVaQTHBy2lBYq8Ji02tRc+TA/BKh4m9RdxADnz2yBBa+0
pgOOlXJv2WLyDW00K4q5DbNtLf+6WYe4m4FeDNZrZRPji++1o7lut1gTZ0FMx3JVgaebjnUt6fPr
aBZHy2aOqiRs7hXwgbDH0Nr2PjfBg9JYbume3HkKA6XoEIx+H1IMByn46yVB5aACkoxHfpudAcNu
I5fnbA8BqtIpDdfwI3iE51PdKdKlgZlxjAPjNM8wHVGG02nOLYknmczNSGDR3FwiI3CHeH3z1Mtl
fugEg4SLdTFMaGi8zlzrJERPeRAOOpwHYHXMnT8xI0+U7Yp7aNyqGj4xIzA7JSubo6WwqeXKl7X2
HP9QTzy1bKCWWxAIgqxpRP4EyP5FGcm8nIzQPBZGvKmErYRUh/fbXc7NivVsD0oh3tuG49jsQbgg
zM6JEbeoCzJVsIVP9mcFgzCVh8V8dpj3RCRG6DJi3JVaoMptdS2cq0qGiZkVkSn0gxiA+Qian3rI
z9mcWxMBSripjlz0l5tdZOPBC41jL7czjyTyw/FiOGNPNLSiqQJARW+xwjrwmm/Fp5nKy15tkFwK
mJR9CUc8LQlorur/h4MsWEXIYhnXmAVP3mCgxSErfoRp0W2/rb1RXhkBTDmiq4/PMXGnq9dqn2V7
HTKRbI6Qbpn0JY8YhOSDwJEsHan7HtYHmul4JTZNcaM15S0hpNyW49m5HWAf+PngemS472Sacy8z
sTYGQOwrHYBXqNV+7A0Y6TRCKjGrmVf5972XuyMJ4Bv/POh2617sslmk7Hi1dMfysnOCWclzTryT
Ig0VvozEEPEVOpbOYpp0+frsMMwfqlkoEuXtk0L1mey3qAXj/j/g7gfpfqT3r10eWf2REEfzJSYC
qod0b1DQxRqXYvsq6Y5moEj/fqTksfDkdERQhhpQGon5SaMOFWdwJN8WDoAH7a7ZYljdaf0D55HF
MK1Wu1MQ6vvvovW+0RMt2x3kIe2P8ZCIjFGMwZ24C7XBr5e05MqydX1pYA8ahOsqQfpGsSYoCpwr
AwXNIgXdqwuC4s2vzI5gw8oQ625wtn/Gg3W44GwctE0x79jbufo93jw9wlmn4fumQt1jdzYnbdIS
qbfjAzzkRsB0P/MgXsk33np0D2AaXICYQBDjCdFq/8vnWJqUFP8wgLQZf8VKYMqg824yVys3dipI
sSHtP8V6KbJWPdqxp6UAs/Z6W5jj+vr23mVKtT7rdwbNqaQdeQcJ4sGGWwM35oKE/MMEx9FVUp5z
D3OWDJTM4yfkimovwv5FvRPl9l+rcV10r5z+l8L3D9UvoGGDej9zurW9LLBACFCzetYuUCGkFjV8
TNxcrTYF3PLb6TS2IEDlM5fjJHg0qV3e0PReoUHf2DBltRIjWHg8XpBev2dTla/Ebn+ksTVVZHP8
kDHIwdl6bK19WJi/EoKKtBSQdllTpoDEF9CaTT+jsTci+d9EVt+V3D7oMmq7UCOo5EBmygVulfrk
JtXttyeogOPjSEPwtvQmDSWxrzNKegVLa/nxYaodpqXYjWqcoI1bJ2WPdlLAjA3PppXfxBrPyw5E
JotPNDWXHUEFUvkzTJjysc+M4J9O4jeVQD+u9awUGms3daQaoYzFr7oalYLHF7JUdJkSpkf89UMY
/WRAf4apd2oSLuzW5BoOLiMKYi9qEO3WdCxkKqTd/q8H2DSg8NfCpGRG6EOOuOrvhnNb4qbJcFYI
bqUBjT6VZNIVO1/RM1fI9xZI8K3LwFT1QwfUZfKW+OeH19Su4E0njn/OdU6y8c8sVlVXcYJsfFMA
tMtBSdNZi7rmODHI5tjOatvxSsECwGpUHASFiqJfdKnOEC+OaLGI2JYH3so/tAieKDS+q0AxBhbE
ajsvaYtpbepXLYDqB13ZcVmFuTNC9Txmk2aT3e5FS5zjhxbA1o2nZQpKiB9tQLS9bc1lJ/J+KaCH
soA+YAaOAfs2lBWwEjXPsByofHP8XXxBgm5OyBF4y4Ofifdp6MS39Z6TlZhejwldma4c4lLCevdZ
1wVN2UTtp3IZRxvxe4XptphFfxqcPKO5c4Xxq6VfJzmUxNP95nZCTANd7jP8s7P776XNNPWB9cgO
qLy5++xUrm5qwm2Gm8Ieg/Mwtm0STj9rSxiYT2W46R8UMh2NHgz75+ViASw2G+UpH7bAcA4o0TDv
2ehZuxev7RB4qo1Oze4Pu7Dj/3A3euwedVlKRyIj2wMmd5O8CCAfln19lPFP5xqczjAwnGuVB35H
OQHqKhMxJgXT/PlI9nQmcjDfPuIvfISrK/Oul7M93NKpvRKoUQSBEZ+T4r9DsmdZd+LgewUhQi1A
uitOgHFDFQhmamzn1xiy0RJrPGbc72WqDJN600QMqmzYfT0suDaBsK/D0Vba0ntgBNchg+F+XAS3
1OTRZyGOI8wUcltPRhM/UV5+z3FieVpA6goJTpl3EiIgzIgSknecM3npeCotyzXL7iaKSxaVWFmE
9Dq4w6atzzi1yUpyjTS81wM3H1GMVUUqPx7z+vRTMgZz3HXpBV1kzlk5gsIfB0y7nthRkcOOrfES
aYc8rG8vu2G4m1/H0xX5Blb0CA6F8QGZOV52AbeYXQxLaUwVR2grP7MmvLduPjNHdB1zgxMUMYj9
8D5RlOwa8mi7nNtW2LzwGx992DNXGXQRlCGV08rAzc2skNLhuiKnqI1g66xMhFDtb9H8gyC7+F26
da+KSfUayZeV420DzGQRN7BvCiOkDQYWn7mzNTGEzkWdHDqKZ5eOs/bd+lhLqoIJZPHz38CGl5eM
XGehkiK8WtLtL02NZh73ixKr4Z9MRIP7VVObjqfuhwikZOEHfOc9NeRqovhVB5Yt6U4gkG+bnPLd
ki1mvxDkSErVUIOFDB3h4/Cbsh0OO4ph3JB32q9KFpQT1LGiikcSxJh+aB+fihXVpCP9rxq505df
Qwa8Ha3RtjgeduAK4hYj3GXpAOqODp6CrxkdR3IcSxYhkiUITK84kZuvfC25dar8KO3V3kOn2szT
55N1xzvSlgLiHsJ06TBbrqAImwVCcoirvBFKi8qkFlD/ZqrmvkJrMzHJBMY7QO96xccTctuvGGef
sjvwYla60iLx37qUEe2c6Dnm7r+16kzSj23hOJfkQeQhA9PPwrdfn/tfarlJVFPqQ2PClpj71VEK
lUbMVe5tJlWm0WOYHogTh/P1ozFw0tHUOk6tqmaj3HnRzg9UCzPNWVzOctwfQrsWzqqd3OOsW0vt
3d25AVgykPcfTfIEMliqOKY1sDC1tnuzcgt7P9JV4dYDIHGXYSI3KAV8M+zf2nOCa3zTDIWGaC7H
6itrzcTfCLtVSl5cigYEq1iPg8Yi5949Y7W1wJE9YvDRs1FLdj+6agquORUEdb9AESph1b4uigRu
anmWeneTyYNFrfoKH927OPOzi8O5Vu0WJvD5MSGoIiAuPHFrKjep3UWhZAbBR6qwbYCaTWP8oxA4
iPwj71aP561o2kxILaKYdiGZmKYdA2zRFv4nnkigTArpcbesaIMRDXA41tQIUxiK0JcAhcLCtzuL
H5Lt86gqY9Y1ewgjSILeancXiMM1sV+sH+XLyH7lXo/zyse++ZgBpTlw/gZe1foU9y+XLlIGOFhm
zVrqisTuIdj44drsrnSFj2VRGYfzRStSIniN3g3cTUJQRW+veMR8o4I6H2ho2pSFvIVyx1fLs7h+
UGtuuNwvReMhc6zJ75ra64m+5ZSa4AAS3LOtMdKzO6mZmjmm5LLkWzVfC3oLNA1N1UP0CunJphCP
fT4GdnvRrcr4ulpb3Vg6cX0kncSokjUoXSMIyyUonOu39t0iitt8kDnYF2Zx5tto7KpnxftFBlPX
emc/mgW2OjdkGLoHMfBbbFM/Y1mYdz4nb0T9oUzOwRJBX38f8ZSBLO9IalHOe0MvO+0Vr01tOz5j
dz42T1r1SaJAw1dSVoDdEVoAhHD8oBL41641McgGmNlw7O2qUVRT5e0VT8H/W8HgnlIbds815XWs
j49RHB5qWknyAeO4YQlzqwwDC1EByFwr1s55R8156ZxQQL8BKAWiTf9DHWx65FoqbDiIibYxysMf
qn4gWwLJw0QOZ3cUU3Z6mT7z35ceBrRc36I5MuDmyR+24bZCfbO1abQn2Glr/jXVwTNFV2Wk3QPC
cRxXwNom2eFmOtlciPlrJMbK4sRnGA9L8fvHi09odc9bGFeHQkVYjL0htDbqr1m4Kk4y1H/wkQO7
MDkzVm5VXwTGxXNbKg5DTL4u1aT2+aHz7At/Zi1j2QymGRbSV67HSd/PTSYobYyPu6/Oa5z/XfES
wQQJWRN4lFrAsG76qg8pwZdOQ1E8iHCtYhaltR2bR3EUyVxjzx4W9VMMCfAw/xR0eTrSc0DDVLyp
GEJDSZ0av30NCXWpJ6ssrXu0SIaJuFDADfhNwD7AjSgXYW5Y4+Gzcd30gJaXyLoaA64CBdQ3uvR5
iBiMuIlwnxWJAkJwVM0qsgXPvURFR0AC5kU0M7JXNj0FIpcOE9OBYagCTlurO662a1eu2fdbqx3U
g0pboFHKIH7fSAqCFBwEGnjtnzA3WZaC/sBPGE3fdt5HGGIWNYoItaVmlaiZ2eAUXFtRytV8IBIP
jKFwbBcOC0bJumX1zllJbzq6T0aeh43qcn06frZ0fYprHzVl5qvSZ5vDtqXQstguHnM8+/6tr5nl
JayB9gN48RJJrMltw+BEdqXnE+sT8teGV0QVx5rs3SwOJfuHHJBmvaqCkKnN5GDOC1CHrjTAlCHe
WY8uhaVvkMCWA+5dsv2oCG1Wy4mXoC5jf2g+CHFQK+o4J2vzvQ1q71eoqS2v55y8s7qADfUI54aV
K1aS6oJXGDsPxWS5uoIZHphecYo91QaLUvFyIsKBnX+E4Mb83n2iKETQJSe5RuA1et5zuPnqtpp+
Uow1k2Kt/DeRHHWHDGcumB3G/aO8sw/8D3cwH4//NGAq+no7C0mgCVrrJtgJt7YnZDsxuMvm3Fzf
vaWssNqlZJgVUZMMvp5tDnFSjjv2K/okpNBsIV+aa4kX/Wt4fNedbJlseCnJ3giY+4LN1VC4UuKJ
NEqMmPZspTxwZGbAbVruQwx5DZD9P4xNToIKnZCTMFThSVVLmosvE1lejRsZoSFPReopWqHZFXD3
vjOWFrp18qWabQdAefljpKs2yVzzs0nJbbwzCwUjZ7CXHVEg5p29nYjFlhb2xVLuwnj9ng1XZmKX
bX/bYlobUO567lfxEJTmQ9a0xplZGAJGsJq+Whm+Dx3+BJHmcPC+xoc7eKLRBIlVWHVP81CuW85E
MHePxLdmowVIP+xUOXC0BDcRP+Wb/XERgshI2EfDPPvdydp2cHFtcW1cfaA74cIXo9F+pvsKVo1l
0uQp2CJ/JoLWd6kOmka+vG4Bz4JdxsZUeYUeQ62xuly/SM4hVE/Ui0/VbrvtTyW+ezPK4y7wWrN4
/1IHGFrWvo9zJa5jhp9ePi93MxvsjpAYDxv8Cl5l9wFfPsyR/9INsGj98k7Mm6m8kQ7AjK545EK5
LTc+TzXca/1DnAQYa2KxUnkPyu+N86g2jVBv59ky+jCLNuKpH5/zaxgsvIpyRmG5CFH41+OsJ9A0
jqRcr2e2PiWROcWGk51hi/pC0DZsnjmF46M2kBSMnBU2kNMPFhjxspj02wzVAdGpCCze8GD3y9Oo
CJhnLuI5C0jQtMTLVvSaykqEli2sQ0CvYlzQhgA9mxI55W48bduhimXoeSllWrWjjrpqiJZ5ItEt
xihmLV8mLurccEVvzHJ86CGYsTQWfQTvlB4xnAMKct5fZJ6TqlAOkJB2b6+yYmQ3BwAsHNh/CeiS
rEvBo4XXBKd696OOZCrs97Hfw8W4znIyRXgzGkdzTQI7G8+yj2nO61kF8Auji3xxfAbL4PxXbcD8
JldsLSJVMkfzEhyE4z2gmLgVuH5Uwwqscfjd+WfFAkXNKaZ5XbVzViFVFjCm9s1vLchacgs9SZbe
QFZyFE0Db096PQUizE3Qng+njTBPxHGmVemlb7+OspG3CC8p6mGu2JIDZ6721OxiILW1GuSmW9h/
Zeed04B+mkcxFL67jmpfZTVDGTKU/WyXbXvOEeeLeDy0ofwt7dIjPn0T14od/10Ne8OVBmSPh2cb
9c4ydVsh8hkjzFYKQ0eX5EfchXqe0rWG5uwFevshfgXiPu5FVglQtRWAdEWQ+b7Qa2uGSoiQXJsU
QpZwHj0QeVsHUx4V3Omua9pgItdFAYCoaoi0rsBiicQqsSHXzFAY0CoUx12gKO2xMb372kabXQHu
uexkbGBriA+Pjusai/Nv5qt/oa17HpD51xkv4chdhJwcJPBCoFzEXkmcEpFfFrL4JsJqP/AxKHYw
aKRCHHPjlZH/ebQRquEFb/KjTXidZ+Y0WRH0bT3f2h9f+7uYeLytc7/avf2rmKGbOnE+Z/xkPL9N
4iljHCsLpKdN42QUZZAHUsZClK5eMunZlTWfAuWe592ej1+Y/R2fQksYemb4g7ETMAVcf8Etp4M1
y7bfMZOEU9c/EUpgVDtt7I94U4sX0N+M0+fmN+dFfkUA6t3sqxEssLafNQ1kbpjv3DF2qNGEgFPU
Pgp0ez8yY8ELWQEYb/T3xyIIEARLjf7P2+Q7iOLFBxqoDCD6PEfSMljn/KsxiGsOU7uDmEp/rcT5
+NxN+A7HqIfmP/UrQhT4tCkz7sGLOU+L3IpHXb4Mtp0kyAONxZgyNkYkJYQpsjvTTr+C4s/bl05/
FofxuEzd9AGBslIlpQh6utDwWq+/pYZk0Skh1fzbQD2eHC5JLZQ3i1U8X8DxNTfz3URP0lPGtETs
OS1R+8Z1H8mbTQagzP5E4usySwEUHdtqSQvMMKo1vovHKEuDzw8+L5jlKxsy4N/KwIkNsxPK3bDH
j8rqwY8VSueX8QOgy6FKKXaQxCrl8heXKvhVKhfo2ydSLBurmRJNr0wvg7zGZtMuaQCIwPLu5lNw
rpcldZC3P+zQ7/MnDILCEs8+pUGq1Yvr2+qmy5vROzJU1uczQatIVw+QgyntR+ukHkgxYd9nZkna
cYPN0qloAFyVqOLoaxWkVe0OKPZKdbvjKabY8qarqMQLBQlWoRJOj+3lo4cm9wbT6cUXrcnc2fnb
f7qlc8n+yXoFxoXtQcd/aqORPgzZzv/oiaTuWGLt2S1FuElCTPIpOEOnPc6ZLZcIUPiIOTAagH/z
AkJfPtTI3e497DxTGA7qM5+gU3Qo8zGjmKo43nwIDjJfeJ8L7VCIysMN2yDJVZDIbD5Fajg381c6
vq5Qv5Vv77zH9B8+kp241sjyK3+7pevvr11tBzLa2EquYpwklRsSAlTQXQZETpV4/5+Bq5nP4BHX
hkOCUT16XQOPPVyJTLvZPdISaY/d52rSV+4sLtRwCpKLzLCkf1TeGYmWbY+oNoOqXFqwl1jMisiC
COVAHFKzvK5QLyIVpHcsXbDs26eOgD7oFdljhK0WVlzcgf1sop4hb54Zy+Q45ObN6/e40zdj/Gu0
SHL24bTCRDVTzIRL/mRGv6Rv3ID+cBWR+Ds+1qYIbS8e0M51p2a/weglEZzdzbIorgq3yR7FLgbA
r5KvsaUoLX7Q9RJ9B0IHxhp6f63melPyhn8e2DBwL62qBcrkLImJU/UoGRCzgNyfKH97phI8ZAAW
mGF0lCd1LlfBrwEeiGakoflwWXdheOCh6XUBK2Ybpqa4YtnAml5jrM2pcQ4gJ2Sc8e+tTt3djDxh
X3+FFIKr/rilz9AKiF2p5o1hMCZ1uB+BoMZnyGv1Y51asyOrgyGYw1E3enA9M5I+/4KtEPpyPVpk
ZTeXqrCNwnDXrIk4olITc3z4J97UGm9XKBpo+Id66ykj33fJ2z0SNKZj8efJTnecvy0+s4Wk3J+v
/as510EdFY/JZ09q8Ak2Ibk8GDKUW4XDKSPeSFQ0Dz/Zao7IswGg2XR4opXkHu6RtJ6T136lHeoW
36zl8a5VqLgZ/syDMvvJZcvSbPa/wTfBuhRZgqh+FTlvkdH+K37zY+DtU1NdanqujccUGC+dndfq
qpoBx+j9YMCLbbjma17h3EYhbRZDl0ytXxOdevKp4kvzy6DTHsOMQDFKXrZrdLQ23ugfwNRNIl2z
jtD+uPuIqQbWw27m8YjqTcpJmxZPyQTEqknnU8rW4lXY91DQLm1Et4o3pBIwJ+WcvqyNcXck4JQ6
KphEvdJ1KyF2x9GrWY/5rc58DXHu27baBGpaCbJGpmlX6oc0u0CrDkEi3pY4k5I6u46C2TuN+vxk
FtWYsaUIwhc8lq8GMHmNA4Aril+PmawqegOboz5ZJfumQyp9BVAGbsCUW4GW/BfxqZX2P0hAgQFP
AiR/rc2NmTuamlFTdxXih9Aa1gTjsr89+gsoSjS1C6VpzUN6XW8SwerMjriT2WIrsqdH6SKjbFxc
t2PzQTBZSrPdec2srv6LXcbVg5kVBCJCwm9znON2Zidug76iqoNJMPCjHXXUuWNXLhkVdPAFRKaA
m47nY0VBuDlCXSnNvYf6PomJi7D10e1wkuZP2aoKWAsolIVeEltPPe2Ua4gib3RKEjBHoNrzb7xc
MPuVRUx1LNo1LnOJVhKBSvty38ECSUe7qPxltgSN3we8Jwp5mJVmAGruQJ80D1z/9cezBPNNLhtH
E/7yc958DaNd6Q5Yq2aFxNCcb4N7VdziYz52WKV1xucpp/sHHgv3aCSJzd4w1FLwI7abxcVIhrbi
ZeqbpPCQHHuz3pIlA7Zi+mgUPqqoEiejSDaUnKA0RpamCENVSuDJjeMCgrlLwqpysCnVsOKFRvnw
kD2Q1LONKx0yEj5reZMEzzKY3U+pT39+jDqA0nhUmfBRb+RjD9TOmpSW9yT7RkO2/PJC72mIP6JU
Jt9IzGM8rkM5SqIUX7CKjHogtOWAhsrlTEepYhNeT5Xaeheg/quVOVdsLkgy5skBMx80XU98qlKa
8FcEyXjWxcE7M35WKjzuCWLhCf4FPVQZlQzAwBIK1+eA7mHU356rp8gYnHtak0aWYfiictIM4VtA
dPqjyRFgStfkwJFENEzU3H6/NNnFU5jENAPJmpTmY8yGMLXnI2oD/jM+fKBYrA1mRh4NWfynhKVu
PBD0w5M7CdlFOVvB6u66dkl1nZUMdQQuTCY1s+Ndj6uSLHPihmYjyVNv0Kipsta7El5W/qFI4mVL
T2C5e/9Y7COz5bTSUrzj9/47H4Ep1aY0DChE+CsJIM9/s44015lj2qBkO9ZnF55GVKKu3nwXIXx7
BHQify4fHSEGiVwUgJyku8cwyNfmccvffPO1wAoCPQYbBMWBjWIUpA+qPQcKbTJyWePiAiRa2T8p
IfQYKjads0uJQoVjmRtPbl+jDvAaQz90CRd2jHy7MEmnkgd0PswjzZPWZ8T5XhIqLQciEx+cvMb6
O3q7Li4KVl+zqbonXLJ+jusPYUVV9Bv4iWgG80goOnBhCnn5ts6DtREuMEy4DTm2qrLLSiqrWmNP
CmjSkFaA3DZwZ3yFNICqeUcOKFjJWnToW+FrfBM6CP/vosFU0nWiwd2hC2stB/4Hk9lCVyMrlcz5
5gouMTBnNmBCvfuaD+S9afZLHF5HC/3KUKNTmsfqC8lNwdna9C5OQ7YWBhFe0+ac1KqCR06SLJnD
YBVI2pqrAB2MK2VpTdUbYa81k7XlKbsxRspQTWEFy14Suxe0yPQlRgWnWrhXvVGduaTeLEYVEyZS
xMpXPUS6h0oFmvDvKsZH8fKh5yug2u+tHJgLGKV46J2aAQadHohYh4j0+qjLcCQ6GfATo4n3+6ow
X3krOnVPNG0q35Mmuf5iCiCZLn8ozBk9s+bbllSFHz1VBxDp8dBgInLpsAms+Vm9nP7SewNPFVtm
J3Et2dnekAHlgdZz73peEkxcvNaLUWXA4aWCaDR7bPWDwf8K5wFoeCc/t6tt+OWSnyVVwmPPTQil
+4X5d7DmJyV4n3uoU5N/VNImfiCybCVAfXzxbtU44BZ930hgFgJns27UvvljAbOkBBQAtVuH3Ykz
ZUxCCgt16J9v+zPNyJZcur1nm+BxBIY8U25ljsyZToFrcERX/DUW7uLWQfJUGmGmj9doKCM/Xw6f
2sNgvCcg5itMS3LHYQd5BZXMf54r48uuPcNfM6m6gwvL37obIzRO51PVPTcQf95UFXHpj0Fm/RQC
8JxegWByWQ5/mREJSQvoM6ZgyPOOpSRD4TAq6JIUHgELtfLWrx8CiRHAqdrv2n8LBJuI5o5JUlB+
0L4mv8vMK5IbLGYqkwjgouPYw9toJXI8LRkQoFV7p88RwSK/NeRMl2pLiotPxHYSMAvGD2HAfMIe
cF/EXqVuGN4y1rhT/WPeich0ca3nS0Zbz3T7IIJNaw2041VA1lnK2/1lGxKW+Kbmju5mXUqR7Lh+
6iLsHwC7Djk4MNEsej/uSJ7xx/cDr8VZGr93mZxUjv0TREXwzR4iCzIKWlGehYAMrngsasssq9Lk
QgXkU9v7C0VNcme1U0gGfQnmFk0r6GzuS1NF5rIz39nqo0ZpLWWkXxQamIpgUfrMYHVhECNVboKJ
Dzd6Ip/U9C/XIkG1o3FWsxyhT8E1tyxv5lZnuTLqHbfePj9hPDhJZN6n0cG+kwvXoPoMIiZ38qCC
tfddw19FIp/w9ccW+SYZ8Ah5OeV6fIAijOvKqK4g5FYotrXDIodCEBK1U2gkioupQnlarYj090+w
xoSHpGdzdQQ3tCKyWGRc0R0odq4J6VdEdouAkLLNJx98miA3UJmQ+9ZXapmtI1MCzfjgphQCtbAq
lhqnpZ1P2aMHcE4oIzaOCv+mNyD0v5ki3ThqVuSuW2nknQWjgV/UBK2+xR/BAYIUX9fLKdogEWWc
UU8mGVsdyuurYh6v57Yt+7q+Rlshp3phAZLzoCCEaPvVu/Xzax4D4+Og9RJj40a5pSICN374X8cr
VhzMryalMQ6vEhzgwGTwdrVbs8pBXWN+GqUCoaUdF2sBe+/eAH2Uc589NnrmCL6g0AtEfcnKTu30
12ZK7ikpGnatjVQC6sf4SOKFORMSug3z3YzQ5QyxxF0pBgNTmuNLUV7dKN0kZGF7xF1n5MypQThG
ld1UXo4olAjaPvgaAz1RI1O8dmKl2I44dwItUXS93lbgkzWDEQdVm6P4CIdECAQIajrU6fzw1QTd
WmIS7vA1FPx+gjBmbIkmhSclS+H2bIm17ft2j4ThVw/g5HnUFWYZhYsaeqz8K/NVcPptr8EMcnK/
+Ao5+w/wW7PgI1HVKgsZn9saIjy1NIQWxeuP7SxtUVAPfXRYXQBBXI8hjDADlDrEhvGkDt3/rwmi
Y2Du30nTR0VejKoFe/DACXvTW1PtIhN8NpplZfotd+EBsJC5/8SAQ16KcZDwHrG/AsqoDvkGgrcn
Q6XEe+XQszPHFlw9RLlgYqVoxCFwsFw20nHOPij+X9esoMb8deIOAfb7UBUhkgqKlYzJ9TPsosuE
clLGu+Jn811XU6Hr3uRG2FSbn/+oacauIjRmbfBB81KKI9y/CEDr2zGwxADCwJAfYljKBTWCnbm7
yQIu0li8ypImJcUnM2WN6mH9pJISEAOHoL8XPS4/CWa51er9fDVIZmeryItJcqu3ZiddhSqV2zMV
TSnt1elMAnA8g0kcs5qHZV91nnYzHJfhaylRejEfoi8j19rcd0vrcM10HUQzitoLazoG4oe2nYwf
nOIoI67G2LqxwvdqZJ3GLxs4DtyRBPylBF16EOx/56MGmsD8Gn9o40Er7BXC/MJTmaF1tgdnv0+i
E4IjBoEFZq4X3dBTLHBdPkXekyXE0yhTJ78zEHuuRfst3CX5i9odURUkE7qkx3Eo7n/wWbL8BhMC
AjMJSoxIvUwe+veqzGaLOV6dgnhGcCDCf8NrdRHNQdb2nIwJuYIkSH4mJ3il+INnF6VdAseHsIVy
4OcC6ktIt7YvET7AxdejaqIEu+6AHJs+D40sot0goeQnbyR3FUQD5L617Akr3GcWr8d4eem9VpLl
YOY3/XEZ4ZrWLy+IVaXL9025fp+8tntGEFxu2EQ7GJDzM/bd1Hq5NI35dvca/QukyvgLeEYUHRnt
D5rTBVVMsOR6fhwUXZlBQS9SY6l0CF4/edDp5rfdn7lzLjo3QDwvT1c6HQwgs2HxcIOWGy/p5Dn/
BqKgpBys5mrDD1BWfI/mZj86iICaLd/GubNt8Od0z8IN4hJadVBybsiwCO3h4sLKxYcpTNnULA6D
6FGYo0Tynu07Nzav5oxcDuqgfInoqGkq+D/Wi/QI17UiB6WqEDSwonHycerx8ph73S+LaDJcblBa
+39oF06IG4VsfUuytD7dxKckSsItcEt7WPXY/riOlXeGk3Jx6DFNotX+0G+t85/UrBMrdpfhubRi
vyJTYaYslC4vpdSvh9HM+i2QRDf6TEkkqGxv1Y4AcfOHp12j/ASCe6FsVhmIfpVfYxrtMwhUigh2
qh5bPIvTpH8IVptmuXcHyGVoavov3R8hh/wZl9Npp9mU/+q2GqKW6NyDaZ1xXIXuAYIxBShrPOAp
0AqwRtLOgX8OmyYB7tOgNcHB3hh/hzNNSpXACtDRwy7paCCPWqJIAb7F+Wl3q5wSgKkmypdVpnY3
lPuDAFaS0A2o/dqr9kW2rvqGfldRjUgHb1RIg47KYX9G80wCSIWfhgIXPMwg0WmM8V4TysnVoONV
3WClOkBJOIwbNkrCQqQ7RsNDPj5W+6JqvaVKZQBj6czwDgpwzJxyTsy0CwlyREY6IIWeD7rJCTue
8AIH4OqosAISL23YgB2/hJBYv5yn74Ki7Zf+ltf0NY7z/dDC6xzVu0fOtCaN57uf+6GIjtAexhEj
yAKv3w+/JSNPKvHnK2XP2NEKUV+FLIdGAbi8eK0dZvqgzU8mzJLmRpScuuxEQ1E8MrLPqdI2Gw0a
0AGfpcUh7qv8PSqaRIDO/suS7vm088weWhk+X8YIzu5ynEXgxhOQzyuO7RWdvvrnl6BfAWmqC0Ce
o5+kH7pv29ZJpkK/7trirfg/Xhf4HYW+nRQTtoD6+QEe25D/171L2Teyyvfl5yuB6Zyp+8CpKWYw
glbUPqPk7JsVArbQh86LYQPQuPAtqNp23A/YoTYfGWF2Kprfew7ObxiAR2yhlQYH+7aWwZeJmmel
IOyhZXIIj9lJFfmwrT05IKQGE+b6g3w004eVZE4zQFAfnwSSxc3IvJQa1aLkfqmaXr1SeWI341Lw
VmeijiZzLJ4W//Ay2v4CYF8Ko504O5bVsdz1dA7OLIQQ987tvsWulpWz2UW5WmcStWFOyj31mg1z
ReWKf1AsRmBQvGz1eydD3EfiBWJPOvZELMHaX+pLCldGT1jHZ+ZS7oVLaQgUN43ovq24cHKyXetV
WUCcwZCJbmJJizu4XoMLgTiSJcMdlE8LQfywCbbfaBAARY5/P3GMzQVBkekkHyuS1JpehlKnWFsY
7PFGVQToGdTAFg+N2X2qIg70LCqpLmZIu85a/qKPEUuJHu0n3LzbwpqpDdHXpKK9z9XUWF82sKlK
Li5FajrdlxL+pr+VTDMRe44/W3TJp+rO/hkeuzD7FzfB6nnQtVXqSHZTVswd4Qldk9l1Q9zMOFIK
+pnGpzywZF+sM/pocrMDp+kLMWeWC4QFBYVFfiW0XBzKWonTam75hLs4GRu15AVz8zUxadRzkoAq
tCqEwxuaRtWwYs6pDWU6PKc=
`protect end_protected
