-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Gn0ercA1bu1CG9iTB2x7B4pnphCBWnO7lDy6SgcmmqkXrd26ubjIb32XsFwm4q4Y
TGm4cLJttIyFnOyyEkAsvD08camNrQCOEW6bThRKWWRCfN7BTGn/4q8abyn10MsC
az63Yc+Q7TOsb+y/VWzyrJe8vIY05vB4vZ/Js24EkQw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10297)

`protect DATA_BLOCK
eBpVzi6ZvrgYAeY65JSLkSIl6TXzJQXjNlm16Z/g1j08l0y7X5pwzTaEdZ0uuBSX
vSWSu2kxjCW9guu2NHkXt7T0oHUAjLkOZztfIx0NsSx/cPfv6pSf9CbOU1CpzDJ7
dbvhJUbFk7hjcmR0/eCIE3zygOG3X0csf/XAn8DSlPNzHoz0eVOPj5vvc1j+vy7X
BOvGX86yWT40s7U9i3U+kArddTvt+cJaNZTDal64gh2NUjvnrmrl9EJ5WMxhBtsQ
X2J/0+8iFem6C/d/i4dPagTB7xEmGPYkaUZCiJh0Pa16JDOOhhHCpjNXbvC06YxZ
0NVH2a8wIGohrnN10sWptnng769ppb1c+qjjGXwb2xTs+xrwDAPIbV7qdA/DUTDr
AFLDo88/d1KJnz4Oe3S5e8C58Lo52lNnpd1uo1QxG3M6FzYHBvAYuMg6+Oenmt75
oyUg6SPJvAw3noS2IpTfurzuiBJxeXl0ewYfPdbl3EXFtPkFyiR+ZQBC8A9c101r
JNYGYEy+2hDISftAQ64l3Az9gfTbIAxVYT6nu7whUtXlkDkdNJGIB4J+OwDhPqiL
9ksvXkjVJUOtgnd6A9ENo3rB0qP+/RKRBuCF+NGzGVEwAHFT5DJJ1F1UoPl7lpUQ
NYaiMDjmAGuiF+S0eujSzTnZBQ73n9A0CZ51bU3jjxncBwQu/9BgPqbm6WK4XVW3
O4zWAVXU1F6nkNJ7KyyBaOHssiUPs72u3wNa8Oa3PLfJNd9zvGaWtMK28yTNnkDg
4EpGFGOwJWYRiSwrMOwYC4od7sfZ89Co/RBlUMqlMxpRyrrXyjl7imYL6iEvGpzN
9RLadOPQTbE7d0CBOrbELqffeQNBcO6JFXFDTa8Iy20nronIYDGPhSci0IPpcz74
KsPz3y9FT2uAgD7W+kozIuaedrAex09UKdL74Pp0/5HM+LNcscE0wehIw1roBcvW
B23uiuxKJXiJ2kG02YbI66d0P1ggt/UW0ZugJvtx12t9C0ZhJdOLjujWoDL42jpe
C1+pVPdbLdK8QKpOlKHi+lj81NEbxuimUJRFkQyYj8XpMXmFtuw8l+MPCN10OBYV
WlpfwSUzPu2656XgRDsz6rruv3idYT4Exu3lL+qXqRT+TSX6u7Kxi9hHDceZB1A+
K2TUKsIdjW7VeYIYqAbsyZAhSBA/NJ5aREySLk+2AolfeOJz9sPmul1CBhnzBCwy
zGAKy1d9dEsCeDhNydVJ8e9xfkC+y/+m0ld3F9xPC0GtpPLP/5kglhJV6+TOrsGI
PQWRRf6luhv6EO6ZCtxGpMLFo2DC0j9voL1y68fJzPlSShZ4TAGllexd1AQyDoyO
TSSt4L+G/roUWfRW1UpLlovpEtJvuH+SDrIJG9+ucwTtogGrm0nonDg9iIc73Kpk
B/6uSDqHrAaYBh/ZO+FC33aD+MxBpktFDdPtZPzEA7365cB8HeZolghpkLaQ1e/+
TBnjo95J0h/6AvFOfZVgtknfj5AwgcM4CjGUFJHrjC5OKzuUrdbir7zrQYN8pxxH
Wy+mIH4qQjs/PuQN+vLOrJoDgJPdiQfV4wd0hDndI7AempqLXZn3gAdNk2E5Yoq7
V/N+Ebcqd5A6nos6bu1pcDEP3AooWlEA6sbGX95HYPyQ/o1XvhtNA14AAOJraFgC
c1DiOvJg8zDQdgJYrBCYCGHWsT4zHtFRAIm9PUlH7bHXj70ilYKvva+Di+aC/rs2
i0cnhLiisI8hF/DdGAtfO9INbIxFYygt/8DcXUSUNzYYSGrifGEQvW1BHzwx6zPZ
Z21yVVkPPqTCJg6XD+tfQpABXWXaId/0/B1KjYPWgIqsp2iFXw7wfIvViffa7POp
TYcewETSWntP8HwnRlfQODe+jzlL/y+ykD6aEsZ9NcAIg3jzXhSakktIILh310//
Xyt1eNvg7gEUpn4P1uT2hUL7wwYlXWTAKX8n/kfy8HbANRLBBKoGkgEmmHw4qO4W
YNyf8WesQyJpB2pT/z279p1Ve8UIMaiSBqAlu/Smbd5HkUwdI2Kicn75bUXavH+7
rkgDQG2CMOujQEIM5Kk1sSyEUcFNNEkr4/f1lyj7CMc6lKl7SNn4bSjf8JR4Is6p
ozte6/Bv0hu55TgwrZabQmU9cJSfxMx7KJl4x+E1svgPPeSdKx4B4jf128PDAjqS
R6szZ2yOic2M2sPDhzGmyPdq7ruk8I7o0p8u74GouPjqaRm33E3OzdPgNNRPHL6R
aUp0flpL2xf8poCTTBL9ZrOTRv1MzpjGwkzx5v624HEr49b1O/pALVSsJwLCKFPk
WL+TS6yj7pP6HCwOFZywPMMVKBTy3zmzw+10vQKYmhF+WmXrsOSjYyfOIIOCnmPo
oFfoTX8IZBdB6uBhoD58b1hOGdTi/DLoUCHqocHo9xtyUKxCxwrvzDGRGtVUBgLw
0vHhHtHBpaW8DXyPDYc0fbu4fHjMtXAhC4HXqMo06W24ZCrfMYcPsf8U9KLRifuB
Jv7tl8VlORbZC5gMMUURvwsr3LgwbzkXPi+RyrY+k+cEfd0RZgXXIWlni64f7pBJ
SqCbXERihcNCL38BtRUBcZOvZdIQTCM6ctiDl/llKr1Bvq15c1k77epoccDqCSLO
DcwRzKrsqme3N7XrKTqmvxpvD8jY/jcm4NO+ilPa9yswMLv9ttCqyEPLuV2UW0lL
Pp71nXyTUvJjMBen+e9GRg1FnQhlsuEjsen7SopGBv08259XvjI1h8nPfD0nKTJP
EsKcSuAyUvmbLPh2LfG2ZOtdgvLEgdVPpQnzZ0nKkzdrwZCMWObV23lcq1vSwA5u
a09iRj8Rk9cpLuDHOeFLAE9poxHJCPDFIx3ZGjJu/gc8s3c623qddRFmEsVcckOa
67edtZLWSm21o7kGlRVNPjRh01pTEi+zo/tUOo43dMqVg9W/sfmXIKhE8q1XlF1J
ArXjb6E37D7WMP0z4wfk8m271ww5W0arIjxa8gdrQ9LPNmN3npLwGX1u4p66Z+FZ
pG/QLUFS1TOoE65jOfhN8FQiklSBDxfsKhgol8PR9CjEZje/UrMWd8AtZrOgLfWz
SW8cXf/1ilY5xaiObBvO4Iu/RtA2hsW6o6HclwlN3MvsPaeYvR5l2eFpCNz6S31i
Af08KhOOqTIlhZNawBGq5XPRM0orQScmHpts7mvdVfl3HqSH2NOYpA9z670mmHt3
egR2V8CJb8NYkmzStBh7xbGgnyIiPc1wyEPQwS4xQVlrJ2atPl9t1lhiZ4WsazvP
JOYQSk1I0bRXtphmFUqndHPCDjsn6lhq5KfZqNFFHG02Q1PwLeQ/rDdE7ZCVYQJr
0eH4vJafjh0yeAEkMjAoFp3lPZgZ5AF2Xn7CuhULvweuhpuiP8ywqe3pbWI0KFtD
xT9ZJaScORDH/KwVjOqb2vwfXcFWmvudHOe4UAFZyTCE+vcvZznc/BFmiLO+0ZVj
K57IwkGMZxBGA1HTryP/wT9SnxwVeJk25YyXZVhcEC8RSJC2AshjwjTfqxDzgmtc
BoxSMNffu9p35g9be2cMisRNabIwwMU8+juHSXkTKnakSdGUbTnPf+lXJ2N79obQ
n9F9gkMvz0iT48fC//9qEhpbPZkm6sc8KJLFkP7DtzN5QtpMAJ8OHNcCv160CerT
Mp+lx4mW40XzwYdRJeOzvqx0CCl9X1jO0a7QM6keFJi63TpVCK5gEHj7ZcTUSV5G
rRwqLjp9xmmjfrC3ExPAoqKLsAwhL2Z9WuGsLT9trl4HmmWSzLGacNRGDat/R6Vz
9teHEE/Vhj3T7HoAMfUhXceIvZb9/j21NMpzWVeSeSS5i+2R5b5fRtgib5UVgPKS
4pQvCUnDR1Dpq1sBhHlJ6ssK8889wdHIKyw/ttVeDIA7oaLyh10PBYwpNinDYTmV
acVFCnHCK2P+PmX0zbNaqD3O6Alr3199CbNFa4/d3h0lMVvlYPq76vccfrCa2nss
PZiFCP4nMrTIsQlJfkpNplTXQnioP6LssOwaTq/KIzGk2Q5gmF5MirSRVKB5Cx5I
b58fjKSJQW+692UeH+XaOsjOh/VSBkWahmVxAOCxSMLuCARE00Z/Hap23ufHYulh
hEbe/7kHf+qFlS+J2o2TF3zZdo+Qnh94p5iYffqyc368GzVUfpJ/g/UfHTrt5L7s
q6ZmRBJ88MRo4mEYEBA/EfVqSZpi3o01zKBhSC0xG3fof3qx1EUjEbgLg0SZRzkx
XfGT2OgOF8VunfCOe40HWZ0j0Mgy2CQkRjvAwC9zuxcxMgynvJGxuKm7fumuPZOn
keUC79zdkG4m/Wa9dSUTtkCxWhP6qavbHUdY6yQ2sQu4MmxKNDm6Z3uFUc6pG99z
cIyfRNcioui4H6n54Vd26He1vAHD8i7S2ELiqF5XLzGKi5F8iUNxqqIU/Ai/vOdd
0uxyNJMtucKJNq7AaRKmHHZJ7LqVDSagP4/LmusFhERH9YQMa8tVuEK1AN6odKV2
cFbDX40+6vHYBaGlng+ROZyEAPe/UEfasM+StY/QsSE/Sns+DKdXFbQAHwLSU0Rf
KPDzYbfg6TWevJzpatCVL87L7tn4/6bQpOMbm/e4xa/6v23AZlCB2qywKpAtDiyJ
u0Yhs55XfavhBAp1eG6xBxzs8aELEzoH+npYVRPt/nATM8V7dAYhCkMr2o11U1/d
LrnnfHr9gA3miNKIFlr7RVsllvvDi114gneRgdHBg+7e7zIcOmxwYJ+APDvqfHv3
rfimWoE2je/smEnSnxPdxvpzjI/CTjqqL/7C/0+gVVapZKrtgUxLnAr+0FQ6+RUS
ZyiDmne9+PKuARUthAV9irNLRNGgGcRvTLJlvTPG7RlDcTUyeN4BaYMVFxmd6CyI
gv9BPqGuYFmahcMI9CkDWCN/tnK3+Owu3MgMY48mcy0+7uXoers4gvN6XU4xypNj
qUY+TZAhydYRPpsIqFAwULN7Vte6/kLkcRL0xU+LCdxStHkdMEj7BWL/3ctD8Cs+
OJ9oTNTZVcBRshU9kN6v3C0M88EBeq/XCrLHKH0B9n/jyop8JYXqpqkYb4LwWbcI
9DkATL3aQv7uO6/nB9CvZkAz38HArXx2jweHAAPsxN7LI2dGBa9t/RNTTjHeUoz8
D62xXZQTua4B/ZM+RayhdPyaadFig+ha5dBQgd/8RcIAz2srxOa29XwIqWBlYXeM
CRxZQWV7/YbPqVl3LbVTXpkIN4p+ruL2sP5B5rzSksRWGVUJfE2FW4qtQ8gh9a1D
TsM/oulxnOvncIUx7O82WtB78lzVveJ96RhU0E7vJdn5lecckeEGUBIi21snmMTm
iyrUbU7DxZbEBZ1hNliOOtCI1JuA/eycshM/FD32rZEAtg2LTzoJmxRhUlYDzZM6
Qr96dnPV3+kPdfPtPdhyVvT/o0a6ZCW7/PUXEYN8USf24JUMeU0AyYPeLC2L2fjF
wqU8MtqRlkg9Bs/8l10a8Iew7+43TU7vCSZ95uJ/tQapcCBwGuj0VuvW8EclFFI0
US7tHdttqRZGZdLhJIoRVrBaTvOQIdTXhv3Sms8YUdX0gALsw95FkqU5fJat4DNz
sBkvhmqNkig7BDBQ+khh5YnIr/1dvIe7P2zNJckzguVmYcQgYLG+8WSb22q5z4Mx
fcg0XlfRrVIaOeC7tuak+cStR7opGa6k9wIFnfq8FOAaUZnS7+/7q2sUgkqTdELz
s/mZ84RRpTzbJJN2JfVsPu7s86p9P28qdFFTk7uNbAH8SF7ZrgCcMw1A9MFySTGD
bsR7KJO3vo2+fvyfu94+Ipy3azSo8rdVClA0IVcfs56MU8miU2S2GhdUg8D+5Ys7
rZbQRKQAe/iFoh7XPjdHv1ZHqrBwqMWd6CV8PHj4OT7KjO51/IjNpyLRHiqJf3IV
OJIdHitK0PD0Htaj0GC9xakKPXEbrRD1D68VD4Tec6WcSQW3FZ/kddRRUbukHEzv
KLHUab0tyGKOuHRzkFvhx8Uyy4AFpZPaCab9M4CBxTO4QIeqtt12UxZvapyUmrBA
KtyKNqHk5qzZpVeeH6ow6xQ56rw076RsC0N+s7fzwGidmet689dNaW30eYOiuVTM
BB96CPP5v7ajJrPftv3qE0j0wj/PJxbHidwgLpcFhAVAPGtuaseIyW8fodkuW6le
f5XZc4mhcsEE48cDeKPm+HxqLCEniYPtqrDuxkW/tiqGuW/epdGyms9KScuzjeK1
Gz+E95w+LRQ7rAprYex1ly2ALt8pmQIkgbYM1u3aQJpl9Z5A4/7b9gLLxoTTGBXP
cLMeqMbp1viT0jvPFe5i/y7922shyV8y9aLqr/n40ITIG176kJuThwaaBozJaCL9
HH1aAxNtMO7xV6ueCoOP4ti7TqGiv9HMN+XzKppymH7bhmVIOTIzpX4WfKjM1pra
6/tbZFsnDbVrJ4H0n8jYI9o+EcDTGPbNyS34bKMFCMGlkROL4HxHs113zg+DWaqB
djzcTsgIo9hWAypE+SciQNw4TKW5vgPT92CBG+odtsy809A9NkxX8NW1KP4sixGm
iSu6y9eM6WTV7eMzuVLxoWBwzrNEgSA4KVkYKRCm6lapFZ4dEO5/Z+l0BF6t/qfj
LE4Jx1BXUF9EMHt3eSz5VvBG82Wm3p0x8rF04zOTbU7mrsK9PuzGmFpgCa12Rc/Q
1V3fgzxhjYIsTaOa2dZKanXUYoy5KnIIw9oowkazBNse8EHcEBA/sH0yYz1x+w+m
oNw5lxlWgz0bPJ68kcqFnoUwJclappbZWjUgl4w+9jv9ydK6pzqNuYts8pW1VeRp
ZQkxwy/8pRwg4XCFuGQZOEQcIzWkQ/5nNIcq568VTVwBYiwN6znjSAcZubzlQpag
7qlWIxMk9yacK1K13yXCw1NVNHJMCiL6EAp1vHLqMfSl3Sgv9RU2fhaWl5W2MXue
k9RpoU1tExYpaA33DTrohseZ2K4bVdHCVIp/zcD9nEj+LKPp3sRUu97vbfY75fA4
bAjmoQSrTb0N+LeQKFIeIBvathX3YTQEpGlePdN86nvPlZG/bxSz7CTW+sBMLBgw
DjeI18RbhH3Dk4hn+9ksG1FnexjS1tKMqCpa1evy8P2z+c0E60X2d7oFII2G5hoY
FtxdG8p3ZTGRq3KD9Ignat6AmCk6cAaMDB5c7ObdksWW07tqPK0hqJShhjzO8g7/
GSxqaweU+sx/T2t3mrpRcsMzXw3nPSwUC78oQyHXaqFpJSoU5fwoj8NYDw0Ts/A+
qhSqu2aV0yKMi7S/iqIJDy0lEj7eXtdJwhEJAlIeySBK/NBadfImOHNxhCKXeNhr
LDfPAo1+kSoHyRIfkLBDfPpzJWauBNmhqX81scX0u/PhF2hDWG99cgm/vHIil8BZ
hB+VeHpFGZ5U5TblQkKwLTI07legxWEudnwHmR0n6oM33KQp97gny1ltvfM/zhtW
5ub5z7gcYi9UVgMDW4iX/XNVQIUCGiMyOdvN9hSHXHbKoYIlByjpNUgUulwo1Q1C
cs9tzzG/bJb80B2XoSJ35olQ1DSIpPjLxrf1/KDSs+PK3WEKWpkt/cYN0SPk8U1V
kQgI6I0YmPpAXm1CbDqF0JfYeCpvJhxT018vCErpdsXx8LMspkhEFLjmbCaWYAUd
tg3aPcRX4KrtPtOJ046SiYKgairZLulOd9+MzW5PIyTQcQtXaICBh8CFELb/jtIj
//RbWDZ1r5LF2ncn4ACg27p6WrDHquv7eGlAYUbrVHEmilVuIGJ0rYKUwlAQyL0v
QrG1PjWrGSVMrF0P5/jc1W1BMg9CDGtQVGls+mQHj10lPnprxX5OlQwHZQvZ6ToG
77ruDplOUIXNkH7kDpEPhUVdYLZ2tVO1Pxtmol9yLDHq8PFzeRHwWIc/5AQzO2Pd
i67XARd15LKKB6VQulI0WWX8SEtk0xHpZUA+AA1HMkmTAMXwIsE4lzfKnXBd2IGM
+vTzNbF4KgaAtOh6LZSNN0bi8rVGEKXK5bicyTT8uJcWqOjbfGN2UX6QmxRGtNev
V5k9Ppml/vcGg36BQmdKWKus/0qL5rsVH+pT7gOINhgWM5JbqXMKj8S6OIg5XP1l
AtfrHXyUo3FB1CJFcxm3duTUBUjrZFlX1NM9/NN/m+AlJLMRhHKa7YkX37pTlEc9
rE7EgGprj5IVF0F02/8V51aEENQylm0fd2fWHVVNkLoZEaxUqw6GCBk6WdrvvYFb
OS0LT/9Zt0M3RlYYB0XUhYoJl72rluFbsca+Np3OFJrInnn8RrAJ8NIvbKbXzSDm
3tuGDcQA/NBuX1Lzwhb+vZu6GZbhiSkVXP/bIvmhrAKMY/TYiCKi7ZyJQ0kX3r4p
ZqoKbvwk02SnJ3UdBeZtO7pqtgUQlPWytr7t1eaFKL+N0AjWJ2g3p9ShZshLql7d
9/G4mGyd6U11mankAC95UdEBvsEbloHMcRXP9b4kCT1a6ym5aPE1x9DFx8R/Wcd8
gi0gg/3THS4NB5mb4ty9vS+eTzjYsuWxSAeaCqIMeIgafDrxVEJfUQk5YQomdD7g
KbQYf27JEAu9MZZWtJ2oSb1cQVG2cmYJ0+bXGmWAZ24K1fCYYhQWTC6tzykUf0BP
CTJnS1y8cyfZWw/Ifin1HXK6LFmOu2W774th3Y8CqWmY/pTB/V5/nsWc10xw7DDb
A+OdU1H5052ElqnNlP28xpfeA5ZbYv322UooAsYq2175EixqRuZjC33xnAKRE1QG
QaXYp++VAXibWGZPBadNfvYgLCnp4NaCXknTfr0r2JJnmRDaw+6r4zO9iSjmldKX
3VQ+AA5vTk2pqc87MkBmQvUVIcHfWHkBo6+e42UA6GV5iUxJC67z8PecsmuOCwM6
cv8Wm8c5ETjFf1J+5zPhFJM9rfUYMTSm83rMNsvP71PpEJHQ90UcyyBuMk8PPM4g
a3l7xnwcHT6i3DX/+ZAT9Zx9Z2ILAd/ooDgbRJErOLVYsKrzM8wXMFrfUJKchtam
FgAgQYM9fH2kpON2sHDkB/4v2Gu79OoYpVVJz+lviXAcxe4mb6hLFmXlUUhl4Mbb
fLOEPhaPvJT10KmtygCQZXbuAu8nOUZjbg1CyTSaXzYrRb31fw/4WMGx6X0bv7JE
Ev0Y404EcQZZnjE/po3J4ImGaHA57VcMPsWmGHz1wUyeya3vdqmtx5cS+EPsJvT9
lJTIVCgPN/cSs1aHCCSs/PjtAi0JWXNvFIhdwfWUB3rbxc34ONJj+XcaG4Fn6HQt
4hWhB7Xr5aG00VtFs+IIA4X9DAv+qJrWLgzmelk6woYs15yl8Gfb4wNsKYONqn82
rVXJ+KdnPCoeU3S+AJbD9USRA+xtbCyVwq4GBKU2bjTnJeEEs990kFXV0bdHxjRc
DTIIVf7hqsJ3dSqINQdIE7DYVdg7q0RL+JxpYKW2p05XoW5qrCKMj+tqDkXIzswz
vyV5OPrCkuFKDwwYo6kDDAc6UeBBWP5JGOai/rrnVVmX2LObWHNM/1icKmvOply6
T13zVTPgpZzlg9g6F1zOMVCy6YfX9+nCMuMAlw5ICH2rBTG6zl2lVl3yXQZ+AV9z
9FRF2nqe+00oEbDsOdGNg+NjTBH0UfKqSwOncq10XwCmwTyGJZRbNmTnaDxEr2DR
6+V+UoOmdNUZt3xo80bYwzKzE091W3fgTyAFl9VZjLJszKdYGS3OQn2egWFwlViy
t8NMaXqq66OECGNUQa9aKlUQrKsU9OgBPexSdkNlqk0cLAxv4Lk2mi8CS/FXT0A/
ah7xl5F09LwtCyKdZf0dZufGVA3l3530WojYFEjn4IGdkjkyfIQH6OHN1SwQ/d91
eYmqtKmrbP47AG4CbVm8u78A1DdLxOtTbHoL6UqVv54pI4Kl7Kzrkg1NuD4MTMRH
SAwd7mzTE/BL3VvRCZV9+nF0GpIdAXlUMetsGelV4foBZFbbXP8mlJRLMV05tD3l
2cmKPUAY/k2mYeS/TCVsDhi5OgA2L9MQsBYCGlooNHrQYWq6IeU2/fQGx4I/Z7Wm
nBL9xX9G53vvGn3PZFtFE0dA2+FODaXrf9NfOS8F4WniJXmyundEVhY6IK+zfVxQ
wOpAcLHBDWlNLU5YuPJ4ex9kRfRsSS0K2v2QP7MtNHlq8jx9JBRIanREMIqm/qw1
8wiYiFRmZ8aPkRvGqtYVeMmmOGt2STGo+sBJ5Aj2BSHnOBkdUARN07BKMVs5fK+J
RWwdP1l3xHuAuFCSo4MAMdrNDHr5niv8yx00ob+9fDUnCdvPQ4Rmk1BlWVGzwrfL
FXDO8fmvfCeW8oTqhZXKX22pbeGPhLKdAq0z2/1t0fjwY15tikiojFBeREy753Es
ntS6MZLapFefwdpgfL0gunAcOlukUhDK8JAg3AuV4022Wo3hh91d2hEtP9I+t3PL
nMRjuApRZLzssfiO3UyKp8zNfjbxXYek65g03KMDoHU6DIHEM0HiJ0GO0X6HYxDa
YHb6pIHKgJw+k8B45oe0P5l1DJjtp0XkZOHT0CYCQ7pnSZuSQdsF9/+P3y22Ekav
GSjEzhu5lqYhjZNkTi9GGNh+OGMReFcwI0eOnBkPdFkvm5Db/zYP7EZATZdcw+Tl
avo2jhQHUt2bTEyay4Or43SKERpQjI1WZeGshAmL6o4wfHQX4jCjphqtvUlxVjke
XObKG2IqxHUlTAcq4vu3AhBU0PV5QqcKL/rUCIx3m+RbpstGvHw7PPJx60PrtMv8
UwDlgHdNPrKHxAX1fPscluET1cRCwFj2HlAhtgaNvrLyuRQVyKjxTrKyuaY91wih
fvud1JUHZvkSoDqiBnRzLDkx8fdaSn4TUi0A/aEVmsFZWt0CpDelONoQuZPq/Nir
4+DCrRFhTL5Q5gFO+23lvnrsCzQabQlcPWUzThw5q1P/d05Fijk3Pi/cYP/7qg4g
+fnye5wKzq3OgD7gZ0QdKR3P2eM8jJOvIU6XYdcPIe8aU8kBObmRUJbnsrn4AL39
7RTIReM/w3DptKGinRfZL17R32zlUIFvjgmKE+Jt4NQe1blT2AdPyxgy5PbyLGqS
jnWkm8Xrz6WE+6OVrpfuG4MsO+onXpkfMFh7YPjoqDADVagWemMUWiuSRcFQMGhy
ChbMCdXX0mTKZNHbZHtOMsxvH6IKZA7+xuIQOxRFaKm1Bb10vLXwfWQNHfs7Lwmq
m+jzNH6w2S7T5pRFWC/XKZ7b4UP4CnKgtochizJtXgbzOcYmeWSE3sLm/6N/WD2D
0ufsr+71Fz3vi6TSFGvWMCyO/A62OCrK+Kt+xbZFL5PsDWQch9WoZmmGfsS1B9YW
dCR2VfT+IKg7JvQESXKZDlX+kdwQPhyVfpzQXHavUq+/Mbh5xGyGVhQuhCPGAhz5
ZdYCPaDDGuiTE0HNJ3XemYwQmHyXzB3mkFKQgqhtn6TjbwcGQS7wZ9MDvK8E902V
GWdcPtzkshW0Zizf001Cat/UZT6hKhajuVilvIaJonv2GRobZvGhTzSfXzTm3nx5
n3ssBY5ZQumExa7afzza+1a6IcEqrbIChBTYbP+BaF/5kSDdRsZdyo8oBX6Kf7r/
dyP3mJL6wJkdJXPmy+biPGoKSnhjyS98gwx3oQKJ+VrAzoANuhKUX+xZ2L6iZb0Z
hSRM/D9E50TLSfcdYmbjZshXqYJeTS1q4GsTJOTUL1bkBPBxZ9J5HJbRTr/xFJ0x
sn6APvSUClazfCKXn3jNRBffl18JhAz6qBw+nG4efSeUzcOx6aPb8J/md7VjVSPq
M4LDUobtAIVPyS4YyHqtPas8Lf9vu9O0qXtD1h7sDemxpwvyKMAkA92AKQcoxETC
ZImm51f71NAp9j0BWrEPMS9VVud9JrGQhmodeOeo4LV+BZyJY2ZBXikChKpeJkR4
U+wuMc9SR10HFCorJNYOooyTPI3koe6f+DPisXGBKNMNix/vmlFmWAcVd92MjB38
J4vKUn92aGiMMY/JgIr506YU8A00rna8UT/6i55EVooJSIZEwsVHSNtbCbCZx9/m
HaA1AsY4YDqqnZ8aOWyJ9SdaMuzjE2anPUxmmkTGfRCDAEHeL2T2A8fDB4t8uYCy
rnygRx4HM6EVcSjRL3cZvFIZJtiSRR+pJ8fR90a+3NwSIxv3HdbgJJPQ3sBokgT2
RX1v3EngdIGY8KfC3LoLkjArG5Ga7YqRYq8XCdhjj7HfalIrLSvTvoISz7kUkOFQ
bvKKs+tmuwKPiYAt7dAviVE3NvCNPNJYBX/81rAk5yuJq27kfurzqgNeOfbS1ssc
4s9e/unTCMR93oTbZ4fW/DluDVHsyC+ide6RjlDXJugs/7o0zlFocKG8aTVGGBzH
aTcCUcDgUd8KCS5uh+2x7Otm3PTqplUYA7T4DH9m2AF43jxzbtlThRdoU62T+K68
sCqUY8a+cn7R3didtQQz/j9LEIaA8OSOHo34tN3Fd/5Wi32FjLNIGQMvIuF6Jd+6
nPrgLbN3aYx2Y55QCn9Fo6UJpH4bXWQyCup5Ra8maDbduw8FDuP+dx+2UGBtxYwt
RdMMwlJH2l+1cO5Ri/TV/n7YnigMeeMF6ZuHaoHEY2obXrO+GDp0DhSt1uCSJ+cU
oBwUAU5IrlnqTPa8W66b5BPAL5Pj3CsTgKJp5FEfb3m0wvLH8EfPP6AGLzOsNXfF
b1KiTXUJ/758/uyqjHMLDID2xyvZGdTSJHPJkL2dcmpDBuNVmoRK3vH6T+ZaS1Ao
IKrdN75YnyXsZgFxwESo/J2G8lsQA9E9cF8stXttv2jzJ6ToKlxw7XCgI1rDifZd
btaGn/YTydteXZU3HYDI+l1pSkO4G6sEwNgtOu+jjovC5kAsRV7/GKSK/TOkN9md
xmLhhpQtU6l4Dvx8bpiXTiPbU7UxazsPZo/znVHqXb8u1crC6FMjHUoevIlj3MgD
u5GiwEUR6grdUwPTB5y/Rx/vjd1ibqwBo5v3qZOrt3/TkZ9nFx0dTXba50ATZXB4
sAjD+s9YEMHRSHCrtNw6eM9m6qaRcDkGwd3gCl+BtPkCeIqBSHz9Xpe9696CdHy1
pFi/lRCU1b8Rv7Fwooav8qUosnjaU4+jbO8CK5bcBkwdSSC7EtEr3iQCbhoDg5yP
lH8ayllNwRg26YgPuKOYpxRYqjINGpn+Aa5CLvDrP1du374ETZsA+wHw/hovvYaR
Ok1/O09JZMIEGqEPJxWtGluoJlvnYjWqq8RbavuM5C9jc0jzrExj81CQsUxyUPZw
qMN0Mhn1/l0RjhEWIG7fnLqwVEJqryxWTSyaiCUeIAOXZGaeBIHTq0W69ll1cjhE
aGKKuUPwjsMb2nMchI5u96w7asPgG0r+czh6eAO/C2q/0nFG3+PA4JuR+MuXJaJf
qd3MBOKs3doKW+NK0ONKJPgI2WYuOFhuB/wd0YGEePFp+1z0NzQ6a1GytRvLgxuo
sIqv7LsXnSRXF7vUBBeKhOAKVAikfM/GCtz3/6UI8dhjwDQ5U1fHYI1a63asluI+
ehnyc7O4LidToPtqqCeFzoFF6DPcOucG8enaefA5mxfI9nP7HaqJxX81zLk8BGYL
bHhG+CIcs6qFT8g1DehzhH8E3LgL1g9+B5mPR+x03lNC0pKi2aaj21XfEMM4S0HN
29zZJGqp7sQkfeVLfUfwx8bSyqAZv32GkUVlDQlnvcoGApcTbcUanIF3dMKGv2Bw
VpxDwCzXaMVA6LRioh6o8cDiJ7vPXLumDmzkoq8q+BawR2+XlS8BtrNHk5216wp9
+CvJljRTHY0uJQhzO7yYVXi4VvCLsITKiXjmkCVzXueboPnBLqcdZtmyBqzJtwjd
`protect END_PROTECTED