-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
PpQ7GsVfSz4rHJcu/WmKwb2IHwKoJ5um7NOGXCeSqXxBEJFMH+EdyOJUXNonZaNE
+0C7oiPRJ/MhvYGR4i67xJzWJ+n0T6vjrKNmR2fD3dJrVo0FjlsP6v0uOy986Gaw
+rKkQEJtnxpWXOZ8eTKiCPZ/Gc/HtPVMo12Nk5sLvv9lM5fpBmKr8A==
--pragma protect end_key_block
--pragma protect digest_block
qAILkkczBlNYQ+YaUyOi9LESImQ=
--pragma protect end_digest_block
--pragma protect data_block
TjaAb5rYD3rEBz1OFoHKcPXPrxgoY/hLLWjupym2vjBj4wumXUY+3JlxZFX315TL
Lm4C5Au9OlzUDpBXxSeMdHNzHaklviow40B8C5M1iX33YdUeGx2fhnuOZyJdCkqO
EtmqpfjjsN2qaEGQj3CSBorP1DW63lYG95NQNyW9nbh9RkX33unsBgohjUthzkCV
t0gIZPmNCivyBB/Nmi+d8WS7NWwF+Gh3ToLOE1wlgGR+GPdbOvjpDIGukNogz0F6
4gZEdNYgZiOScD0XrBT7LE/fnU0aA5rgAAmQFC3g6xqW2jNKGTCB1bekymp5CxDi
6VeqGJ077Bzaod5TNcL7GO0eBYQygfSHXHMW5mBkJJq5uVOQQcIz08rIpumAC4zA
v40YjvhsyXiDTcBBR4ikOMpVL9VAFvPgqgdUq4f0IicwzKCr4Z//zwdEw7xSCdxV
I7kfXmMqRnkfEboNhgaMatBWJit7k7ehyY+Sz4Uo15lSXhmQNfztvnEpNUS1wHhz
KeAkspokfXanhhDI587VB8eQPE/Dc7Tswk0kowZpI/nqVCOuNwkGpEaxO2JYRvtl
C7kRVTto3vXxj/TjVJSkPlsmvgnDqJ19ONaKn+U0t2GgDV6lQW4SoyeugygF9BF/
zOMJ2nm94+v9z1FQJfoi6akAVkmyQ0jP9+7xbmaHBu7K1t8l+h/hwZ3VqtQlDCq3
3gCZlmA1SPfeTm04Mhl1HXqDzaxQ757NG/FRZ0I/f6O03+lXBMonIe8z6imLLHvi
gQ87L+R8L74HoRQ1x2gRa3pldeR7qM6lJDCE9Ez0zfpk82ay+nVkNa5OPqeyBBQ1
7muH615dAhC9bYkHQWFIfOQqLveg5OheDjx7RSZCxA03FKVPIfImE0BGUBkibsq+
ovjpO2088ARo2Zb4eNtT4m9IAU1/IAxIlJjsp2pfHjHh92/uIDVvnw2jEj3rAssG
/UuTXNxLQimv3TutZUuZS8sxz5YuO60TxnSLZMuqfAfpesFatmKb0OT/WigHtlkg
LeobnLuzQOXbFVXCB6N11kFWKmkTOSR92ipUzAvadfXoCbZEeW9lBawFdxZSjVNh
628n+N1vOr5Pr1df0I61D0GrzvgOns+AkVR0DqJ1n9ERZHxTpjVLe3abrxmgkGUb
o1rJssZejbtZTUllVDfO1jxrRxSY1Vj2RUdSN0OfSn2g9S4jFNRDPGSJm8KV26K9
WyBQ1Z2aJJVdbzZrjPoDPinRGht1ZNIsopOhmHFz8XLZCMAhU8cVoqPbK0YZM8dZ
DKmiFqAF6QURiYfe6hF8K1Q6F25QxspHNfMAUxlr47ggFKhdi4Fap2cLdSrgOXlT
6EjRHolDr+eYTQp04BloTnZbLRxyTzrp0eQTYQbUcK+nBCEC0s4/NUx+kmRk6M36
u6IMQQeaCfIOrQVylgRp7GcKjvrKHKDlHs/hbXbwDNQIuFRY+K+iZRwoMjvSIF2Y
dEVRU7YD62Iml+W0TdwOBuM1Q5wtPO0g7W7v2uVgeKE9sLg8q/n5HTcZOVf77rG0
JFIucwY8Qj9mFvB5UimEMaozadigq5rN/A4zuZLiQfyoC65MeElAsxCyDmYTQAa6
YW5ufcQAOqD52dkBJ317wF7JCCmcdzs8e/zLglpB1ZfdfvB3i2Q/IUt8tuyG8yos
ILPMFCxT8Pw09ch5tSgaiMDhngIdByFjVxbWqH7EZGh0lLZeUa0WMg9/jbrBX175
zw9XdGfgjrEsrVnT+zFW4ufgVGH9b3jkIXS05P1dfWBUCEOzdRNMcpIeq2VzIIO+
vNLxQEDkFAfrlUeVy1Tz8eMMfg2suuYtnbSVENDlirhqBnvhqsxcTbl4ojPHr6ps
AtoFF2qgduuXmS5K4PpzPr4liROApWRJTFEQ398CoJzubQcupqf8qAFAP0QHh+Uz
aMsoGgOpjF03K7dn9w2NHyR9xNaBE4a0L5fJityF2MThwo6M/L91SZRfmKH4+TXd
FLXjAJijxloT1zncrAPgX1zxNnEY7C1E8FgdDKKU2wrfO1SZi89Hp6cVxZYqC/4B
FH9xqEwA+yAFNljgKcqgL2JE3bvK6gqo0tmnd502epqe84QuEw4vzlVX2m+zc376
1KHiaNnkU7jKmpUHUBO+y+8dVm9DbZzZMqAGu0lExn5Y5N14wSGQ8QPv/r18yBOA
bZ5AX3/fFkA3AsGcfAvwvraJ7tgBhsrPrB3BKG4/OjdNhxGVsfA+Y1AarwULzomD
XEL/kS4sOF0+BRWaNBWdt1ZiXDEywm3yYkr1Vmd4Efx26cZmE2U8KyUvtAT7gYh6
DhvjYri0dD3rfwsoZqrrl4luugEWgaB/32z82agqBY8+77227O/qaMFPE7GY90Mk
CbsAsYy0XslYOtqq58BlKG2oU3+fHvWf2PnFsHS+HXVGT/CwnDB0WMhJse2rzeRK
qVJGUlrgZeFRnBgIEJZZtV2cIII6V/Vjy2xbsy7S3y8XEoGvcWBBGc6CDR9iDEQu
5T6CQ4WzKT1ZOpCQMkCGCQtSKO5WliZ/YJ9586cx2YEQnJkoA1JWqN8s6GbjhiBz
/SK+QaIRUrl6ODu4sO9yQYbp5DYPSJ6yofQB3AgdMGNH60K9NJeaKWl0+N0NGX89
kIIdDIxjPTz9J4gb2erNF07NDbp0ktSrXhahem916sGdkYvJyGE/aLpBmVyXTpZd
feVulsupg0i54xO9HOmGbPCp8fuTGOLr+ygjhbWJpiNPYsUYuMwDIRQbkvQ0S3jf
XWGJZOQHmgFE7uywxeDF9ZCwCTCIDWU2VIf/94RurXx/NMrt5VSra+g57SGM9J0m
ZEyXdfagWjxkydY8r1mAZWSDJwnbXCYanWlfU7IdeecfKMO4WZzDXH+2AYzptgTq
DDdHuboYmXbyp+9zSznPysUUr0nhmgOzq+jK1O+zAJnjLu3ill3SyLQNpeuUo6mR
M7X3FvAApnFgjVpX72Aj2jxwydeGbgGANKLibR6cUweU3b/cNV2ANIQ1epPJbGte
1lVQCiFBR1o3grpH5R8mf7hH3n7H+kBHMeKAFIesa7IoY+f1XHQ98/YgUhnYdbM7
IgQ9PqTJ7IP51zgiv+dRheHgHtTsCcOQoHCADqzRJ2LZJIAr1GN8G2zTt1ivBztF
H7Q3sSGNJeu3UAl36eXdXC9HReJIGyg/l4TTK+/S3rAjqLIpLooWgqTe/o/beZCy
cDH6aTftZoeMiAj6XAmTLCqSaWYzx1GzRfTbt9vphvBPrFA6iQnORQ/UTFbf96kD
MgkGRQlm4QOQxRDj7cUQps5a5iTdaqUB6vaFdOWjb2SDcEo18Cfdr/xFkF0iBslt
1tWS0KO8m2digARgEmiBQnZHew5ffvBh5MeyLh6KexoZK1EmYHAYWxB9Q9dqdVs+
wbWtvfFg6Bs0v4kj3BcjI3PyWRcwQEyk6M9X32VGUNKeNnEdK5f8wA1fgNcSvLcF
nsy2a+bHV/xTZw3fNOnjpEDQeK86e4XICaAhc50ZTbek+gtrvaiFmuiOJu9lLHrP
0i8rWrjHM5i3GcCYhNuiMIgLSPdNGRC5PvkjV16zim24+vQuWU6tHlUhUWCpc2DT
Bg/Q5SHZ5skyZaKvZnYYWd5+4bdSzKZLFJpRsgXoZTLHUxZTCqe1G1oQTgsrjm5K
mJ9Nl937LbgddESzujOCnKAJpNOOQ9+SdAAOxBQ+3izacoZRwNhPVymtxW2W188o
JLfscYyNaKcLgAPQ4cadNRnDaz0VCtCmhP/DYlgPVLzKAUKR0QeqY0+mXIn3SZg7
W9QUO2lkmm3VCelVIpN4qE8xFUqTbxXyYJNRd/jLxqccrYowVUTR2OuNOe9nYD7/
LMPsNQeF7sH/ehAPRGY59aiW49KCXhW3SUVtuy8iK5y9lSiUlWU0Ia5zNjdomvs5
O4G6lmy+nn0KsENCDaZ1paK3EWIOJvRFMZ2A9AaBLOeDfGVDFPLdneKK88/fZoA5
kVtjIe2Iqey6R7YD3CDJSDE7jWbKgJINSmDp/3pCbRUg25SD/Rt5m/tXQgH+uaY6
LYFtREYUoewMnzAziSHcjyFHdrGbRfk1mOLs0F0BfhjQ8x3Ktcx6T0RZqjVQcsFT
FJdXQ82Hynn+RXBslVKglN/wPcuVzmouSTkzTSJ9wsynefxlIQ+CgD3hBgWSPLOd
47OZ3OV+q4+cAFRFOJN0zLvblZXIrlA74BovKZACm5AeAMF1CPfxIiwp1yj+N5KO
JCAl4x68CTckCD8g/eocpC7jp8P6RD1mWIXGokRVdTZ8IPuCvvCbT/buBJGIjNN7
9TJ8KnF8SZ3OJVw2MB1KLTFJPHjPWcgvwS4Qom1DDG08BZtBvgr8mwO4V2RxtW/G
MM+yPxjNqxyUQ9nzGnyqxUTnoCb7NP5vr8AV27fzbJ1ax8mwQBM6W5NPavA56gtP
SaaLuf911yzu+ayky3nZ5kNlACXtsYx7rwadLUE8HUwmHCJAUf/cISk3akUhSgxb
BtF6xAzYGLFDbd80fxmGjkNnW7khrHYymQkwf1Q/qfbvMIe7dIYQcRxn7rIMzYGh
wFfLBedVbqB2Ktv/Y08si5yt5p77FTrYGNeFGkEgXYP47V0v1NSj+4t9xwfl4P9p
JLdhASYoHX11Odo78CcFWieEuHMvDek6NGRoOuLfA/lP0Ylbbj/pg/v672KHehGe
4uF1vYX0ta5OgTO/3ywLLW66O7NHaMzg4AlsRQfXPt5BiDLwyhx771YPSO3vSpbr
jSb/A7r099ug5Kl/J82tXkmSFh6pBKlyuwEDb4MIFn423r2IAHWulMMZ/TXdfpoO
V8KD0wAJo+WFEA1f0BpR8AVG4lBy3MZmy8ul7r+hhJPiV1D8lKs1MnoaTjhYRghT
idsE0fMlFptaIH0dUJ/CNEpSFyqHh7IsVNBo8SwYAya12kT1D3UUXunDWWmI1x/v
fjd4oen6QLsr6V0UsqwYr+8cacCbFz9jPr5MZX/JeSOaf1OUXranTVYAtTPzOWIB
1pYDXTBsmFOeGjAT/O09KvAvpoak7WRBI//hdGrW7oKUHctguXurkFCatCghxbTO
Ls6SsKJPv3g281/FnFbLOgrLD6CApGK+0IMNXmmZG3IxNnHABFYkhBq5wiUQwbNS
7UrlVebXOk14QEOaRAodwq8L+i6busFg2JgQRnk+3CJ8EM952oEyxXQBD9VQMljx
h4B+10c3x12FAFxs8DuyLVRMhXLt5EeLA3jAnLfM/ak6l4VhUKKRHgV7rG9MtuWI
Z5tiJMp8cHU872yCU5ZAgiiBeytZWKKuREWi7izcs+ae7hHJ1iyEYOpGqyvGcX8g
Yvtiwb1E68ezykWkIm7aHRtoUb41sVIpnin/fgTdsIpRBPZHDP167H6ONpLc58Se
rBHtP/WhMjz4cdEWpHhGal48ztqbZifIy9mobxJYNMdcuW5AUY/aG+LQ/CRIM5J5
Lpccn05COxTombt7kn2cBE9svklox7znNpFKKsxF+Uj3WYGQDumhlaKZtAzY518/
3tBdZmuhDe36KXyhA6F47e3X9YYdmHxPot5ymkZZ4ONHTxdRKuzu7XAmbaDiISFb
waa1frx6UAL/Z3YQrVQyozWBvnqX4MmNQMqL0vPCm+OB97gOVR+r4w7u0PCmxNxT
FxK4+pJ9LihH3Gg0iTU1a+RnqLdQqp/V6qP/BHj7tBUk+b3lMY0DWtqJHkh82HRI
XyxKi+tQocrG++NWRNAEsxAvYTQyq4dj2wJOU78KM04o9uRI6fuvR5ke2zXN6obq
7pBmxLfVAudR6DVx/BuLDc04tSp9jNuqVvPDkT+VklMvv6VGYDlYdnqUIIZYJ9Pi
zAcIC3KtyGujZDKP2W5oN4gKjJRmushOCTeCbSEFrsZhGXQvMQEVoOOK92auBzJJ
Xf0az9cBuIV2fPR42W+d9xvmfNsHmaH9yn08kdG+JYr5YOHkB/BCjuMjtrqc1C8c
L4g4dYmr5IlaztGbGKMvzyQ2wYCjsMZ04wzH5IVH81wRdud9ril9QNg/6wtN1it2
kRU8mDiliYvR+SLs8VT2XbWqPkITNMTSxzZu01XC6gcKERaOMB8mzxF2Nssd8x/X
9QVyBPwdsFKmxJMrqCAaOls1g7zCdfjD2b5zcb2lkUbc3LAqb7ijgolKAeg4FTIL
+3Wfm2G4iulpo/kPVDkM9MGFA6AcBvhsVTAN6ApCpYxiqi3ylArGr+ktQqYMwjW4
7tH1dsRIO1FzgB0ozCZ/0qVMxAYavcmz4Qi2E4xLyUAaXLK8/iAbqwQoJEuAg1PN
qz3eBgEWjdGcHsA1GJT4hFoAbNKZOms90dCKTrPgy1cqglIYsoi5oU2wXO2NUYTL
MCv2jDg8mXFTOuYBxfr0GE7g6ODQ5qqG9WWQNzG8NVgMVnglIcbZTmVxU8UFMRAv
HeAeFXF36GNcN+vQenSd2aGFK51p5p8IcdeWvp1j/X4dFwOWuxndl8ZHh0DsebhB
rezHHL7piE94ScC5EpLFDZzTke7VKEMRrN0IvhoiC2yZRmVRdd5DLN8EW6OWtkUv
uWaeVcga2yDTtxLD7Y1sgkqWwcN4vCCNQYM1zN4ehUoPkHAmGTWBU6OmzBhjh19z
OHgHkwXjE1nf0naXUxEB+m24C4Vc/vl+vSXIdXaYe9APapCkdcfljBF1yQ++e0Yq
wztoLLVh1WgLxNKTV42TwT4r85VysiX6bHY7lk0OVMveCWBoycysTeOhvFU5eLMr
HFtxsPcf0mNNI0oe7H5tQ9z7f6iea39bHglNbgA7d/ZoI53ylsd3cVmA8BgFEb+r
Y8aTYqXde5deslAmkF65/MkCpjJ4nUWZ0R2eOy5BU5ofClmQTCajlpFK5bGQlOno
IaDWMnU+rlvTK8swZTyja4gcsQIGYYP1F9i9wIx4VodBs2PeMakJC32owXPv7YOH
S63gN65dnRpjBa6wkpJQDyFx/otRuL79EvSupn/gDWoWLYQhEvIllyVPu+OWphBm
VhN0fCgxcXetXcN0xULJiVoJugMAsZfR5ZwHfMcX1wVbVYctakHy+1DkUCG/94uH
lhTKcdfsHxcryIuzzCF2l1eLJ0fys84pe4fJgk6BwKezfgTo2APXkjlm5j7okc+C
rwuyyKfh/11SuNNRusNB8HZXWnaUCfwxXeHp1G151hhmM8kSsE4syXxEerK0GHcP
Bn9otWnFIgCOYFGHqUOkOAyTZAOAdhpSb41LjIm4ByD83IqyIfoPcfPWgeLWxDM6
mTfl8b8Cz1/3Jav0dfCm3DANasLYi2wXtwL6p0E9MdKjo3bHnupvb46g/Z6/LxJ/
/o1Ca4AQ47RfOaGcULWW72CEAqjLpxUkdZnkdoHRHrqH3N4281lkt28t1RGGjYQl
sZeoATUkUXBtt+z/XCBB9dt1e77CxzGZ5nMqbKBVCuLQLx+g6hQQTYJ/GAb58PvB
6xBybteSEB1ixZZD2opZ3qF7vdsEMOA2HVNoW+VLUPuMaXSYy6WWi5x3bLZJdMQY
3EjAon7s2nAowRRTodByx6Hd2dfM/k82xRxr3jPj3L9x49BDAK46oSGamV3DR/Fb
AwPIiVnYpn68A60vWK3+1+G+JEYexmbhaEwGm3plYibIeTDV1QUT1r6ZbvKAa9QZ
muXPCPXRTQhKwCSs73Z7IfrCq1aBQdVi5PNaSq2f8cjOAYRdTxAgXIylGYIXtzoc
lU2Gil9S2fRP2nqhDQsXnGOID9jaBrbox6dzIGZ8yecA6IywsyAajfvCVvoMaq5L
ClbtOu2woU5z+puDVbgXYr/auOxcDWM+YknSiFFwfAjP/IC/woYylezVAYn2vIMG
5dgkMq50PRez0P8i0F7yqTeN3vos2wLPVE0aobpNJ0SRIAALip7u0JO3dx6LRS2q
WSS2AcKCZajLq+kGSN3/gAL1AdnxXnBcJL8+0Curc4zk0c9k0khYsV2PTKjXy3Wy
8YPJSRwmHQdP39VFH0lRmIEv5HD6e/H2W3Z6rPnCX379EMMGMTxE4soKDg1xPaBF
Uu2T98dZry9Dz9VT0ospqN7+g7ukmch97rGBXRklzpcvW1D8nzrAIxVVjuNQXR2s
Pbi5N9NXIjMI3BcYBJV6QODlhIrZoCzN/QGXxqN0JzX2hbSLALBlKDalB5D8GbYJ
EdIy2k8egn/2K/cW/zmyRnrVmAPmFWUJAR8v+JHvVJocq4tDY5Rb/pFbTRkyTeTQ
lyrNbppstp0cShtlfRn4G+rpITDNab8YGiv8cCCLimZuLxeZ4Bdk6seAaVge/Nxf
R+NNjPse0RIXCmTXBowS69tqS3tHKImOE33mnPgXT3yZtfgyC+koEx6CxyfmNO3b
sO+kgokl8PGjSZ1qo6nmfAZi8h80auAO2CH3Dhd1olOuKMCWEfO5UV1XOtAHjdLU
8t6r1n6phbmDJfjOz1DaNW0F/VpB1geqjl3tJ1msn6HxbpCLxvnJK89crGkIgX4R
J1Lrhi5FyxZeobeECExm6cp4BZzBwunvWUtv03cJDwU3LgSKeDnJBzz6081oHPTT
rVng4uu74eoaOFJ0uy+T03ywwma43JCDdJe/K9Jl0vT+GhwZauOAMvd4PIUh8nAG
wQjZVXJFPtc2oi3BlxbcD5zZYCFmTJ2RETHmQcZ79urKhP4qrHvW4gKlDTFIMPPV
krQJZ2TRKlw8J0ggW65Ip1CNulAbjd2NWBLQbfVB1LIr+rPIjhXN7pMi522Pp8jX
FBnoFi3ioCaRt/3g1T7jgjfo1nb5D2gNVnPurX35DDsIj58MXsFgBJNEvVCCexmx
O4p2P0IhB1iYtHLs0Wx5vhly0b9PXfW02Kq6VLjHkCjLu+NxCBj2oexG/EHSLoLT
oMPadLLmfhsMBlBr+56MmGn/KXzTYFD6ZSacqpLn+zlQn2Yhulw4DJ99LB3YVo7R
GUcX6MbfWk4StIH4Y9JmT9NaPcUj9ov68auxkNrLZOZSWSdambnPcNwB/K/MXWjr
JFoiWsNkY3oAPLvZJFRRgeMWyV3kwkIxN86LShhXfsGgC2Heq0E1ZNYDO3itJpwf
asYgJn/y4FrBKzsDk4EqOAzxcwNwsToVRz7CI5BiwEXeQ+9o0rBLRkjkRedsG13I
hdMvM2i+n6qBzi+32TOA3Fvs1ieFBFCLq6gGdUmK1MU0MqzGd87wfv4AUGAhWFk9
j/pJ+mVabQMnclwGpyA4+yzxxWqGzP2Y66RpMstzoce9Z2rL6AGtZwTZWVmHZHsJ
H1DN4Nwj+aAj6uS1dCTr/LZITIButz1zxR+txhX5Yq/YRkPdYGeb8ZBGX0ZNhSuz
4QeZKfbQ5V2j+YHiS7i6zd5OB79MCV1zCCGaT0P3oErFuF5srhCclvTLqBpDFfnw
4+mWtLQZbD4I3+yrREo9MZIgjEkdL4sZDZLddhZYKMvybnYTLo8o87fa1QBGJSOf
geBzzXjUcTCHfvZfvXOkCqK9FMbpjDmWNpElm9Uo0G1UtU54tH4h28/dySVFmczP
1UBdZMVJaJEHHqaLS/9wHE5JB6Dfp4/JV57OfZS0uDL91GR6MzrLhlkeOasspMnZ
BCHzzGnfamerSzH/Y7FrBVdbtOnFj3l+NiDyFwnlInUGvoQbRVMyHsvNkDF+G8WT
ldejpytGFwVdgLj54jbfpYJ6PyE4C0pIiQ2Bu5QChibqDHaJHNN9UR0uko3LHucd
3VtbVLAsowEy0q6KvXLrutLDz2lITXnUQnaeL+RpsN4MzX/dpSH2Asfrq8U7VYsh
j7edkUOCBYqqycWW9vWAzDfWk4A7cteElX/TS0u3MlFmH1dhiaNz/C+fa01vvrEA
SACdnAtQMyrMhV9u4XGWGVp7YjcW8jZtRIEL1xw4r/3m/poOHXeeApFBU/rN3U/Q
8goG9q00c1szDhqydczTgqwo+Lt+z8e1uOp8cG3ZMN+RCb79iq6ow5pXcUPnMhQN
nv8V6CdXJfK17ZL9eABBJTaMWvW9XOeiL7GJbBpF3vwbmVgUlYgL4R7wxK0WsqY9
nSrBbgLDIzTrlKYoJwPmPy+hy2wEYYEfaqDd/3/M8cGy2wJP1pfRvLyOPpridKbI
5m4FCuDPXFIuqa6hxkpou6vsKAxX64RuB4q3TOmU9rNOrc3thGlFsjlHQrL3q4DO
9vXkgPHqbtm5JCgCr34RPtnHClbtkL2uVVQH7s6Moj7uvhRE/SmV3dVwQPsCr2yM
SoMnRMvqlStGXQfXHA/qC+AntcoYutKZZ8ut9E7f7R+iykzsRVbY3xcEf29mk+HN
XB1KoUF5YGvT6OxuaX9DSp3fNEQrmQYVfgqq2dJTF/X4YhIae2cyNia4NznhkdeL
uH0CCCf3n6OfyHs+QUZGmHcA/QdO1NaiSERTZ4NueeXrA4FknYZJX9xewIJD+sIh
eQl5duGzKTwYuxJMW0Hl8v+KFkknSSHnDFzG9rHMgmqS+Z2yijWczJ+aco2pNKmN
OWRiQk36Hnj4U+ZCG9jfbF0lkiyVaCCNKRdrN6Lp9jDVwQYcqyq0LEnM0JPtd5C3
AXMnh3EcipryVaB3PS9wb4ZPK8mLInVDMw4UQ947r0Q5BATmx4q1t4Aby2LLc+RP
m44Smg9lx/YoM7ADHFHM7wi6wOL1WZKSSFGdX+Z9bV/QdqyUMDa3X6wwpvVxs28j
SCgrANJV6BOUDW0KYcPSGcrxO0kYCj1TItzL8ULs8YETb9BsYoMyz9VOlMIy7U8B
Idf5zOot+kbvHtJfm6EveEO4G80KWVkafl5PBtTHoo867QhpzG+9zZN/wFf5VeAS
CzoFox0A/WVbpXAwViy0S6XDbMkCB5iif/Z2q3c4xYwTQeefD2/6a5Mejl7fp1A2
crTULG48L8WMHD6ttQicYw4bHyzCNjcmlqZMIHQyWmomkWaHgAoEXZM3tuscZT4k
+bRWIS+NGYmDlBiPmcdyLBRFSxqoXeWTJ6JhktAKgmHKXREWpNUmRgXi7xSRim6P
hGoGaZD3/7bSF6KXo2YBRiINw0xMe6qwMsaMmvFhHnzPfz4EfJDA+CRHYx2lJU3M
fHGmdLxlXg+xeNlhqUCrsDw2ylq81UHsN90emAq6pr4AqhhyUnU+AX6/0Zd/C5Dk
GTWCJkGe9JCvrY2scseVnm6+EWv8ORAYNSv4c/zW+nTxSsNYauK67OsK5WxGQ+cO
SxJY4WB+rCN2a0Oimf5l9oTfN/l3DAKoSpuMd+WCuqx5rB3YQjg0ISolqNp8CoW+
c4etIqmbsmpcl0bLqOXyJTyKbEiR/TCSK8LEm+pbcGMZhcNrRJssT1Rb+jk9lUH0
tw1y5sLHf3wgIPwFmVtjzEsSaYCHU80aO8ssMDcsYddCcjba4hO0LZdrTJWaw+aH
ltpuhio4YAB74gguCWaQ3oJ+ZTnIvsj723kAhjnMJmqOwpD9GujW4G/zvqSk7iFt
yNxDPQ4yMO84qh6IU9i+YcrYOnTjB/zeycmiuf36q6JsuRbcYVLKHd2XKGa6oJ7X
TrjQWzYxBMNJSn9Qx41eMjesh85D4Ngs0SWigvJZmsMdYGq/AcPFVOyC9Dxv2ywC
TrXCf7raOgBJnHqZBeyq7rqkJtK2ty5kQufzqqBsnJFtkVJYIcbGI0lI8imcSElh
rW8lv4fF5j7NKtOGzhuOiV0KqQyUTax9EMLYPJ1nZXONpN/QV9BBuvC9d6R9Qvn4
3L24uirN3CgoawjxugPRaFsvLOBlFyMdcUY6Xke11IzdQRDxvzBrlJmIlC+UDBQy
CstKqauR5eb8eiqqixQ8q/EFBTf0xRPkaXeShxYqHr3UrnzNGBhgHN4su/FgrfyU
7JReIBKrZfsW3FkP6dvy/eMLJsOowU8cteB/d5Fx0cG6Vc1o8PdrC0dxZmx9u7/R
4zMSSl8dQP4M/FKkoizFbii7wALHSwBp88ptx1mcvz5kH7dqhw1ydamYaFs9ZY84
pcBwOYQZfHss4GSAgOj1yEXL2LjASz+NmYD6MlIzxlppn9MY0ZNrZymgwaBkP1mF
nfRdJ+JRWjF+0MQ6stgbJbnimwxQFDHu9e+e/MGwD4l/UfU+jY1ySDWRtquwP36E
e1OVikVtsZU+RlYxZ1vXpDTZ3UZtujnsbMtR2Qxx7jg6BSscZ78pyM7YsUu/fEVK
z920W2kz8uvA+VRJqnnujLGc8PqW1yGRQuqb/MJquUl/EW9Dn1vKL4INuNfBqaP2
e1mw1rA057dMquxGvo3s+HDlcHcAe77WjP9UVLR7uJQPtPSMHFjX/F3iOW30gkGC
GdKgv1flLITGfcxTPDddW166Pf/KLCLKjdjW732/anEGyQCT4rKKnJUGBUUY+KlQ
WvWtQvX9T/sRWIPUqY+sTO7CmyIZNCZxThik7a5OHjfwWPaU8RYIs1gyGdnfn7mr
x1BS0IyX0t3o9umcj2nr1bCtbESjiT010aJihl5qny1kV3jCcGBqCGwNRnDdCXpQ
c9ZHnS32d5B44I7jp1sxCqT8W/8ZXOo0l/zSDDCd1oCBezBYCOiI+vk+l09ysFwA
1jVSL0z1BPuG/8ScOktIMrbq6JtCXgeWBU/Y1+sfkw96P6mYGhoU+SYe/Jgmj+za
zXVUL3clR3kieZWcBPL2cq9Tt99Xaa0GORbdU1uH3U98C3Hub0JD3FQiKr+gf7Gp
nMjuiP2fyTLckdK53RCy5A==
--pragma protect end_data_block
--pragma protect digest_block
XHa9e44YOyYkzZ8lQ1wtz7CZHRk=
--pragma protect end_digest_block
--pragma protect end_protected
