-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
d55TsRioo17vYZod7USxSGIv7d3A9uXKXXDJgNhJ9J8MLY65e+W6jlQSJzu87ojs
KY1xSM8we5kzxDd5T3GeyNxjTRgTJzWSv/fdKL5z79o6d44RPwHlHOpz83Ou6Nl/
DveQZwAo0aulQ64grYvi1uAtP+xNFRKDHvK/hLXDVqmfC5NqG1aS8g==
--pragma protect end_key_block
--pragma protect digest_block
+Khtb8vFcS+LzW8EeBH8ts5lSIg=
--pragma protect end_digest_block
--pragma protect data_block
aojYjONw/em0nPSTLjqn8MbfOeceMtmmyv/EvHqDYD24o/K1AWbUpH0uMv1dtAZ5
F973UsNt+N9tqUR61omKa6FNxOAvNZ5alhrdwqqq3IHJq6STFtFs3SnAHeXuTF0P
ogbphSjdpz7Rt8ZiC2w2+ecp6/gOG/fM7Y90NyvC4pr0cmmjcSKFCh20FWBmYje7
5uGTaezTFK3DQrq8xRV82WgmcPJQmt//E1qSF1AuV4dTtffvDuOkyE4E4smnQpC4
3qCtlWKwQLKBXJ3uKfg0M/QCXz5xl2kXG+f3OQ75kpmY5ePZyLxeVGPTkXjKsxn+
N+u1dLneAu9YV+waXuXKhwekCjwLDAsBKADeyZ7GOph3utjmXsPbgB7xINKolDIC
Zau4CKJUQmMJXtZgpUqMWign4BuJbn5dw/2pwarexDeJ+4XHk7KSz9h2j3yZgWJ/
93egMuki8egvu1rqekeyg1UMHtBETbuCUrFq14F8qvrF1js6ygw1vNEMY7BFnqZD
FBuiOZOrzXEnIQFQcCBF8wo4RgUkW6WO3eFdXHrPkvTMfca1MTBBRnQIG35Zdl+g
auki6tgjXPFgW0em9t6HGFs4aV+SJTJnc6jHSkkOM8XQTf/lu9pWEcVNA4gu8/KE
BXev7mk8zPQIxZ9lHB/GWTSG8ygibvddWQsf2J1UW8OuGACdoeFT2xUXydEbmwXF
li3X/ZaHh+G1HBjATHrRkf5dHyob3UFOeBYXh2o4IKT0cY6kAJeu2gAXbvuQKmce
k2qXGgTPIDuc6B+S2T1bpU5pI4/KCzywlwW9yyKNidOF7GBu5VHLb1AK/OxJN8PT
bFhBd0/ufxYN8SOm/h0lceemOZMYn/GQY4uScu0M0mKEx+xvcq8SiLtUdZGqdlo0
hfiNhBM2cL33OSbbd8vrrUDc2XWYJ+oiBHDBAAGWYarQnEBv2glxjWpH/Fkm1y+b
jyculIF0F4pXnETPqvbpG+otTkM7fJF1e7RTOmyscQL54deFGwBYIDu1cTyola7w
pDEXhSTs8FfXI0+Gjq9y6TwhuuSKwAlRZhmDfAaiClHz8+WGsOyZBFKen2at9RlX
ERoshdZ2xwsKdOapqPL4Uu+8OtXlbCttlNQsrSuZd5V/YDhkSlglP5EJSOuK4oq8
vHAnRgvfnbk9MpRibs1+Xb/DGIFMFmBDQmBz6imKz7MSsxwEZeYZu1qQadU3U1qe
7pOZTNHuHjPmUOw38zBSIcvBxFIMUW1ack8FsbV2tsAFt2x8tfiEfTPYesJNAwRD
PqDknXbJJUWGGN+JLTb3TimaLNRIFzlx3Vh34nIXVHLpT1m7Tt56x/d/K+LMg6tG
3RWmwQd6gLRPBWZEJn6zDjR7dyDGa+Yr4WGuhB9laDwx/laSAd5NYekS1BFYlKn/
nv8ilTE60M9tburOMALvbQSCEKBvq7w21oW8u7OxefYM97wS1xkpOW1++6uWA3Uv
PSJnV6zTYH7HGgk9h/VEWCdQUkHVwARkiETOuXcHQopzOb7Ql+cQwgI/XbG3jaXq
at6OXvjy1U3+zA49kTkG0o0Ujyig/UPyhVzZHdRRyLUiGko4FeKW4ZhDrZnXxC8A
SICNI9+8Vs9eaM8PgshJzERHzWeTo8vli2R8+qQLPIBVWiKVmHofZjeCj8zdtzGt
ds73w7wl+JT3vPiLRZCwteMFBf7UaFd6dJ72AG/EmgOw0EMXOD+yVKCy5cg2rcts
9+IbPUu9htznapHmYKJdDWGO6RDgpRywyCG3r8mVo9mYksF1x7gwvwmWD9puuP4p
wEejtOhfLCvzQYBRme+LcnEELJPWWT5XYvGaTHAkXvm1ynNTuFwxpHwD/f2m7J8G
RApoBTkioC8X7FLFuDSMxhAReobe27Z+UpSgwZGQsYZxHzTzxDFlhx91dGlb/RPV
oWm/WBJNbuDCKHqmteuZrismK/aOmismIrw9I3FNxBLtdR+6c3h2aa58NkKXPryK
J0pm/3kmVN+267jEAXqeDj/AZKWANxp9Yr88+DCbmI03gNsshS4YmPJyoyQNgphI
s+l0pOB+BJfosRfu7m8qO1goL8fwTsT+R65up2x8oW6kThlVe3TJ3XJeCD/0bLE2
M6ZeSs+opXpT+kU+s0VJiFXWbrYXwk77k/6MIaQDhXC4+Kfwkjp+l/74ujKXVH6N
vLsFRdHZ3B9FYvPbmKpgb9oITwE0SPCPQPoM5wuf/qfDysdDeXh7d3BnvYGN1Qqq
ycEpDVf9Ojz+LS/dN0TkljuhnSTwqRw7+UovWyr3Ng0VXADQBht//jySFzTc1tnH
YA4YL9Jn5kfXH5YPMXNwPEym3+BKueLhWbXOXpeZXh73SR6TUx6Mkly3Ak/qsYyH
V3g5C4Zu67mqiO7gnLd+KtANuLjGOP3nvrWluDLwuRQS3cOnvqWmLqwLKcVqFCwj
6PEn4UvuDZDRw6+tHidPBVlpKoCGSnkhVDG0NJJCuTuENorxtepZH5vY0VYAe909
8qxTlroke84HtrTYUDa76UENbjYDLiE5VdHUjToQK3gvBGrMCCCOD5qM4bsep6Nh
1T7TlB+AbZwGg5Rumb69qNVBquAZsDqKJWGlDPfvOZtMNMl63zj52AJuVm5JDl3y
5IMVtdzY0zKQ1zbr+QWSlTICj/EeYn0RcrsHLuYQwlw5oUzW6bM2/N2G0Ikn1D7A
VaiDWDlyvdHdtM86rV2sDDv/3uiEA34R/bp/fkDCcN1FnAVr+6dJf2mSI/JoL0NR
BlTnRK2qYV+ub4zg6pfomxwnesD8x0jVcc5+98kmmbYgsZyTAXTmlKTbCC3zg4lH
ZpzQRQJtolifV3qU2ZKdTt+oTiKOCVBYtqKUUbr2oPa1Ex6u/7AbEycrqGfHniM5
RRkN4/8I1ZlpeDK79OmrpoSnd4FBmoAyjxxfXyCjVAZEogNkBYWAi7mLblRSrIlL
Jal6RK3xS0f3HpJ6PLkMlxYFz5fVSN2QeQ66D2ijnkowzhk9LKUVghp0e2A3SkuE
rRoAiMxW2A1gZk/P0UiK1USmAHaeqDDUgy4Y4fQPUGT0dv3WakV1WOEQcjJghsmR
n16SfQbIKMfiAUTASR7kTX/BEu08mp50LpGJnhB9cveSxX5UKR3Z+zFGJTXLx9N/
MAJ+rnUYWg7cIjR4dqWNTtbqCZVh5ja4hqUYC2pLM/MqrMqvLJI3tvjYH4QNmPT8
IstnQqEQoHOvI/glNHnC7KgQFl+VDfVMHQPjfrynJXXIFYgH4F5Nku215TnOI555
BGXudT/J3JHsvvjsq6X96mqIfLqNeb6oBVeMI7rBahmVhYAX5ElfEDhffWQ52iGL
0C+vaZDgKAhN7gUDO5aPmB5yUkOs/O1Oq1wxKX3kZ+iAfjA1PBFyVLe51pWDeTOv
IMJIazmryCQxHaPVUR1S4mExeDJ3jcGo+QxahrSjf94TGTl7QRvEQLHXHjOz6DBQ
fcXj/khalyJ4oYnMpzQN9fca6yLdb5ObrzNZlUU7KdGu6txKaTe1RVnHyVKmDBrb
jgxC9oU5B3li40uz5zzNGTIH2pySH+15sr9BGT7fGYAY6z7E6iug5g6V6qouGFiG
bPy76jTQolzIQAYiIhuV15UlTr39m177GyO8uB512fFewKfSVDzwF6KEH0b9HVrC
H9PJZaCoyUna920SH3QgcvM1chN7Ee0L/7Ci/UEOI/xjYLaiArGv/MySJM8Q9URv
v/0bB4YRffkNo0iJ9wJReAgd9RlBqNagBecTgu2TjBFGmpC3cq12EUwXwxShYRpX
2PypOfq31WqywK7eYVUEecDBNp5lrPP1xrfrlenwI+OZp9ac+XypSwi+pYyzYPLd
cVnw4nLwuf1vw1UmZNLJvkIQ4XLmccQ/9XkqF4bE+QTtosTmwK+dr3EHEZ7uY9fc
w4Rwlp75DW50nSCmJbANQpiaE9m5clH8TsTuP3pGX98g46/Z+GwUjUf/iRszhXW4
qzCfUPuN2O0dT8Grs9sT/vG5RAlyvlibyS9t/PQPf+1oxk1FzgOcU3aXfGfHr1PD
7uyC69HiMBEkU6YTGQWaAfeLzAei3XtjC+iEVQFczH9tlt9QF75cWWwA7HBQIRXO
bU4U8z7F+KWpB5lezox5qoRF3faRQyvXFEjaUYiPfpyiBDv1Ul4KEy9GNLxR3dmo
L9rwjbs+6NUuTkOCGVgDleWknNTKXBatKvVSO0zGoxwCIUisFu/gPY/cLGvjHv9N
jiDagHxX4mgnrewF4hHeyLorR6cSx1dlFkr/Zauu1A3Y/2I5j+BPmHZrIMhpd0Lc
CHD9CIn3IY1NnLpXd0smqbW0a1Hs+Oc2eKBl9cqX26WgyBuExOsmL+/R1v3zz/Wo
7JYEXgCmIUkgBN+ebJLR052EM25Hj/I0S8WuYnfDBf2d7KM2atRwarHWz016XL0t
5JwdwkQaMMLEuyGLT96MVii/WlHpma4Fz5BqGj8HmAbsAckBPGbMb6SjATEZZD+a
fKLWFGsSqqwf2M2+lh+JS3UYbYyzZApo7Bk8SFtgWO+ya7JZKYovkhYafERaeSNm
onfYYEwyGeUS9oEhCDSP5FG5srGqZCdteMIPRPiXBPzrsU77qQ+706R5LDVQxYjb
XCnMX6QT8SbT53axte6xvV6rF1fPcLq/UJ7ARfTinFVrFDHcyXrZFKhXfPec8fDS
CGwnEUJ/OpjIcuJezNkXGyAy5EqzHl3mx9t3NHFuDeu0Fd3lOhBlBV9qNvOr7N1j
7elL/utqnJuI9iHM8sp5+/zJd428+lo9P9/ea39AUsknAwvej8y6Sy5hcKSFJY4U
r7lV2xrjvCva0b5i/OhXOtR1nfnpSkBFbQPa5nU28BQwDUW3/DJ8dyBypeiLjgFe
p6/9GBtxvy7U85WeB8jGFrx/FkWPJRwWCSbQDry7XXGidIq8Itiw3LgTcWP6QTo7
xIwXwD/4KaGd5QKy4s9q1TH7qCiiKPUB0vDBX//p77vx6rizTbl3454YoCFzSNWm
BRJj46FnpGzw8y1Rvs1A7H0rhLnl66506zliPG/RCSFMqbBY7b3HjpkFcVMrxhgg
lpH4A8xEGvlssI6wYrB8DZQKQ0vMLrf/XIk78XJRlNuPnV9WqeoExCHVpqarnZ6b
DaSWjVEQwa4PVOSK7f81T7/VASVkbrLN95siaTQcf3I31ugmeD41f9cMwjGLMuhE
hNHgGHMUMHSPTv2M1t3G9Vds5RfaWOVXEfaS0hmT9d+8RySjaQwXbdX9013jodAb
9crtFZQZlLhe1+V50hkVCVaD5wNIHCSWn9+DlNw1S4XyuP0haqhHApiNA+fGZH/6
Gn49531WKMpsC3dByKWot59JnuxX0X14tptg2okSXTJy1xyvYEqyIUvyxg7sENgI
ge5PMoLlsb/ksn+KKOyr5V3UotPaV3T8ZhW1YAp5/pPBazyiUBlc3wt9erjKAJA6
2EQ31MfJkxE4CN3A+4JPGmwMZbfhmfQsI1DTYnlQJfv54Eh6etSijuWcb8Q9lG7W
GGj0YQkuImLafcjBT8gFsrRI9rYdQ2r1j4KRbkyAkEP70/WE2zH3NsaZguN29ppZ
UlTsjYH+7B4Ro7Rrwr/id8BtTZM1+fZtNJ0Z5c2xfWI7IFsnA9LpVl3j622IhJdQ
T8/BmjSJf09yCGeFRV4xcwMZareGw5DNjqbJmC5SXP+8iWtIsyCKCfc3Az6y4Kit
1j2Of8VTbj5CVXFWgPGIkbZY+MjIIy4YjCRD9e7fw2Q2Xj/AYc4GvpA6frSaDjyG
2aVHTFtm+bScdV8kDsFjdVm1w2OtrGczhfelYlkPpnrnxakFlO6MeEN4liM5X9bF
t1XkBRMtARjQO7d2R2bLTMI2xZZALa24oShG3sN5qOZAdMCw6eB9mnCu7oMP69UG
zoCecxNwwNMfkP+Hi8m6YRVSlTIdrIV36JU17yteR9DN6lsTg6liZfw16AWztIpV
/M55BBcTxJTQt57fuhnkZi/8LsorqiYF5O8rF4gGCFwJ3V1BlEX3ORA8UOH0QYTs
rLz6b+lXfUa8IjD5dNHITCIlFQ6ZuEkipsuxU3LoWSq/BL8vlI7UP4x5FBwbk5zF
lCS9oPMynHzGpfdzu5x9uhZFepQlUF08AWYJPGhih5TtTa6BF9oDAZ8hPI0zwJzf
9d50RJqlVPMFSDDqMmFdC7EdYccj7MuxbSgaBybuRCUQhIGmZ4YeURAhyWAKlwXQ
+uk0OkVXlYddmeUJh4sOe8ik1DBtvnxAOGlRB8m/Ocm1ZZDi9jXOk0DYIijEXbKN
EATehWD145PYQXYuBbz14EvBrcA3/z249w5lc++v6yWxlhtWOBi+E2Q1YsMvyWre
kIX4yjm5vsjlhePDnXXvQd8TK1khWfmfh7X3YxXSHS7Kf0WGGfakdoFBp30Q01M7
tKYdhN5xJo+hUDjRsz1irWXlEEen56MQpvMMpuo5vbtqirDPGt325XVvIdGsUbeF
iC33srzXL5xN4yBdm2FeqKC6KmZRsc+OTJ/3yt6MvbMEWs8WvT0qH2kpPFZ7IiWa
uOjVYpvgeAutPMY/tavMbQLlPWnZV9sX/vaKKrmJa+N4Oo803P/gBWJJ/W28RVKg
thXoE7x21oWG/sWBOz4fv7q00YtpFBQfvDzXWyF/ZE328bjJJgX+KHS5DrFN94ck
h9ONdshSzKao4ugMGrC0JV+A3y4PNcN76GfX1eJYifT6kAmMPhwMVcSAMRV7A2vT
ZlDlvMfGIfM7403TndoLY+dq4iHyJeatyTcJbjFGUSeUmposNzp1YKVbmRvX4HI4
5ik6gXL9kZP0OpVQEdc4YaKbU3i2ho+zInA7vlZXbiw4obOQcPwrP+TA5YeYpqNs
B/Uki5fbRCbg6wu3GqcLAyqcUTij8SZ/yZ5eNbATpjajAXfoj/YDrG3D0uY6tpE+
WH7Wl9TelROOCF7Vg05hmaslRjExYNiBx4bvQBBY5T7+ih6P2H+5uUM+0NbCN5Gr
DE3Lz4/+G/eQEo3qWW6hqZ9g2QSr0F6ohf3eBJuX3jK/N2DbV2CCmCNRpaKQ8rq9
5ZcL7VcqNs1zGzKKXIT9ooIbpzTMyVxWivoINoWWicPNxf4qNnYzXfKAuDnZYpoq
aWDfVHDFGl6FdMgGctYl3wKJk8ozTlvkTvR5U5JkF2RawDc/VURz5qmmHC4BXTHZ
U3+wonPzOXlZ3p2jNv5MPdrWYJ6083SedI7QYQEMKGfnAw047H+Ypee7aEz6GG5v
uaXS0eEIdYRIYyVq4GV4CQDuIcE/mgvqPmDdB52kdUBUI6x12vOhu/sR8Tcr9sU6
l/aNEOkSKNvAtqiVNDdTjItNg0i59v8jBXytHuuN00eUZ249JeOFH8XGnBMw9RJj
Sm261J7VflKL5DDINivdcZQ7sGnd0bSG+Lcd/nezWrBMp08PTpxTdtmMupWSrA69
29tkgimjhGERdngDbxeFaxY5GHqk4WhZs3PfoKRSHB4+fK+XRGJmr+UKSW+ephmV
1Kh4ya4BFCGhHdA+D/M1+7bIt/E/JZLgVEdNRDCBpfJg1D7XmI9cxraRfnAJCUkx
EcdSXbXDmDuVoijC79AnRk33Phx77ptIig8jkzLtfnb0Bjg1gz1p7Z5g+Ttr1QV1
HtkXNlQzNLHLZqyma9h0/AEqnsYygF5b+QEMuaFUTRFfV8/FWsgRHH/OwA++cCzB
VwLR4oVm3GV2F5YXCDvdYhwcn+n/rLKLSJgoowYGHIBxuy4bKZ3ditt7rIG+J3CX
kDIpTplVlzdxbASkwUZZIJY+t8PpT0RV8Fb3cNvDkOht0LJYBz0TM29PSifkC4XF
9oB5ZdcBgf10gYTKWNrI4YUKy2Y3hXlY1ifZPViGHt0IcL9QDVkxaUejVbOLes+P
Flmhn6KVUaOvTuiBleuMX03V7NXXOKU+fWrJF+YbyshtGBV+cPcxpW93WjAMCJGr
Vdol13fK1GMogInftTjJc2dYlwCZ6sYM/VSMJswlXZllSDaSCSJliOht9hosHr0V
q6h2GpTKQEpxGy2GbiZ+Hd/k1sXEYpVJovCJId/fgNRZOuxfkm4xQ3SLprwycL0G
sJoDq/wGiFMCHBGSVl1BemZN4aE4eLn9QwOA0T1d37geBQDW1CkF2m53XC1KHQj0
uH9BlsR+FqIIfuWj9lWWyrTGjGvSOONK/damY8mACD59W8gnZ7wIF4eVthh4sn1/
rs030JIP/h7d3isyKNZsDrpFSyoEyHKhDB3kHKui3Wy1M+xOTWMj3JFIcZRl+0aM
0AOoQvBwrRxf522H9BfxFKF5nC/qMJSOOkxjwjn1HdvCcI0GTpyYsCauGHa/rqo0
AnOsFjG15z6UBVNNZ+VO2jqjipFJKFRW+vTJTPOELKEURa1LCxEASLf50TMUYsKG
WzzLmeRKzPiVbCBc3sAlIIVc4XYQlVMp1EuVd46txbeaJQLWdR53wOqd6+gWYmO/
4dyQBZJcgsjGK8uTUoVyx/N4IOS282VeB39o98P/e98rBf0vZQ7vRo1Y7N4uv45l
jx8ca69MfX/FtFQZE87BFH18wmB0DqxKpOe5M+qvLms+ZigU0S6hnh+jNsLcErwS
YbgWnL7WASCy3JiQ3NGJ1G5/SLbNbFQ1wdJwv+qxdUT45pfesvS22gf7x7RjhDbU
whtaHNjbrNuwKvfMzRHSiVDgLGgz7V2LJifo6fK3eJfevbWjrg2FbN43YkXZ2/Oh
o+Cxbx1CBoqqHJfQ8pq/SVCn10e35flsZJ1zpODzhaMq8UziXmWfUxYPgmeexm58
uBz3VaM9WBYfZJFUVNDI0PZrEt/5v9DVQqszrpFE9O2Payz7GV0U4aHzEKrFBWg0
BTTf1aYdApLd8PqcBD5ifybv2zP9UwqlSbVVn8ZERa4ppjZ+r5QBOBBC9BAaYvdH
Hqee4mfBVZ61QmcHyJ7c1ZxX8i7V1QPTV7jSs122Ex8RsXEyidm0PDsqLUUHeZSF
hYH2J07C9AvsxZFWm5D/smUaNsn0ZwtdwOhS2YGUVuRzGdg3LIXi9WPriz+gb58J
rwqnzKuXtu9XF+2KzE3FssuxCZhhBKjfsGZmnHLJI3sVFaO3EF3OFy34/Mbd7GWg
n0nQ0RtnK8vkvt27iF4XQcqr48WQnobRsYPRhuY8qE8r3O091K7166oEx6oalfjC
3BV9xlD6WxCCFS1bD6nx+ftd/KY80MKBMuW/QwDr/n+9iL+zRcFu5Ovg+2IOT6FT
jg/crhCf27HEpXR0Qv0LoerYShfQuykQqEWdJimQXA2YuLYGFUoqWjPewAkUCDor
PPZtLVt+MDfbkj02/uPPi8rebSmZ51aMj2fAhB6cYPnabT2K/522Y1Jn4yezIYTe
RdmruGlOXgCGH+xMje5mQJEIrTbDhIxmys2VNEoZkL39iJBrQKDKaRqA8AEVgOBL
LUF3zb7VHsKlsTnhgCLUeC6HUz9RZdiITEgAYKWxvvJy0ggryIML6nKCZWSq+nyO
iwXd8bDhaWaVWI0bVjK/fVxzKKw3kehACyt/Ncx7Vv5kwGtEZx/tFFlej8W5QvOg
gQrwcsEdSUol7cBMk7zFnuGOKmLeZPeNFfgHWI9LQc+DD5SsjEHQitVIVJKmhTH3
cAkjPwykRJjeX6wClQlSM+WYWgVDdO1cgt5IkwJpfHcEKrdUmX2H8w4r7aNYLLxh
6IHjpuSAXn81XU7sDuZObBp50Lt1FLKCnqa9nGNXi5Dbs2EQ2Y9dp/dsBpVmfo6c
Fjs9+Xcu9OBYcT3ZTcAbfjkjebrtAvERyMMFxmjUmkX+DksM5408fvkNH1q0TyaL
I9NGeLoufXcc06R/wTiMYhnUNMYl+7xtiYmCgiOtljZmlnmxPTVcQ82Tt2ulcspq
eU1B1zDSti/Gav5/SZgnxaeKLXDkX4JFOhBUzqbgyAgM2U7R/QCknbjojLzju53m
BTtGivBTd5XuhYMQjodm3EnmseU6ltQ1AuEaJ6w1Cy7vjI9xPhGzM0k8k4HpbtvY
DsVYeeA0PyP2GWb/8nHGKmBmnoKoAgF2/QciTBq1tNIspMoAFWWeVRdbjBh8YzJ9
RpoucaHnbtcsKXy43eBnh5WHMQwzFiQU+AHh6rd52uInwR/q5aDhff/Tz+buRtyM
v8zFMEhAM1o9z/2sgrXfe/qdwQxyuYxoLYC5DQA2yOJcnw/fGKC/n3nWsDbT2DDh
6IesGfGoLZpkC6F/Gxwk27O1Jz0E8o06EqEexdeYNb1Yj/1pE7DMEpzo/eF8hX2L
l6dU990oaCsYZB10i4GEdvKM74BGz5gjbDLQ3yWetyCS126xypLNBJ7usk/nRm1R
Eh5ytQwvsJJJKCA/ktfOTZiI5KFZyApFojf+/F7Gbh95Y3hlR83qd5GkUgh0wVbY
eQ43wIRifMn83CnUcSrk6SZjrzVlY8nH/CCmBp9PCWcbym4UGybWa0/A42bwWvUo
JMPBN+walr1w+8z8shSJAcuxs8oQt12zoz4BjHh0uAHhjKMCEBXhjEVm4i4nlPKz
X/fdFYrcoL05mFzYvV7l/18IgOylo9K8yZiNlbkYnJUcfEIuxhRQNsPZnOo65lGV
GoA5hUmlOCAx80b3h7zfMqLJpt53lQt90aF7OL0UnpJhFqBvd1IGhOEC+ha2cWyf
T7R7hN0bbD+uXmemjzWUX26fA+QtwhOVmSTBEviESt+rJ70w9KTtuTSEocpC0u/r
hnUCvVWkFft0MOe7WhJlK5keckiNk7xiEzjN1eGNmpqkoc92QI/W5WSETBo1lUqX
L5XJuCPn37+IOjLcSl2uNsniyAYTkIG+VMcaKTVaAtrtgogFdCQm6P0azMiFV+8q
441vHAZooltbBsQw5Ks8Ut75s4qpu11cK/vF5AtUyBYV8q5FCYvtbscugYM8yQaM
GyLxPF0jv26bi9qa30P36qHe8eMv5k0nX8lOdYZHj4RLIGwhlwYbOt1t0mHOBEPq
5xmeij94B/ANcNTpSpnVyhlZQPV2ANY0INkyNBF60sQ/cUztO8ByF7xcYqvqQJYf
Gj0EG1KC8gOKkcldtyqUEwSSZHBsMWeuFWVXRCl5jBimUB2RRLsrq23D80EiPqok
x8WrkzdoYV9O2CuD/HiFVWGzfh3FD6zMpQ0YyesyLEEpSMxFuUvh60U4vY1ClurE
hZSGuNPtkMe5AE3dNY8F5e8ZiOm8XjL3PgY4NMxfQ6k2DjCmmORnQAVx7N/UQBlQ
YaaUhVouFpGm4WuP3gLXywQPJQa7eBMuly4L0h3VPZDZ32aOjq4X2reBQ08Ax94x
xouiWvoEwgDNjO6gwPBrHKyIw0fSSYfqjkd2ixtBKIcyzoQTlvzEDizzrykRERa4
/SaFNx9oJ5ViMUWl4nrVVd6M8OF6y41xZDRz0PJvhCggBRnDNueHF5XvAjo11wwD
rKDlgD9q3J3kHtGmE1nxLo841d/N6dYVvCYkjUXZKPWgi/+ZfzgaiUGjZWfDD20V
TKK5hQXKI8XFdHHy1PLYAoKUQfeNkN5xGLl7iaoTCm9GutQziSH3tDzLc7FX458O
m/fdwEeoa2AnbGfrLXn3KccYrUkZ+isUWhZK1B5eUjmZ+sHmAwnUgQ3N7B3Gjgyx
2DM8+AnafqtndK21ty1yh+RJIyuItm5JG5i+3AtvSOgpc5hKTUbL7vwqJztHS7u0
XgbvaiJHjIVorkm7RvZrKP9AdaS8FC+zjGlwMGqWM1zJutFEkbvq+H7gjHHQyp/u
KZ6ou5icUABkj6b3Kf+IZ6M7dTA5xNoe0y+1O+dL4PAeFHVTNTx/UEHl/g/0rSGI
ItUdkTA4uhXCnUyTboBl+TLIecu432zOApW68q3tH4bB1bGDsXf73UDg0wxtD8e/
m34pFvgt724Cs5PRsS0lEmuovWV4iQfPDBfdq4wb2gGYTgYhD8jbNTOUScc9AQ0u
ZD2Tx4Z8iRWMhejOVYBNxh7mDAbgiJsUYtORIVLQ3kKNCRvin316eCtQRVFhCzqP
bmmygcNAhftOqmND/8poT+LhRAyuDciZWykYPjL0/DZHZI735tJvQ6JdhoKZdtQs
s/hX73JDvgVs3TfcG6L2zvOqz2F2AR/7HdpEMC1fdMRYCsYkdad9XY6+ID3fOmJG
aBHgtd+YMBa+AdDhKvI22qZxZu2uBdUUZFW6eu9+FukBMFc0W2KxpqobgIY9O5EG
LQwkzyDshPK2jQjgwDDvZHbPrO/hS2LmV7tAaWbAxc9itIc07Y54BXnss18/RHee
431KA3aHw2+Q27fM0SMHPuWFuhLa52wUTKDocZjJxpVb4z2NrUMZqj3hU7V5wQft
dbKU2W0WuRQ7snJqCk6OI4MnBFEyiBCJb0WarZ8DGnskYwVmstqOYElzMYM78nIQ
lKfZgojUqsFNotkgd9uhmJ1J6B6mozY6prOVpBdsOq8pD3tuekjaWZt4IoM3bkBS
d5I+LUGoMMxqjnezWL5UWT8nez9AwTgz+rK9uAp4+ej5qSizfbJAjGUV5cdZHz9a
A6qAlYN2BumsrwP9aKreZ17kdZVhd9bT0AUQy3e1zKZJbNrtNRhulGeWYWCpjgHG
YnA3i2QzW7K5M2s2cc+lo/4sQQyrXPgeh+3vHVylG+xcMUiGPKHi/N36SCjOl7fW
nVBt05wup8470QfatV8rC32b3PsFmlyxZkSrT6XRmhyBW8pCokUlZtMCEIIFbvp+
mXhWJFAnHPqpCpOQCjSP0O60Hy3Qgf6T92ChNTjLtQ9RJwo203w/LwWh70iZyZVA
Qvd+tgpcU6pT6MPa1mfYI5d3rMx/gpWZvMclewt5GAnK6Ua2RwADr4vbjA2W7XOQ
d4SVLZdQO+g7fvYb+DAPKJBKxOyDBi4UxXL1pu9kkHgE1S9jSmMNQj4GFERt0sNA
/Pm/6DOvTsAnTFpN/0xjJXHggUn5J7+y9j0wHDS7qXKEwRAI9ly9TVV6Pss4/D5F
2lPc30ueBEX7z9aNagVCtCYLds+AhBqNJNU69CLC1dH6knvEFtqwGC8EaEDmtHSv
MrTsA2Vb4owMlW8GKteduXl8lQ7p5dTdF5FFAVibk7iOobqn/x65PWYc/ThwyBJz
coeiLdml1dM1O8VWVJJHDFl7sWGKpRQjlQ48vdYWG2ZUvVY868jgPd94A7fkE3A4
RW8sjHyAI7nHhixdbzl5kOi2ER6IslGWA5KzjCamjgwD+3Y8piUT8QB3eh01cYE5
+v1/YpwvLPy6GJSiX3wlMRGvnawr05OmhayBzkvhq/1eyRXKEiDBSLhbkaWxxMe5
X5KoblpsFOFKL/28hc+w4PZYXuofUIM/O12Ln0E+vBinczT7av5XCuZyl+XHGjyP
I/dts/k3MCsHSzY4v6Ky4tPYAs6wSYAT7y6sDLd04roP7V0W5/zYvsx5vwKDItnI
KkXoOjb7j4gzxLPpkjL/MmFcyXFlEeNSvdz698MxPhzV8q5dRPv7HpHNj4EHx81T
ZMk/8/tLwGPjMyyngZI6bXXYIITdVl/FqYyMfFNNM9PhDQcq1nt5zgrKhsq/kQ0w
5eeMuj1i+Gb606YvaH1tTy2X+vhaqlC9qNVWJNujkdaj+13F8HQpEfmpkNs+qYCi
dVnwxQetOFF5yjZ2jyuSG4paNB1sPgsrX4TR86ljtVLsCidcNdCaB4MRpQtp1nA1
utls3TafkomszNWAhQoua9I0K4SRz+TqH9rSVsaxCn8nAki7EyhEoui7hGnY6U2p
z0u7fD9jbERCvm5m0lhGyaQRbPvPlVGeRclYNkt8Bby9NQ5h5jjNekCts0ZMccx4
o0BQ7zxthgEZf1Hqeu6ofDf73YYzR8D52X4NXM9SGagQJ0I1Q/0CVniaqweSut1q
hGTiCte5UsdHyjfHUFDPH455KzPcz8EhYISiaHHWqeP70JYXmf2+3RZsRqsgxkAx
sMb9EzkZ4G6ZfZZpycdMvzzxeDV7x8ZdAfCadiarfY8XqbSDq1h78aKx7Bh4KnlS
F0HkFjlw0VnIJV46CwN+tpbdxd8E+Tc0AwsfS4dyJD19Sul2nAJOxkvJeJ4muF8r
QFxKJlUgNVU7pcSHbsWl96M1u8UZK9rsQk3iCn0YKtqFAXj9sp/I/iLzhyS6mB5z
Pr4WWWawo6Iu7iTXPZQpraXbthlOSLo8Vgl4Bl6jUWH0h9i4IiOx3gpRgHzSgk6m
ADMuJBZB/1MNSLo/IjK7HMj+srXcC0Z4K1DTwRetJjnGmGGyb5HbqxrU9JKRKkCe
BSkdHN/q1utyQNg20Ua0JmA9+/y1j1k7eP4547aR6fwiYc8nxfLUwy8KnKiVgJlh
lsqAsuNoJEiZRxJ+Z1qkExj52ak+2ixp/hzfX1UKweEOW9QB+GmCzvFjsFw4AySl
fCZM8af04SQgLvt95TMuNd81Pf589Bo65Eql3tJ8VmzTwjJb9pWduUz0k9TgVHws
a6p+FWSwK5VxPVX7BYG5U+aL0PLi2O5NBPKvegdKpp/ZMOnyMRtcbQ9zuZlJXDio
CLIQmfg5K1mFzv0HiR9nJ14qgqFz00n+OwzeXEpU7u0DOk+5MyDrkND8bUSMt2Hy
FUIKUZlnzsqJK2h9LbktkZPcfrALHzWrFEZE6ywF4809vNpTijR9ePIQ/aik0rTD
Ddd8w5k/v55E7K69aOU5ug3WpzOC8YZaS78MgW5gVPtF3TyRlnNwxd/Wf4ens8nY
AX3cQ2dUmU3pWglBIUSXIksu2vBHBYhQ4pyxQWmyWx3UW5qpnN13NmM+yjEJDaKv
qFhxiYIe4Xh9CRZvNR8qa6tRGwusG+eZWjspUl0K72frjebTdbg+v8jNNDh1wT18
68zi82Fkbf4Cvnh52+F0FX/R23jATb6fp29HV5EPsIxStQSO5Xm7wFYJvudKE6Re
BdMz5jkN+RFVLpw5LYkjwfwvmRlvCm59jq3CTf16pSj7StigTeYGcB611npb0BVa
9ovLtIgDhHV6kfiuJK/P6Og9hdpMy6njIhzk+vX3R/JkjVGRtRmi55JujqpMnWGn
rrtW77/vA+cz3kcxFsPKuqTEI4fYQItP0coVQuPiWeoI/gga6mLV+UGhVzgIEn6M
Bzjrw8Rppdbq7dnBMLPjRwV6mP4xpsXdtApeGT85149MHhye4jitCCjd8Kzst50K
JqJDapbUPLq/9kY8ye74IhT2Zb/zgBw1fT7jNLcXdtc6iB4TGIM/meavi11dN7rt
kCyF1S452oG4SsBkMMPzxPES42+EwyB+cremwUUSDA1Vb5zQVpi3/qpblyahyr+z
cKmrLB4HrZUUzqBl0J7uD17XQBBnhfzmAVZLcSeEUe3qBum1XNCwD51nK4Cxt3YA
1w5lcCwHWf0KpTusNqqcM88OQkodbeVpM8RrMQpvRaWetDr33sFU/EfwYBzllARj
UnDD5scbKyR2IBdy337kUytcIMk225mtaSjzb5yNtt5tZhQ3aZ9XnXgKfnNCO1vi
cnnEv28o2AqKTzjNDZIx2TytYodvBWyO8pHlbTRE+yg8Nxuw2YkKxLgAkScwOv5X
PhcKTXSLABjNbyLAqezW6otl2zaNCM1gLHlG5h4fO61QjkycZR9zhdgXn+t4vWpB
1eU/tJt47BK23/vR8z+wBz+pYNJr8TFrIsMCKjse3f1Yuv248YwKPXDzx5pXNNro
17QG8/pIgc9gszsnPizAYxI9jVzKX/Jt7pidbZnUgr5LBS49i8AMJehn7kG+RZog
CNRI7ye8CnSEF9Km81zRpLKoIFeZWdZaAvxgd214jaMYAjT1VyIKoEWmyeG9dliZ
Xpd6p7Xo4OFP/OGMPirN8LMkK0RJuq9bfFPfkMLNFRQqZNFUlnDqYBbiPJfj/TTT
bc1Xje+Jf3eeuB5eEkBMC/yLfW2C55nU1RzXB3A93jz2oM3mr9bCTA473hKjcmiW
2yq6lu1lsWkP7Sk2Wzk6mI55LqS3Gcqwiiy95FtdTOfbr9kXZH/KhzFh5R0hPFws
I9RdUOB67Uelx5fVOf8TInW3IkIQpxE6LaJUel80+PsOa6bh0PzPu83gx8DWAcnu
ERuWAky4vPDzGQvRS4t16IDIHYQmKpo2ZZ0tBRdPEuUXmvLiukwVadKVh+nE5Ivy
6xOLlnBZWU3EhHCj2v2d8EzUMDjDiXDqHu6obFhu+nGhjXDwegp6Pc5Y1Y73UJ08
FzToUvP2PJ9c59HLuvLhCr9P7jDrq8vl2Hipb4H94HJgX7k4HMuslgghtXrmH7BR
dk4AiC6iLJnLy0YFJVUqiLQokHS5roGgok3ulNwEivZnJ0hcCt9HSRQ9FaEvHEKz
5GMqip3wml1qp0ydmZDHH7vtfLIeR6A7/FgezLu3zRVkvmLAf7+5p+S30bT3fxrA
QjUP/YQmQFZh5hJKdXOYOvgkJQky2AYd3J8rqJMQhSleyZaC69cccXr+XFP79URF
tf2RREzwKJ477DDVCx9rTiJ8oXYbBgAs4xZaAN5wc0S+Dxy5Y6VJc257fLJpxasi
lFsdfsDQQ4uJTpLiaPhe1XPxG55N9/HOb9reXF3b7m+sAQGHIGBOEB5A/xMLjhV1
oSxdLBxXGA9Jdd6VKefm+/6CnWk1rTop4KNwhrWwv5V35OzZky0/boMbbj/tSuOp
zQuWoRVe9hWaDaR/aeUGngzV2O5GLPNS7PFsM5a86j3ClAUtfjCGiaxVLbupg67X
xi25dKtxYzWr2L9NZBqrPUEwLp/LPqJwHqeEH2s+xefUVptSpf/Rb6EvpG+DHO5j
D2UPQwRiQJXy3WW3shrFzi0Lzql7r1sguYEgzyUGps3tPu4kB9OqbCotOxlQoI+E
INDHu67URUAAE4LI0o8TMnCdNgvFBeztusUCrRbJm2tF7p7xAK6WyeDGgs8sqhJe
UfJRsmlqI1q8LaeQCS/8CTLNQ7HiHDC+uhAhaevYa5Gu90s8gCjx3tz0VNfVo0ah
1gM5r8MQr2On1lH4lFwq5YHfayK/uNEZjuLCUHaA4GJJvflQECgXejQVOlumzZiy
PWZgQN4JNuuuGBdptiXxzGgfP2YzgFP6AxxfzU8UZjtzWLP/Xf+vFLPPTBQ42790
BlY9TtEJleYsNBJ3qRU2lt20EHiS4S/upG2fuUogQLsqUuy/nBMY8kv+HHeOzaA3
oH+msKqvuQL+dqlyCyrXYN7Z++8Pqnv8FdnvfuVTxM1XsMbLlPf48I5Ak7ncLobX
s6ccnEwAxOpg5NVkKq7f6UOOsVGnP5OKuYeFUpEigA/PkSpq95r2zmhXWeIadfUP
8AH0hznUlbnxyt4Rc5AjfkhSKKmNHM0ozjqEu+jKR5Srb0eCSatnbIkNH6RDsTnE
UMGBcWK0AOJo6AieEGs4sBB45yE92ZzoJtaWUtXTZkJm93t9RJnHY3dR8qRhda+d
tfL6c7JUkWrTU6XcBzHGn+CrApMWG2uxZceZMjjoEu2HuN23VZsKSMg5C1gEtyHW
EF2WOH3CGPqNKTv+UXQEo5NfvPveQ8R6Tk1cYpyW2yev9aqB2H8qy7sN08w7PpUy
/2EqHn0rE/OxFG/xdsa5hTA7l6izWzTFRtc4aUynByB1JwVmnYWdUqvNXKdbOjCd
RPiDmhzAat9cZKK2wWSj60g728zQQC6yvRSZ7lxPGykYvve9k0nuqbZ7nIkGdOGF
HH0l4sM0sEM5Hu93Hp1kzbhsJEo82H+Y94hyWDFlb6Fjb7yiR5O6mrU4GSINYD3c
w2DGGEvTEjaC710j0AHTTas1yaJ7gf1P9RV0dg3TK51bi0hQHhbYSesA8GnmaNIC
kzNBddrhBQA6rYSsTj10DE6HjKGwH4q7ZXajG+UQ+Ed4N1i/lPhibW0eMKzBq2X7
NRWna8iO+57FzG160baxmDdjRyQu4b9QSdlIhqXI2GA3ylzWpzMkbRTHRKfo9jRF
LwxPPM7YkBQvUzldu0kl3olSeFVBFg5ESle3Styk6exolmfBoEWch71hIS9hNnwh
N2MM/tK4uAwv9gyfYXnF6Qs4+4ZtPTYx1Es5zdRa6BR+HEnrlLGNR2EX+dAPgZAW
l3cchx8puxX0NDiE9e5kKVgpFktyq1VVRF+p0NGh4MIxyFgJMw5HjFrMB0tuL7Ui
ZxTJcWnY5oM6xmMjN4PhD78AKfd/b+edynBPIpZdhz2Z+p5omuji8/ssiPXtGVMI
sLIROpSj0sNRR7GYQXt6NwZwtqTDqV+O4bCfHZAZcpvJabCZu/V0lr8+kCLI68WC
RR8EyghigG0LHbeT+V2GFnqg2+lur2GvnRl/7Y47qGVLST/kIGLRNWqL/l+7HqOL
uLWTrb6QGovZH3GL6wfXiajOwLDxSUdNpibDVJW0kgj3pt9Ywj9T4eyNpi1LSwAP
FJeu6P43RNv/T1nlvI2xK7vXJbkHkVNbsbnoGCNRM9Rz42DJKFlsnSpVjEW00dHO
KOna5/6ICMyMXAz7V6IBcBTlWGo15FlO6H8qYZhY5K5LKc0iY0A8gIFx4GBvmk4k
Q6p/dpxmjiB6DLWBQOnNjUMd/eiim73G6Mwxtkukm3e4YDr5r3BL4IKofO7/Yhi8
cIgE5p48p+D21JQIQ4LhFbEn+HEYZUH7L6I3fq9MCBVuYntQHw3dzfBQSYo/Bqf8
CvSY7AWIEa8jMrBbXBh+mkCxCAQGQbwaNJOFr0yRVDXfFqLiptd9z0eTgbuZpaZP
F9IreXGPZkVN5Eso4qrYUIlKx8RgaHquqH0FDkWw53v+PSNN96v7PuHI7f7qkvAd
TBfwxaMjTcSVITRL7nUorfeq+xofiGInTu/8FORsxJPmPMpbX6DEUv7/gpxw4HXm
HPzwipvLdowbpEQHbevAvzOJwfHbiKno8FjCLXBqfRYxb92TMh3iKsYFuqYUc4RC
B9LULyPf9/X6SVpg3ezsMMNbCqxSLGwahzwJD61ur1GMzD0iKfY3WX8eGenoTLP0
SWnb5OmxNpgv+xLIHdaKhRI43sh1S7x+F7H7MdBbOsDcesTiw15vDVetsjJrsdO/
LBQEbhHJd632YDroAPgWxn67L3RWse9+xeOWg1XBPFFaMuKq6s2Z/KcaSh5JJEGW
i/l/BJD8YCuNDpdU6HCDDGtfuu6/BbZXU2wVdaurHe+laijWmD22KToipCeDDtGB
Z24nbRJHE0vAjPE2WSNDwiRhcLGSAg0m2oLhHSN8hU+0KMu11KA/B09BASpxrm8q
iQARRPUU12XSxnH4i4+DOXvZ87i6t5UCy9Ox1Qp8W3zmFo4LRHUG14qEMw2HResc
L2KJtiC8E62PfcmaXbLZuc8A6o6rid/mgQRQ6UbJ+K7w3HFvn76KdRc25qeF4fSt
yokslouXq5+HimI9MwPrnF6PZwzN2v7szrRjPNnUwGA=
--pragma protect end_data_block
--pragma protect digest_block
a4hoMj6tffw2qk+AFt5qVL/nDcE=
--pragma protect end_digest_block
--pragma protect end_protected
