-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
jT3/WA5/Bi0o3CXcSGZZpDZxTpeLGxLPVGIencE1Mjoz7brb1Lvv1/zKrWvwVehW
p3RDPSCcNuMBmo/nx7mhA+4Hnxiy72RlJ6a2S+nbnxfROhGjZVQlU7eupJP7rXlU
VPbR1Qrn5O4NbShXDqDJI8Q2xObzMONx8UfrqjDp5lw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 2848)

`protect DATA_BLOCK
6EgMFVsGhIcxsz4QTWTJfUFiiMUNMmTienM2YpvwQmK9fLZWks1jOpTDii6ohibp
3Z+LEkmWepwrbrbM7rxBl0EWIk09AVQFeytt8hVuFjoEEG+8grlgPQ8eXJ1oI/bx
3pqdbIZdDcp9/otEqVF7x3dAmyiP43+9i3R/3VbVY76S3LrYOaGasHeRB2JffniC
Sl2b9QJRiLiBG5RhM+jd+l7Ho13TgtqOzuiTaCt6J6+0UFWzw6gPB4/SUz3MwgDd
7+/0VHkF0FppZvnnUvY0OppJNngVPPG5rjTakAb8GeneXpExzstgS0Ym7xwLKl77
jB8wSrkpq98smYPcMHpVMWfatM9Uz7bdLIC3ixEiSHuIsAcs//Q/Ui8VQtuz1aoK
WUgpLjjy+K3krL/dXJEmzECjIqvprfKYhJqRTO+CIBV8F/zveZxqIS8dFc270D86
o1vwWn/UGaN9H3EBHX5v7e7RqybyM1zntHV9SW3u1O2QZdLh1tW4lbgEn2ue6EGe
9mKXmRRd1Mpxhgt1UL+gwMcI+WDRQnmvPN/MLxZ5evnigjd+OiuDBu/X/KJyt6y2
mopwa4+mpUotoL1YZerVx1wkJA2ECnuyqEnJXE45CKwe05VJPzUZoxeHzEVJ6EQ9
wJsUlrNne04IxnOWOoYNYRFkeswm6/IJIhXFGurrNVOYjOSmB4Lea7wx4heiMkza
X3+krVS+CGjNXhnyh9GTwm9u563b00VB0fmMMIvrkotNAJrZDA/3gEp4DJR+Z3nu
VRpWMxch4WI/WDPRFUB/88LXV7ZSwzxWfi6+eHmAvFaDy2DJLSFxJIEKZ7erDR8e
S1Os/lyoZo6tVAEcCpj9ZCGeeNhS+VNPclP6oP6Cun+SqNxX/uz4ZplASUc1dXrl
552m48Ddvju8YsvSdrjUPfe7hb1ZSKtjb85oF2iUxKZHDT0+UmkgDiW8VieghoVj
I/btTY2KG9lWrAMJ9oTb411pBMPb9wUZz4f+Es1qXBUAsK+4Bax5ttUfLlrL33Zc
3zlZ1PoliRzdrQd92N3V9MRGzP3XJfrnPoQJ3flrs+qvM6fjIZmUfrp6Jjhe3Dkv
1T5t/M1jrnUOAgHhfVqNHgPnY+PA5srBgPs5wlHE/kWAxNTv+VN+3iBl0qDh0l7k
t5EhSwFBFyk1qdsCBXSpoc1NoPHXnM8qUvYqwGa7OG7nTBedFL67KoStV5BIaxap
4XbSQ5IJ6UelqqegXI3NvOJ/rBaRQ1MabQ9WRuZN5UY+XHLewY17mN+jBTNEQkbf
6oJnjo/TRrqrchZe7xRLdZiv5ZGE/T2xZeddFscquUk4A4zQ4xGmOkaNyYGLv2Kw
aZAZX7dd2rf8651WCww6AEp/hTHPe/OnUnfvicHkp9BpH9sJzCUmZif+qMjXC8Gw
VjVfVdBmhdS+3qse/tlBdxHHrdKL+8ghK48h6hZHKdnoLTDCmAodX9hllS+u4bc3
JNffpSszZvQrpRxTKdFiOdsKW5xyOhFeD/i6ppx4xQDRM/MSub5i5tAwNttaMCWX
qAYdoFjn9tbw9MgmDSqgsRoDZICKwBz08Vg3rHAD4f2oiDlftOOFdBcquPfoothu
b1KoJ7KfYbGrwOxVvXGEgyDkfkIiGbk1Yl6MA9sMhmJxPfKTNF+wTEGvUDEZLyUF
WoehlHn818GkIl78qfsmTKKfkGKvbz85XP8PsBS+LlBnwg0DZ20NzIQCEwvTx5QS
VojA1aRv1xEGHCTxBTgaVwcOcYwY9l6gZKZo8fznYCzN6tp5NrxN33xVgoXk3g+s
bytChyV3+98Tg0H5J6XT9GWw/27L3+w4WVEPsZ203gCujX0qy7SjFspUGtfH76fT
1OvID6aIH8rOlhuiBd1hGXW9xYND3wnGolTQrVfDYBQtyAnW8qDc8WOruLI2joDG
swVGFa1WNgOUuJXi2+9g6nwMiv8iQKHjnwn3HJ4MuNRkfPbPcbMgHWtGlRXLqGqq
psb/8CY3938KVvUpNf35X85oQN90e4bTJ9aOyfHkBjO9AknD0l3PrcAZTTNNHH2B
WJuep6dgKpPPMxb/0MQoEVu/256dUKOfgCbuSmIPLyEq1KZRJ+FdiWnONvAcKg+9
a5nPGufg5wQ/FoQJAuLex3qou0uXE37k0IDH+L2MNu2GUCFnu4ElrVZb1ZCy7xZU
Wkv+dhheymlqAq8IAj9n4gv6VeP0wverr2PtUqua6202PWr5LUv+nxVj3YbD0XZD
pDbG0qQqckBC8sHCZDn9zJVitqo1foW44Yj8MmgOyFfZOmBh2mx/EkCshCf4spvb
OtJSLTODmOOfRK1u29Nm5WfS2U4wy1BOpwUchL7tPAjbBPENk+dqD4y9KKnQbYY9
b/ekfjWWYSG/oZbfg2H8Gcmdxl0YflRcnd+RnYfBPjWRC/lRVUCv6+ZxhxtW52g3
CrlARoanll4Ep8U8YyVTxU/j+L0ggzllvtDSm+P/4ehxjPvr/b3t46wr0G7hpzLn
nqCg2daP4OoPKNZB1SOq31bvVqIne61TB1+dcoGyzRbK11fCABgtsjEgzPdNYAMD
CRPhqv/hLM6g5dImOVEFoyjlG0+SMXF10kXWPdJApLenTmuFLQxc71I8t6sM1lBw
wqo7pP/x1eo1hLDydRXK0WSv/Nw8tyw9vXkwMJxtp4s9uTY7l4q29EfpobrChFoA
xbQiVo8Sp64hLgTsKo5fopF6gfY0rTfiv9P593ErB4j3SX1h2mUtJSV/HSnfvj1P
K8xb0HzaJMAZzlq0GEAoGF6QFrSbUkhW1n2fMmMefz9VuDU6KJyMaUN9O4cfFAGj
7rEymlqa82GKQn8G4cNRkvlJmv1df8SJnVhh0F/bSBn8na7mZ90vklxZAT4Co6Pq
L7MgeQUIPSxhaOBxkWqluptgNTgiXa2uhYFJWlfpji7RqBIuQkiaYi6LP0mtmAOT
/40vAD62EiCC9qGiwtKq2fTInurAnS7bBe2fVscuD7hxFfmhmqyw0HLpGx1H3LpZ
+0GllY3n1HIkvjhO/Q0JB1Pim0AJFpNyYz77VnuyjsiO9r60ZzhYOzyezVcBFAtA
0jc6UJkjKDzXYvamOWiIxj10UD7as0M1ZbKIbve3CqLUw+N6Lp0/7ZRIfd1pGf5g
TbzezZz+Br9x807R2TOqwRo+b/x/gQUsXtlVhesucEYmUwD2uqB+3yEq2oqvUCDf
T+gXLa4ylYKdrKdgwI6ZmGHWAkMT9D1Gq7xBYFF31b3DoRST30J+kLwTDq+UMyek
SrY8p5n96tM+00pq+NJ6Coj8hcelMJOLItWtffqcs6a4ODOMoK1hxzQ/4zL0oZQG
wgV/PCnDjFakXTWmPwflrC+i9otAHQNpD9aKwkzVbhq9OcF8WN2WUkafpvnl291a
s4FfpF8TDxB87EGWXQjPwZNaqUZfkJrL/t7KLxq18Z0xWOwUx3sKWxWJtraQKZla
L+4i/iFu7Yic1Mmwaa8KvwJIYKURiDkbAjB1TajlstTWrAO5pn9o2uSlCWSfpQ1q
T8u1K7TD4ax4Tmq0SXmoa2XOZqkMsYvQmz7vr0hFziYhMMvF9zOFiCA0FFm8Qt67
QAkzbec1wfD5hEU7W0wIAzGTNIhWrW2Xax321UZ1Rz3NrqQVmAD0aVYXr9sF88mr
33KAh5QErH1r2AivZz+9UT1uAq0gBVr6LPfy8ZMKIZr4oxSA45MbfTBt207/GH2r
igyT5o3fK1yFdlSwtijajKyvJz7nRnl1PQVq3xqcGzCL9bB0VlILtDSCl/+2xwwP
Z5cZxQX4GyZRBtPBcXXRLguNJ//4A/97VXDMNUtySR0//3/4FHwHAol9kbpQQ0/U
`protect END_PROTECTED