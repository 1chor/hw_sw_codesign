-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
HvyW4/3t7IIP+jESCvxT77iok07mU+UwuqdZEjiDfm2Xb9IRM9L9iAnmPLaPpGqH
ytdRMfLPS+xKAAXdP+TCnnC8GTbtC6zt7Op4lTr+mS8C4Y7B5ovq03lMMeBUAHTN
6WhxZDD/BdWTmFJnLReTf1RZnGEmuUNkOK0CSxDm2tA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9510)

`protect DATA_BLOCK
sbM1jUCMSsA0971ha3yKerWqGe0a7Z0tegCr4BQKUKlc6Ms5UYW4LN6WqALaQFV5
Ef4RxdUq6ZzwZrpKM6XMzB+cF/y09IGfS85RRJr/nE8ypK7n5cAqoPeDQsUD78Xy
yAnmd83dnCpLHKMyHE79VW2k/Hzp6rfyGTey87pLoVvCt+BEbxDvsCCQHfCBKHJw
UzKIDrMEQALti1LUUVVnvho6paGHBBfOyLJ1dBQGAOydkDfY3fngAtUT0k7aEsJV
qbjH5jMcYAFb6/X2t+oxXERHngVgmW//ObCbp0W9hBGPdsKWPNobIX2VOReOcUTU
YpTSpL1nXxSM37y0vS/hO/fBy1wWV9KwRw/qqtiTCDEyTdr3Iog6WgGGvNdQsaus
vAxCRkx7NFw6csvwlN5P9whKy58J+4HEblwFsr/PWTkd0iytlP756VygVyvbjbyO
tJXz+J56kHmD5X/DeSqfOxKVojQ4syB10LC7MT9AjKYhYEgtvzZR54hVwWuF7KV1
7+OxwFxZBmFk7xcZRVPSuKG4NB7ZCLsU5nyYTIIYZz7pNIsDk6qK6+/x1aux2Ox1
Mmh9cplhS/IIQgQGjTBSjzWIcAfw8odinAZFrLKWZw4mA975Pgm4c04Hq4yjCT7B
OttFpom8FWuIWutrHJKnth5Xa0AN9FNfeG3nP6Gsh8ccvBHwcpSu+SGt3h1vk0H9
7VkaqsOeomDsCalOZLR/TAHO9LF0lm5cAPbN+kZP7RkMWCWn8egOgnWoivD0YLpt
DE1E1lZOJwfvDeE5dJB4JPEDjPZ+baJfE1XgTsd4WVQWACkg1smyEQ2WIFskphrF
xbaw2VqdTD3y5wJHhDukJ2104y9jYCOLtXTBsCgzdMZiy5M459PRdipDmQvN57Cz
BmQy7CXmOgKMoAwe0N3YRNpcCo/zT0sxeb28a4VPgyipH3fUKlgQL22EL3t9Dhsi
jx4J6Qz2rctMD2Hcb6W6d94aEjhY6/a2zmwrtT+Qha2g0U1YB/cXh+DERpk8LDZA
fiTnzHusXXJEqCQcRl8jxDcnVgf5GehYstC9oJG+9X33BXd6ZScMDFwdcBHx7koe
0jRmTWK9d37+XW1O61XHzPAYpNzt90ZskHjXfPluO7QfWCnbHJP25uRJmy8+Ngdk
inw7cOwLJumqecrvR3rNqxiYci7E31IN30cFsdoPrrJQG/tLsdy1uNgzfP6vxCGd
xJ7DdmapFLmdxKPL1ujjV534H1l45v7rg021ufujvMxH5lDOE2hE3IUYXNHjvFxD
oYoL8oyMO1ymJiygBbt5U4kkbtyPgiAFOLJcdkZZu3I25qmqeuCMaAyhJLWLcSwQ
24hUGzAvHZTBAamnKj/Ya9fzEZLq1OE7K2o/ya1ORF5RkblZ4QWqihuSQWrtk6KM
aGyNt2stLtmJ/xrMPS361z4n4bPe3Hg3qXmkart4pQqTCbDbCjKoZou1YGizrHg2
4VkuMDV2bcsr1pJBXEvlA4nBcBkzocwitOEhmbgHA7A2t1j/hLo0lCZBzqSSaulN
vMQV3LJayVxBIBeZ1Cf3uunMecqvHD+WF/Jy1VX7y8akc6tn6qnYiG4mn9Sk0fSL
d1z+Z3X2gaQzjGs26zzDLsI3WvHFHX0eQq04SWGXnfrsjJoqDFXObzenY01h6sT8
1Gjo3GiE4yklzUGXoHVQiR9h/UUndk3KWAB3SBgoQp3wQlKhKla+GNAV3OzVICad
bxFrLj6oFN92TKuN4qqv4pwrpC5Wy5rFv+/AwfuHx66a1sAZvXpJg2gVnVb6krN3
OmwYdi+uAdulZtSx/5ptd3ppuYVyP7dTQP0gsRI7P1uldYzMIiuyTXepm7IE+5Ge
0Ko6ozr5V+L0Wl9EgjTn2onxhW+ifqujJlgUK3238lphfX4Zmo208X65kosmZoGV
edNhgsQMsUVeDLpoENeOhOtR7wpcDixiIn9nfQxcVh3PQnhd92JCZ07qKrUe8toG
SbAiCZ68+xFJLgoUjaWPBtwRxCPMvLt1WhW310q7bwJDtrMCL+pHZk5zFDfaG4lU
CMVqsXN1GtsXuwFOolPfbwhPnbvbhbg8IhiVsM53lOOjjAetQcAXKv/8IO1RAWOW
8xY8d3g1NffZ8zEB71pYXX7/lng5+I5A9N1tdrJ2SPjG1wzzsV2PCj2YZwFp2X9l
MvHsfFBDXt/ZkCS0e6hjJdUyL/jK/55U9y1IQhP+N+gNJFUFt9g8hvmAhKQtI9mZ
AoDxqvyKvyMkwSVc7OljweFyWXOakFpQCUmyyI+fNRXMBjKl7T1Gs5CiknIfEHfD
ZGC8+iMSX5IVov3apN9RrfSuHaOGMCX+3GJvF9IsR3j6SPpVWwFjlPC8odckJEm2
J0s8tsABJvMrR/goDiAptXbDp2JmP2fiTgnXV7SvsL4D3we61BGP9inL3W4iHZSr
F0obBsEQCM9i06ah6dZZ945VrfLGV3o32ttYqHpolMwmlMtajNAWhge0rbRdSO0x
AhRb5QNyWB5Mu1F92lxS6rVsJrI6qunq3rRT/k900+pZ1MxD4qqkMLM2UWZIBwq8
jAkPtikjAIhxQHdtQmDxmwEvP79aM9LgG3s1BWAP64RqIFsKMsvPYP7p4jr0v+Kg
03ukgVhYDn14k+j6u6XvvRmNfZfpM3FOKkPqGycQl5xyq1VkyEdhR4XsdAEiFyOU
KFUW+G8lc1sW+hllhWyXbcbIu0xf34+L9EtrPuojFPeI0DM5LEm6PmpvUKtd9gDC
QRUCUUgl4+AkN22jFgUkmGqfqAPX+JD2ilSKicqhsz9p3iuNvANmvNpp8UUKKchX
W2PdZb9TG68j88jdMRGCfAK/5YIXfuGvBuhu32K1PcOP74vV9t7mT+d7MRpmLsQ4
qUB6jrmwOLOMhD5yL6Zc9ODc3ZRfcRdlHToH5OIM6S7xIDN7tBtrPAwcsoZqWc3w
EZ5M1aoie5EwnQgTh7Cpmips6IfW/t9e0tv+/5DwcyrNajPFnspwe/1DoZYqJo2g
NHWJGYO/l80Qfc1s22LJBB+mJnCBIQmkseoN96VEjZWlfRVhkN2tOUaknkLm8RRq
HvzrqDmVdeHHRNJrkuTh8VjTDIkOJ+PHvovK/yPkxM1wILHEk75GSdZBkLnJu30x
To/lUfk84TpHqGMydqCugJMl2/KjcoQG5svHDgpZT/EQ4WwEQOKV+CgFIzFyw4kI
LtSZcoB7cqUt0wuvHz5hNsRoo5M/jNz04LIQckJSS2xQQhLsVNJlrKTHaVj3Rpxb
UPU8uJSKAuptelCkNbjhogprg2pm1egC08JSrq8czp1ytuL6daKsB8qhxeKL9HGX
vYZ0POJhfR4yVOnXyhtqT+g15PcpGYMaBfuunB7Du2TbwsZa9+TZJB7Yu2AYs0oT
C5T4Mh0O7vbVt8lThsr4BS/Xtk630RP66StMFE8o35t2Tc0oMquAPhtLEuTl33ob
eY2Vp9PAJgNYQHjgpu/B47SaRM4u4O1YnBVAw+Ocn17xgc6AYEWffn+hI7QvdEd4
ivTFG4pOXRfGVb8FYvYE3c2A6IwZOsUQgJSZZ296/imJzpUC4tM6D5pVWWhVt863
FiKspKmYs+a0M1ydu8Z8tQAE/nXymhb1XIXw53HpS/XkEvg9fyEDFQ15jNCMlFMS
tJ2luBsovyVbC5bE1xDFjdQ/xx3JbLz640nAF8Ke7TApT3yUZMJO3D4wL0vfZEOZ
1boN9glYwnvziWfkCgl4STrKf1vvpYxJT7XFOpyk6dfADHp4nCoxNEoTS90SgXkT
bGGHoatPRmWm1b+PaxlYwzJilT5P57xryXt/PAn6BR6bofr7M6qea0tZUYqQqTZG
CEWV6xmrCXcynbj1nGhbLZmmQBeMUDX0Ptd39Xv6MPEnx5vw6yw2Q0txEOUC7Fz0
pSlstwZu+WowMNUu8fmXMZrfdy5Djv/prk8EeTB5V3BBWXdgZdiNrzz45HXwQSXy
pjTdECmBsyUGY3uYK4aoqxIIar9+ihcBRNEDEMfKXqx9WWWJPqQqr462tNP31Hg6
D5j+wUHSM9d5yGTzb4vQrf5whB18TnIvZUC/FFyDathP201JsZSpdgt0V3ql+NGg
aLEJ+B+5a6Vds0PM8MwtzNhBXblp2rZtWk2QEGE72DpE0w9MpBWnpfUnua715JFJ
cYs1YTJNHyNGquPahbqRsF0not2Muh6gnYsmAy04BOZvp8gi/lYq/ZZODmu36aTj
QNPJl1BFt/8Ev9X0E8D1wlM5LP0LT5x4bJ89QRfaqKpcBVIJ63jLc2MfOvpUmGe0
vJkVItiAcOKmO6tn+qa0Th03M6tv6oVPgaVQpecj6BttxZ2b47tBcnzdFvn+oCe4
d6Fb11RS5iq0Cn3AQxF8EyPRaBDsq6sgdlGftZ2O5PBwNeBwJhyzDl1MPVylf0RQ
fV8AgO/nDcnCut5ki+y1nnC+Sx+WtUupHsfcLcgulxUD5paDErH9JX0cMu9Tehk3
bseIhZ1m4tv6YtSqdhJix7KER7c6HVQZa33ixKtkxUkPBKH7aVLDUwMT0T82ycEx
dM2jlwghmVDRW6I156DmqbTlJNlaboHqP4NjZJDbXK0t2aYzTul/HfD3y8CHeXaJ
ddFhgOV9Uz5coJwnkVrs8Vw+0W3eo8NvO2qh9M4aj67Jf1Ha+akQQViokHyhqpgD
HN6QJZFKqXRXcBx9Oel/2JlN1dJ9fcrSw5XS0BHaEGkqsCo+ZhBeiWRFU8QoIvsk
Jn4rAD9iaBm1H6/vOKJHlF07KGIsb9gnb0UlMh/BIf0dAilUASVs3LnJ1YmjxuR9
FA75iw2FXBXd8DmmVgxJfXnTdPCI+cY1ze+ACfCp7fICT5X73pVyEs4xctrQGqV1
GnNz0RNCiSKaz9unqujjJbXweDTrttNDaO8+LvVw1JIT2/JBJCvuG9mRiTxqtpMV
OOUKhTZ2ovSS7GEdTwKThlIduHsSoNYLm1ApAYWd73ltnHAPr/CKcWrlgCUtSGOP
bBCI/H2a8bxv0c9ee7XL1VxmGskHc1w9npqHFeZryxR0/SQduhoUQ5jT3gCjvyTW
pv56oTkC5XgNZ1hMJT54Y7UJDMG0SuId3MPBZApDywiD9CMxEorgzqtBSXmQ7/ZC
bCIONz4NXIyOfkNLonhtdFfdz9GBm9IagrMx4X61cEH8eV+JeZgCmuuoDjv2Jf8g
vnpanme3GlUndq+u/Wana7qK0SLWgBcAUcG2CAYOvBXXd8g/TsMWkVhXZz4uk4jG
AECKh7wPQrpveqERjeQtAN6u8C3uDdKGmkt/PUTcx1M7yxDA23x2ErYbFH1ITT3U
zal1edpIuysf6Pcq0NwgzBMm9NbpgfXaemJSjt2Pkx2jG1WMyfBC3pYF9LlMgf/j
ee8zPJBsvIP7O1U+pohKjE5nPzyniZIbZU0ffF06zbHiIXGqZc+RQdgS5cXTEAfv
P1q5dLmaxMf8eYaM+m0a0nv7zDL62JBdFS8qGlwba70GZOStUwpupNwJKVWQUFyd
ErgL5IceYoif8rZ/csFOv6sctqqxLQLrstPvKYlnfKLA+/XGbFZDDChEcXZPdPmc
nW3bqfC311tbiYnXn/IeR6chyofTSvCZ/mrxqeKj5QTijN9WScsVuOrxpXJsCj89
dpjSnH1jKys5xrbWxITeGRMdY4o9squnVgoNK/CsluGfwGfOvKenYjcpdSPTMNDp
dG/g4aIrI/ZpmaEiuMKY7d4AZUpE3yRSOgKUBaPB4KcY6S90gn8VtLGb82tFf5vz
gq266CSD/dCcHJK5jQvMwPdEPY8IEl0TSBZOxiC8d1aH1AVpy680lROcf7KBvIGw
lpeH3M6+LyijZEzq9eohzgxuTAelkdLZ4CsZnrHLPj/pZIn/jlEvuSg5pdUa9KTf
Kyi/cFMz+WNJEawG03fYurQ1rp3JGa9VEm2ubGgHpptQ8LF+nWvtmnNxCgQRUfSl
vTxNmSlQ+WLNNhImvzJFEZt0j6z02kWB5XUPLDP6NpV4TElv1ER64qr9ivpidXU2
cmG5ADY+IP1Jg6R92/BnP1v7adZjxHQKzxs+Sk9fP45SRr6B8VxIGkxiBkfSVnpG
LBCOV6WnticMtZezkNFn59K2nJZUvx89EQWWWwgsqGgT8OsN7hVE5Xt/LYjl0UHj
/bSGczaZ2Qtp2coFYPvmKcTlRfTBrDRyDGpaRMW0FRzTJZiWfa0oo5qvtLyr+x+8
KyXvUk/Blk1r2vf1dsBNOkvki9uRb4eSI410xhc8Y3fendk1CVenWefUi5Mn6YbA
HzWsFTWt0/O52UwJG4GCXCvu99dvW3xEzXuvDnXw8x95mqmdUs463zMfNRV/y2zr
uByhJrGHoFGYzQ8E3B1v5sbMv4RrC+9+61+aZpCCw3r8ClsRwi4iSkyKLN+OLQjF
Vgfol0l/RyRHKpAvxaPvRQSexp/BV/04oY1wCo739HUF1HN3oUbaBfvjBEA6HyHj
iIQFR4zFvcbtYwiiftA/AJAYFuYHK/A26SXV+IXpt8he6AlABiLCR1jRxdSSgUJh
fa6/oni7GSPjpFAJ6BhpdkuQEMSeZiiBdufmsSFWhuVUGCkGKUPkmHli4oebxRCc
2PESBGlXpi8GUXHgfjLU+P4cyBRWMwtpz2+RD8wyC6rxTgr0Kscp5kabQJ8u/NXY
cOY1briN2eZ/6ogtOb+8UQanUHhdj/XCqiVnkCJD/iraL7xJSGQwZW8vy/0jfvg1
C6lMu7Iswt8MzgJ6qsmO7AtJX72FQIZ1+Q0gnkWFZnTyPUYf2R86yy+2PuDsmA/g
TX89p86xgXKJpmziJMniUcoAgOQuje+M4ILBNUNPMFfWayxxzFiy0TU2F3AlK51z
VM3rRp0nOtD9LnVueJhyh6T0P1g0RDizeFh7w7hiWg2zKrSYPij9fbfIrNe/pI3j
trJIahr1sbF9GL5GIw7mNvL2ya1UOD4glOHyI4Y896mNHY7GJERbQJfu2EL67N7O
t8N5kqZyZ5xG8+MQkBpnDmdbY9X6TnQ+Y36EZ2W82KJ8AoaGSPmTnpTrkhy41QFc
+6JhGx6IifwgfUTGESNt0kxFbfP5aIO497jWFoNBplHULvI5ISU3dL01GSqYkzsN
JRnxzyj0qYuwOIbC1SEnXEYgyE0NsVaO9p1XrbXazM8SNhHpTLOfkHcolGEqhdSf
EEbOobi+FNjBQpD+gEm6+wk8nGDlY4C8B9+5BZLbZ0ndy+iByzcDwktPh+zneI0T
C/0scNi6nt1ngJ01VRTbgWaqnnYSMmnrwjV1YwlzOZyEOrvH5DAjZ863TzuiLE0U
4F9712cUNnLeRT5KFr5qOf1bGD1G4Ab0Qaxm8RV/8vk/6BT1DjKjD4MxYBIfBKHb
5VDorr54denia2JbBnp6sLHYaVoBVwPB8xBkXyWG5JJbPtJoxEQM/SDxaOx6S1Pk
rKvk9NxMXKt9N0IqHLrt0EhMUO2bjlbGXrOUiZi6lcwSS+7MVR7dpL/M+Fz9wIRF
USaKsmWjLXGvWfU7fhmdDw7DZ8aqWTFVfgX/nP/H5UuJmnk3dbicPofDq73TV11a
ONGQZFsQpAiAETAbZus2TwhqSWBYS5gm0hNbLGvnSTM0am3J0LFEe9fGReh2CTg0
FsDYu9M3f4Rzg4jLYwKzC9H3bk1H57T21YPAeyWD542cNGHjGMngUVskgrGO5qWb
pG0Lx70vFqXY4Z6ryNGP4XRmljg4yqqiXaSauIfIpZEfoZBrbOO71vIF2tUn1Bin
lzN/hm7bJQ4u4pBDIcGfa+06aPKIIc508i4xqqFRvJdZlS3RZh1nDeMWMJtm4PVY
vLurn31yfAsOCQfHa4oFH2JpcFanuoSeZzOjKygISbX48wLJW0TzdaR1MaVhA8Ey
/lK6KGkltcmECfNyxiRcPp2+em0mNvq5JjAH4AEt2pbFzhpH9tWGqa9ghOr4UtdR
h5folGy7PYp0V6MNGJAIyMIUPYGzdd1lPeqrOq4skMl2/CO06O3hnKi98+75wb9o
fTlOus6bRhFGp7gZPuSwCKF1tRZV42lakEINhat/HHXXEkfnePwJ6PyFl4/L/HXH
7orjSSSbnQDJWOprywuYeYhZfeoqaiRBVqog8rJVuvIpZcpC/aOl93aEtFKrcxYh
9PN7pvfry/2kDViN9KPlK0kk3G9Zu/3lq9ixTAushVDpOMASrUnoVn3VafSDce2a
WgqTcwtn9TOF54NfYuO6Tj4cvW8z/0Jb7YYi2h8YQQrznAjuoISJkFHBC2hZ/8gC
675lsn5G2BnQh7JA/LvELrxaOaJeH90+WyiAYqvP76PbZ6Z6Imx8VWTmfgrG4nnf
Ovh/NrS469nQ3fzy+9VG8uT+FredueM3rqZW4XW9P4ix40W38J2WElSWQMpUMCZG
csX/iO0a6n0qFxvdC/+iULnnv4oASMel+anifmQw9qPcM1sbNYQtvYvBf8ggTFqL
eB7cm+KAimGN7v9FWFJSFvDTMq6EVlgrlPxR+tYkFOHVpPp0N9pBQhOTiJOhafJk
GI1CRL1jpkJSBExUnaJIjh9EFkK+uijNq61fij5RvGwkB5JnGd6Iglj9Tbe2R4rO
pEyVCv5XHhx1JSXTX1gxKLvIifOvmWJ1GZbZA9HLUkN3Yz/3Q9R87zu7cp+jNcxW
9sbfz9xfhuZUM8Q9jeZSBqzSpIHmiKSCj7S9TtsNS5u4bhd061qgceLJUPSze2MH
W7SQyKaLSjIGFClXCVXZaMvrQJjsQNLF+6rTZstB07Y84IAqgBtqq+mrna6RjkxQ
b4sZEGzn7TsD+UnpkfRGg/0hMpG0fK+Vx6TI8v+e4zEucGkW9SV74R7bYXJoAXgP
cFZxsolBOw/T/A3Qjlda1BtU7D3iwrbibCnrnlYMiXoMXtYSDaQJCIC6StX1RbyQ
DrLPmxKammTmbxY2DPDgPhAwJy5bULazl9gB8RWzIPEJvof+LuY2R6Bi9G6x78Bs
TzOcGMEx0vMOma+jy814syx9rxIIJP2p8+DlbSt3cm8Spp/5QTCZmY3yFOg/g0dq
1XLFJEDiivqOwYkwPM7HFRNzN45zebRCKdMYEx4Np9H3uRCqJaoNja/08nJ9HNs9
w4mNozltNtz7HuX5ew/iLB5uuI49KbsH5/okrbm6KnT2IVhol7l64I5Xy95nB6Y7
hTJ/Cmn6DEr837Q3t1Av0Ae17TTn133CDVqFK/kftu9fnK/Vh8qtDr9qSrngo8a4
0L6vva4D0BfHH7O9f4hxljcepeRvpI68xTjQb52T4jWZ9mYRd0kKXzl/rRPamqjL
lOaroO+UED/nYpJQeJXxY3Ay0iDOlvrBzlAHnTfPhltNv6doldXfdgMuz+XwEVeR
L6MIZ1ep56H3uKAhXqtqEaYd2cVfcDsuA9fuA3ohVLYkWS3bp6RPIoqvhKkIELnP
48VxEqLk89KRPQjgjhCHVAa8R8dU0wfCggEGFgN0sCWm1VcR8xgXOELMF1DPum0m
JOzGhNs1wBM1kRYNqatD6Dx/Mvti+DIA1Rgd+hHTA8QFiTO1b9i5s5Veq+T+7I6q
dyIcmMJSO82cbXHV3QqyNpCtiP8+3TQSWlKKOmRklza1fOg0XrBUSR93VVCuw/6f
q9PYqJH0x6+rG9qOu1xjFzl9WkBe6n5T407wPGCRUa07ktrn6WqJbvWsRyuOdjYO
3mhTLdUPg7qeiKHT70+hmTDQaKs1f2Yw1O6cVk4AovBKUqypV9onhkuDG56BPXVa
gBCM/3wglo+uBwi8m6r7F8lCYzXUPjlNHLpfwO4IhSi3T8oBhqcf5W1114U6xDm+
JqERTFkOAuZMUTU2NQF7kLgQWwultthIri5mr3ORK8s08BfW5fbfUGSBplS5/sYP
0pqJB/mylqv4eSvNJQ/o23Nm76FQ4Wlv2ByrPPKhHRwYX3PDRUBur6MYYgSs1qW7
Qw0JLtHwgoZZmc82c4dehHo6XjpOaS1IZGckZ13Ob2yYeEKBJQ4Mzol89jtKgYKk
p0l1IW4Fh/V6WOW30yRLP1y4fQFfL2ZWNvt4ahufJIMCIhXrZncRfsr0LbYzFeLT
Snb6oRfGt4BK7bUnS1yROHyY0ZMjsu3rBxrrGetapa2sskVYQN+huC4rH1qVVWWE
ESHmY5CXgxsdi0FXZIKrSuMlQrFd3mYGC7Px9vfa65H2HFyq6QzWxT1G8VroUeix
hJpHAM/Hsax3yHFVXjUxnyWKkRevlH3e46lMMUuktrjlTB9ueF1t/p2Z7VHTr+UA
Z4MydIclhWX2hWkvU1KDPodO53WspM7KXTaHnhLxUmpjuCtwlE0fIZxviA0K9t9d
EgckitTSEQlEAVNSMJwvna4nuUqez7Kl/mb0Uk7L62woPjept/JunYC/qp1QsKao
Q6u26lpVyKK+ruZlQo8GIeA67NULRfJYzMbTC2byVc2SErPe0kY/YUVwY1relyIn
NvDRE0ZReqk3M7iXNvJttrV1o34ToMSgELDi85M5dV0g4Dha33ecQYoK/zeUs4pd
ApYg2ZJMive2EIBa9wZN9GXHbMmWjWEPhpp4n2ZP/CgbXZt+whb6aHZaZYyA8f8w
v58A8hJEtk1TN28JB4+pBW+XF+nxO/PqzFpwkDBLM7epHyCuglpqk9ZjXCweQ0zT
wTW0/fv+CykluZPYWcQAqsJ1RfRR0sLeOrNkWe9QLRwPbjIKx5g24nPOVqJeskwE
gx9X3UuenRnjepyPHPgzJxT76rhviNzbixMoEBn5BZCDhFYD1SMvmYgPUQHUH4Xk
XRT3N1zxPrqamvYumfQdBJyTgpY4lYW0rRYOUmWCI1x+vfxQwJochj1EB81WxCvf
0GfwbIpFAzkNveUnbEeHCOsoVL5GgvjSoi1CvakZVm6NWf1N5LFA8OXGGjRa9iyq
64EDMBr6FC7ZECnxYgnBhlFPrTrL7YzRHPLXCQSDkpcp0L56xKPAMwSR6SYd7z/w
P0EF9jdbMk8hQe8d2ZuXVQ5ELS9vFSveUTWH1Yq6+yu8lcZGVRpJpGASxmAUs1KR
wH32cjhxQKI5O1snkDC8gsUt7j+Mk+oW1poC2lvzBQNWhAuXi3ipGRjMfZSVVBd9
G+zTWzUi4j8kb1UMFpCzA4fnwJZ5YHBHRM6f51DLV16Ddng1m6YfplD/edFnqe+k
B4HiEUSq9Uf0qQv6GMhRaRz/jANiaFMAWrE6qAK3TKNOBZ5442qiz/5hyc7uUZqs
GdWKT8IXP1aBhMfAM9bxhZounZLRC3quFIQTfX26XVTC/aqQED4273GbYe8tAxue
pGvDWZ2SjRSwI/t1fjcgEmzdE/HDCTzYIoZ8fr7Eyj5wf6yUHcyWUbmwKyXci47R
7JrB12il+43Aw7jZ+UDwhX1gJwuLVXW9XHU/CpLRRQxvE6Xb9OX0PyMHO6EqJxUD
AvVtZU0lYwjXQm89SPcT7zeHXMy3Y95XeGQclVwgynVg+fI1L/kD0b9ODwRt7EkK
kGplsMB5JR8TrlS4H5BmDiyv4S6I/1B1dnAb3piEFvxoIYR5RDH/hWRYY/FGgXpH
GJRR0I60ju7fQkw51EohxFxBIYfgfmeOxlhIYUsIDRnHc5XPg+GBd7crWLrq1fH0
qk08yEVQaAKRTvi7uWh8L2MG0ITssuQ/4cUAMzrs1W6AMimlcdAO6a5dMDeE6YXj
kNTe9cmeDHCtcEpLfnbYwytCu2n4I2USSyu5RwgU15a1Scy09tyI+UtNf7Wrs9aV
SQuu+hiekHzqNU9a1Jh10rxMX9ifGFDmebh+AOIyNje9aBUi/Y6WGfU741QsT/UH
jq5KI2W/0z9SOzzx3HwwkyIRYVrfusFcyYCSyHl9hdUWmp3SfT+8TySBkPuknGxR
Ls2e7Mb6XMIQzAp+x7CaXg3FytO6SolJ/+WvPBq6EJd1WGZekFitb4XaNKdoqEcf
NhS/YdpWxZXilkK4RgpBl/D6as8IWoTVNS2SG2z/GZMydgVH6P0ZhJ0qP6tccDAa
OoAtTn6JnLwznbIiIqnSZc+mOCfGMtsY1RoVsZyiCzv+CgsREMOcG8QZilvGyTqu
Obzm7RBukT2Denk1TEO6GsJesT25qfYMh4WYfPaQWJ3T8fZVwHdgmhgc2Qhf7/kp
CV8n9tK2J8qxok39vtQFKxEyFiiUdfmqZ0e6ZjeTLxEwtnsZMeZL5+qvLRvaVOwf
iBvtBG72z8VOy55nZkVhB9K/AIDPh0119QofnZOGBIq/meGJ6N2cuKItlriLP2yZ
e1rfYacJNUd4bpd7fMALQaN0rdcaf6HJO5ecjiaj055mqG1KCDisuht0qPRNfNms
xda0ZJ7LTpyCpwp7A9SHRb6pWEgw7PrAbu+sw4hoMEFjTwqkGAPT2ukzu/q0RXZT
wY5vTgpoxbyTrSXfDFxD0NC+yZGyIUL+NWymNiFmtm7IssB61n3FN4uCB9vbzgCY
Ye/f3ujeuUIC0nbkRLtDBh+p4vRAZiBWHFGfgSRUCXObfIwK7XHz6BkOH74xsA+q
JomPlxWb7EvgLDm4w439uiEkIc5EMIM4oEHKyGQmlRWNQ7GxrBCC3SKegIbYjaXR
wP7Zg1ZCQWp0eiEkTeJ0+DoyYHF6GvAKXU8Kcnm5dMRP6342l6ysAL09xOBiyytg
MUE8/OSJ6jXH52/9A0TOSYw+Z3K9tQKnp7+ZAGY7RwxMuJpo4MZ7WSGmde5tsFOG
+Z54Jn3OZx2JHnjkJhR37sK65L/6aXjTF10z/u+5kW0=
`protect END_PROTECTED