-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WpP/7RMHGuuBm5+LPpRQrvup3m9OIZmoh8Jks3H2eIn219swvmjpYkyFCRlWd0K0u8Bi1VadCh2z
SMPdu1rlIfZdxKqZ9G43w/DnwS8owz7/quC+xsxSN/HVOZfdqf6kic+k8+YZE38iBR1m4dDy1iO8
cPqMVjosZAuPIC+YtEkSWK38lM3RuMLa/Ano22+nWjIk86+QACFVQ0mWulwcYEqt8n7ziYYSNGpI
HbvPoHhPBLTS5EdZGYB9ssKnwS1y9Uq6SJF13MKTEFVvJBPER7LSRGLw5svsYJ765FLNVAooeCED
4hnlBjyALkqWx+3vOmTxYoMEQ+p3ihqfOdUItQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 52288)
`protect data_block
lOOxJHXinX7zkrpvyt72ls2/geVjcz/YrFht3wS6vNcuWKjC+1w16nrrGPhz53XFdLAEZLHm3ERT
FS2uaavPaYglwjwiYoA60Nqn4LAK1XDKlTixLOfQHzNeIxzzHq3xt0BmBT2cbe2MPgFHAuKnNKoZ
s4qu2oZ7lB0GwdEfaoEnMHOo0zoU7w2ALkeM2Hj0BcHipbgCSkckqxd81wopTmALIfqgToHLR970
TRBPtwob1WrhPJ+keYEmTcweau2LA/zKn+2byy6ADjVmLBp3xzQxYffOMfP4CCuO1VZbEWP43imP
40cKxm8Px0m0GNV4IFtNJhl8o8/vspQi/tDIEFUF4l0961MfTTcy/nwrmtkS75fIRGv/F5frkFQf
qbrjcm6mnGxUvs7iTOmFLEHpGI7vBmZOko7ackwhnrgJPN8CRZxiT/jDFcFCbjo2VvrOimDcQVku
7fML20hbArQuBfNPc8I0evIKcZOfZiUMCK1WFD47SIMioN0Nb0MqH4TktCIeHCVvlg6hSdHYilLy
aJ59fKPkaNYGcgC4PvLbEAH8uNeednu61+PTtjxzNrABDV3mmnNGnaN13ElmSykdER6OMh0ldjdD
5/hFWtk86Ak7IRcWCb7mBuU7pjuelkYvB31JQ0k74IFnGAP8dt/HXhySm4178LH4MVQfg95wEHaU
1aqQ7fwg3gj6bRuS7mKuwn0MSKCpHZAG4HYFsyPmtmy2APsrWaHVmxe6FrcTxdugg1Fo4vxgPmMn
zbDY2B+cp8VaY3+4/PLv31jyxJrVUS0qzKHTJRbTlZn0kv71FThvwszRA1hnfNk4yzLf5dEeKmSM
iPNEyPLy0Aq3F+3xKZbiOM/ATVjT0I4fY9MqDOLkwfGRE26guq2fRROCus/S4psQgN8gXXmmwgpu
wAwFmHw1IrBiPzrUTQoCpDqoYvGS1sLP82l7vpL4HKrrYz9SejRX4OIH6ASJkChp6KSm7JtHes4y
qKApq9NzZbAJcPJBEvlzMozbbKVpXVEa59bN9nHHN0AT4uXy880xH29RQSzS8FhtWb7nUKBGe26d
UKogXGiY3fKqN+MwIIpkjkEiBpIVENHWt3FNYQ4YJmLEwfIHk0zqgfvtIBESqLzUiy3Vp9JaeCIC
FbXqDTObKIbySHdMxCDWxc7jahwVkkWrYFT6gTa/a8V0UcYJPqic6BjIAElSyw9XaPCMSsf53VTf
H0MdAgq4FeTqG/OeDzsmgDMiDC//ml5SgvQneYm8nyGLFADDRERU8UStb6d2oac92I8Uzi2bfcTC
TU3b2ZsofKmtM28pb1I/uCjB60DgY/M4BeuJPvTnfsdyFsr9tjuoXJI4LBaTcd+SyOPvu+fcPG2a
4SgYSnstSLQjIAYXLtQTXuv/Sd1gD9mKxMFCDEEoscnfhguLTw746P2+604sjPzXOD27iZrPuBn7
yYWh48P8yurPUPSYib+ac8DdkGu+SX3eWK3U2cGNQxpRbgr8ozN54HdAwu6BrXoq//4C95c26wHu
mAvF/9PtoRYX9xGHkUQYt93EuT9mSXnNEt70+/jk+0/aCc1J44pQplOCKZgqA58GGw9+uMrrP9fN
ekLQmcgwe3ZnFeyvUt9b9LbX1TLAHu/Okoq4yODmZrrQm+05Mi/Qxl154wIX+9QXDnD/leQ/VKgN
Rsm2X/zPW6Po9Oa6TQyYCctCBsnzRGrzfZ+u6LtEdcqooIHeJwOVM3uOet2JSF49SyHbnCv906tI
Mr+5lfCS/IBRCVP9MzxzdIoB+E3pqFdNmvrncAuKrqHnNUNu/6On93MJ7KU8hDGj7FRYCE+wXz6f
NcHzHm5QO73f5znoUxDbPESPPrZooJEQYZE/sEDVmkaUP9xPB2t6yNfri/kkcgPSxHriFQ+Dujq0
sv8K6es2cQhTHrlhKEtF3pVaJX0e1zmLnbO6J8jbQynk2K86mSK3iQOzn15xRu+who/GdacBzDh+
12eKUr/QmM/+jZW0XDtXIRXMbie7FQsznGnmsmAIsEiTE/9zNyg7136eYtr6VS6SLtgyMzou3gvi
g1kWgmdMH5F8vf32GnmKwqTM+LDMLOx4cxNC8IhZSHC428mZYDZ/edPp2h3OXSHSG4wmjJmuKEKe
S3J65MrckMSnUPbFB8Amn6doWCmrg32/47tfxpTNdpod16KF4rKFQS7MFLAOLNHwTsVncAMLmR7i
LxKkoCM9VkrIJd27Sq22nD/gWJtc/uXpd9z7GbdX8oQwHMUoB4gGaJy2Xcgw5GWIMulTzxl3hvYy
u7x9FzgiTKZOjtChervz1undC6ukQnyv1XVR7IIkfXAKwm3osQCdaUpfn262BT185d+ZjKM3lEqy
aLyL9gpdYp1b5KspVx1sHaTr3uYzgGPE0niUOWOqsUzwa4XMFnvRbzK91yYLOTw7syDzcZPN/dvu
OmYLMvtt9vFeY6cCoowAhNytdlvsT7CJsFk5TIr2sgB6v0adkP5kOfGslJ2XjJmHSLXAsWB65BTk
jbvDMCTqHDw5xzfScSJtV/1srcwH530UjBPKzxB47ua3m7OWd/GDq0MO5qoLbKcSwOJron2nHanR
n2rQCowJqLn+GFCQ1AgObdcvnk5T3+TRQ0RbelhGAfYnLQFiuRdR8KARpRJmLQHLQ8rx0vc00Z2+
uqdWJEcoGp1c8+X9ALR7U9Ua3dJtyFpcwG+UCmd8rGePGH3WBGd1nvvfYHlDkLfbJewr114LH1Tl
G08oq3ck4e0LRzJMXBELBPHAyZsCc3AH9AuL9awbLHyNlmFBKC5q3x/duC7bqeWXRs+uqU+6+ula
05OA6pumdScHL1Agv1Fo4C2pwcmlnhc8Bnh8X8rBU8VwpBudypCZ5puOOgZsVy+15f33DK+JJFJJ
4szswfAtjXW6gzvYuuthN292a+M9fPYlMg1KLhmW8vfgYjSgOeGiiDpeSOcYdGtJoehJAiKVjRMS
fdscS+DS9nAX3UoRBG1rA2V7hPcGlAx28PDZHQ60UMx4igqx3h58QU1jl+lqr1thmOh864VX4BoI
dtm9Wbh5D1V9qVPMaBi9toPAbl2TLGnm5BfE0leHp5by0s+c+Xp7U2HNviNERS+UDwYw3rhs+Gfk
/VTc33VbZpOTInlksJvgkKtUHKk8fM593SCXuT4JmhJyUoIOKeftKVfz7H+5+SzT1Mp/N/eV9Iul
f1HA1wQG22/7uvAzM38L9xY0zVWB6uk+qZUN6FSIudSYxZmRnwO2HgLzUWlN+QLCl96QeE+Q+7RP
SC5IL7wB6exFGNDyAapxnplanNSga5NL9J/Dth6JfGqGF7fVzHGAiCOjcnSuUqnbFEygOLuPhR9B
iqTiFfFhFJBGcUSX+tXu4yzNilyi3j9l3OIGofB/AJS8jURe0/WPDYb7cRRVzsTaVu1TFJIZCXm7
lJ0vMiqLWvUkRkir5+aDw6jTYg64qrvftm2DaxlzaRHu5UYDWgSgCBxUB1ZsAxZotre8yRov0LT/
prOu/NbvkTlrzy/jLY1WnwtszprgVkZXGOZCuYgkQiD9DfEOc/zsN0QalcNIgs0wHsUfOg7sJE2g
wP0JZ8AIx/itmLrI5PfImZHclj3IbHcYNkuTo87rmHbz37jNw+/2j9yu/BRs/yTxWs0Qu8wGjIz8
nR0PLhf4x3l5Y0ZUKz158TUH8Q+RKrJJ3HMHy7PmDR32uyGzOefMN9V7Nj/7RpBKC9oxr7hxiwFz
D+/bEthqpDep4W/wh5W3cqfGw2S0pvyYAiKYGpUiFXN+wfpI1VXxsKZgg56a8LeIOJQ65jlySdai
0blmL5ygTuEtlkLX+b1Q7tZdSnEiEezZ3ZMgz7rlYRCQrrM3pF22TMAs4Rvd40tXjg3S19tTjNC7
jPqcRtI7oyJ3fK88afV3/eLA2EfzkVzGPZFp2dbgELVO4qPYSTYAZA5OAiKzdkkftnYQsDeshcaI
oqDIbh/+KU/c2Z0Pf1m4WMrgPoNvvmjL19Bs33S6mvJNXFSsdGpd0aYed3x7IV1AKk9e27JlX6cb
OjS4/ilqGaZw48FxqF0h0OsLhT732dH81otfMFjoCkGZ/+GqRv3ofCDmxpS+fHWfBJm5FGvEYHjq
Zor+ZW7JLFiRs2IQs0LS5cd1yeKClP+f+yCxZTRrhL2eesjmojABQzPY7ll3y2y8uYa+s1HVELU/
qrseOpD6culhSvYOqNF/HWgkXVUUfEJsB5cEbNQJ4fzQ7h4kqa7NWxMbOyjlS4zfXq3zLHZwztok
ZecgjDPUN5ZJmfWZa04RxTS5qDjRP6QTumwqHW5QSr4NhiJBw6VTCMruuD0+GR/IOtm46o4Es0eS
zcuUInZF7vE2r5pp3E4rRnYbvNoIK5fN5vfEW0d4u4qtlx4dUMcsqXVSIWeSEL7DAv1fLWx1C3WT
dUcX9l2xstaze3lmf5oSyWQ2CwKPPwcz5jZe7bBazmXmsLonbNyU9vaLmfX3lvkd9Iz3NlcPB4Vx
IeKfgiKE14IZEpMKsRjZ41gXZDRSnHIYc8XZAsvw4HMVaL36PDuHJ7ezP2i10Sr2XTnjhfv+JcaG
JWZtAZaD6eFVviDT0SvCZfUo4/jS68dyzpX3bhqa9Cl6TmAlleFi7ongG4DBQRA+a3Gf0I0Kxak0
n0LqyhbHrNC6kIxgHONQV3kz/vGDRqN5txsHsB6B0O49jJ+nactj8X+iuW2RecvC0X9xXek8qZ+Z
W4eMm18fP12Jwth78zIOi7S9pyButz9StjKfLnzMtbD098FXdinalXBui+XxnyFBThI4vmLFuToQ
gWNp8GiXZLAgdvsp1LVC7wSZKvuQcWC/A8VVpeNlmTkDIAb/HiLprbN0Bou0SX+df6JR6YXqMlFQ
n8uJHFDdbdrtC0kDVTd3hYx6Amg+0aiiekA68X7Klk63Nd+UOMICksoqhHmHqOAxxZIoPNHNHMKb
KTHsu2XLr7DO6p4PdKBgWsj7nfOBCM9SSXv7Fae/jD5qo1LZjN6XYlhT/+SvQeB2OgMBx9s2yZPY
5JQEjgz8NfywLpXw9CXssPcHS2pN/67v9rjaAbmj2FyiKBz6EnWS4zG9GDkeFuu/4rvMdf/NkGhZ
BWi7Kx8cckNRt8DgJsWCbU57Ob0BWmkR2U3nxw+4AquUBo+0Q3dEOTBblJ0mBV79lGac3oFDwhv+
KwV0Dos4FF/Xd1uF4iEfoUNYi8uIV895GoLEmPX5fqS2CJe6nvRwLJwNFr7fFDWg9kNiEcJAADoJ
yY567irhiHLtsTcwHE7jFiWOhkuOLrbDIsRA7JoID0WPFpxzJ+TmVO1tHVx6WU2URsL8A/MOIHIs
FyJqU6HsZokibldhPu0R8iV5blrmxVqsd6UCdQl9qs/C0C2r4tCO+BrR7buWOnX3zgm1OESWwj2X
cNdVcDCDPbezY3AL7bSUrR9F07BYwoskjdaeRobx+pG4zGpFS9w/Vw7jfPaHIdRDI0FI2qqj+0nM
gB1RfNQY4d+TSTDtD7BEtjP7QGcFM5xYHQVjrcq/1QR+2rmV1FoWm8PDOzjFJ9/AvoQ7pBfspd1B
QraqN4m0GxM6+CppCtoTmhR7kFGGY+uzN/i2ZsnDeqdxAvAiPgSNwiU0vgzpv1R1cQzAl+MC2q8Y
SBkyPsSndsVS4qBuDtaz2M+mmqe3j+O7hhNMMalQKyxGW9Nj8a0HJ3PEmkj4aYGp6mOJTNq7u2dc
vZTJUJqbQKb5rUl50R79px+OO06+8PeF8tLeOuztQHbSU1ynmiSEVjKDPIMbot4V/D+MqZM3UQqs
6Cmv0LNzz3bQZwN7KOLSbfJ8ETUT6ojzBNcGet3OpwrgEkkCoaTvVEYBv2YadN2Mvx+pwyD2twpu
+vY2S7vIUYECndd1aiHU3rK2qvBpyHIKSvOf8LKP3BBtk9dVQTNg7HH7cUk1xhUTb9t5nFCrxfEf
7ZbJYDcIuGehRtKTZHY+fmKfL4p7GY7OqR/PqcPPTciqJLQ/c0rEScPRBNN22ZAWmie1NeBKTVlw
n3CEvbe9pLcbxDRZDeUK1gL3lYEH+mxGMcSTHfQBU0Tr23J7q1smviOU+YFAdl0FNSVSs7TPaAp9
Bptctc94FDdr3et0gAPRyYzFV8G+9cvcf0yH8lw4WvjZ9g/N+dKPazZuDPhKuAEvC/7V0fp7niYE
F55fL/0t3/bv0RVWWM2vvBVPgvVILvYaPUbasYnce9twXssNGOalJAdWPrTJkm3j4Kur4MGVadCW
pI9bVeBQBTEwGIX/sjxEwi49AGJQNucAIQQTv+yVEAvfk7iUX30fmEdWlieOep91bv4aStNEJkCw
CzSCXLUJlR9EJc0CGppbZAamcu9j1ET+bQHTPNhruJsgBCxv+myn3h4syPO5sv0gh7on+JTicZc5
I1ZwC7I6GjLazlW5VN81B6eMWfYd5ZezBfBt5ZvVxb7VpSvcV/RqqVLpehiJa8fWEy4GVrdPG2cw
ZMcO2p912qEqi4AdKpLSdyIuqxDIZWknDj19y+PkmQpxDeos6nwEL/6ubqfPWbke6BJZBDCltvi9
aNdmkEvSXJWjIYkS6DGTYzlzRMftqzFbN0JF/ULeE3cYtzf2FVyENfBWkhnTM56BYVd6BkFggoRj
mDnUoZ8IxVAgSt+5KnfozRyPcACaq9/5TikLkGoApUsKnqU6kZWEeSzLrPeko+h3O+AnhBMe1oxp
Ddi2ugRLISG21bt98o51t04mVJLO4Ik7Kxd21qsiGrHrtyOxdYSrtZZSi2b7aeeOeqYNeGlWdNdt
HNHS/orvvWB/sS9kBgHUqQN8D0ZxnoCjTc+jXcex6UP6+JJ7UNl40waMuckMeNhWlToDq7YCzv6f
ntSn7sZ5iwVV2THIw3Uxs9IMt+laBlPhNYz+/rYEUH7Q9CbLEEEe9Z5dPg3o8p7+rC2qBjaz3U+g
TyHcuDy5jSzae+6sSLnLUYfKEDUyLftwL9VjyGbMF0g2RiReZfm5EQ1ZCiWE1Kl3bZ6rnhbZaUp3
HeyvCg7kVl0CRnXTHHQhZFmvwZkX6wr7rA+/LFis8VkoMZYXIkk6P8Lsu0c+4iFh13a4BIBoheDj
HKeIcUX2f82SR6LeC+4xziCURZf1bwAk/O8WIk/Dri60Bawz6LQRT9hs8rauyysyBSbSgLxDuM/B
li3CPZFQa1If1QvUA514CGZkUPqYkElyllSfuPk9HSDRDd25/VIf8h8zWSOeXfN/unuv4snjZpXk
LIYoyAH/Ii1RmMPVJJcrgGkH45Ij0xXmJJNij3hFeY6icBEGsDUkmh0k7hiUF40pjYckVyK3CNcY
LrUVLKgkl8lvyAyeLuo+YANsvx1yqU2BZTH4tVTXnvZYkzKKvnAKU3+15k1em4XeVNENezzne5LG
q18KvVjA+SOow66UD/mPma1o5xd46znQl/LUlOxPjoL8vGCbzIgWi/UaznRsDjjzcwKMQGmC4Vav
3F0KERfZr/mNkJqnDf9FbOpQUdSf7grcRy3sOStOim8C6Jsx6eZpDC0zhDgXoXQWABmvB+m4ANSh
39+F4XBnBOmO3syfcv4zj66SDHov+qe1LdBpQZw9NxX4azsy1Tvv3AVGT0/RbNh2XrqTRTmHZwM3
xR4cbfXX3evrG1zXcfqDN7o/V3hrgcO4GSiIZgQGs5YslElejronxHw0vqsL1t+TsttyhC0BLJTP
y73BcVt3+rBgkxuo8JjRlviY3buX+JBP5ojBGoXkdAdURWtckDnSt0vE4InbDeNWYY94lgoCOovL
DP0G2K4stzzZPzfgUhNQYNNP5deHkjtmBA63Vn2ecfZ7joLKxzZsMrKNO7+2Soh8nZMNh16C/KFr
Pb23R9YDrrWzpakTFP+YEtADOYsyP+qysVuVvRk/5grCDURB+J5puAg0bueOpilcbP2tPyEaDsyR
LLXPv74mGAjQse95LtcEKESrbCTlLR92Xq8ibhh5RgalKCDNhSQvWWns4UMuG80lu4hJQPlQTtOh
3WoHt65AJRXdlgrQ0cc9CMbQlf3CKKkUD8SpJsL8H7rbi/r2PEpFKabeyeJG0RsFKzmGoJ5qY0Bk
sjBH9Gg7LYTsuXuRgLp744BxhUvamL3JYqQmBzd2cgm02lqg3sEhihR4PQT9Q5zMYYaxvXq6DsEC
qTwRC8rmY2I68T/TqVMdSh4m8EZe6gDev1Rps3ozkg3/W/hFkWPaWzSWTiKZKPTVvJ+PWZ3b38Xb
QOXhlhfzwDM3+9wEN3atd7C2+abZs2ZEHXRQEmH8LkxpnfAdd3JUO3xHd89R4wFOFALIl6lmyiOl
BOrCSlOkPKGPe/U4kVGM/9wtNMBLpOw7gSZCezk0ZAd0n2hRvFSNfcQQndSHpuYPHbFmASEyw5J0
FUnk3L1fB8Hk6CRCJEEnqvf8usT9eoxAWaeT76N0/iHuxrv7uIQ+Y86TQQC0MygmI+lvxYcg8SGX
viapSPw+c15zMyxZ7a3Y0a9ppcvE9WjCeDq9rgnzA3A/GI6BaSAwVfqTKe16f3D8Tr1mcf1pyWi6
crzcKc9TRDdbne8LwJg90QuPUMeTNOq4DkzKEx0Ht50wikl2XZJTTNlJCeRg7vqOn2wMZZJ9Sudt
LFyYars+8OV1utJ5D96As807sKLxHQ8qgwEREInyKOx46xUeuFvEEDSCQWiRxD2IDt+zQGG38zD+
KQAVC7CazIT5rTeksbs8VLiPDMXTMQfMOT79uMvHpPMozYUe3YHPPcf+Xh6bfEpXNfeTkq2Z2kkT
ED6QqiAMjDIZKDK+gScW2Puy4zOpMuTZkxgv0kpzSXV3NvwHnWg/MzxbElbi3/kXgl0HIR7WAHNZ
kef/UOh7oSOde0Cxs/i5q2C4d5J5SvyMIS6qhkgDuz/SLKcPUEPwWONmWiHhF331yWw+nK/LFyZ6
hbcKrMHheuY5GXVCEJOWpFntoSWtUuYQ0cLG9TQS5qVaDRT7mBfqxhKTlCkKCL5jvxaX6zciPrem
xOi8lSkME16ASnYsfn/xfFn+njaGrdHTKhw2Q1Kk+cdLkkNxvIS/ywllS/+RzINpIDdFEMyP7Hsa
noaoE+Nsc1rWOd/NW269oUfO5GsaMg12HzScBXKJuCxGj2VsJMMO9pm4vHDztelnCx8vGue7ShQn
1qkPuNXhAm7zg/MH0WSejMXLV/epkOi3yPgXC6AJTYyrwn0tXMnlQHAs6B3bpXpj+7T/+KeQhFoD
wpXvwAXw/LzT0g+qcS46/cO1DM3Mcam/OGRpDWlo4GEKlaXNwsCFwGD+suSG0apGQPuao0ME4HXy
g/uW8unnIar5US661GBKgptNnt5p5Umtyrg2zLPC2/vWYlrbCfyM1kQ6Lus9wotdjYodDjjgiSF/
N8jdT4PtjbLtajPDUgARxLhvTylqlGcTNJ1ANYrIwtzuPcZC7vvH/oBwehIKNKDrHjjBpYjleRLN
1wqvpXCdypFegPVeW1QOR3eXDAixj+RH6LsK/cfdYd5sX4KK3Ed3ZDvJqBUG7ulMkRFZgX+c9Ygj
q/qP3ExrAKJVOPEhjzvzmfgTFEOBW+BtQe+bDZwD/n4c6+3Az/41kOzxTYQIFLIAqJQC8CFzCYNr
/bM4BW0+p9iau2+91IX+TjRVRut/GwmqiJCUij4sL9Cgbz1qMo9eHAkXkNPFXRTDejNkLgGCoIT3
AJ12ztoNB4q462oEvLDXAGJ2hxDwPWfvLxHRQC0HKiHGoYgm4g4OLigdIy97o3hJgiKoRJJjl/JA
rtTtreQhwapPnsq06mlUuIqk8hkGb3YD5X1cbPXZNGf0RU9fFQQ/Hn0saKNcBHuastWRS/78pVSs
rVXsjfmNwQ9JMX1yeTtWUkg0kLi1lag7NDgTE8gHg0dI8k1wkee6uG1lYu00m8t+DP73xJp2UgR6
mcIHrSMEgTQoEIQOnpaJ4J9VH54Ajz2PjpypyQLtBxlshYgig/MkzQRXOimtuvS2D59+rbuw7zMW
MA+x3elYgHeSlHlhYOYUcdcR8cfwQuwA3ljHf6O4h4kQPi8P8H2u55fH7SajTbULfWTu9YGpyqZf
2+cORAhyXG2xuePKeqc8ur65j+vyFRx39ChDmu9ghbydYBDfEdykFUevHM4hFgQmr7rOCPbpblXt
HEwZVX8/g4H2WqoSh88HuUqb3fNHO8wbtcTqhh6ml3k/GGa/qmOPt7EuLV7Je9AjFe20pNP8Ghtb
y9O7v15MMGU00l7VhhG7Yb6rPVyvMaZ7RCKaQnKeH1hG7Xik3HP4sAo5/gCU1jMbTf+Bwd3IxFkd
G9OsjcYwUmixGYXB3yHYZ519kTWBH4t8MjSwbbccYRMIpWHvAHRhTaQRJfd2f1IkVsNcKxMlp2mQ
YOYORaxAhGBSx4S3p7JEARk+HRN6sm+tzIDQF57N/w8NexSk0bwKGMLRUcaAgMC/NwUWPaLCI2Q4
UQh9DvMLRXmYg00C2m1CFsaoAxCrMuyfBNkAajF8oWE1RD/lKIuk8w1dVKy5AQg6cE35KCeQ3Nxg
OG7nGliuPWvRZcqkshkK+ajpE+tYm6TcLDCmNOI87ZEhJfAr+oR8D3UUuPUIuELCQtEgcTTVxmgC
JnRw6ZhMi3SQ8orGnSQoTEEGc2yHvZes43afBwH7CdCUzLPRXshN6T2Pxczim0DGf1zZoUElWzmK
ZPrU8leBa/iXj9y8Ukay8YDrcOj3Aavwitu5dZcPbbtxv5Cs3Ry14v5v0JyLr7+4qXMBiqi5K0oZ
znS4a8MyRpYKAywPCZUlCEmpLa8Oo8tmc5Fq2hrNQ344ZWoS2B5C2DXXXkS+Fb669W4SPgWW3vuY
fZw/syY7onsLLePODRglm2lDLzFWVeoGuxL2BwGcxpzh/hjO/yHlvFRBCCdWm7ba6aZ5M3n80J28
R7OFZFLPWwPpMbVpkYjGmnGOi/8NTmx73X+35TmMu781CVC6wLaIwL/fGwWydMEsD4mr9OdEecKb
Yhj2zZ3wo4AeHwhWdj5GsobBycY4BpBNz0Isk74PIQ+WwzgnqbrRfeLfyLYOEOuCxcydPnKdZrpY
I4bjPSAPioaaK7vlhIRFToBGLZidy9lsXDbMOhUm9VX88vq0hEQLfk4UKvPeJGKCUZGwMRSYfIE6
o7q+rr3Tdq1ash7aWzy9yJMp97nSE+Ht/oKMWtT5L54mikPqbv0QMO/u6XHA37lHiQNcSwPzzlAC
4/zkT5sEa65ACooR78zSh2X0JLg/Hx15FHmnCR9akrE+mFY6w0zo8kpC2lvlsvwbBFxA4A0HIzHW
dlbhOybhhxThDjt1FT0qzdxsMfyw95p5Y6pwKgzoDb0HCzL0TGKuQQ3zjUESCY+S8H7DwiokXvx9
QThpbOBCIj+55WS936p4p6t1I5UDPgzJLRyMAgMjg9/Bc/D2+Iz4I9C7/T9B5igHinVGrI0eNb1r
5mC/LJHtfNelkUoov5SpJb/OzvKWE7MBNrkMCo3KyOab3dG9RYFlVsDacuCKnskDcQNobh0XeGaz
azmKE9C3YdMv7KljcPFXrMmwzV3XEvr6Xp7d0saqs7vDVTq4N9VSY5EM4ww5XWu+j5zqD60/sgkA
ebgUjWumNTo3zXcFdMDuxHzkZt57sNHNOVLvf+pezqWAjmv/tKC+beB8NQxWcx/nnFnZrk4jkNyp
AD+GJgiTsdv9ThuozaYGWcAFTPnbiVgCTLbMWSlwGigj7gH4827grErk+elrs5MZ68OyGe+Mn44X
jTyi1x2lFJhDhYing6GmKdpgC/Cur0WRHxeMUuXDNgK8lXgsd14NmsHEqZ96lWf11EORMjzxCblu
uQiDKhrEmHH3PwSZhCQAv23JwpJaVJT8+o/mXOpFMSdLpOA4oEp6JQxw+KwBZFoHzVSClUw1mn1L
AN9BBh6OoFK+8Gw+pYeTsssl8sqPIpvthQTSs1VebC+7z5W1eFTb7ZIeaFGZPHHUgSEfTMl9JhPj
3NR15/U4wQrSQ1YCe1TF120wkZ1/NYkoeRSCGTpPLetHyOcIgoUAkyzWFs5GSFUWoirlvx3N/CQi
6J5C+h4X74JzGfuxXfPoH0lQCZu7GcVfX7QzoVABMN9sjBx6KQKpn7Be6VjY/ZTN0jQlAjieaYmq
kvmH0Nxace7ISx2fVED0uMkmtTDusMLXwcuBueTlOQPNmir35O+1Ad48tgNXcypN39xgv2i4gn4+
h3HkRXtPPcELq8KHxIMF4vVCKop0gNhAJxp2TnjLcCDkIwyeswMUMXAOxlpgfOXYgN2fUUniN0iP
1WaaYV8N5EBTFLAB9EiRBFVy4OlWQ7F9g+w5QFRtTIwsINA008SejnvrzpJ4BguBEGASFMzNStk7
tex11hSpW6qrJecwMPXuX9NWWkKI0Lm0a7bfcUISK1M0Tz4T2uyqDN3CkWFhsGEtMxYc9tqmaQAV
Gym0Uz/vqbB2VxR9EvCnOv6UPAt8Q/KOolE1Eux+frGEa23HOR8qFoXwWuBUZfAwvFySb9qcfSNy
pR9VQ8zahmNgeVxqG+hVbXQYpj3IfwvTIRXRSO6yb/qe5QAowLFE4JBck8ifhMD2+zypCXpbsn5x
F7U3COdIeycB73mbhx1WgYQa8AA0WpOyuqAhJVUIYXS2QIy06b3jFESplnHEUIjrXnXnMsV0Xcm9
YuWPlSLcnnKow3v4tLNikeG5Nv4JKt5/DCxYYPLa6hUbCPPqn6M7eeDL8Dp8yu93+bZfcTa6dmaO
BtFkg7iFDKzoC9UlHPnsjvv8w0FbeObSGwYD7d0e3wuv26ikhmKMXl9YJIqHeVmYtW5dpPu4XavU
6d6JbGm9Ejf9Xyw3y6VDnmQFr6lA/f2B5k8Vnk8KJuXcVrjJYWghLwwl/lNETtHvdnzgFJMDfAea
N04tmfCrA5bwTanGsGAc2z+excR4GSjFVPZovgyVKV/vtc4fIB1+vhVwlgof/KmxXNrDecNpxgLj
c4K6pmAhuaDPafzB1BwrN+EgOFuX4Uep2+deeiBU5tNBnfDfyrR1oKIb328WcvG1bB6LA34Qjkbq
h6B0MsyaiBvwpDeBHEAChXZ8L9GodN932Rinwt7ShhQHLGOkCf+ZZp0eHi0AougD9iFaqbXxrpgf
KlwghpJnomLtguQsKaM2VyLprlCUxWAWbRJc6jYtrjq+3S20mc0xUFoPr12XLrox1y/fnr55ZL40
MTO9w+PYr1W2vESp/xgZqKHZy4xTGDNrxVXOPHg3jU1ZSx1BafOzbUXqjOV3HJMMLEXEtcli0u+p
gyPe2NtA7GmZHsBb6ZRQ4PO/CDMWkU76w2Yyu3DClT5PGCE+15VZ1E1fz5Im4zhEga0c2NsGzVyW
edzV/Dleb95Qunvm+E+ajm+0P6iaLg2SouQSxLzXH3oG4OZlkesPo5cjDKoEizVL7uTdMsDVRF8n
KRLc39USn/MGy0wsp/72cL17ECeUTrbEl8E9qBXdZFGiz+EGTPgwyrJ97q8Yf4k/AJe7NBfIihqW
xCtjcwnl9gHdJVs5V4BYmxb/T4bdIr8zCjLfv2KUcYVVApOEEm6hctQUoyLzQ2QOxFdHlOkcGzhS
sExg+3ryxGly/1lMvl/Ok6FHlsvDgSsI2pSWYQ/RRJduU0kmIVsgvw1ec52jBPJvnNxPJ7cjsITf
HBghb6EGVmdo3KhNrAvG7NL7fN0Ep5rGMBiihT3IIe56Is9moVdNAHxiyK7kjHHRPxfpnMNcpQfx
WNeU3e3tMYpr3qUCE9G3I+brGj0YHmxvbvSq1iJQ+KC1V1pJVHisa3cNz+ZmDC+rl7hZZR8VNUqd
8lOLCmG/LVTULwMlhiaJL1Z7Q6Q0d9U7FdMZJahje8ZUojqZXjLNzowRV6B7lcApg0omkApa0Eje
Sh0W6CuI0tVG9IE9oqpRNhiPc+cVtdTAwMrDP1Zo6SSf2r7NmZQ6OWqYOntp24MHVBRc/LAWMehK
saqZVDUMXj8OUNrtxvUfVTIbobNwA7AwpMg1I0r3VobWdEu1tZBwQ0imJIfRkp45oKIVbzoogjIP
tEzowasZDGfk6jLcJ+HSc2vQBR8zRgMzD3hNQj1HAolhZARYhAeN6EI7SEUZTGBK2z7Q/SzStEB7
AbKIl7MZH7aqglyHwhT/TgHRUBmSYOeVo2r55wX6ch2pddbZsfDDmV3ZfY/JIEKWrJ8jWTaGne+z
HQUWtO8MXo4ETzMyJaR/dFtEXiAdVVbjcxPXvcsiCIG3HYPtf7aihKeeeFp+QP7cNi5/xfcosPDn
tS578hMHX5OGZAgCkQC+Hw0M/Y5YJD/DYdPx301NpirTcSxgue/VxtHV6wH4SAeZ1MFjS8DAf1xh
W5ceaz5vs1gpyW2MyqQ7nDTjJaHR2kcxEerx1Hk/M1gVjYrS5PLsY40QcQ61g8OLtFg/rSAhDHFl
6tatydqF5yDL/QEk5OEcC8+6yX5ds2yPnT+rlussJonFxAU6nJX0oGHY8SsqzMsUQy05hmSOekYK
7xGAvcVYtCVYYmZbSCAoQzoeFyqMHEjKEQ/Kt0aiDNAjPJX6vspLAGvWpA86AF5RRmbTr9hCTAJR
/vAsmgRD08nUVBrmxVTmLhUbPyr/KPzlolgUciikcwR9i7dPx5aZrOZu3ysY1IYNZNAp27xNrkWu
rjlLFFJGyxsFTaDzVQNBxtETOvuijBOJg06XC5ldHi+92tTXwpsgAmHpOg+h5U+fmO3LicSwFkg3
5pSL+sg0QusPWLZjoNwAdL3ZOBB/oV9qm4suqPQ671yqBKkglk5zfKWc7DGIfbQcSjfTszLLdOAG
G/HGyebPLTr6o8CnhRvIJYqD4Ct7V/G1+zSc0rV63qT8DZXn8g3ZpUYO0M/OumSbNHH2zspbOXkR
qcnPud+CeAM70J/QR+UutpxXznWrojUBJDmGYWiqPMrY+CqrE51ISLzIHWngONCS27fMxn8iAHe8
Wl+ZgzyCeFdPbD92CKBKUF43FCIV6YI8lCx26GwQVENNDdXGYQuaKabvDeYUQ7q1I9m4ZM/ugpci
D4ihtngEpkHfV6yF9rPkSSYi86xS3Me+u+MXIaRgPYWCOZh8awnntm/po5wmHKZ2QQWd++4XFfES
HIrB7Ce2WOjYW52XT5xlygvPlazmLW5t75UE7cawh8WVQYy1GSHPEP9M0lMBMTts7B2jQ+k6Mvsp
XFWrJrcpeZx6+2DfZGa4Ix629sVD8fYPNyniEQTk03I6N6w28AgHlboRVUCMwloVGVU1LFE3sL0G
ZB5EMCwKR/kp8sGEVlHynjzzkKhnzbgaKncpKCGYoU8GiCBVLAGqVHjnhJKAXvwLd/pEEH5H6YAb
HQjXTkeuYGcXj2g7ue120wNkelj6X/fJftdVqWhsOlnSnTtdr645NjxNX5Chvmq06FYxlhd3v3EG
a8Vpb8B0MOds1yS31LFZsdcXMBb/29gw8J1Zls6MA/s/rLGpXFgbX/By8RL4CplCMgCLjVpg5UJX
s5Xuk/K7wlc9o4b5vbEDkkupy3PCgsoh8riAdTuUO5EHhiSILf99kcTYFmQ+mcuoeIlWSZ0HSWJc
6cxZtZsupDqAlwb1Z1ORhCuPjeKBmVW5c/CA/9fDKsoPUOUyL9NRNR3XdULTXtvbLJpqwj8+yzU7
xhZ8zpiqcsKzH/6SXsfTXfApBaqcUiplllnP+/cxvZqjZfPEVr9U4W6Vq0fbsyYbrvSkhrDigda4
Egt96NeLNVxs0zigjcK4rDjHffnMjZ5bxqrwVGzjjdyji4GuJiP6W5kLY2CbX5sOk7e9oHWMclVS
Y4L0f18jXPU3buTpjhgi6NjP1vv7qwOZBKLyH8k9uJTKL1w+FK9U9X6lX4qUJnDj1p0GfcD9a4ev
RqfuFQhKZq/xHME2Nwei9F0WuXlzI9jNwOomrlfjilp9R3b0H01rT9l2ZviBTRK5zetlCxCE0Yos
ciBrO0AhIJeaNniL08wFHRmSwgfnDJ4F1WkD3A+CC/bQ3fjIx6khKAGezp8GnyHHac0nasRHKaGx
5xHYW1N0/zHMNzNuJaKOewu2QBHnYVbaaObn4pDsiHcCXtERS2glHi/53qgIOvc0LZ5zkUjvxUsP
wo1Lcuuv77PpoEC2HIqt/Qp+IXJMKqyEYVeU389REhEs2ZBktKgeIa1kDlUc4zh+qlsvzAdIc5G8
6uXVjVtgWJNDOzI9Q5kTZc8CiAYMsL7SDEq51PvZl91kFgvMG4JJTi3Ve7631RH9ENB5laqmjzV6
sszGHCFsrWx7O8/O0QtTPjhN0lUywomiAPQ5GBbQnvyW0RRlqgqkDyjfEyTifXmoyQ2kgG2wKhDF
LLpY3MKQvFpEi5vM8LRCoidkhLMA5jjqEmvuB/ZDCVihmDeZG8v70FT3CK69hsglpBI2ToZzoGWU
NXEv4pLwCb0yV+RK7ByDL5Ch793H6oHQuH9fSDSdj+XpXJLUnAnDzEZovzhia4TZWUbLUdcZwjx7
1iAyUeBqrylU14M2S4nniYV5oAmsgQ36tvsnCAHsZTTtOEJwYCIazGBuZFiu4QiixR20Q0Oa+cTk
8ArI1svHzooAdxpF1UdFYb4cktLvS3ED9RFh3+THbyJN52L/Y/XC8QkTOPNcA3AHzUJPSSy8eoVH
Ib8OcO3HUa8DrnJBP8Qg/uvV3DYDeljIsL+1HBWy7Hw/DxYfabNQrEw5EzeWE1rhnd8SnSuhAnGL
oF6yBcFoKRXzjNEKofh6iKPk8aBCpy2l1nNO/y6CF+uMj5oh+1INY6pFAQgS0EtfeXPE/y2PCx/y
+Mwx8MCzH8pmfMvmewkJYKQln4kfP2bViTXty7vbWVX/yAw7ksYe0D65bHpj1FEdZJpUuT4fL5bF
PKTdQyUZF+2dQUP+CNnjUhwC0gtgrAQTUb9quMyHzvVLRZNDUuMjVd/95tfkwxPex/Naq2UDuvJS
DH6FuIFWcsjvPSbiJnjO/H5IU6vrD/l9jKWredGq28F7SEd8GHYYrEWOqSe1elgDIR/lw7FRj2gU
EEQ2gycQuzuiprxhYrtSRY5rgJaGUVPodIHMY8FLZY9g05BoQGPEZ3hNqXcypGV4cI0gCd7oZ0c0
g4hMri/DffGTEdAEgalsMmlV2OlUZNcjme+d5jJoq9UDJ3bcDlOuyboajLA+P3IZ1N2v0qTi8/Bv
X4+VT6VgJZY+QVVOJ3Hmp+9GlU+mDkVdpPKhF+I0QxkmnAwfYFSJza4n6ZOsO89kKzGjoZGVvgce
0hbNjF0YciFaUY0gpoDU4bsXdHVWm09K+lRz4qW0Cw7Vo28rZwdzIPhdmEtDnqySmBSZ8+tFY1jx
wVIu45AantwvBkT6w0YPyzgtWeuumllLs1N1Dhov/hkLwFWd1MosQhlnp7a6ES7zq8xl64nTg4Y5
FtJHkB7QwwkzC1sRZWyAMvUP9xXjYqhZdQE3OQrO5+p+cbwtuSiT+V7HaoYbrSdONSB1iSdbIRO+
myeQ+YrpiIUIZo4BY22IRStbqGyFXVxneDNtadZI3bzV+Mrpex44D47FPvpBcPeknAK7M4GAdYFv
Xsj8IMjjldiP0ndwsEU1p9eLu7luMojcsXJWTMWg39bTBGC4F5q8ijUQgc33FpaJyk/ZLqQpQe2O
ckb7tmWX2PJCDypWkjCMMZL8JSJjWoZzz8KhNV9gjuFXkj1uKybLpiVfnWGEi4hQVd6qoS4/FHjr
kkFT+TNPl3QYEHAiRwNaEhpM77tpMBTow5jLyyyC64xVhnsKUsMSqfzcCOP20I+YbtIr0Dw6EsUw
vFUDek9iMkCGO2FR8gz8ArXJskQGUdReGDp4Esw7eKdZtRSMZ1xX0WM+cGba3QdTYJ/VebdUlH9z
hBTvOr1Zb9dtZI9BUprrRF+Rfqv9m/mr25fLltn79kzuEVQQbqL6blX8imXiiPyfShfciW5fdYZN
n2Clww0T/wmCaT2S8K4gsO01H1fd3QP2VKlDo+hHbPODQk3eLxswTDzRfvBXb2aJ0yvU9D5ZQzN0
4bO62C1LqRlXrBKaihu4lWu/AQkHcTYHyD8oEqDKTWJBiEy1dqlFSjhJf90wsVlzXHlOsrC0Oj8u
qAb/b3bxpyVUi/ay9c76+s7bvJPkoW40aLsS53eZNUC9vYLB+asUMmPoq/W1d5kEc0Ko7tLee8+b
S55YA3rkebKMFuo0ZAUoTPAUjbpDxezq1Uh5cJwUAbIKnBS1qXeAEICfuUhR5DW8ykBZ9dl5dsmn
ZXuEdE2swCtN5OVr3bNzJnQNNLsCoKgp+mYH21KJSyFnN9hwhpHWfO80w8IZK7W+eQf01zow5OUx
vRcfeXz7w1ptnSwZYOdaVE9AizidE6boucTWvWMgwlGcNyzntIBbxOxEsCvL8bmLHj+9BDruItxP
h1YcqHum9DF5Oun3PzONlBf04GTQLWw+iFIZW7XVtaD9RCQJ0TiQYnMTlzrYO/yd5TXmNnPrn83j
S3OupkQHgKWgqvWFKas2ITSkgNFMG2VOsnZGQ4de2eHfT5gsXygzaUCQd32VSa4AINR26HRiX/iY
tmctFyC3Zi7av/1xoDxXdSrebGnizupN5eYQwDlMQ33UzWoYHrb4n28PZesYppM2CbZM/sY+LmXa
EVNCSYcWVhGGaZ8l0Q7v/QzJ7Baw/W4blBhvqd6+Sg8S1Ijnmw+usw/MDrWd6+1sITsfl1sxESFw
TUEFpcsy40GwYlyPNtBYtYDKmJgd2A59IG4IBfW34v9HljdkcgPoNBd+1+obP/EafWU0/gXFEeJX
QoTlGDZLG9we5aDLVKJhKaOoBJil5qRA9NNDAjWIvDCY2cEmeoIyAdoVgangHa/cgbX41hSgY9cP
x4bYywux76bhB//4FbRkJsBKnBCW44XbkJIfIrAYUaIcLeRpICRDkDjsGbRg4AAjAzaGwCCQ2Q2+
CQU7oNdQeRj0wDIPqTS5lvOm1j+UB/nlHehJbyrz06oZUl4tyrtZylernjcyZZxAN31PQQsLnuQ2
NW+eoKUb2yq+fjSaViIWEOvZRi0doGvUXQFLKWG0SAKSxjj0BxqE6piLWXgKx+h+9V61PdtiMcVO
thZnq5zwkwaoTSdwvp2t2M0gxIHqhCxIQLQdamfhytcWWyuz5skznQJTaDA8qtUl+JxMpHstKHml
V0ObpTMZ3mmrfAOX3GUnAsJ25XP0Vf9NcdtutT/lTwOBJFBeXAWgUsc3nBOhdBhZlu5ojOSiGWz9
dOhFwedCC+y0yM9K0NeVzJcee9diADC8T+rNUEag3H6ti3jusLBmGQNknRIvxqvt85B1cheSdnRe
TGo2u6/Cja4AM9DOSdfI/En/sCzbb1HZ9twPqeF/opZ7h0diZD/hOTdrPQ9AyuFKDJhqHS7kVZvs
meiQ2eyuxahMWtJ1XXejVsbyk4Kem0DSCZwCJTLrVdjRQO7hwbIOQw92oUtesZ3XC8CfgiymYdJ1
eqqbhRuv1kzBbwT3IYR/eP2oc+zSoLz4FUgxc8Pl2CNIIz/qgTM+IivlDQR3HEqla4yN7SY8/hqR
IymK8VNE9YswmTFHDo51uRsZe35KT2cnddZ1DvpFPQgmIShGwVnkdvc1inicFIr++xqoXX+H7n3O
WkuDGEU+BINqQ/ZVoNfO8XpMLQhN1cK7Uce8xS6wVveM8RjGSW17onTsKfqxhl3xeZJOzva7xvu6
CijZ+Z429hwFsr7CZjSMcHPsNJVhfQMvV6jMY6iHb9ek87CBatckIXgGZRQLZOz50sGeJtjJHDD1
bG6ubD7C2wb6byM3hT67+4aiwT4m2KuN/XYXpk42qEVwm245JA6vH6m97jvimjZBHgEaAP8YRE7D
9ep59ARAr3yOkspGf3G2UJQN9ukus+Yix3exnP+zlCM8l9ToAih5/VRQmts1TxSG+blaqE7/JPKR
HmDtCfXnaNijPnjbvyB3Zyaqlli9ApZSC0W24MY87Ee0DLhq7lHlDsDOOcIqJzAJ+tq8x7X23yHB
xQ0ypbaKy0TfcxbwUAa6cJIIOqqTjpLa8U8VnUtZ2aEopA6PfLuIpqFlwpLqhXEPB9bHQ14SeANk
gotAknq6zLemF717CUtsmnO8abQKiX7qwrSxn5o4BhRrt6qg56Xn+zTbA+/rXUtfqBJZYIhGPls5
0l6Kaq4EmNUOyALE8NVK4zr0W/habvirq5WxRLdlmdQBr7jlEftDwIcvl9Vy0+DSR5CeiRRs0vMD
QNvQ56z0WJynjYhYLjtzhv1VcfoHta3LzCmufELsem9veywnoYxNiqp7ixK0CekPIbss9kAuOiaZ
drC1IJb5BFYtBFjcjMj906phEsVSRxR0D/A+UMwW58+FFntidTVAwat74oWRr2gnk21fUuLmkIfd
rz6ym/cBCZhLiXvMij7rAHe4p4zpjV1PCxaOMDW5t2xVRGGBJnueIHDQMop73/FugxCh0A7hwHp0
lW3M9gesmZdtAgZBKjVOgD/shQAAuP69a2SUy1eP9wDStKn/LQMHIcF8qiEGk8A1OBF4WPTZRwrI
whqzvMI08hUVI47SOl2NP9jYmiK0UF3K/EwjU8KMWzDYpxzp2VCdJTKgpqcONrS2cAMhq/gXcPBL
3sFmaDv45oOS8CXBF+FCngHVCk0W8Lv1FEmSi7KkhcH5FUkazzhS4Cy/K1b08JFmgqPGEtIYxPOm
I+H2nNPX2mPXuNo8J9HvD/YOrz3KX2q8unMos3Y5QE0+Uaa6YOD9xlS1xdpuAFXERjSCadJPmDoh
QU3AdrDMidSgLBifQjuHEreGR2sMFAHkVxzE6j9xLDPVZYHjKh2Mk96cnjPUy9gw9O3r1anHOlct
N1daYD5OuSoJ/qcIIaVhR7S74lVE+/BggHfMMf1he2f46/nF4dcS42pDs/PWIKp1Z7k83BNLf8tr
o7vUMDRFwN6myStjcydSwq+ozpq0OKkDemhh50qU76lctSSJINpoOcVmD5zaPk+eXcZ7VyeSDut6
3r+AgPiFyJr/PVAX2aiswaHT475kK3J2BeDvaCDK0AJtybaYaxGAzwCi/UQx507CnHkW89e9ym+H
SWIixDsQ0dWejadoe+gow7Q1vv/yxRn7YrlzAbgisRA+FDq2BoXV2mPtQNANZhaG3LyOksRlHSAf
S0csPAhKTyPH6xadfzBDmGyYxwPm202QHF0+lgjAQQfZO3llWCPO5MEjlAc50uCrofyQKI+vkSY2
zf9Cyqd8S60+0/Xb27HklvFzYF1tRRPZZcFHheV9Rd2z4TCwJynxh/QLoyFfS+y2r1MdyKDt+0nw
gDdCKgiVc+us7B7yUo4twbwDJ7M3U/WotHc1HdBrpDAkrzTH8mqiemXFv/Ym0XeNADX5R7KX+YDZ
ow7JxBU6pMxHg7OjjFX6TC4XTwTpXviwLcEZJbzwLXv3nVybScB4jjtpAiBGPfAKpCBgbnZdrxur
8Z/0fG9mO1m8SrtuHiBCG9HFPdgpB5zWaa3fSD+q1y7rUyUzSrM3mX2GxM9C1Mb8WOsE+obJ4pQs
Flj0xXORiBITS/W1fXB/nBVYwGUsF28tNSQPb2KnDECuut2s5u6MD/9zvgGzaAHuyksiuyFVk079
x/X5UdJv45v8S+kkWPzla9hAylC61ZIARZTXxUN+zPa0wwPZRvQr9fftBTfK24COv28ecsjVAOsd
bKI0PTnbgF0EdEZ7ZYIw5XwK2VSpa6076dTB/svV0efAl4sbh2PBZ4A3nVIi1Apt9dJyiPTxkxrY
LSgvBJ+BJGu5aFcFg4hqVVdfT1zo4PurfKGb94Gv5FFp00t17gQDdSt1mIqoRDffTfTrarrkukEy
dafZQsuLxMt7dxfn+y7B6lDJUhR21Iw2QL8Tf2x1gdAkdlgUaaiw+ItkZQXcSsMvmylM8iGEQM9e
ZCalxxpL49BFXio/0oW+XNjk+hjmt0rSq2P64Yp9MXLTDoABsT2B4sYyVbPk+nF3MWV6lPgmtuUA
g3DgIxgYrW2Tz9uBL+zLTYC2vPdAheeJCb9YGc3zQtQGNOmlZ5WjwgOdVWrEJb+SwrjTZKjYvXMY
3UrwgqiYaPYEs7UjG4aCsvzsRYUSUUWr3FXOkhnrLjtf8gVy3e4V8zg7yojA96BDmbeh05LXqDPq
xAFzNgEz+uGBOLx8R4NmmKy/tanf1VogrQjCjeE6/R3VxnZvX6vZUqD7f87Y9t3rfRa6Wf3CPFor
sQhtioox8ie736nMg/nYqoNrN8YeXExFns/fCrzHjU7a/kIHQgwvg+72cFOvzrN7WXDJ5PCsydvG
4impm/STElznWDG+AXklVs6lnXliY/rEDZflFimjPL3vt8Kh2pMwLd0NEDaq4yvviA1aUKONfw1f
MwMhxmvWb5OWyzPNJoL9TZWe3tWysQkYqyhD8THlmg/ISYnSr/ohJfB/uE0QIF2dIJhfUsN0Ntxr
3HrFhZ4poHDg4Ejh6QsyuZ8m+EyTj/WX6spBTF1UC30ky/71tRANLFLQRxbE5IpoYCBjCOmTWZ0g
qlLb/I3M2yOCYdF3bKlKFYg5PW2nWSe3GA8CiNhwSszLJCPOyKcUdMIlLL7TBU1pn3HPGm2KVk/9
MIaK/4llVH6wxzsfWbb6zWPEiVZThnyM3XKlqUnZXwpTphBhZ5yQhWPNR4GsgMZexIlyc4dMhrW7
/Iwnw2umNSLiujgvwXGYoAkl/9bqz45wdFsAavkmdwBoW16p0T6aO29Zs314kdlRK0WpCziEY2e5
OeEMzN2x6vjjzZpqP8jx/7OyXfCH6xc8UiwJmyNK9LXVRXOqxhc3RtO0esAz3uSyhRjrtHG5/sw2
F/aflLnju2E4DeGnA8d/o3d04RyIE6RPJeuM6mqD4VyTdcQUinMzLnPMV/KKCq+EDJlicMAMBt+p
t7JFB5si3WW80FQFlWlbgZjRIitbgP6FlbquFeUPtR731PyFqQr92+0hJzBtaaHyKr1UnEYNW3z5
7sQOlt3nTngt/Nt3EUMvvLEIEPo8FVR8KLLV3coIOu4bxi3gYhN7Fay6xqLFb2/01xg7CvqmsJom
59q91X4MnGBxcJuo4KFi2zEOxkdmdqfUj0T9bAf6DUhf7uq1NisMux14bJC0MrI+k/tZbRF2YpiW
fE0tC2zqOc3x8dIwBGuZyCXCD6h9Apy7XTcCrvPAGVTqp+TSlE+sYk5yRWfG9SghgnqDfs2tr0N4
eLfMjBIO9WJ8BKihgYfWxs5tMPLoECal9wg2sOGgwLjyUgjs2wDKP0v0YiWrPdbnXLkix9kKkIAP
qrNiJW2wY3jQ6Ewe7+xS5R9xtYyw/vaFEbI1nUKDyB7RqrjtkLU6Sp2P8GdFVtOQXIFp0I7zkzgC
WJIKbYL64D+HSxXepK7FY/QOILzZIMBI0uqYqIgNtDY/zuB5flEaod0TIX8sVVCL/9u3saEIzZef
AGrUDt0P5eFEs0Tl7Q6uCpGfNWcGXjjp2esLk7UeB+gU9AqM86MWjwYvJDD/vU3hlFzuOX0lwsh1
RED8P4T3hfb2bjs8g6fmr0YEVluWYdau/tFDqcfIvqO/ADqmk3Jm5RmDQtqu46TjkoeGKhdXnBmm
KoU2NGXHQYbkelQnKqFMn5rADh+++KHFg17lKRyrIXRajH3Y/l4DVM0ZxhYzx5jY15ZJT4X2OHy+
/GmZ+Vuw3TVXGQfsj4MaPY2cExm5Lj2KJfUToUjPeXGSOH+JQOp0Cwou9iq6MbCn9yq5RZbFvIxH
tGwP9jD1l2zP2rVIXPcDaIohqZXZ73nUQdQkGEEJ0/Ul26WRhc9wKLNHniOi4quI294TRdC0OGLy
HSLcBAvK2/y3j0rUbH11lNbuQkXv7O2cwib53nGXGu6TBdBb3g4ofl2Uc3oTSioxIx0P3CKLnXcB
0kLOIKIT9S3R1fxNQIxcGXLTWaZl6kSXAYO5sCh7TPJ8Jy1MExK9bMfoC/H7bhiiPU7rm6SJw5ar
kMQFwmrhyjb+iB3kjLXQo6B/XvBeyxLu3sXoOn9rVGHke7H8CBH6FdCc2sofztuz/iLvIBipKwCV
bVoXf30+yGBnoIJyxhCRMyZKVk5aE65uk4HZkcEd7P4XyS8tqksX2jiXh5gsjSWYAqQCn+7QGVX/
NqK1jPltE9g9bPLRBPfoQs9Zwz6Ue0y5bn1VPWexEaIsOSnLckK1PtfyUeYoouP2A7begv6vwB4R
Gz8sf98O2rTyfd/pRXhCI0NzmqjDmd/eQffc5fH/u/RvCkXoX5AdzUVgfOmxIBuFeTrdjk/Svi2A
2Xe42FPo5pt0mfgDExXfXBLiOg81fPcw8oxoYkFJezjM0V/6RDGNuDe+meqTKwSbY4xQC7ie8Tev
NVzm+Iv57hbo702xnGEyngG0dzUm5ho4t60EjdK1FjCpPZooxYErAEM/r1GM8W8Zr8RMLLfcqOwc
VtVR5aCOTKlMOq7O37+wZ2LzX5tr0Ql1PLiVetWPP6HjXxbfpssgvMSLvUMW8Pg8krMtYzKwv0tp
BmI/Zf2jWWuW9y88pjanhdGPJ1mjgultK/ipbhxx2x6pRSvPdylo3rNhLNrlW2q1O1aiNU7oOJvn
y6sz0XkyB+K4jEoj9oOFw+HpN4sx3SRLYci3p9q2qeqp6Iuw+uoAX16ade6JN457f376ewuUdw7s
wq1658axAOfcwroew6tVivdgj+yO0aLg7hXFnCcRdk4tAbM8S7TXChCVLJqqw+SShN79pDnKKY41
+rzizdeGAXR6idlCEMOTtonmenkpsWa9PJFWlzilhZ9iIuWYDQpRKqqiqxnalYFKDWJTdTPftUMi
vrpWEyHiHXnbOij1ajPpTxlb0BNvGsstUyoM4imuuHnOeKrnw3abSLiH2Yc8JCzwbXlPC/T0pTfr
/E9aFbbWMz6CPZ9Zk76Ni9n+qOPLv7V7K3fV14v/GZgxv0mV6mxSa+PnHiJrjEAzu49LD8Q90KM9
qT8ncp3byRIOEiIjwfH7/KgIXjZNtsg4aeqLTT+xBie2Q6ydET/1rmfv7V/zYwC9NBCiliXcyV9k
FZRn1Rj7Ni83D2ZByiG1jZSH3dqgCBpyVJNoKBdaerRBiKVb7HRc9Ya7rLPjCQX2D2yrFPvzwNmp
NMZPRmnOTooQ6rbAwYdnfX+34BzpFPcXcWf1Ubx1angsIh0fvDkO/5H+3cmuDsJT1fRfb7eUigOM
sHyGW59XC3cDsGj50rxh6K7vbzkyVTssVHXALeUhxqTuYYluMLP6GY6Wh0xCr2VorFtQoKFMj6pP
GNGR/hMdC5GUzKlyT1RTXNaOMCpY7SyeTs/arLhivCWFMfX62bFFRFbLBetR9yThd/tr/z0rbUFR
2/W/VJeAHdS3YpTgAdeqsQnPSiAtN//0bSN38NhRChocrZfOitUDmfkOpz56Gsj0EQ/EMaZxLDSy
n92F9acQg4Z03MRGgJ37/FQK0gm2z53EYUbovbHXDbvxIn1Qxye9iIilXsIAbjMjTEz61nG05UUM
R0j1bj7TZMZbmZI2jBc6J+m355aG5Nwrqry/zzr3aTPbsi6i/BWiFMPB2bAaUbwmWpuHlouqxzzb
7cK2ddbVJu1uQLRKOn50fjgL6JYwY7yB+HEYanFOpUodSwQzbRsA46OtRKAmIFtGvt3R3tjsJPnD
BZZ6NMQhLEP22zhTGWDbyR1MTmI00MDB0YknXoWotGFIOuh2wFO4aHzUpU/8ip571rrzBhGy33Sy
RgcOvYu30F1QlRx1uuTeLwKblnDIuNpWd/uTmx91DhYwqmCifcW9O98v+M8aG0nJGcx/QSq9J3NT
m767sUoDBTaMYK99W8qqgsl8gSKwESPODdb92X7mNQleEszt/gUV5ksoS3jq40ZiUKNI8IlqMnLR
R0bTd7VvQB1RPfkn9YHRLgNz4dX/B309IRacRZCxmTU/5351w+tm26Ihp93UAw/SdbbLxT+ANY++
OjVZuPCDsLvCVSfd9u1eeU9q3XFZIZKOxFrXv3WeFGQRuERvuQ+b8H3EPNiD40gX3IrLwmw95zC3
jK/yEZ64Yy7+OAmS0gFOFNGQr/uTzYnweF3uZ6YaF6PqLFCb0/52yTOFDPZdzUlv6hhKzI5l6AJi
2kIejzaK4ctoiK7twXNTU2aQhh/N58L2+Pfac3Wrt3uRqTwh4Mr/yFN4ae+SfMN2zO6z9k96akmh
2aXPIVjPYhO1k2pPql/ClLqj4rMaGShyExiLZIY0ATHAB5v5151c6xhogeTsmOnd+60A1lwHDqRY
RV7qxWxgn/c3kAnBfLSdgyHHEuauuijl+VEuyTB0Tfl4xaHcvAenPXDaLtQv4B/q2izRymuGjb18
kphhhNKeK8xpvzd17XV/FETYQiplIpsWM2kYsj7YvBBZnxsFSgoSc+/Jq+doxpVT1Sti74Pz62gw
ZHDd0xqkou63R/oXS9QYSoAR9pp9Ncf3VLtbyrraLAgkbSyUt0svzpnMiCmmZtG/cMzOV9gsBfpk
9AbE+ky36O/ed+liLzn1GA1YWy996HJnk66TKbE+HUU3KW6mNuyn04UwHcQ1h2PT5lj9BeN14PLb
EZP+hp+PItJgBfTVRr9gDJ8J3gFOTgtu7zhUe6UsTQR+nv7WZbWb5tkArV+IitbDa1Pp4hBefv4h
xPP+X3VkV6c0fkZXqVcJDtXAoZ5n6do13Dj88nRQbAZldrLixIk//uUl2CUK7ZdvDRWuB9POl1HR
Xp0Ro4DffuVKJSr5oE3Zp5Zca8s/moBA9mUEIRWkvFTubfxY1Yq1ztVAtkK9kq/RdTg8e2JPm4iW
3w5TseXCmX0lkN29SOUdyIcc5KwGnJpCWCuZEGAjkgQXFXbxetJTtSiVsIi8boaS67slBILBYSD5
e/NknZsSWpDULvtgkIwF4N2V9EIzDB5NXe/gJfXDSvfr0Y2ptdtFSb0TsT4QirKB50geUYRs2MV9
WRXoZ3C2wcDuQgTXXsq2Omjl8Jp/yA6kM/poHsw2gfUAunSQ3yQKN3wQIsx2JC8Xszv9nnFU5X+j
OuKFlLL0Utr8gM1p4t5SuOC/2T4TVYrKQezXK3CrnP8g7QRRAH4lowO+eK+50HFd4gFk237vqtTc
R0cll2BFHENCwWqP+xKzpXmuFqA/NbCxK/lWNOWgvS0SMHS9ThsvZ6EPdrOekPkiAp6VkY6HvZF0
q/xT+rftI6yVj+HQkGxtXJa8mChtHJE2VtKueiHIXU8KpXmZhp7R+Rc8xJbX3XPAbXvaINUGLg+A
+gwVbyI/64Sk2ESMuYzf6ArXzHUGFjcIgS863DjqWCGf95BzdntkBaGCtHYV45YDSM0P+2iNMnmH
BpieR9oMpher/P/tf+tasQ3lE1Sp40pwi+rCo6GkS79YwyHncd9B2z6zLV8ZXQ8Si5WizmNgqL/Y
pnc4RdgUDBYjBwjmJmmFwNMdTEs0GjHTn2BfwLPRlhoNOOkS1xfSsHRyTjsMSCg1DpxFu5Wh6E/2
UdoyKmo+Uwb8euoEZvAU2d2qfekS7FXJEhpmSlpGqkBg3wkiOoxazopsEdrf+Mi6MvR3TL55PEn8
lRzcSbGCWbE7U0OgHvGIP7h3L+z5ilzoqx6L04TsTk6vmUS9YEhz8oTuuV0BWemOqTkxRpnIPvt6
f9l6Bj9SNko/ZJ1UNsB59qF8hnahBXcme55ktUIWgymc5nrnomMQ9SxiJRAucFMQiEIRgydkx3Rl
TFZe0fOxXaFA25dWVFK5aXXa4NFNKvNFfMMfzK6kCGAxba50K08FQlw/HTWHt3VrI4gL0FOevgWl
j9wm6CvcZ9KS2qHhFhsYBJzpkadMUogMXCuwOvDPg53xyI9EN2cw7Ae3t9k06Q6isLGwUFP7Kzmd
sBsCJJnA5oF1tJJQ9KOpowrXJ2Z/V1Io/SbwCVcHpwh05Y43/vGvnwyTBqTmqQrs9SIIsaXcKOAf
ILe1+q/JcwHnF3w8K9qX/tatd7dWvQcBIGXob1WOzt9/sBZwOq0VWa5/b7Lvz5fqO9iCiPEpbKRS
ej1QwpROZRWDxwP2GFkNSbawYkjCK++1wO5S+hfYTYXOLD1D1VqUq4XEHMDFCCqSKlSc6wfAbQQm
DIPdDT0SD35/qJ0dRcGzXyG25E1Ny7cV2kU7QUZQB9D8/wU3tHqcXtvLZuHUe7n/QLtow1Bu8Gey
BazMT7VCUVF7F4XfVrtI3Td50t0C5YjYxs1dO6OGTJ/J4HHBbxptMcy7/6QWkaGmXoVJnod6PVOs
FIeqs9iBM8MFjZOM+/U+EE8ciOtAaI13s2jrFc89mWBJHWlT7IVg6UO8V2WDnud+Fa5KczyDsQP3
2SB2+XIVHoVDZMFf6o5DytI2XPQYC5r9LhAqHJu9GIG0KEi5XkNFMNOjtnqf5qXLN3coXM3cXB3x
ieydUqTq83ws0uAN0qfYYuYn8IR60RThE6RhdM1h7kAm2TWhr1bWSp3/2q708N9mdTIu06bzjvZF
TGM2ekT6TeEPI8zE+LEtdivtA0Fn0Z4uYq9nyqxfAjfFLl98VKGroGcXHTAFMdY12WcMPXIEPmTt
zNlE/L3m0UKwFcq3SwA7ldFvfIoCImqWQdGAY0StOwu5+2Qd04R5xG+JAfSNH9I4JVxX/817Dr3n
eG2QRex4FBesZhGti5xcumGAEVtTk9f1P6U9nTnoF70NxTrsLEBwWMC6i/MkhvEzXDprFhzQznbF
G+rrJG6dl0QGW7YAh5zk+b2htjsEvHxHDImF+APh0lSS+3LdfD6H/Fu9xd/iwkZzJo/oVSJZUPBp
9QN+tWhL4X2wBRtcKjSAhNsZgT0ee8DrFWxTqme+/9i01xDvFbApB1Aer8gyl8rkH5gNWoHqAp0x
wa18t7KUQOx6HHVbn2/sIHrixOIufDcOKO70QBRH/hzd9fEYHBbBkDoL6PSUfCb8hkpdzvzA9wbg
QbDsUASFd/cbjiBezEy+CkjpP6ghNfiS8ygUCfc456wNoJJ52ESHL7xFq84Tg4ov1LWgrdvDD/Z/
yglLORCCJxqQqjyNF8dLxQAT3wmpjzs1xoLxQBqPN28hbWe9c34MGGFySpUdpCNprRXW+ql8z2SA
nW9eI5+Hulb7SxVUp6D3rGvo4JuOR6yiXfp/UFBt44Pm4pg4nPpKBh+9MeDOLOUJkTBdUm66rVdz
Cl2ecOsK8FnifBPOjrf9IvUMEQWNVcQ2Tpoi86PMTHoJkgmrLrct3ByaGvmU1BddgUaWpa8t8SuD
bf7Zyw+e3RRTceRyPFNae6BxHeXi302clGTjw1zP1n7o4HJWV+9nxO2V9TZigAhPWJhsG3E8Hp+Q
Nl/a+qmEOD+VGi+thMeyhwXzps9ukiLodqh6CESQP1SawKoDzXvge90uEdTPQBfROK/HJQyjisGS
Yk6nBFIRupcZwPc9+WVnAjFmVdbT/zZ5uMisS0uYNJKnm7s5HNM7R+FrVwnR3cJ7pWgbXks+9WJA
g+qCUZQUgnciFt0N3Bl1cGvwnO723B8XR7rqdz9uZANWCvRYyw9dB4De9HulZFRXx3pAJIPtoeMt
wtP2SGpeaqJ8GyVTSNpc2HeRQoG3Yv0Hsc+OOrJqNUTq6d8UvVC3Mr3dCD/PqIGXgCwhUcI68dHy
kWIJtPojyiqpiravKRV+SrIlLn8ngNwmLQHOt79EtbH0ICev+BfGw7jQNWbmsAOcAtUsTC5D+0hD
Oo90VoN7h1qqPSoVNRrMmb+00VovPrKeN1kigw0k0Eg7L6xiQi80R+Q9tON5w2Ep7e2PuSd2r7ES
EDucoXdujgkF9X39I7Sl9OOoF9ZIusrnxJkUpO8f/V5pp8KGkdW2f8oxx5ft1M4poCtgYskOYOIj
sVyOsO6xcN5P2eM6D43Jrj2B5rWirkwbPMnw5KeeujSm5VJBBEM/fZbMpHHg/0YRXKQsWLLl0lKe
gAhlLNTit6KXKtnHngYow5fJF58jSA/TTHagMCzMFBOCO0i2VD8WJzj3DJoHcKvvBCrhiOaZ4zRB
IzrWEKsWpVwgSWRKM9yIZahIysMlnbTN4rw1wyGJ1xB5TBnwtTb6zFPipR5pu2AKtA00ke1C4I4l
igQizJbZTNyTzynNj8vOmIjCiEghS/QlB2P7ArSnIbW6wkbmBidPZQumgWvi4VneqN00jycqk58w
7CYCwWn3yCw7tJ+QkoexB5vzvCNAQegF4dSXvA1PoUa21VmMh30MU0E4QiBh4y/eRa02SKsF3PM7
5ODw6J7VE1HRAmz9jwS1TrBuHFsHt/jxZKnXse/3VyHdsgT+nrHEyIBivLMID3ku6SCV+l3pKJxu
cSoVuIoYeLe7Y6ET4lXt/EIqBXN2BrRL8ovKVuLp1CBO8F2G65/aBEY6Wc0tNfTwQAZ7sVbpoAyw
7fjRRCIMgNQiG6ZRP6/Zav/ErN813zaUXHaS4Ptl7+IUNO4zA8KHh4eawKiQmYOBD7v8hkZliijp
fbCn7NGIplN5Aqd2fget3Z3oT+YTQWWabCa2pPbN7DX9kQXnqfJ1MoHmrR3dvC2zD4SsK4qGrBRh
Z4suJwZxCro2X51birtx/6yyMsgvXNb3nCKJ8YAgJyMol76z+rMC8eOVJsJ1JlvM5ibHkl7c2xcd
+s6OmfFjjDqaj/fRTOj+TXn/DpKi9gC+x/l0JiOOnJFp4xFebcgM+0K3vDtGsaPld3K+bj2wuk/0
emKbqQLWVcUx/P1evgOpB6CSQtj6Z9W6e7CoLesdue1fbVyrvJtBpqYlIjRirGTbjH02/pYRluGH
WwgVb3/A4IXwtXWxnvgMn7tro7xxG+oH1eZEOsvZ/XyUiYrOFjVRk39yoYELo+XlG0uQTApo2T6/
V1AvC9+g8hGIanla9/FcxR8Wf8fgRTxspkZEYqkx/q30vyyUURKMhOUyW01zdTnLIHQZ3AenVUVA
p2CWLVayIq2R2xeBJHq9HvA3QeTpgNnMqOKxlC8GE5SB2XvV7vuGe55fuT5LHPN6KPQ+Y6mjxtlw
qPOCLtVg2UOW7bFq5v87Nyr7PW+GxpH6rojEHaMAMw+6/J3P04jEOa0VGAehV4UwON46SQC7u17Y
4m/WWvS6nrsEPa4qw/5gMWvmAV2kUkyVP8oSwEMAvIs8q+x2sIybQkOnomfmDsgDjf0tIOpkoi8W
c5ID/nc7CQOZSbVzv3aDo/aKQqfZtSEMyyN4oBVy+/jr1aFFf/gI3B20qDkYSSJrnJMFybYfr3xh
qH/nBvF2LFlzy+Gcw+dMUOeuMBzFvI3MPj34tGoLMmTiqBSFQ1KFUfjo5/nRqQp9KLLSIuvaRUk7
SORjpF8VAY5ZukzklVjVaJ6J6o3eWkSPyf6OdXSD5iVKjhgyjM0mgtOB5Jp/WovFoZ1J56Lz+Hqu
0Qgvb10pTXAYQRQZ/p+Hp0UAl9WcXHlH5LWi+2eFZA+OCd6+SKJM7m0m7lGMcoHxjkqtUR7bsKYl
aVZzObBZZWjeaAg/RhvnLbhoxMCkywPmk3v0OypcZM/X2PJX9MS8MYPORyWZ1KumSyEA/5l+xOn0
nNKE6Zmf+v7nfp3aMXUGinmGMgfksBZtvjmpyY3GSXE+SY5s8oWZrhgn6gU9TLk0wOVlK7wzR69R
MO+j0EV8K6QAiXTP4WwXXOOOlefEzPL2rWJffrDY0GOknao0kYS6cSYIch86xamLKNEeyNHG1+Dx
RtrY+ZKO9SGNh7aatzSUXJ0L9eHrloLjSYaAENotf8x7yfDwMx92KQin99GOH1wGR92bBlDAbCrq
HK9cuAKCdqMk1QsyEtj0obxskbaGJYzfABDO66oxR/Dgr0Qlh7Zov9Caso+FlQ3Nvq0ygOk/cuNB
y6hgpj1EY42KiHcUR1ZWr4/XeWwuERn/JoQpMeBMzntOV/YAoomRmjssdqgqJgYgB5HaG6fBRD/7
eMsNw5cz4aZaf7ZdqyYBBqBXbQueIKmq0iIugt7Ejh3hjwlUwx75C+WYP/+y4Zcxy02FD8GVd1fG
dssYuHJtVv/mL/eCvrBn30CXVZjhEjv8onpL+9RhkCNiOlnTbIKoEgfvE2hf1I3k4K4DVtkevbHW
ur41EA+Jy48MG+mlCOQBPkBZkOvs50LPklAbzL2vD3Eb9Noy8Twy8y90UcsTSPNDR4IbqsvaHZa3
MIyb1xmbfmyka4tLF9d9OLON58r3uSM8SJPGnjBVhpYRtrB3t4JpZjwQ5ZWLoeCR/siI00cj3SOQ
noraRn002AJ4fc5Vz1DzAvU2I4lXrwj8oOsiilBkEjxVe9/NZd/GNgLICpuxU6iPNU/ESI7nA6em
9q+92KxUSxj+DMWdOXJ9EY2C0cpdNWjU/btHhE3aZgW2rlnZOIUO14XMPqKL+wRm+D5QhDG3yA1r
0AwVTWIar/lY3WXU/d0YZ4UOZxyozeRIsR9zJjQztEKVL+nvf7TnXvc9+8xWhR5xBsxlQ/0uP7Bi
zfPZtR/3rQ9zjr177gEF5Z1UDzPtVW6+dg1fB8ienGrCtSWV4ZMqjsgxiAaW2QrMPFC1XVyTd+l0
CexDXOfj+xvT46Zj3VLzjTc1KKRoFj10HL1uF3kxdd80uNnljI2tb21bgJ3XvZBgGfPIdzu/NF3K
ML9fB4nuCCFZOi8j81bvgRh6I2alRzl9FlLCB7o63v7Jc6siwFHy6C50HV8fT0gmCZe3l+hMxD+H
vDJ4EvBZL20qRFp+Q1LUJlCQCY4JS0EH8sWf5RHMLus+mDTKh4z53Kmf+tBxC0XrmLYVExXScPG/
R/yetykuOMw2xMPKaf/TQpTrTtP2dCQYEc0Sw85l0borKoPrxkh1iqRxYbNNv173a+QCpJfsF4Bm
OO1HHlxQ52Xl+4bunOjpCICjxPvs7hWKL+oOC5s/uomA+3pcUAKtZQrhx0kymSZPhCvVBHuEqk9J
bzMevNKsR4pMWIVbl4zasyEUVj8oaxB06GHPicVQzS2j+lZD0DizJjmNYnXNoK3G0QH9tcqIpQ0u
gzLtxfBBI1F7R6eUA//iyuUSWiaBkaNbkxnls63r4/8jiH9Pw56jOaS6YUgSukF0Zk/Q3Lbqw/j0
xtUTEIlL5mAwKUzb8TzJ9jr+QRUhX/sTAG3B3h1cbtBRJGfmXk/wQ8Ih5u4pzBzuAVarWtmQoK6Z
K78gpNcmrThGn9WSPqfB+6gP87ahCWVoHmD5RPh3u8bXawhaRpsFv1HC2mGRJTjDn2rKHpx2ryHj
EUEQBl9AqE9CYBvyHyM6FwttiTiRRssyAeEABa7uNUUc3ULYidnVLuYAkDM2Q/ilgJ2WQeN+sg9f
sH64F+AfFowLWHzYbruHCel50SiyV7NZT7Dza8SC2wZxzqBYl2fM5GcANHmOlFR4HrU8xgJ7+fyx
n41dx1n9SuHNN18TJc/vE/zG7Pfdr+u6vZirlWDU6rqcsTcqCI0gUQp5Fe/ROz5lFG6sWx0ZmEku
PI3pJTNRaL02p1a9BFdCwnLFvslKjHVxQAeM2tpRyY1j8V/kTYwh4zJuwgk6SVzoi8SKNqpv97rc
UeX36oZOep0GPfiHXgTDKz6fwo3kOsP4SaZ4n6uZuFs99mmquF6tc3oUqsFYw5WSLRVZNPZfeJ/e
B/unfJZSLBh9UPZnYTcBtC8A/Kne8isBRhX+OHq8ShxSMuAYju1SmTeGDhXb9u14Px4R69FBl41G
L6jI+k4tDwAjHLnSJ9ZZKeMsldA444WSafFDpz52SHl5GiLSuPI39rJ/MDStQspE0csbrf8sDK2c
Gz5Maemqu5P2JWGIJvkfkosQ8B9w0dGKhKTWJSl10AnyQsWVW1IylQESlLobwXPKCyBJoxvtSwFD
5yyKONucvVn2NvlmxsXi4bIMP4Zx9GOYmAeGCoNHOVi9ipd7pTAyuOnzVl40ZQrZ8LZJV3YBsd22
E0BuVWISbl4vZ5hp4fzslwGqX6kyn7kIdpqWAv9Hvchumory14UuRsqfUIj0VDF77DXAUqg2gKVg
cdKmV1Gd2SB/Wh/XWw9Mf0Q+1SL1y+Qk9fY0NhYtcdkfWS270fFz8L9vdq6BSP8n2oUEUooMbMZW
XEQ8PycsQZ2nEtPBrbtdPnr80tHCfz4m0KHK6HUfGAfV9RzfXC+3M/0mjLc6/Q/cDDk8eXyOcD+j
3ILeb0YRaw6AtxFygUf4Qe7n7EAq+osJPNYy54bAVmiaq2p12Hfg9Yt8zLFGLKlGYVIZ1WrDR4DF
bl5qzRmgLmD4InKIhMKehW132bQEtzDO8vhAgwlC5B9oLTbqBtd8Y7CbB7xtkbdmZqPK8Ax6Qkqe
9cytgztgqAWkeOLeYnQv5b8XFglNvHiHQ6Jirn7rbq9pSJcfACvqDuQwYNaH2xpDZGi3Z0cd0Oiz
GGSiQK7Y+6KsFLp2cHdXpa3TLuC2ratvJX3WkKGhpBKB+mYkQlkB0qpgqb8RPe5btYORMK5uE+L9
pSNguyAkxcnjg4YJ83B71Pata/VQ3N+CwyxMZsSZvLE/wtZ4IgOv4CcXOKu0wQ+aiiF5YXkVRMz9
qehm4jjqc1hfwwIpct9zL0dTQ0VnqS0TYnN/v4KnmEyfBO1lQm3vj8lu/bE67tf2NH1EV5YZI+KV
GWcL60GvDzad5wt003dy9sa7PtQRKKFfhVzoCdpw9r7cqIOxQPS93fKCugumKvHn85h19fIUa30y
KXnBSwJAe9kkE5nGySOZYSPmW8AEPqO1AfD5eZ7gmn06qT16sTjG4WFToWH3oU+QQX3n37Mu0D75
xWzH+G94OIcNvgj85uYYFQcxL8TdZP8y+y35AHCjVWXbD4PfhKxcHxASYZIe6op4IFA5aWtAiYEe
p6FGoGs4W3YCpJAk7vNeJqo3alaa4Km5B6wCiUeeobQTgiviwzgpeUaJDcMFcBkrjxTa6SieKPCg
NpdUNPZQlC5Lh9hENGdnWZskQXmdk+RPt24LdnpZ4ZGS7sbv4cla5F0nADoxEQd30Ei23Cdrc7m3
g8GWElJmAQa94Ybngku626S0qpdBlJnSoDrkSX2jxzNTt2aH8qQpyWdCCb6GEldg+t6qI9QFxBZb
FThoS34vDM0CzoA2CHos3h0qZ5pY10OZ1/AGohWkM1oyWcNkIMW3IvgSk3haF1wepksAijhfHqCN
82r2SCtXOR74lVmaVRNrIh1E827++WN85jwb1qO06dKW3iofWHyzNrD/ZtY361t5/sPzjFQmvsJt
0lD6IdwHWofkT2fLITSyXr5DUZ1nYRh/5jx/UqKU5CuaBbS9kyW6ixxri7OqxKoC4Z2fzD5e9CMP
qFmNKKghkztYKapWzMG9Py9m586fFXEB5ENRHkQs1+ZwF+yqSR317kqvk3gk5H9squQtnp+RrXBB
t0c0vO+JsFPHO9P6wywcwwQBgW2chjGXYX+sL67gfsar4CaL+N1yeXE6NG4O/kmnDf8gvmroCLaq
4j93scYmhZliVLITuPhDu/0T3V1YIvgjJ1R1hvyvkAMdN2Kx0Bu47WlajTLY5mR5OfPLu/q+vp+D
l7rauTi9vEthaG7D+siaUio92tp9t6tqmv0Ri5qaoJgns4yBA9wJ5UPR95ewbqjL3x1Lp3BTkCX4
Pza9f+qs3FxJsYXIfWK2OBmcAvdI94YPi+VdJkg8jvDK+K5+sViYQaEZ4WuItSLgVC8Yth8wQ6Kh
OJHc174IXMTcw/Ab0RwHJ3pZbHfZ1YkbO+e1S6vnqKuHY6vJb6qMF7kTYcoSIfrtsesOfVnPFu7L
GbmC1FgHo45rN2jqChJsB3W7+huY0+GmvR7fJCTCLFa2znrLF5pst0UZuRtsTsSjgaWtMK72AUX+
Q3I4vtP0uSMVG8Vu17ewQ5CvFZmuMckqZTRjaI/TW52akbMaPw+Zk+oIjxdm/wFlg0pygRyNYLz5
2P2Ypa2i07vxP8woUxZCLb/ZG2pveFxj67Exnx67TXNuE+c4mH4AUCr49SrxIGBlefuuzLQ8ULyY
P88jmG763XDpilFAQAv7nNiXzL+rgEhwJSJbArpfyVO6f+p9zYPzmBh6yqidGRBgm2OAX+Phs7ta
yd+YgYwl2wm2BQUIXmwCfqDqyYKYx7661Fr2eReJQb28F4iR0jrlaagbKV9MSwiasqccxTFATJhX
En3Bpj8mf2uu3KRIYZao2u2WXVVdR0HF3ax4pTg2afs170yHxe0odVTX4Vi+Mf8Yv7xR/VHZZBzp
p6jpoZgexUK/fnrvCZbQGtFncFN822+9qIIz52XrHRGc7YBkQPUgBNGujGL09XVBPiVoC13W4Gzl
A6vbplqc1Wta4utatvmoFtBEFnQfqQ9L0GoOm34hXZh0L85MxC/3ffdBLUtrM76xc5gqb3wmsuP/
81OaOCwWAgqJtO9F6/UtW6PUnvaudt5ZuBhfquJTeeE8IpFONK/pNMiufcsSC+4t+d2dhCoqkp5L
FURQOtMSnsaL4MoU7gn7wm5TN++Ku8mZjy1zPpudhXpChBRm6bFEelBlBlqFJtauEFaPQUYHhujz
SCjIwI0PvshXGl2MbnNJnYU6Za+gaI8tYptI5dup56SzKYdoG07ZJbE55DY/PPCKqV4Bsdbg1Cy7
fXZRHMFF5Q5K5DIxnckik/QqOEaBqwvrxEXfCqWgEKgy1UlEuR5HbGT7JLQfcPrbRlzTYQcw8fvM
mGPvtCMIIqapAi4HIswRIHYVKYYi8BbBz+BPHloc+0QAFEXnkBknrjZaonX7mO3kDwgVMzyygWI3
1ycKCuW8+Ka9K922PGAyrJIhzQZpJoct4MOuRXEj1j9svcSJQnWXViqa7Ih4vmuAWxE6awDbrbzA
vsLXqHJPnKcvodPy9dz51pYPQ2tN93uD+G2Z9baesXuOsBA7OP+8OIbM/oXmwh7w5hmtqnMIwZ25
IpkuzZOQn6OfoI0v+sjEgracT7YihSstLFMFNO3WUqimN6UWEUr1HXelPm+kfYhPx/sOmgIgdxrZ
OWAkm+CHmhWY4JdUxj7QivzBhbn82T8SZpYDRGVqkR1D43NX19axpj7WRSs0p/dPaCV+VVq1hvRx
k0dBZHOBT9zdl5epmt++WAlJLudRvULn/JXmBiOAp3jjQIVhQiB34hYOtLtlA/ePbFQBu5sbmwed
V67y71S6DWx+5WdXh25fKIDLWCcXYp6qQfqD+EkGA/RTGumlijEpJ1kgfmhDhWR2GQ7vnu16fSYT
r1An9GjgwjU1nXU+6dRFyoFJ219VfQbXBCBgQtcQjYVnij6dte9WjAA/2d5tPuzJ/PpF3Mt2JqoU
D6auQ1L0vwFA8y598fe5zmhZhIl7j8S8cPMQ062unrg1+JPGX0FCRQswuApA6+5zHsEnLLlnqX5Z
/GxHgvesPn/Xm1qwjGoUPHQ709DST39PNYNQjNK59Qm8SVfG0TFVTmOQjXcAVOnQWmgwxLCeQkRO
ySRQEIea79bHSPmiwWb/33jl878xK2b3UwzsfXFF9djEZFJnAD4hpvwakZdP9gZBcSL3ktz+oTOU
ibcjH/O5srAAeP6E+O+fLCwAJVS5hJkdnl/zMCxpjR5kdvp4mko+waz1zehca9up+0HuDQHHgT6m
AtOZ1rD1a6wZ8H/5uYVAPs8vKGt+8UIrzn0rySaWLYGOng1Ipp0DS6O2L8l6bGQNz1BXo6uBvHab
9xePSn6HBtcYl/DVVJ9fUNwwpTRPkT+dgglt57htXb3HftjRxg3Og9iYsKLPK2Kmbi0qzBiEADlS
bnDYT0+wCPeFQRWTZrK90Y1HGpaJJU9qTCMA0oR1tHvLPKXpyrB68ynBjtVcjTmGpoNu1XXASTly
M2Xahp084hbIz6wwhDBo9VT18CyCHJDHF1vL0VqCgOtYNvWzg8AXqc+t7IJID0Xcg0V4dvr8tvdw
nXdi6NudBRQc/IZWCct3ma4k9auD7wAgUf9XaxPOakWlHsCiWFB0SKZGRiolJHcEqANastU0G2Ye
8saD8Da42PXVtaKjYeqQkolq7+XsmzZhZgMtxDvZ2NGnaBz3oPzT0x+QkVYZN3GzjE2dRYab8H/d
cIXVX79r/swEQSNRaP4DXeIuP96erlYZ8SrI0KV3sCfguYMP/OcVlu1BRVl8XgUzhgzU8n1zdGqW
GZn1rdxRXFhbFjQb+GYLU43oqh/1wTg7XAyGY5cGnV5+ARyL5x0MymgnRabgOfYUGYN8BxCg8ISc
L+MIZiZanA0XGLdrfrWYHWUKp5yzSLfAeuF+e+cIdeD9z6234emU0bxkb+24djTOgMKPgfHuODsU
bIg/tn5NlqBGVr2091IFDONq6mnpyzQQmgVUIo5+JttT5JLATbBKm+0z/XHCwUupevWpp0mS3TXm
bmlKwTlfWrPTjBD/Uj8yp8rKajPZSnydC/RwxjFfMdcDe6UWfh6hNMgTsHRdqvPNtw6mejkfIKaA
ehuql+OqSTJIFtuqSY/UrvUZeGeQ1Hi+5YSUHbTPZZuEfOfXEa4gbqm1TCMAfJOC1MaKtIjNyIU2
I2+orcyzJLpiRbl7Kir1benxZVz+gj0G22E3aUj8ia1DAcMvvga2Aj8EhuesJ112GgBM7xnQgwTi
X8qBej9ETwRlvPChxzrKcqOz8X9Py8D/IHZxN6z9nqB+ju1NfMYDlcPx7/X8cSMcGLhVvfdN2KKv
2oq/Igds1RvVsJ8KWiLmmE/0iMWMbxodcNP1+Knh67ua+/4uZbqKLsag+73CdMJf8viy56L3OiL7
kykHlLqgMxLYOsB+nhlA+BZ7Nu7c+fmGkarcE3yiDsr+x0vF4eStJ96dgK4FezFv2PZDzBwyLcEI
aAFMI3T3IPUxq105N9MhCvZijcvc4QQz9sGekg7BkRIoRbyu+9PmCbdqOrKJjSOBDiMNmhkWunIy
Hx2a5QqMoTGB45DvMaa2/jWzacYVnlbbLfdOPPsJoF56wa1gCgSJIidspNcznXlXofff+hkz+ABt
LVZW4trB/K50Of/eO/+ZKcb1FNJuwKC2GF4ZyfVamRtzPue/Kvx5L3EA8OUjV7GptkzhFk+nWNGt
GCdAwyVuUHsy+dhrIFcrH0/JDFBJLoPN/I7HVA/WEaS5uPCp0IdiefDMy0N2aTwhuXup58neYGa9
+Tf91GI2ZEG/ntR9TYEOA+zHBOTEgQ8f9OVXN0u2uMgm6hoqi4+o/VzljtUjD6IwFk13D+IYtTZa
DCnce0hUGJKm4Li7WnF4D7GJ80iYul/KCYBBeac2AcbEqUj3enI+A9EZub1OAz0sXFkFKP9MEBuY
CztRlFyGNs123gBwGRtzhBCJWFAuQYcJ2MXm4lk3dCMq79313Zk9b7HGEIYu2kZP9KMXzyvcZ7MH
sMSX2HThbdn0fI+7+JEGfFBgupricKzoqWXYlrciGIgx831wtmjPtKT0tkLBlITl4cpH2x6ihUcC
fOmrHsi4RT2fUxI2zOdHNpMqsFSlrz0ep5ibqJsEMyUJWpCCSqyt9QOhJUx3SEU75H0flFA46Gr4
6elbDxbyyKZvCjtCVUtrTgXryJBQBV5U1FEbu79tdJ6jM30gEBbLOEffGbSX0V7cn8ai87vjcbCA
gaJxXlAMVoEY6Osm58KWEmhtvKd6zQjxr4jpnS2Ws+bQUY2VyIoBXcj5ujgy5HLQs7Ugg7am0W3d
5MvPpk2plBWbGYunU4ut5/mvQZPamtbnn1rD8zU/8kJlU6Gg2aVTCw2THmL/j0IIo3eQVBPFw/ir
IAfjL+9pRgZOWCCLYJXcntIk0sNfawU4WhQRW435kf0GL8rXXFT583h6xqfLjMzurPCSpFDvygOL
j5kPvU7/t33Y2Y5Em6EC5NzkKH4+PY/8sckq+1sSHwJjie2FAem7vr1ZniU3Rr2NfZZ5FZKzf+l6
BC0hT+Jv0fzcVkzTw2coO/n28YfcH/HsGzvL12uERnbVp12nRp6NpHQFVgU3GmCuNGy2JPuNwRVB
gv4v+Pe45CxHhLVJiNtpOdjA9/A/xGRYZ8tnOduqbzjkok4OcLbk3fk3fH8yf4z2dMrIT6IeEh0+
kTVTIyOLI3weFgBwp7HGaoi/ZuH75S1yqr06vQrzooEJNb+l1Gc9OfsV3zLZnhxF5F4znzNgsg35
1be4VKb7i93RMYObuNx/gS7CaFJfQqbxUJxg27Az8qii4+PhkZJ0Nkq0DvTlF6UcdfDb1bUxmaeD
PyKt/JJnH++m0VhF0I3ZqSGCQWei56rnE8dSzonM1zFdGOv/eF1hqKEbANtnQ+Ds+3EV6waqGdBz
F3rw2JsNgKTHaDmrvBV6TdqW5+7K8JO/TJyQOgW0i6x4Ub2UgdEmJAldWbW2Z2VxYUUh/nROydxo
vXeABPRpXhikOzqvyb17+wIxjkseLlCiWC+9Hkg7ap1dI7NC4JnCvBe4vBKbHOyeXMPH8Mmgzpur
B1Qn3YhvX1vm4Lyze2aPJ1WekIc3U7Eufmo31UB/HkCGWXIrNz+2iPRGilcBMQl9qdNFZrWR9pAR
whPPbBIG22UDh2INK2ZeIubB+E3E4x2t+/v1eaATPTmVUSfxT+MgT1MGUfERB6XW4A8y323BwS5R
W/X9R4EJSag21s/rDXYcxBLlkH5is8L0ITBQ3ld76FzmskJrgXcO7p8b/6tYDlIvgszCdfrDjx73
09G4AprtjvNd0xHmzSP8WT9e5khaT3DbNvQgw5ZJIk7XbxiMg9cAqUco5RNAo8vk5TAHzaw3dRfn
XikS1V1dIAerslwmq9ai1RvDauWsT8VLY/FYbs63zhcllato6hocSNjSd49TuIK6hx2lzWG89Chv
GduIkXXKHabHkE0hZGvkflh4qdeTqZiCs3HUvEspBIYWkO1x8IVe8sW7pXBBjaqRLr8D/l8fJjNj
FIHSewnFSoplv/yskP3APJF2nTY0UJjxkNQejgEkpHmx1srPxWWVpWIspZK9+Z4Cf8lLBiKqvlWf
MmgMU9G3bh+2l27TmBwAZK5hK+Fs1+qxdRfgDuxv7Uy/G54Fanlp7gUg8SKR2u1ob9dSRvqNS/lO
pOx3t3LlTfcMpq1nsTsqXT/FlroBJU67ugodxmJzswyxqXBg0z4hMxa8pPM5sVX2fhbimpqhp/xS
YCREfI03LDEqA0Ro5K8kdXPNCVo5+1gG6nNalV+RS/bKnYXIXYJB/LWzxeabDv75cgmkJ6K6NVcu
2sGeaImxzDQPJROYO6lGR4LEJ/vN4nOeft4JwLGpfLOPUWbX6pvV9GBs8SdM+Uxs5htD9gdknNic
AccgAKHC/JoJ7iVWL6fIFDuxJTx7I3XeYtzDM7AEx0Mbh0ZPnDa8CL7jvOnmUFRfSanj54/up3yV
zq5O1RMAACQ3jtrGPjdBlylLstnmllmrj619DHXEUq230fotTfsGRg6iyRd43FPY4jSdT/3SPdSn
RjYkN1ULYMtFptzudVKQ9vdYm0QoI7icxz5UVakrigCrlreNMEgBWzZWadKVSRuuJor8d9Hobjj8
xtY1iv1GwkzloChuE66frMaW8AFHOv76CKpgp0EowOEZLucbPtXmwJe5w+MgNS/hdei4tCiSc6a+
zqckcG3BS2qQNHalwDkrT9mNml995CVH/2n79UvShAfRwIFeSLOr6javKxzPf/5B/LqwEGK2lCXv
q5ydIDIKZ9j+KGnfVYLQAKMhEorEWGTKnBYeyvyvVD4nvGAOQTZlYNTKBfbj6qq1uXE9zwha5E0F
e7JumeQ6jPRWZpn/oSSlPOSNpVdVTmnmipz/h/kzvxEoWqv6DQ7Ppa0RwLJaPtuQ+WYtjJRn2n14
aRzab7l/5H516En63JA8f1krAmQ51uG3XbqtfW2dOywRgCVWg1ayBUblnAAaqzi121zxeI+A4ril
NStmrF6jOJAnIrjOGbLoH3Qnca/GQtQGPPwC6wOqLDCIzyYpzyjVKwQpIOx6IunqSjjZRe1CP02s
1gK5VYfh59hdprEWO7lHHHXgUb0dwRPQcVmMYv/hqEZBYTe1oODohTJD3YvMlebuX5pTRyhWe8jT
yNUHpI7jwfQL7Fy5pWySHNv4VUUu2MRdI5xsb39bbr9xOj6ELfGtXVLdQAon/h99iOcdN0NX1aYo
ohDohGHBa8Lxr2SmCO7DS4RJr1dnIBWfaxo1dNEEU8/ScY1qbnDDuvMymmzpJfIrUQII4QqnW/9W
jEkcq9swxj1qdXZXagdJiM0dWxsidwuhrizsInri1SriuqjCmfiGcw862s3A42OOniORTWTmfpjt
DcjOn7ajVowqRI0GjhKCW2hrdd07HOXIUhmcuPCh6I4WYWj2nZTgBEOo/8pufKafg4lr7e8XZCZo
+JksdZpEDbR8T4c+g0Y45KlwwfnRYkns4HedIu4KRjuIDgfp59Ke0lfUnhVXgpignvI8umrnsHqd
mtbDKsZxWFarqq1nJ7uhdt8i6qvRjbyXcEJ4d+msz9UjDsUzTzDIMYD0qiQnw9k82aXtAPIp9kCU
3vrP/jgtGa9RnUKVwcooZKyCWp2dnhXOB7NXJ3RGzQ+9ZA2+rePCxwyDsQt1haqLpyo0r++7F7tr
QNGUtbxyArB4orjsqD//EeijNm25UqvSjka0nrNfx54GKkRq6KAjkQMBiIbD2NuFOGaCuFdcoKYf
jiJ0Bkj2n+R8HEk3qjbmuKPg2fcYioBcL9W/LvkJKwnI9TlYISNrIrxjRjFBt2oc/snjY+tlfzDk
7kqnYcrY/7VOxVYtoPiuJgzhWMoep4o5TMuBt/L0tj/UDBKVspE+k1N7hKALpGUHHqODV1yXttD0
XPqoqZ1iKneKUu9rHKs23sPHxeTEowkZ7xQhj2VUmPDvCfR4gEY1nLBMtMb23jfQJ+tuKxG2C2S5
uJxLhVAVyOPKQ4BjQT8VeNVVE3Ick8+xi1+yNe8r3ZDRrHt29VO/ildURxuWbrZEY0Ep2KtvTtsl
d16vGD4S6D4d6rmljJGXZ9kdJpNoDNR89eLqkrl6b82jvs/xXDXUor90eLPCF9reogC3TeIDLOO0
4iZFnnpdAAFv/V7t2i6vTNLBbOVSGan2AsdSXsEJraEoc2TSQevvEfSwNIubmF9acORdiwm50Fxt
yh/JrAWarHI4iFdCfN1OXjIBjOOgHedZMxyLMZWZYRKtBcigXIwO125k4f1/+3kqKJFwjJ7+TeaC
P8QQXDOQ0F2yNyD+a89RW5Dl9vzW0U0fE8aRmvEtsWc8Q/lnwtsaZ9Q18+jGnp5SKSDF3PNNeuLB
XWjXcqwci7ddbijPsw8hZ7+yyKxSX2BgAogaBW0LApP1lIH9dsGxBJVhjhtE9pH6YRIIKAm1JsVv
Ph53XYTiIEdhkIHRo/2Zdw6F2niFn6VTqEIUh2n4sK2pL0GeQr4q9T7JG68ayt92OrQ899hFIxfj
RO78u9U1gjoL9jlGT+CojjGGN+Gn43uceKBD+MWrJSjofIHq13Op2Buj5pbTCpchYHf6ABDguooF
4nHoTv0Ya7U6VqzIlGbnMLuZyiIivyozGAVzli9RfA//beboByO/uyZeI92OH2hBLPdL2QUABDtw
ExcY4eMcxzk+oQYjSji7XkLECtV4C7ue5bTv8EBZf8L/G3URQxjTRzTyTv8ne5eIabLVpuYLCwtb
k5X2qZ8crNuE+Is+jkmH3SPJW1tJfu1GcN9wIl9enxyrZUNKhxUaTFZNHXI54PTwVWUglkmWXwPX
NfJP4Ov4sTknGfTaAfGToS4ZAG1qpfFqSJYIw/NAz8COPA6k58vPd+srbLsrGx9dzHdZDI5MkkoU
zmQZPK4w5aEqvbWAByLeo13wQBpZYvr42Zudu93DqqSjuH1TnD2Oes2KoJaSX+Mgk5sHJwjlZcas
SikAeCqGBnPgNnaCN+3V1YM1WeWixBc7+T7KtL7SwqZFAByXJYHFTBUhoi3NImAqAPK97uLc0wyN
UKyTMMRVCabDU2KsZDtZbH1Wcb38olfe0fjnJ5cVzNZFF4mqTj/QkwTPGnEwDFkpi6jABBbGf/Zv
9eeTkj0flYvDD0du3j2w4DDGIc+dF/orowKUbL0kvr9svIAlDQGPnRvKb4C45XuOWs7fYBgSyJ1N
4L1q+BP1blKy0US9L6SPSNrb8vhR0sGJtUAyrBAxnk74EJMjAFdI4MsJwsG6x02tsA03VqNng95Q
69VHd+PEnLQW+eJGVvJR3Sa+lzeM6WJz2OUuLT945YpGaoLbNKymg4UiMNGSC0JvVNaJyW9c4xat
JygiMIbiqrr7uTny+wy7zanor7LaHgHigkYk/6zxtRdjKRtZeZOQoa2NcrLYvuDkOjkNez0gDJ/S
k1KroqXt6rqIsH1mEPa2/pwKr+egNq6kmd1HFeopIxXYVLB+GG0/2DXrIqb0JZ+llUyrGPvvGKY/
3r4fBwon5Xj+Ze91S5f/GeRDtOoVGjJUkrNj9g/dcmMpChYCSi7jV9DbNaVOWhlSAs7keRykG5fS
PD90OiFkxNmiX1njPU/Wodhp8aUZn0VtdAGKf25twXicUAaxpYMt3w9FPrEp+vAkg5sG7Fm4vvQ4
gxTtsdqufWu5Xe2mNHqSryP/NKUX5legBTe/bKc7YWld7aduDE/F/Nu6UYCbdYiu9YmZ7oFRZ9pd
som1ILuNxtmOUiis9NEsSvm0gf6Dsl1UaB79cJ0rvbOMQ5ECI7xNDFNl1a3Ru9SI8FTstUxWBHg6
gFCGBfvUt9bouE4fW5gsa2fFsLdbNiDTaUOu3IVo8Vux4ZNopKFWPZXgsPT0KxZr8PFAjpVx8q2A
4jUECSPwIrzlvR7p3aYV87rPlXz7pyxZaSKiwuQdqEnoW3xevprvJWFg1/chsNW+PduI2/UOlnd5
bbsHGZE6wZdx/Mi//Kv6Uf6SM/1cPLhifj/gEobVeGQHd2/6ABqOYPZzzqzWT5ZZicj89EbTog4V
Sp2pKxy0x5uylCCxcX069pU5SdcJUbrGJOMSz4btYj8rl6BgYWK1t/Qotp9rWUQAyyJsUJD5gpJf
WB/BKaXyxzzfV59DfERL0CPuOD5sLDo0e0jK9Sxy5ZlWD/loOALjwm7UDgZUGOG61NJ03/K8cY6o
vC3KCO8MKy50C0KgjG9sojUjROAz9fyZQzLWcQMtlgKWZzPaNxJnThQlCh2gsqYvJcwzTEQGVHBJ
yo7/tz/LO6sa97QreGZKx9/ZwSrGWnzxUBvr5Cd5EknFeUddlSyzLLSARpLd1llnE72Vyz22gPSM
3Qh+HEU6meP2aGF/RdWkIPN3o6ZsuC/FzJpDNp92xsW7qO2y2rUA1oUdIJSBmPC17w4o4qo/o5bS
+dUDPGdMmcALln4i/VvjHnPju3YDDgp7pzRW6dhhU47W0VaRAzuNAdZ2XW7dRnqDP0bP/SCP1M/B
7nvOIos97D7i8oydlLigvgMST5l0nF4AwHhL6V/JLIx0x92bRezgVD6U1lYEiHCOhelm369blIT0
ZwwLSwZap3PFvY3OpjRMaTv5VtYAORQVqPnX/vpu64RcCQxtgPjT9xixYUWwZhxu4BvOCLvTnSv3
zW3iUGH66D8mt5iIZJz0byNrdXGkrPxMGFH3s6lTHyFqwVn5575VlVgqye/5hnZ95kJOFhBgzmcK
Qd9rbsIE1UJGa81L7javqu4DgS9IbKEY2/w9Ou7JIUPqwkgpvt9R9Mc/F5K8k1KYG8YPI7pnf2gn
FYwUrvoo5DTxs6ZtGp6PFnb+IjL8LviN5JLGuIqbJRlppcWsLxEd2PpSYKOCLKeQB/Jov4+zuaxV
LX3dGV2+5Pz8i7rp6qbgWtFwR0ULByqRxoF1uCFoxSmP4sMgPpf1w1qw0xPXIBwXMXZiUB5RD+pG
uS58AHiMQnI+9KWUu/bqEWootbQDSnBNykB7jbckC+LvcSGdW+Ybo8XXon5gQAo9OAePdNMF97cI
w6+hbUzOwWdmIlEerWkz+Jz4iitZeoXaFo0FRTaCv673pvJfVf/FzHEu/8IcK6T5ABvdgMv+MmYL
+bEZJ2twrqIygXcSojWQK4IKYS322oIqxDVc7/fupfcbU8SqUGUoTGe+GL+pOLMlCHYWWoejyP68
2skxhwc4+KyPrISDPJRuuwKag9dER9Y/aWBjHKvzjAWMPWt1DEkYXXZjLHKqtvJqn6Dpb1NYMCQG
MS8QPXtMccNo+DxsS9kfbZa0Q4FEmKMZMO5fU4W0DW2vAB7XX8TVH0Pgl2+wWVGL4Y79nbKCr3xa
YiUy0/wX83iI3yaQLVbqg0iHCkjBtHsC6f0DwJfwUh3+LCx0b3ShpXoPMm/IXB8P7TAnvPAJPYts
2PeIpxZJpZXKOgSuz/rkyKvj/otkKddYFafGG5HpS1+bfq0R/wSSeaHnnl6Nj3Cm1/+a7gqcliE3
rg0DCFhXCzxVCW6sWOvQRumSWzMo6kqN/7nBbCUbrHInKOS+kiDzo/0vDXOWJXiRwg3l9XGESxrJ
b8bp33ebQ/mWRVBfuu25goNuLp6OFBSiAr0FJYr/nMA2nmgWtKVFCM052f+K0kHeN/wXid21d7B/
9N1Z2FCqq36KZ66aQQ//N4rgtZIhgzqbk8Nj0C6fBBXo3UazN3Q1SEc69tK7YRFHkAxUtGzA12Cb
4odCfXFID7kqgnWrhuOKwrYYrJ2Vz3eMWbxrzvosXvrfB4OsnGcnpdhwN2D5BdiSi6Er27ucpVjy
y/g7QvHZjbTxN64PU9tREV+YpmAHWdmhhbRvtEFA/73iuCq08S1FYp2GYvzg2a3Hb/bbM+L7sxTh
STiY1KUX3C8sBWGo7iLdU/ry+h5/yOkTDwIDI5shMJ2ZzW8hAk0rJgighQGVhO96Mr/UrIVVSy7y
1USohHL9j2sFwBO7GG3GHjB7JmJHWz4VZDDq1Ic7wnITzePMBx1Ck+rM0PNAuRHozV+71BQfquBJ
hzg9BXfDrIf8khoT3HIAMK238D0p2Am/jxZNDjpbDl1W/ahEtHZRcWDH0gva7onyUPZUho5zvVa2
RyxYaoXA2bhpqbW7UJ0qZqB7p83vnHwTnWye/PM0Xdy4DHSUO/QRf9nWl10DooHKlto/sC8kGspZ
VndC+XIIoJIOh6VvX+jt4/0+kFQmoQa7qWTqyhut9XED7ETYLK3T7QnC+6xdik02LBruC+65oYfx
z5H8vqlNpgR9+5Itvamtw7S6ehIX93yFRTxSXLoKh2wt4bzngGl78yihT6+PblozM2LG5S/gSKbw
68M+Vo5yJ7B7eQss36EQtQAjlMJnmxKWJOTt87qwvf8WjrO48wnMozNk7cz9DG/GAf1l7dYoOLWF
I6IjKnzmYCitroN36gv0nwbPCPngX97Qx3a0oDSf8OTZm90XglDroruVkcR1GJTGGEcz99kFfZR/
VAatLWARwNPSi7uSBqNy4lBLuS0jzfTRxf2Yo/379HxGSR8/EaTIiYcj2uXPCJy2satXTRUtfU6h
6D/h2nLCsBQGNYCGqZRG6vKSqEqORGqNH1kOJGV+yj1LdkVK0SOFqotKST5Vhcu/3MIpjnBm6LJk
M5Azym2FuzGSQu8SwJ3hgOiXvAcCFZByIjBN+PV8aGkt5F6nVAupisQiEJrRNKX5pwqd0QBfCLke
UTXbKnHbUkNOMVVbBeD8vtbn8R1yo08RqHdrJeFvuJE7aKvlgCvxu9zREksozcQ2hIl0Q78mkqgK
3kXTtR69B9OKvtOPA0C8+Dx+d5BdTsIG/DYNEVwWE1rndFljegbUMe8TC/enAnYo/yDluS6aH/gO
0XHbxdWiQXmpZGYfuYcdcUnJsX5Ft/D8M88FC6ZEQA5OAMFJD2JzU0umVr92LyBteoEYH8tD59IH
Kt6qjkduV6G5TCsISChqSulgC4LuUvQ5E3wKEUIt971VvZ+B/1vyQB8RcoguT6HJo+jiyiOG/c65
yl01Uw7Y/imhw274x35glIj/30EpcO9CCChY66xc/tW2Y6+Klh91OZLGSuboydni8QKER4qBXPlh
IorNxNoCW2cdrrWF6ML1nlvlRweavBukyOEvE7iibEba6FwC+ZEqZmg67dqlEgkp2X0Muwxosoub
NfvpSbwVlMC33FRvEL6V+9RpuyiiJ/Epmu+nPQTghNWYq903HeClQTkwbhPoDa4vUOs3QJri0IwJ
SZTkmk+cG2MPikbBNhu+wlbndOfPTOtYb5CvbgjsXfdyF8/5xrBH82BEj02cFsapKBhH7j0mDohS
IBcx3jDxzA+GEaq3MBHynNUpkxC01Y25F4z3kO9iu2uhW3eqUh7xkOFJYrUMXLBA1wd/mQr4xtP2
lxJboG/SgWD91vYTMUgyani/DNprR1fRVZ3oA8aVtBPoiUtSGgb16nAr0kraOTKRu/i8rRymbhq2
vCHCVIA6cwas/vLytB8EjYBPZ6ONOrFTD6F/ehLu0WQ+clVI5nvlC3WgcCD7XRoJ9Rw/m6EM1rjT
5Oc/oTspENRHjWWSoOPcjPo+J+SkYYHrF8Cf+MfqDoAP+bWkV76Wzt/1Dbio1wNsYSW0Vyyx+w4D
GjL4w0KFVUlFYjpweJIX11wIBEojLH3qscNoKVMWyef+vnNJXqntDRfk3fJ5HuIwZcVDgFPtMgfk
EqOE4UI7+fPfTjOdL7D5g0MnKMravg7ZrRDTjZtHGRRw7T0LNx65Xzadx8C93dnY9foN2rF/3+eM
/HlWA+Ya5RPKxdRv94pPIwqd/Pb5/NqxUv2pFSNSruQEVi1PmDr7RY2z6xikMjXP/QKdoae+4LF+
EwBc8bQV6UPSMC66r1GM/LBMnv1gBLF3wsaJYqjtwfiYeh8E9M7A1VDQEdUibfATgFctvZb/JFA8
Qqpd8u87isEgiZpKurpIQWCTDec8a/T5y8bV4yc3eOalBgRmILvNTfht5ENqEX1r3SEHiZNbjeKs
ZmCGpcXMC9By3Ql1Hpr27svn6M/CdcdTmn78vHR/QYDOoHRaqLv8DstsHhHlKFBYsQVlI72tdG2C
7CKCsAdKPE11/q6dGhH8dsfBDrHtCm6NOpWDBCb0RD2mz7pqRKpcKe/8bU7qbEfvwm8K001ssvXH
CRtmAiRw16DWpQn8g52neQ3RpY/Y6fe0jscTVFGAh9dztz8NRdp2mrW+JZd/V8PZzuQnlUNhAM8F
9+bLSInmiNcNt/Auq4EnVP+LdqrHoDUGQ9JM95RFzQdLp/EozJl6yljP8YmJK4Ynk2CP9AOhAfla
HP2Ft/A2GQFhyloZ2ILI32oAXIGxJFUw1QkWuQiNpgvRlQjFZFQz8j7yqfpvJQm21qP8G+oF8zR+
RIaPMHilvEQcg6g6CbqQ/gN+ils7236YTGMuJsunUN0x6SGVAoTk1kmC6/L0S3EyicCSQbEHT3Cf
nwoGA/HkidCDjtj7yPCwVxeHaFYEShnR2PvaSd2to86lfAKtTlbBpIkTY34Pfq2EV08e91c5FqlU
J4i6SX3BscTvJajhvslQPlCMICUHukRMSOXMfhAk8PE656aDHsr9WI5MbKw7zz21IeBRCOCbj/KJ
Ae9yz5Dlhd7Iw+th/4izImzqNRu5oYI9FFMGVqlRvdulOohyzqi8kILXbsqbnLypu5kKwt0QImKs
v5nS3IimxjXTxl3MW2RRIMTCL3jEYeIEnx8VcOZ1MFmIw9FF6Ey7SPpM9tuQb3vFuHFwQHIWLQNJ
65+Bhte2EGm8QhQXvyCSPfQMYnDcbP53Dj1viFWpAmTS/QVyTLGy0zzXXxO5yL+wCJm6+AMRlzZW
IcMy5qrcryRwvE6By4pRFFNYv3QfPBT5v07IhjuWA8RVL+8jMKUic6culy/9o141gW/tU6VwPdNC
1T+41rpS05fMrB0LBo/Lei7CVJhv/axxu9cOJOhkjqRKiqcKyDaCiOwfWl1q1E1Aa/5KotY76Urs
HUxNcBpBmDrJKJpEAZj4sN8LFUtBPnI66ddMorm/DSlB++o9bwFdOQuBY/7S1WoVhm97d7Mbz4o+
d5xaDwyfEMF4spbLnc3ElzCgslknmxcjgN77hJGiWO779DMsNuFcQNkpdwU/wN9KcLztyoZznptm
IKxy/VRFYsbP4ow+/FI38ilUO2rT0CMMg4bfQRXHVuFel/vz9Qi/5Sxy6U8nAWY/a5T8vhD+PBmN
1tb080qLA9swDM3ppOL9wWKQANG/yytwO2HkBwEWkpVSDvnySrktjrNfuqlsTWrOFhIf2cY34InT
OHu7CeqPIJi4H0pJ4SNBIDBmAl08ALpxq0Fwtwem/vZC8MY4amDBjH15klgcAJFYZpqWb8nkNUIP
Hfope6iQs5bHBE1TpEnh/2zilKL3NKrBjvU7DXQHrkp7pVjTHYH9T0OB7EDTHnrNWQVXC0a+ezHO
kulSFN/Ipq5asERijIs7lD/mouNiU8LVfL3g0Lsj98M5sBK4KoSYaOE0NZt+ALRtn8SAJmVAuoRV
m4evpdQRB+Q+9eR6w4UOsfhRJIIA7RORAvE3qI1t5uLWLQaEeReN/NpBhZunVxB4rsBplwN14zq0
Mq5MvwamRTpPS9GeSTJ4H84hiQuWCSHyPqbKtRN5UQWDKwslcnEFO3yzW/+Sc6/jFvmE01+0cBqD
h29Dc1QiPN55ddoByRV3NMDI9+en7isdprTaUCPn8W4JpdtFqbbsB6YS6RN2VS/62bsHuKb8f6zU
Ph+kR6WtRfIyDz9QNl/SlWK51To9PklLYlO5fpS338Ga+8J4NqtSutfZLT+iEnhGQORrlAPVdgoj
FiO3uvNtYFfC+oyBn3KXxiJdP6Rw8aXIJV1k+pE3LC9FO9UNB2Za96z1DouqQT9xO2+VYr0T2IeJ
LcJahvAMgI77rPQqHRPbLB/DQmw5VBqDfCCciFNNaU4CENyEuvyCjSe13B3NJpr4aWcrKTNRX2uA
zMB2VYiox4MKx8gx/Qek8ZpM/cDVYGQSIyLUvuCPQTNm6G9vZa19RyDzZ2Gufx/QMWHjseMXhtTl
jv4GzDwu9Das3/7+oAJoLCOL4aACa3wBRbW05lafA3FVSc0rzRqqNSHJJ73kB3TiV34cfNOkLkqg
8oTXbCntgngIU+DFAjvYXb7MCqte2fNt1bFjlU20qDM1l0nEfEZI4e3NRmbv9ZaElf+zkZotqRpQ
HvuHS+GbBFnm77msGuHzYYz9yy7AHAT80M0xo9YSxcXZxuwlB8kAyBV05EivIV27qwOAi79O2po0
ARZju1LgyUKsxL8+GeTNSotJTTc+n/yY+unly9EARrbR0vkwUstK7cOx9OBJ+y6JBOE0E83oj/1E
niy9OqjEoIWgSFdpiF3ZFqVUtqOdIXiXO85lzb0+SBddTAaoOt2qc9uhqA43qKmTx3Gg6Bj/0LQ2
OBXD5hUIVx8WvzgBuZm0pt+x2cPIZjpF1gVWQfKePNn9efsCscGXjcClWqQXdKURZcYxfkKC5qM1
O1a7cTbv/fA3jK5RDusAWmYliPeurfX/rnhiVHyBwYZtMRbQD5rYpnY+77RwHBjH7eEAHcU1AuDe
P6fq+zKEbT0wvrCKQ2RUPRsxyqO7aCsfVUqANBQf1efWi667NFlo/N4VnYM7a9xXMC0aodGvAdwt
L84pEoq9XRr/qKfldCpmkzuiDDfvmtPfr2wehp1iO+qp5cMLjg1WBsyLpCm9mmYo/nLh8IovZhGQ
tolPOT5jpc+pTa0fEOinzEEVBWzFyzKxjy9eu8mlJ0RPTzclowA6/JQAyp62ckVDWQ9sjhX54+zk
tz9P5J+gdZlprwW1TjUoTKR+MBChDhbzvZaIpdnWTc2TWw1jiYRw/g7YkINSEaXzpLN1kRGMuDkI
AgoZ1RsaeH952WaSE4Im2lWU6dIDAVqowrLh6u868kCJBtLoytxYAqj1oR0DgKiOMe3Kib0VBalZ
Z1fosAxBIlw+SjGTRfMgdaHSU7it2+9qSD/tZTda6rFPyyGiQcAaAsrSXnyD+W2siaIS9TOw9yai
xpp+0LiH4lhfTJMB+XX6jVebpniibJnpd4djY0vT9bKoocK/TtNNQyw28dC1OrcF7q/B+r/0RfT4
jEGQRwSKJlvee4JhY4rg2+5nYRsncKBYKM2FHaejj4iKOqBkaAIkkyaoInAPri42TMQlBKNTzfTS
oo5DYjcy7W8pRNDuzsHdZiiq+ZxNrOVxC2rsE+7931rGzMybN5rOy74IxoFZC9CkabRYdXEdH4Us
+IrXOXHvKsUeT8h1b94p1Mm4uO7OurRzH2cSh7Z1xZZ8pHJRn1R3mkwItz0W8NzMzMdptvwHEqs2
pjuq0E7pQJNeqMzVGSnC2ZKo/GX7frPuZ0tpL36DP+z1H026DXY35aIj4XEF3Y+hbaTM2B2b0r6u
vXwssPOcNaK7bATeqqsEsZ2ckn/uEgIjSxjP2TCSq3QgxbJHf5PoPC0A3RLsfv7X5EegLJuZ8JId
8M/PvTtd3L2gYnhNL+5sXMr9lAlmv7g4fsDtEKSx9eQfp7/gPAwSIGUip5bPCWFZzrnltalHAIDj
F/iaubVmUg84tg8dF6VOUM75QeF4VRvudgYzo9ajiysjMjGTOysTJ0GxUJE8HiRY7Z+kAhMGX6zt
ZJ+kNp/S4rEBP6yNFXUFuLocN5QpM1o3gAb7BAsvIdn5aMQh8+h9aU/dgW3gtm9BDKN8qMKBVcLp
liwMeNT9E2IsCM2zOq2vdp496xDHg4MmrwtXB2ppMoFjlCdOWBiPiMviX/GT4pSAZSb6JdCsiu8t
tEIk8hgGw7MexnSMo+aCgcxlhYuNochAaWggja7RaQBV356Tfmzy70G4UY1HyxbSDyTt5wSX1mTO
sry45qEVqkp7Y0mGjHAiS7s+5norXQai+0NP+fb3pTU7nQJq4+0ICMmCPcyX36YKMbGAUl3znPzG
vyYhe6cvEOVPJ51CNMjCOoPPjIzQAt0UkY2CngI7d3ujX0h6ei28KVBDyFc1S2xWPrJ3x73/bQz6
yM5AoZl/rsS667sM4/P7tVCzo5svTA+EjfJqmk7vQOIYbZQBA47kPD1yAw6EhS/wqLRC9eC870c4
LYm+zzoSr860KCqOOYu+WZweunhZUF8ydeOsVk2LtINZJnsiv+T4VYOqism84A3deYi8Te6cRhsb
GjNFSmwJjXhA2zkeQ8ZLMqu+h1LkqN1s7VhKq4mgDQkdccUPkTZsURJaggBYPIkTxocM/mkerxHn
CwFILfZjaJiRkxNjNzXt64jqrWdlfFeUSk11HtukbTTun+gxpkS5KObm7rhkanh+0OjeeqXBXPyT
apDOYtgrtrzccesmp7PJOu9UvcUnd9SJGIlMiuozTzsc3AI9XGKRisMo3R2XcSee1Q+cKpuSqYo/
xHEHuQPswwxc7hud9h9iVz/p34s4fop+cP8mwFn3yn9SXf6Ly7EmY3JCJdGORMdYvspE2Q8T3Cgt
WL0rlU9RFSN/sI5oLUdIVxzAcWCZWqU0wgVjg7d8ucaFF3DcMw9kw0mi9YzBythFVWaXS6RuqxTv
xeISu3kS0/+BOuAKs4ALVBOCDuCjUQ+l4dOCfAB1zwImKnd0JiphkHAQ3gV39cMjPmv0bOf13EPf
Ef0GALCGEmkrqHESBkxT/MCQYnESIQpqXsRVkDlIVrU4qVselDBNhrQHsz/I4xkY22VHqxqYxOTc
9u0sRHAfSjzkhV6fpihbjBwz8hF5zDIP3Q/9De160hPSf0KRhbPOLdSyGO7hql1Y1w7vmSSW8yTF
3vgYgSPAiG6pgbz+J3Z2OehlIS3U1lIrflCVPohUtets/jt8ATDiqRjqST/RN0AXvwtd2wPD2sNs
AEpWYThspVHDL32TwV3Q4cLOW46sA7zk2f9GhXRrWvfpXPvTOMb8doCyZzTj57+6VGTccxFOtWs9
l8ESiHfmHqyxAkb/YlDXby/owpyDrofAYlBNTV8m4sy5fXi22cOQ/YH/gHZ4hanRKedeSbS9XqSr
/95qdcQpOulYACAV933evcxSYutp5UNuYyv2gK68FA8fO3+rxtAHeWHHPyJ0umivZStGmYOuD1S7
h8+2+ADlYLiABJa756zFzT2G/xcmk70QLX+eoa63mhLwPKG6tLBzo+ZjPiaC9Kkl11Lghbs/AWPj
0/GpJEx85S6rjxv5pak2KOIpQaqQjnQgV2+g7KYuxKe92xw36BWj3RuLHN+VJfpExlhuCCJqJk9m
aHbqYKXdC0wJrn7JEp4MgEFT33jej9eh4pNVy3rlV3ykUKar0TXWQa30guyh+uvVmLAs1z1tHD12
H1vGQ3deqCM+y9GCYul/UOGXtvZb91HpbamJKtYFgBlEJnXeAQ0o2v1oHhiNeH7D6LRBwjGIi9GE
5cSp+XJcFD2Ea0thpz5q87dGXbhXfAdVvOl5Pzya9r1+uZXbmNvpBIKsTX96m2W7Cys0TE5sMoEf
ftqbnfgjVgi3AdrC++X267zBx5OBqpjtKKKD6iCvM6PSDMOvb+v8b/Yh+7fCttbsczJ4t9r5Bn/n
qczItGGtFRPieNFeQuh7kQPgXOf0ocYNzzq0KdQCpVhHTOO0WLywYQ0JoKZy17npK2vIzO44B+jm
LICPI6SYOYKo0Wuss9cpRcUOKvLIVzAsmdHihWd/jKT9JnAXzyWVvSGeCtHHaevvm8odJ8KNVH8w
TLCZqKYmhVn8IGoaVu/kXodfJnq+MzS/hZBz7yzWh9GYv8iyzvGGn9lhNb2FLUXLJIH3vvuaRRq4
b57nMjzWpXg1vhYXKKwVuV5EstghGT3yU+eqWKQZKiqaoPc0DV316d3b+mXtXGnj43uqt9Svdedd
kPIW8tZFqW+t0XfywId+gTgI1tVVwimJmdILSMrr1k57ooB2+bHwoAxdlzXEx5MsIkLcbkyFy1FL
R4xL2LJ8t3bU8OVwAnZxgv2GJFDbggliPTDkT3UsIDyPpwc6HDMwiOeEnxGZkYAscIZYuE5Kcsct
KYFIoxf6DBSZEpaRdpvBkD+ChSgmemdkM1MpnQAcxZ2NpdTShdwEQIuB6Q1oRotQCXgdsikD7Y92
vTKuxbvmbN5WzPXuEugyghcJfuPfMxjOZQYrvOInaksXVKi8ifuf2OGf17G18XAJkg9jzr5Bozpe
Sj4wMCwSy3TnS9vreDpl6vjTu3HHyNZJn7RcRMOb4yIAgehCm8kW+E/BcpUSg49JKpEY0OaIY54J
0l9uTZoPLm3hwLUFk81evMJi4Ct9r2O/UINrS7ywc/7123B9AxSGPzpMoGQ12TgUipNojAqCfOY0
KhQCAw0JTdEJdsEoXioLowiwoiXXMQ8AdtXde3nm/Ni1YzuhtYwzYaJmmOkw8T9PHWExrSULUZji
i/WquILrJnYFxn1Z2Zf6p7uNqFRBxEYEDksttGFGzk/L5uczF/W/LVx4v2nW8F8cB80C4yfs+sAu
65SDbIRgQ89fdjHwf3qV3CIQvANdI/0672z5ACjZgnCneIF/G9GI2NdFlgowfVr7PFgYm55A318Y
BQWOtodfD4rmNq08UI3LinRciucH+MhwvdlD0hEe7ZBPLSn80na+YYwO50+/I2BYNnv7VH1mo6d4
DwpllBmR6DbxQ8lkiq2je/9rNqEt68t0EC4resoS/X0L8ouj2sCfFA9/Vts2pdUOg4SiMDXJgvJu
TREWCPxAD1KNkiv9s5DPyM7CTl2sU/AwRI5UzaW2S64L+9eFmBxSErhBk1OkQn2YYROvQSg/LE8w
ZscBaXvtIK7iIKDi8f/F4oCdvgL9c1x7uLwNzp7VK2uTE1XrkkYQ46wPlaRFXdbthJChWgzqaGrc
yhNmhYO4nx5bte7z6TYAPl20ULrt9JP6FMd/BkwT0q4TmLlfvnQeEwnWC2BuCs3Q8sjC1nSDIfdU
poEuz1M1cMXbX1dH3SbIJ5V43npe7Bt5P2pmNvgmbt2RHp7HbjiqCscfLWzmZJXuEOLhptsTJgnJ
k2xnPhld9xNV1WYf2fxDwEagzBGRyoH8WFEHOsfgbzIAJZYg7l1y9+K9wBUdWwk4P6LH327ZOiZ4
9twKrkGpuhwq7AKEp2xi0xV94b+tzT4AXxMgKUX501JNBGfZFrl5nazpNZ3y4c1NMu3GeW1nVCBI
xK3matBazKtluN/zj1JOPr24Tna3IxOgHRpeLtmT6VQ7gi1jz9jb7EJSnmqOJlFbI6Z54cs/6Nvu
ekpdeIoxIkOmh1GtEtvYkdZUCE9Z2ISWnTiVF+KrHJo7iQKak4+686irWpvISOMbcS2Z7SDvnPDa
2/jIw5r01k2/LO9cbGb4DL1Mda8C0UfYd4f0JoHc8KLri2h0edQiZ2UcyVIgJhcEPlS5nc60flUr
958ZHKZ2gK6CWGWHRhhnvikYJoLYkfBAvmwnWb7fOTy0N8pKO8jWh1sqbSoHFC49Ez23Y1oudnar
Un6Ib76+zNJNNeAOB7Nk12YWL4ZqmP3LV2XZbNWfdphhc6C1Sq1iD43H8hCqygWdT405ZZyyuZKt
2e+nvPAhMxUX9B4ON1AUkdLuyX6PbR0eR9KC/0eNR7fqlRNxGtc8x5KCyjkpWfsFNCgsHlopO1yg
FcuQv3RH9jnmhzMqCW+Bja2rzIFnSnM9gdSUEZREa/UIo3zTBLbIyLkKh3wqkh9aDWeJWj+0fui2
tH46fzjt+ANde3IYmy5e/nugX1ABS9379zjUoq9r5H3Ux43QT0M6etqbYeCeT5WC3YGC7QzGOrcb
WHOvrEHT2JHhhHQkaz1p7lr0S+7gDsFkWO3jMMskT8Bl110YOoaxNuhhMPZZjH4uZ8UIhFR+rM8I
hU4qXrgnPV0bT/OWiZtfGwMiMeE5sr8JDJFiveGmg9say/nCtzVhNK77bBv20NAHPn+iYxD7cV7l
khsIFhPcKQPS3wRhtiAuj6QK/KZflvWptcOmf+rm3LSJFTJ3s3EjQyO5cA8tF67EzzH7IUpfnm+M
XCEVUbcneOq0UX3S76mfe188LmW7wsDGpkfW1H3dLDblcM0DPJMBuC/1w4s591Ka5BFUdCIX1jcb
7/GHta5NSzuR9DP/Teu1k8z1EKIXLc2l97iJs9k5Cb5ITG6CkR5PJjMAJHFEVgdEuWBOYz5DrvAG
H7IrYGDJMejxqf3nlxk3r+r4DuvfjpY/lkZ9OVnuS61fUFl/cFQXH4Az7Xr6iU9YIrAYZiZDdThW
7x1ddTM5yczYZobVh7cWf1A2ft2pNQx0pR/igS8l/I1uuwWzjoLH3fgmdxVZaXdteZsB1nf60T2e
IQRc7JOdLeZrvwPYLsG193+wz7F4dcr3rcze36FgasTog3YW1iUBVG3Ms8qJF1n71bJSb2szOtD7
6OMK4SDeiupqb1iT3aDCFEnGL5SPXgIzF4aufz69S1cygdGOyaceFJQGEiEKetf0PWK6fKpSs/BU
bzjfzEREFGifWH5ITv2RJbP2zS7Or6afOVKv/tqcAU0adYxxcA5A5zakSlJgIHu0nV27tYcv4BtK
uqW8VmgJ0Eh7WskR+dniBpAlJQhqHKOLdshSd6LY4X6IdEsHORhQ67Ynws/MBsuO2n08ns7OKWa2
n8yeCazAFzH/2/WELbDLUzeZMZWqqepPVOgvI+A+OuEItk6HI37uRGRgf4jV6SuPj8BNVeKa82JC
H5N/yX/FLFcjb1/VrnNfB+MVTl6Ozo+BsL+KhA9WUZyPY1OOkw9xGJ3yP6kLHtE15+P/WMRAwApV
LS52RuCi2EKpLnODY5i8PRjrIqi5rmsHaSEShZmKwv4pJPYhEm0Qm6SGIy2szmvehMNinvjiL1E1
JHtQ/f8YFsPaJt7mO/I6O0xdJ0AViFX97OLTaESEEGyohxs2qCteagJ6a+CtSKmbP1I19/dcQdeq
3+UpU617pwtiCGgjkB/sIgBSziXa/TAXfp1ST25zeBaV5w50Y5UFNQS+g0623Ca2IF3MwQlgnfor
Ai5XHGo3yi7jTBo+DtZPvtcuComzH6Waq2wq6dgpTPKPgZb5mkCAuvd4mV2vZtEeCDzqLE8T4dTv
dndj5TaSXs5XshyyDxCgm8zvU0/qHo9V1Nw+VdQuQtJ076vw6k2riu2OL+qo9tni5jUdSrrWlTPh
SB0h+1SlUGKae3tbSl68ZF5syR3uNZlIkyJ/VubjiflkXGO2FPUoB+GIbmcH9Z7IqIE5tWL11fI1
PdmEXYjMAHNtG+0MvtqPbLg45KIMVE3muhvAxyqLV7JQdqgNa5GzgXjLN7p4+2Jyqp7CChbc385D
n0N0VpA/bBLhRpDQRlktZ7XagZo09MeXp47KuK/BcgexMCHgb2ZW6dkAQzYbZbZiS8l1R1wxABXz
HhyF9CN9jExBG0QbL/vB7+Q4iCls61i187hzQDW/UM7mzPOHRZa6AlIoUuoQrN9ByUCHUwh7iTrA
0+1BF5UVAdhCiidQXxn2sEHXb6YSu0mG724tiVQsOnwx++36RLqyZP1iqSTBTz/leVlII+hhhlkM
+rRPSRovi6C03KmoY/0sIP3gXJtMrANsgRpmB52SMC9qafDkDg2Fh1my3N5OHzy4tx1pHywSl1AM
ml4pDxj2mgixfZdUII/dYxe69As/K220ofeiLsVWc2UNrrXjJjY8E3x1H/9MXtVnjqt5jPKCwNNN
nU6lEwfv8heT2n4/YZJOBFgf8xGEmWparZ33GR2DYQyd7xZl3VuAxTsmReeTHIqtpgYbCv8jf5yA
FRaiOpiTlQsPlJgoI5h+K0lQvTw9SUnifH8QmGAqBuOAHwAuIWzTF6FxINlXG4zAPxa1JK20o3+n
poT2nvy6zhpyS7Ts9YclhDqBa3iAPzXjyavR0GOPBkBPPX+ZKGNyNOHgffImcgIv7lhl7k+vbQL0
eJhV4MUdMSdmYEVN6e/wqxUTmsw5EJocDNnpHpX8zsyiQ+yyFYtXD3iCX3YiXseqOSde+a/xdhVV
vW8B2YsCT7+v/RzRLJmENe70v5Eg7FVL1XTyrQGiBPIsJ7BfhfJbZprDTEF5Vd9RHFSX6s20srRc
KvHRRZIlqOnI00EA+cuEAqiMf+OUiL6ox2qZwKlmChcI7CdaRGh1fXv2+VnB3znAF8AKSw7QiOoU
KLhVebU3UwuPL4WpC8j4eNf+4ZmOHqDDDa3IBeRIBMjIBtbUeDK3tWvXni7Y9X++P+PzQtUlnwry
g8fMu5iMhSJh5RbVOyrXA68zF1TB+CAHAVEspK1GEKVDD8nORuKyIUhkSt2ykE3/gUawNib95AhN
puyMKLAZCLLANPKeY0VqewyYwfCsBzQ5I0iLd3ZbMuirZzsILIU5Zu5LBvaturrqtlOr57ljA2ZO
3J6bJFIqW8moonkEVAHvvJJaTSxCQUfJroWaC3QGJltxMqGo9YBgPpEw03ZsILrRqnT3f7D+X3E/
6ciNdaQYRkUSm+/JgA1xdPI4jOejLeZs3v3HOVMBsBS8BdfdDyJrIK9SSMUNzO/kfcAOmFGHZRo3
lZKusszY5nZt4ITIS9fffpXvrN+ccbvlk4+LI6Uk9A/A614YWo+e8L0I1AK8IWnhOa/IrGCRl8mc
cvNMTQE5QgAfWxjWonDZLuTxSgpTK44unBj8rAJAOAFmknFb3yAC7+90dadZO3s/IQg4PT9tq4CX
VUSY/3crmiiYsSoSoZrrhhZRZh1sSXGZUnAYqTLxFtN/l+iwAspZnf2iNfnNSBgut5G6+xcLpzUR
hfkKrxEIJCcPO7j/jNy25qmdaCm3mYGC4IEyBOY1TItpha3Zt3PBMik9YPrk6P/Frp7OkHlUNFoS
vAHt0J3ztVxM6VmiDZCxwKHolq6mvhteceoshYNSoUL+F2lfm7RT+v0J6FW2wmhcu4xVwKrUkj9p
prYBc6YojLf7fsH2FaciL4XkQzbAvymMDGv8KKXE2WSuJsuVKsSDBPq8Y39pMI7b4wAT/zjp1z/p
wacaioA+Y2yy95un0lZG0W/8D28dRSujdrAiIvPhTR6Y5ENuo45V0Gx6GIMTISZswEuCRDcZ8c+S
G19q2CqP3GU7AgdkCYuX+5wsvkrmE3UjK/JRIVOS9knt7RHl6QSlbYr86FxqJCztS91zz2WbccVO
12kPkoPELJ2kbj7h8BoJTtURmPNBwSWP/hD5Ig4cqGX4cCLDNv3uZSByhT5tdVs7mM6GxxybMLuy
8PO0VbplgF1HmJDgCBN4x3wufOQtfX+4vf/5/c62K9T+I4kFzaJfIGcJyM7HCzSGk+SvgW5wsWC/
xixmwRrwLhAOXlKkGrZ8AgKjlHKVqPEA70VEIMir/xx7M/R1jyEljkMu9zwt5GXfAeuMabcO8n2V
EVy1jY2P8OBVj8nwGNvQ8BP9ZyMnnB4f1Csyrub7B5NEF1Xb8Vb0UHHOu42AYNAP5v40Tfbd7fJi
/2pRq6ZG+4NeK5tCijhfHyaePIXJu2vroGjcIm7fhGKczLRZ3ht8gsnAm6DGrevQQDecnABF1gJd
+/iCwjLyllysBW7Uf4OhxDGamLucHgBfGJeqLpZfg4U2tiHm1f/qiHOrwyOYp37PyytP4qgS8+V9
JFfMo1Vt850OwzbGQaxz6N7q2yETkKctcQ/y2farwHk55QjzMjoxU3hGyrTgdrEWT4MooKKpdUaJ
t7yUkGW6X2leRjwtNamMfah5r+qEy006o/9Fpw7bavhxenfjsf4Ea51UBr6M3i4SlB8ZkBa10Nws
JRIfMDrk1MjsKbU5R6ZpXTBecwhYdYh/569AqU5g/Qs8dmka0DWJrpSZiOO3LjCCE5cQx8jwGJ9V
VUoKgQA85uEomcCZt0aOHPGiVjgaNSoVqyA+Nh2XrF/IiPC+FYLymgm8pUW+NrFtuPcQ8widCJR4
yEa0+++vlpq8Xpjw0tnWi3WQDHsqmenXSyitUoH3q9F3sRyoq/8+fp7A1+W95LM1C2By9lYHSM1r
ke3y3/AlB3wyev0xe3qoJdeXeRxjT4AD9AhHWzOB2NOukFj2HnsjpRVunbu2eBUTJxKYFjYg4RqK
Du25TG49WKVJof1GuL/PDh0ftD0SWG8LvWySqgQI0EZPVvxgbx8OsD33SwuqtllaPmdi2mWNlwJg
LPobZsiLXJzW5w4OZyAnSJrEPTnixfUZeJrG7TGKlU/7Vn92f60GGDLHKGkKrgzYMzcEj53vXw7U
cCUnysePAFNm9tq5OH1a1+FlwArcz8xeel/oYbDkUwB4SYFEUSfCHuK3f6bl81EXbuTFcXrIK7K2
h5KiKkfn72sNyD0t3GRv3B97ygLldCh5EIEj3ct+UAnhwbIp0nQcRyshtk8Ava/um7iJMp0vmHvQ
4DXnS82y495gHxTkJf5KDDMNOVVnlTAkiKpXaYojZ8RKnMPdYtuS3JsSKHzeQ+2DSJvxziBqmwoK
S4XH8ikxcOShCLiRcP4FngqCESvqgVYDdFTWAxFk2oQPR9vAy3KdJXNFFdH4C2A+7QNDa1UgzRv/
MClsTuw/0wVLwhoQ6QFakafXoCoZ22tlspgKnhrQsa1W7AigGzjBA+qQ40JUN2HrITn+s2vMdHWd
+7bxOi2L4wuEx+5u71ljY1pwNV0GTbWKz7qUSKpXdYx5Fs7Qz+or6cmP0hIdDgS+PPjVO80j3SEY
D7mnuec6zjsT5DTtG7XohZ7xAYO2PMeq3dr0nrCa5Sgsy23gf+8/2Wj3a4Xn3fPLZnBfEz3JJChx
fln79CymoPn1k25s8Q12MoxCjQm5tRkfn3zWJvQE6Oc9bY+kHaATi06x91pdw5lFeNlBzyLN44aN
YzAYNPu73SDr9aexOI9k5jBuhFFAs7+QSM9SHEV8ycIcgSwDXst+jBKEztNpzpJHIGlQ174ZND2W
NsjshFAUXG4Bw1C47UUfTnIlmjCr12GZgPsERaFUlScIN4O5cm51ZAEsqdTLmNFCgtK7TQy7ydIW
gKN4KblKrIW2N8UT979Ru1FfSXsefnINH5xFgTCdDRjQLN1/ZkUSICiKkeRjampYnZ6G7X8jNvOZ
+DHlbnZjvu/Of1r/XENrgjdHi7HqvxvLChXuyOuApPzlEzHVTcNnvx8bkW2225qDAbxUKayUSCD0
CUAya128EI6yyq2imiv17BwzjAJCkefI8oyZv4HTt0SdXSH2F6YtetTh7aQ5+LAGrXq9POScF/k+
1I7mXzyxIZNOElzgnVrLdaXnIghJ2XSyDFUqmUgvG95EShtwLcPz/O8SNBSbMKCAE7efLmtjMxc0
9P5cLmMYpPVhVQkapPFgC9s/CMpM/Ss8jn/cIaiar+vM9omxmcquVyJ8+/DklCe8UVLGeH6WruKz
zTRNjI4gYQGNf2vBc12A4/poGPSeYdiMQpdVgbIs7elHeLgDm/NhP66sCVlFGgLeyklAPusrirQ6
292YLl7X2Y6Vy4O/rQMxcHALWy4hkuBReml9qHOdj7PUXQE/wGoGtlIpuhm0B7jfdsCUKzIgdEfG
bj8BQC9nk5RFY18wkhoXItmBbaOkPsY1rAyZL5jM7NlXiU5vWvBU0NhzLz99/riuDN9xw3n/8BPe
TTJkjn/40mDn7dB/atJeJ194Ny+Immc0kNFht0cFi+UihyxNiqOF5TITn/dLKfjcc3/9IwG6QqLE
qGlY3BhPruUecTAz66PCJ4v+o8iUO26pvSz+RbnsXKAmSR6c206uXofR03EkOiJ5TkRcViz1Cbmw
r6HhZaeltmOk5L/w2aBRper2EWqhTPqQmYDpn9e19lYHbEE2h9ACbYRAoookuRj4Ddu9IAl4/S57
tXWlZDwTWA6Z/1QBV2I207zKwh1luxxWJf27YaVKNvb+lRB2G+SelRBPTtorMfoGj/cRDf5b+6S/
/or3t4KJu744A1kyMrjf755nfTc28Oyzkn58g4EH7WOKMo71zEt7exCPndnfTkzfhEJ2VcAr59+X
RromJHy/qSPvYJs/oC/JIJFOpwXGT3+NAsc5Y89pWsDsJxI62P+cLnqoJUDbmK70HdXSHTJ83Ss4
MvXBVoaQHbiUHnJSbwtk4nXGr7kHN3MpetlgN7lh2Yplw+aW9jbqlbXKnO2Swown6xfd1z4HsmKF
W0IBHxNnmYwYy8P1YyHLUok0ONIrgGfLwaLEoWQRczzntPEg5JWyNZEGbjLYCBl9qqFaBlG9lnUv
zeF1BQo0VHzXDExgUu+Jk5ZxvMjtEIXJAkJCS857cXS24TnpzUBtahSWfX1I719H6uRjPXBtv0Vk
j7aZVGI4BkHoJg9WFMgLwUifraUVZzhtRF98+zQU8a/l+z4yxAk50I6P9xjpcZA0mNMqqiBkmhGm
66L84DTZ0Ap/1i68SyuKxKlCSR7kUMv6lIk0b7SKIBiP+4VcEJ+Y+w0yZwYACgp7X1Qp4um4pRHO
XQl7gHGN1rPl3V13H2EOMKErDaZFTfkFWVUTWHyV4nSjMLS/Tg5C1+bETj2Ln+QD6Oi/m3am8wp1
nwPfBdRIQLcGFFhx3IEWtVjIXM7va1uF8O+Kis13l8RGd0tG/RxPjLCwZL53QIq4tbo2prjXrOUg
a4zGGJVGz/ezLStht8tBvhx7AWaf27TplxaQhsLXnXq++h63D8Xr10WdpuMjLAL+oRFHsIWSuFlX
fZlBANX466KDiCGOGaGcJZIDb9ViXQACvKVVMbN2mklgUK1KfAKUbcxmwkiFG+FvJ2q3VDecaZL9
Ccs1i4/u3uYuxqedcoKgYl0d6fNnnm9ose/Mvyib6e6Mc+RqNudBcRbwyi32yIWwi3EGcfawKVnx
xp2KeU3Ajrp5CmnyDR/eHGJfK/3fmStqlrBGkmEppBa+dD4nd+3IrHG3OI4uQ7BQ1Q+tFEsxIJ5g
d2CHqDRCjx556ldgkmOSzhdt0A0JFJElfA+IIieYBxjoHoW7SakybO9zD95ZLPqY0eHRBTqDXC58
M4DjhlEYpWsLql8Bg5e05dGrC61OeG8NBHxYdYeGR8m7PYUOcvqDqtZ+f1KNyleD/TSBIw7EX5JI
9AYCPHjxkX3FxPwpt5fYRSM6SKOOcxl7UEL9GN6cuuNXJSr7t2Eu5X+Okxk/15+o550sIWr4yRgD
Z6T31Ov5/cDmo6BYTCS1y3XPEGZXzeNuAJj6HIH28hQAOknDIfV4hKrpO1yR/g8ENZzMAMEaKDCI
mKDu7D743oM0g757MeT3JLc6MCJv3bOQ8FU1bxMC3KMGEyjouML9EgRPcnBHURjFPNvb/XIlJz0G
rRRzMHs2qaDqnIHu0gUWz+q+8UG0IzLx0UUKIIP+AnbYg0XU/qQ3Uq6r4dLJB15T3ntMkpy5HAlw
nJbfzXYH+DE72UuAThVCj7PvhvUWFWCoKXikdz91HifASV5AzGlSIN/s17a3hB+6Dm2jH5VdNcWl
UA67TWGkCgucpflsScfzuyOB7b7Jq32JEgBIWeu3XtJFE4B48yOjJ0O7j0AQhzkPWvT3oJpmX4Yw
z6s+Z/VKRlSg1vOjgMv+oTjoIKimnKHZKjCKuyUmKpQrFyyUSdKcOaHely3TLM9mOAVuxxf5ZO/C
QeN0yatjV2BP1gECf757rV72/Ybd558Nw52VWSbI3Dh6bg0R4jvAdV4VHV0e8/jpLRRFlHlDPKBu
a5n7kbFueGrocZL5+ClUcHa7b31VcP14Isch6gYgKs/10y326d0oAvQX+zyRZeIXXTRCkBi7ZTnu
Qkj3cZmV3eUoeHydtRp/l7CYHFN5ZRXlPpPQEVZWQfBwv2ffxaqG7fKvLQjHEJk/NNyoiGzAb9Oy
WxbEaS6lY5Dr13NPENw6b+ooaTs8KrVWum+3L58OkNVaKx/NzBmN89aekeNP4oNzQgkPUrYUgEXY
/BmNBO1RQhLmXKiPpOYwWIkCmNwcTcSaqorTMb8jS91k4sOUqqSNso2VK0X7XlvR/8A9kVucUJiD
WiP2G7Tx75mMupg4o7X1/Lhh8W4DjyLKDaZ45Lqb1SPPM8MoJQHAoq6jl+K6CcPJktTEBr9+tQ2c
0w/s5ca8bpY+NR20DI5SbgaxglTbMeLYYpwOBmV8wIpOJhNc7SYSvSYVMOzwlz/CF3IHq8h7YiL3
lYZDw+DIH87KuhCTUaLJMrNGzeaUOS6kymmnY6zJbllPXL1u3P5xDzk0BRairwv6FUW3kZix6aj8
UkV7GWf95YxuzQGmVG9qV+xlGWEpZoUqkrGnkxKlgbiGAjyi6qdjRa3Ss6QnPACpSwdVCyC4q8wH
1imTcC6go/4THfMq2BnbHVYvP+RbaZVfdbfGZqDGDjZUz7/YcjkiOkcpTgBdcx99gEcp9Q3t5G4U
nrBwr5eud9IcoD3WZzZJZIQws57yuvtkYb4hpDVMU/ZoorFTN3QA3TZb3794c/N10CgyhhnuOPAB
hqgWotfxd3gnLMnAHoDXFDwR7PMmTc9zjA6rI7XtUEkFENVZXzIkZ7Y85wHM8RDe6p1Raolvs1mz
QJWUUyP76MrP0q52+rpB0HektimUcMglpwjPmKrYFhmg6wYNoBn0k9Fl9nGi++aQyZK8UzYON1HF
mhUEjxqzpl0eY3c0/10YsS+kgzUKXDUI9Y5DNS+GYHZE/0GnWg4b+dhCaGJnqvSgTEVoUkw2llvr
EATHkWjhCGh5NwO1E9SEknwpHrhd4DNPqqJvJY53DCXiS5sth6XxT4pFUNrmdEMDbprNuwpsszoC
x4sloa+iwxItEr9utQxhnWnACM1Pzwpy7wXrUujY2M4udE+Zyq5aGMtBJcRyA4LN983J0QhwlueD
6y8B1AxQYK4gcYNbSN8C5Rn5dO0qwLAHKb23KZQtwzrG34Fc2w6/aTfPnfZ0YG6liVz4rLXD0E7r
cM2A/hOciKr9oTcvL1s6jNVbhWnHWZTuVNHQzcd6XZxeuL/tOSTY7yZB5LhDABMSYwLejz4FGqh2
aiCPL+g+gnQgxzzjHXHCXtqZFI2hAfEopTeQr87gwxmVhZjoe5lQxcuJR6ehfDclYEUC1Xg4tAa5
ytuPqujRMbHscnCgiiq2u2IrE4xweT8qFpvJi4ZuDpqxhl6h6CsnzLrVloinyZWj+sBidCGfrJXL
E1pM06WMKd9xQuhQ52Az6JXer3Cv9oSUFLPsi0/DFqnrNYQVFlChSjNsQvN0FlwJ+8czuzEpg5MU
wZefjG58K3BAadoHuLfYde0rXNNvc9kxtDSXJofDbN8EnyMbMOnaHFDQyww5cuZtjGvp3ouCvN7S
y0/wguH/NyMHA9MXLu/C0+GVeY9dqJe7OafRpPUZOEwrDiuWcrxMg5hYz4Xr4WEJahOpFu0eLmyl
H+9RUlI+wJMSvgV8RzHygOujF6SJ0Om1EZycGp0cjq0crKfaIxNIppY6AxRYtkRrKJh3gbNYrSFB
m0ZagSJUDAH6K1zKr3rjxouPi0ZuG+bMl+gDIaaUCaLbd4JxP2X//1u6+S/b7irD1EwJhu2jwdJo
EMROsY9fN5iqefLGA9C1NONmQMr0B9FwexdaBGCxSpNgqylZ21Eloebvm+N0dI/sGTv1FfKBb2az
0U5s1rS35l3wcS26fXAwJ7VtRujIrbIrydUv126+cDEwfgaFmpgIO1FHfr92nMFV0XXMk0+yKh9X
ZkbexZPP+zsku5cdgfjsJJ5AmIvU3oZ/DQfRVhfxfW0yL9toujfV1+ao9Kx/KXS0ZD/ReVIMzQ8V
UloVCLxHtgQFjUNMirNYckLKH2Od+N1MWIs/Rcuc1ipwbQgPSWSooeXJMbFueeIWrIENuOUc97Op
wxUeaxxcjQISWYjSCz+cvGpP9wE8U3jJJ9Rr5A7RAxfd5P3guvfF7jEppCexNXnWDpDQu+lWZTKa
s+BkXP+VgCDp1Lc/ZImNAwAX94OTLM2lgd5ZsWCVkJfo7GT0M2LA92C089DaeTKVEly2AHB0pMHy
tLLuSsLLpJ73gd+uxvFDyvzLrhRkpuzvhel/iVzYUcjDx/YwJf/zpmF5GLwddIDnRhXFJ5R406fm
AW3Fw7CqLf01C8o/MC3QuHN2QYgVLE/WTJvRHpjBaQeeLW++EXdR1SAh+h33/fzDH5e2YFMTA2Lv
eVOVjTJDlEh82YcnfEzrovnFe9jIG8MuZIFUKft+5OMiMAGVNOeKFC9mkAj5q6Pi+OwdU7nPVOZ4
a9mUalkkjKd1sHUo0vgwSSRBms5eEVw8hciYQfRJubxq+IwXeXjw8KrWE6/G4YkSKDva7bZubSVw
hbANc+BAzOwHQKC3GDm64uLj8fy2l8vAW5m4YzsCXvtOUJ9YBJkYPxG2jD94iKAq1asgnwWAD1Id
XJStiaxAjcRfKE+OM+1GbmS0TFQoVnsyuCLF5B4kjGg6g6XQmANHKxLuPfP18RVDdokxcUpXuu0K
FAKKTPHH0Dk1menjPHdLAtxkYw+QEpH3710FlYGAXdZIHpjO0nmRONe8og/qxfxG7MQ0DWUa//O0
9FWVhxVvNaNPpu1RyNYl8SXAJ4kSgfzhx5rPTGxpO/mHNSNdJsLJJtgDNMLdsitQ8QzYUXKy1MuE
C+0OqJU/tXgmDxG4f1q8ZB4sPkgX7Z9Q+nO68BziC2RHVgZD9Lm6HkZwVsZyhv7/4q5+QRZbx8//
Nt0i+3Zrv05cW3KAZYPssR4l5T/SwFKOJ2SVsRFMG4z3XANmQO8yy2bjJvKCfFCBBWqNQrvR3Wa2
WnDZcD+gOrSBa9yhasBchEcLsZQkykoQfZTIZ+Pxh6dRqLqi4FXm18HA0jH1OKOV0KqewNlQ0QPl
7HFuU4/xfvuZBNDGuwW8bRH/B1+Uzz2uzR1m3gimnKmD41Q/Bf3ptvI94cmnAoOfyMRMX2NReu+P
Bg7YnMVv/YJZ9JvOd7G+o7w1l3EKzrxOuWB8lPhTFB9vqF2QIcb7AGzGkL9lWQgFo5iDgNsbaMsr
YohpJJ1Rm85btGH/pk7PAs5F59J2pNth5l2YWkAhnBA+kO9sRl2olrgr7nbgVb/ruolN8rY9XgIl
XDI009GKIfagGQvIKrnvKikJSBeuRXYTGtFZmXe95J5VI4X/hFkJj6jVnUGMnLkA6nIqp2cuyVeh
wyERc/xkGZQzaH//Vs1ym0Xpzk4PLv6PghWSEdsJKlybtwOYIQTrnCaxRdKq2gttaUlpf/OYQqXz
qzKnkzeUmh/Ncdjtgxbt0pYdrG+PDVY25d9yxckihBtmG00ObvWfVk7rg1I2Dk/1Q+69niCtEPH8
O3PYEvpSH4WmBRGwDXc/geP1Obj8jy+pEVFlC1sjWyPZTiI6UpA+L0nkxjBqsEWkZm2vS9r83x5q
HQFdx9H5l5a+pLEK4GEWzF7kaSTfzTnrY0MRHQJ8PbkodPnndRlZkYT/kkmb3N81FYAMPzzTIMkt
7tZWUets/ZlnMeeTnKYHY4ErG2lr/ay/Izk0psnlQhsJVdn05ou2MM724qoKa4nWdmaov2OSl0fM
HxL0niUmZplZs0llsZmcPuSXGy8D41jxoriTw5dNxRTMM3yRaifG7B0ugCRd7ZcNEKMkZLO0dUgK
jvwTcFFJWhpt+M4PbOp1E64jDmvYbhiyOMk+fxbTIWvTuGTcU4yQlbVkITRvtMT9Vu0ftqHTqRuN
SzBthao/IlZsRfu3/3gh1BLoKdXBBvdUvNfjvZmGOBUBPZD8H/83dVj0ajyug2DYmqlOfav5ZqLz
I8vGSn34esKFuNyamYQR6Suj8r/eD+JlstkYxgr2dW3b2ykoyI4vwtDSnon3ly0pvWSa4BJVTa4K
wXmaPiirsgpQ1BLzKQI2oHMs2eDW5A4JRTKFzVOWKCmx7G4e2Ac0b2Om2L8lIYppRr+qXvsOVQs0
KQvZ07xHplKipv1NQOQmxheRH0asE9JwOXGI45Vyo5QmbHQFi9G6OZ2zSJTUFVr+h/9v1UrLKsY/
vWOoChSM47BqLxNRDoLITEAqtciJK5Ed/184+X74ARwZbfgfOnDQQkRbSOzaRH5Rj82RQQHUtFnp
m8qkX27f0IviaG8AiEyPFhPcTqYq+zJxwLtssPYXdivfjQtmmzckzYd3AXKFepurjGnEEeW1ssbU
p8zJKEqni1UGHrcMmzXWbo5EegQ9em7daAs723y2P4RwSjMjXO5AkzLT+WiJo+hY1oJfcz5fh7H7
bHtniwv47Hkw/eQs4CxCkYXak6X0rSN8UU9SVLwm59vWaZ871Wa9Y1o4BkDTUy75fEjGmj62Hl3n
kUk/X1KBvrz5bRhdQdENBlq2R/CYUFAovqAqopExchu7GrEvgbY+ZbR9Buh8yiSd7hArs5bfind9
ruOy677KvkOlyk7WAIxZUpsrhwUSduw8tYdn587Su31i/rgLhbI6d3IpmmLfrtIF6jKCUkBSG+Q4
6A/49r4k/GvG/mUU9AlA+DFHHH5aHtB+F1qpnsOv1Wi7CzbyfHzeQ5F3Q7icgFqkQVOZIs9j89YO
7z+6D8EFL1etsYltzAH5bFzSpJvouLuTnMxiNtyABMH3nqIz7lVnXkX5MlCbV0xYFVpxE/HlFB0Y
qKV2AUdErY12nIvXb4cLSQR9rYbnV/N7XebTi6WSxNjM+dTgVG+BezeiyelJu1reKsNh5AyyCWXA
TCaYZAtQQdzMq2fZUe/2fhUlbKjtLxBwBaPuAK/OaSXQTxW6he86yGx9elppD0UmzSVlgA8TaBRj
XmNKTTV3VkSL23zeeGmmZNH97d11g7uYKfDzgA/3+4lDzvDZEWO5rHdkTNtiWPtlGP6q34Va4StX
UuwirC7Hr8PXWbq8zl5tR3V+KTAU6+QPppBSsaDpqTVTjxvfbvCXs8CF3cmx4OVKnstAGMGnmHqY
fSNqpLwSC+Iy3FaWB8rtQPXg94tAmIFmTD5a9thjOTUNgQuOS08D428W9lR0MZYxW9NHG9WQp3XQ
r7Qq+DBIYlOhRYPOXT6krbCKaVZCU1Ql8R434E7uTpw2In3zFlfj4DFocnFYF0Y9FPpkvMml/Zk6
z4VMgyx2jKNo1bkJQvS0StO7IRQOtWEQL5QJiTXtgXVlRM+2MK11Z5uqjQ6FjNDVLZ4VxcU7C1IN
qMwce02QyPKCufuuV1nJPsByuaKPKWbZMqM/XKSD76kUj+8DYu9kw7wJiQnKo836agDIYbFe+F7S
j1Ws3MJo7uxVli7/LQQeqRIOdw==
`protect end_protected
