-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
RlsvfqmOjywYA4+ZYKw+BzQnW/IMAqEmVwRkLLlwOnPCmBmVpkuGGPF9pxnKGpaB
u4ly1qmtm86Vcaj6tEpYS2szn0oNHJk5mTaHmfgYLeXBVcGCgjMZ6Rs0DZJhBpbo
fruvt4ye4z/qhEolX/UJgTjAMoLdYpp+Khavb6AHO4Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 99863)

`protect DATA_BLOCK
mMVQ2LDbXZWxGsHlNtMt9yxq7i4tH0uYL3SDW8UzOj5vom2B0QQ5cT+VEMnSGJZc
tVqP0Dv7B1LZuT6UrIKyB/fX3OOXT7+dw105q44lpOimBt7wuREwAb14fLSj/kbp
2jAJTTupvKDQzIygPwBtUhptxnwo45HgAg/t0T91O8VfKUTNErX4G/9t59zkbAyn
3ZGaq2e4oo0ywvSLhhvPX1Ff4AxecPxyw1NSAJcQKZin8WLBRppvM4eQIvB6KCiV
Wi6Inrq+ybtyiC9KR5wKA7h1ouAYh/bRe1qMBo3LrZN+8lPfmq9QCQJWeMk8i1lp
lLbTa4s2nfsqG8uBnClGjyN2hFttQqxRlLg4qCX174RE0C0bO40wiRDQerzz5OnQ
5EA1pRx2icr/WoYk/8NNQuvw/witNouh1M359cnFdVJR1aY1r9N7TDJUBlRNBeyU
BQyQVXIl7YWHY0FnbIP7hDllaTSIt5tyz9G392b2vW8wEJEVcXPrNaOt00WQQXdp
jkxxHh/96D18wAhqeDt4fX1jq3QHX4/Mt93Pe3bvTmCx5n2zl6etWUCdMWh2kfBi
FRt+6jLVCCRS1G6iANqnyiahggvtzuShHl6NekaJwHnHCZme4G0/deO8x9RnJ6G6
dsPD7LlWhocDERFLAUEc8PQqpcsYdfCDTSPyySDPYyBWuc69RY2NyYRDqtIqv8Di
HeWOmtYZfVeFRttAGkZ2ILkFszMfQtINOlYZBboXC3AaWIkqg8M0YCRl9C8Xdz4L
B0fkhwYsC4BJqT8iVyFDCgF6Ra7LoCw8HaILSu5MTh5RdWPuJ2hvwrOhY+jgGtQT
W69whImz0NGzh4ZfidC7yVGgRfF5l8S297bSyzpLlG2xLjucmeh8mh1UWRCDM8Hr
ATRdpcjR7lVeYO4y9usYi4gbRx2p0NpKzsjFiCV8EuzO5aFX5H2v5Y5rbTJkJKKT
2kGJv4qiOFL4l/17iPWjsxx4smp/pC9w1Gaw3onGhHgByV0HT20KVy/KMUFhQK1i
i5EK82nTu0Y0qvAcACQ81dCXLNUaBKaJzPzDyWH9GAbdxhXh0fZSvKXVuz1ayQag
mRJURV/xX9NBIQwIN0eDWcU90/eSI4mk5rWTSWic9N76Wq/2UN5kE+8uScVIUfXY
LgUEYaagy/3hRq6VvdNeQIx9oA1/qbidpVw24ud7pQaYIUSsQyULSGDvTxRMsFT9
QSzO51FxV7/gPiD9gZnOhkk8/WcSQRdXDnCHDmIQGKd3tI74oFcY75XlJLMglq61
hPtCNBr1A+/8zZx54ZSR8R85MFanJg8++qum0IcujR9knzZZt0bLpIzobJeEkvNk
bYvAkpdcdo2EvXB8iycQkx+d9CFBXMaGxo0aoeDSm3u32q5mgvc85X4ThEfS7D6p
KFjjz0y7t/G1tiPFOWehO8dhDgIRnt1MofMFhUGg8ywiztA6DgAcMHAm3Emg+VH2
VLaV25+YaR3Ei8u/ZRGkLyE9guJBmF5rYue+oYpCT4bX2sFP9keyQY4Wh8zTuLHw
/aPWZ4v7kXQA++qsz++4z2ZG4w58kkKFcZko3lzPOi8rlWUqPPYPfzyF1G6ge/72
fh5em0EoU/C2awfjdHkl+c9apjZZ2vCpNh+8t6SatPbg1JcuOMkxkrB5x1hux4O4
xlN5Jn46TVLz6L1pWE45a5Qo7m3UhN/V8MWdgl6332FXLyqKoRbGKYWn0VRo8Wg6
dJNlCr9LB29YzSAWMZlqgEmJMu/+0FQpMfbnD1UtoYWYmkB1ZbBJS5zCpu1D/9eR
4WzOSs2pLl2Ap1v7+D45zWQz3qLbFBs5ikkUwoDfRilXxqcjCeVkt+ze8+ImlfkH
Ea+F3oTs+XYWCZDEoWhik0avZ1ju5rLaXDpyRQp+Ek5s3zGvjJexl6pW46IkzyMi
/+U2H2+NYJafGjPNx+U7IUV+7k+PlyaiJ+WtcH+cuIsN2qzBmByhomWghxMBtn2y
XzM6VWUZUGHw4Im8lSjIAbnXPUA5llNT2gbAKVjJe4iG2iZNaFCt8/iph3TPUzXj
UdgiGkWm9mWTUHX0mpk99WKHE485lUKwGmlmlDHHNAibZt7s609k+tzaA9X+//aM
JBQt3GqC7UK4XS0EXwMEP5N9uAofOxhozsnb0hNs/Ax+2EQolDbtil/pP6gAdzNC
IBEP7olY479Z6s6lzT2Q8+zJpYVsTXA+/HqZljGt8NKitTlt5hvN62jJbE8Ojz2V
bMtebFLXlYSV2ZODgT6/2I3T8vPZtAgY8ApNrTYjA0H58UIsYTxUWc6yPyEjfGj3
f6nNcKNhXB0X7ngslQoeS8nKF4mqCrmiA6oGs4aCvpZvguT2G9tmL539RtdOWpzT
fPQS6XFwz0FilFE2k0+jipreKRSU/BfsrgMCoqW9pHzRc9vmjgikqsT5wYr4MWyI
irIDvo89jD3dULyB6Kvb+y9nXrBuCNn36u7SXG/6s5jcyrYifF/QBNeqpo+7YboK
KMAz5BOhkGCBkQSpHuvyMMSNTf8jYrlzI32c+7CEibmyfhNzqKDlYGHspwuixKNP
7jS6TdsbJ+Zt0BfCrYQQ7hDstfF5jzFA1M6JI9naEmkbnoIx6CpI6CEatIkCdv0C
RFEvrwooU41LSpEDgXzYLvqCtntyB/ffWF6lXrACyo39lEJsx+FykE3GRuqWuTmK
cOQxQpqRdvQNBdXUO8842P0zjC24g8TqmNsY0JQ1thn9xmDVqLYdqOXuIuoxjqk0
HVYpXqLGMiPpl2/2CWcd5w/ZiEK+Vc92K3TgWvqmgY3mcCgoawbHpljYBWIsUorz
h9BxDwQrMMdomhYPlM/dthQDMkZGqSSlhBTxd02vmVyrUH0sIJoHuxcvtC/epgm3
zS9lds15pjZkibW0i14MJ2u8qluihZ0073WPrm/qWKDrzUuroSViScWfoJhDtSDO
87KmaP6ecBLK608nJqu1EwvkoWnY9gicwu/mOpf5fhAVkOUIytANLR1UuV4Md+2K
QvI80d62k8wnhTxSxwsVDxENvSybdLvJKvNDdlOYtneg4p2P236OBgI8G9AtQo9h
VJ/6tF+mDCQ6HMwgAEaSS8EjKoIZ995O2ayxqV9J+LdqU3mTP8bfL3YfzpxHZ+tU
y1fNBCFGj89wiUwPGdpMaH8k2wcXUKNNUeenp+edRXJ5ix1SdLOg0Wr3t/78vJkP
g1zPQ+R3bxIOOsUTjkhoQ+x7V8LuInZ0jiY10Ci0Enf2DmREzqgxbnhwRulVyqDE
Ek8Axf1nxOR5Jv2GE+QZP09yQkjX1WM/H9lXOuTdOnw63NUiq9wQBjZlyUM/fXgq
aZBqXVGZpTgsEudPVhGkMDrz2rkAHVYWZiZQ0JJ/JJwaD1//zvKGJu2zHkjEt1hj
wEjI5Vcx3SnqcaOBkvOsk+BPWwRXlTXXvV33oyTfkurA48o5LSfrPeFfK0C6bMvM
/TSN9nrOXjDuO7TO8W2gp+ihkEmwurJ+8hFqyIjh/U5oO/LZ3bE6sSPLtdmmkrLV
U+87MXQ2DD0fn5qv5vjwvcK/EeNpRBwO48W8tKKXUMFE1LUKHDQ6B1SV4rgZmlwE
IgtJW0kJW85s97eb4ZMgghHIN4XB2eRE41TuddAKAjUSUT/StiETbD40SyRwqK+X
AzFDa5uuOroMSjtBK2nJsd397HmimOFytlmjIli/pFSYBOoEeBxIz38HR3yXWuCj
8hW233syL7UlYnoZybB5t31rwlrBMpQZ12bw3Mmg5IeTPwiZ7/ameW0sSGVyEk6c
XcGIU5zN/N3VUITbV/JWuB4zrKNcr13j0P9Lwb38hAOD0aCmQ3565voy0CHO6CZY
Y/6CfB/u7RqbhqTfCCdjr8iYdP4fu4PiS6/cE8a6J//b/vqbk3gLaRWLZN/2lXhQ
Qvbh64Cr6DDkVG+/BYeCbee7blmC2t8qzn6XEdpGKxlraoDfZhifVuQp0SxiPJFP
4mZRcX60rUqBdAVD4GtyJZk9scy/i9L11QJBJCGcl/ZtW38zNh5pORXQnvhtSi1o
wwk29IJvvfBnAmtk2vAWL53WJUUUIx7UTyZS0LgN4sJJ5If8WNkR98rVjqqbyRPh
8+ozMXzInXibkwuRdZIYiTTxcJf8oFEzTvVYwe4xV8rdo5N/y1HC4ua6pjk5xNUz
6gogxW+EczM/2WuS3ZuVCJ+8boKpizbTHCzl8VmcT2A0uJxgQFc+MuCxcvTIXq/Y
c1/cwM79pCC5es7VGI/V8TTxqAhC4DA0ipQn4nbspPXS3XY7ZbQihdfe4rFjM7QU
vMw6jhR1Yae5aW49jvAS6peewDXsGNxoQs0hQ50cJOaPW65I4SxSWc4nkBsUtBR9
WRCoSFc7NCtU2AuMQl2TIX+f9WWosvhtK/Q5WhtH7nzQmHkatuZwMC4c/4SOMt3a
frtEc65Bn6wBq+1L0i/ZrQWbr+YILz5rAxtAHX4OkIpBRSiCpNRjhrJ4n0EDrGMj
F9BeEkGmdHBQoWIWHIUlQaz8c0I9JzrpXSwJmHndPj1NxF7k7IijFduzN3ST+xaE
R6BS/MRAsLqhWzjFiE1n6sBw1etMyryw68BsGP6N+vOcVwFEkctD4mx4/jNVR4PV
RtyEONdlsKIfHJkLD/gOxBIlwt7oLvr19By4HoxOqU/47a876eYz8PpYt+G8tN2Y
F5nzqFsMsnzRuFkadA+HPB/0cw4zvcb/F9dIxAX6sbKAyPZPvsAZImghk6p+HdGy
nunLfs4nzlMCxePOvCfIuGYQ3Cfb3+MNM3tFMiNg5HfL2QuTosF7LSONdfKrURXC
/6URruN16a/obJ7WLBCfCCFPCp4ic3ESEJD7O0tvD6fd+Mt1CmHM/7DKBCrS/lWv
q+b2jim5gXv1pL+mGbk/VzqDHknnXQUGvvwCS3Py3O6jCRD/KIUODdd2vR72qGsZ
0VYTaX+AAcilbrVY+0j1DtclGklk9i4BkmPz4fTtSlNKw0Yyjzk09C4Yjd29BxIw
0P5AxXwSdrUnT5u+y/7rsS4ftAdLJJRgAIkun+3hZmQ5OqH4vzazKY37m5JQrwQ1
abi6uRqDx/rWH6UWEXsgBHPji272Ffb0rF2Kx3JgcsJa82uI4616qH/p5FQaUz+R
8Wi6/Z7g9PbqqYzr/Ip99vaBRuo0CKGrJeVUozaNHN8z/DvxfvDtPXhe3IUMYMAI
Uxq+6rFSA7ifC+TYN0H3eGniv/G+DXE0FTmL9nknVoXXUGcK4BgLWfV7BuRe5huq
WfT3TXdfTquhTa0H29i+iLqh3gjvZ7PcidjqYmqvZxPupgnPUV4YfSMCtsx+JViZ
eWLDcBc/L8ovtlg5n2m7dtBtQjrBeJifKucNchuyBSOVfAJK1AXknxg+7IrUZmbd
wClaQSkxW1UAxFlA0KzAr/MGU5QVtIG9Q7ga9vyraMcy17WuVMTtM/jkOo3mO9v2
LqyXvpJckhMdcqkntlp3md9XNrmsZWR2U+SMmrxlMhZ27xLAk8cl1uDX8UEujq7s
avjNWxzrPrsUfnNn4lOh+oEEnf8NZM0EhMXAOVYAXCvUK/bYjDG9tFoEb+g39cHw
yk/DuFeIgJ1YW2wp6bSVFoFIkWbckkBq1RUXWMhXe1A3AhqHb1pTzobqaTM7YIsJ
EDVl43HUdbgowDccflJLbowwZ8MJOlk3nkq7vdt+roQ+1U26wsNJMUF2Bko3ShLk
EhRBkadKxeDW/so97cIV9eqnKI6oFBzZ0jNz8P98cazarrPTx0vJ9UOvkmX/wPli
wdGpRz2tQKhc8gU+srCJrNoU02uwlFFOsD6dh2kfqztciI5NPjRaAdD4ZYlM9/c4
CAhRjC/hBfZ/A0yg9S33d871GWB2sgqmDjG3rfRjmiRg52hxsiixFlAcYHZjiu1V
PejRLq5kGtCD5xYz/Cx2ozF5RGM4vYKJmg4pJiP0rmioeGBFVXTfkBDvcqO1+AoO
OASvCA/1GL/NR6dbjtrl4MNf4mAccs0wkS9NzgfGQkqqewNgyQt3KsQTjJwgCsXn
eZIb4H4JUFq9EPmOBUltmVNNjZwnPpF34BTyZzmQGjnaUHMsbzSlCQbULuh9s1dj
w65k43+TgSlj8t8ePxQmAuqHldSoV8nSUzNwb8KmffYZoM/KaU0Y5+aOXkePkssQ
xqfxbZnoTFDAMtdSZkj23VWRmm4yI426Jcl8pO+WdhSDqqyUSUNbYTRkC+O4xuad
4EIHnYWYgBkctGHk00lP8UxgLomX4lWL5t1QIRjProIQaMYSrXaZ3XB60GkOo77j
SVe924TJIV+ApoX3fjieVOktpFfe8y5rtnecZZCvcIg3eWG1KxlGY4XIv2m632L3
YxJDJFNCSIjpVWos0bye5VUFg53rs/DeIwPvdLlJWmEa0KKV+euDmr6b/1Q0bsrm
yL/yRNrFDklZqNZGkv6tOw2n95XkGswgbI+zn8ZikM1tgsa/44HBkyFOBDjFZ+Wf
Z2pMMSdcRiO/qh5VCWdhSusAN07rG25pUTjnQMA4tq40/ao7UWdZ98y/rAQz2Zxe
wNxKfVe0rHEFUpnU7kLkCBe8dONoxNYRaBwn6ep36u4332Ttfakv8/pFd5HGA4wY
w8jaO6nMIl09466dbo7ZwkjgotjUUBpDx/YMNGUR73VNSkB35l7yBqVmypqxVeAz
AhcFSKkiyBPpK7GT6kKDqWX8P2Xjft1lvHKb0ut4r1/2qjaTtqY8uHMDSXyBTSsc
DXexiUswEmRLkqmsvKoH07pFJ85S90fWCl/37kWzHkSMoWqkQvwGMzhW9TGFidKV
ItGbzrLOuZVh59gd9HDx840DeY5edRBZxGW8Sa4m4hANiLhtqtKPrH/KKNnKY+Ma
xTPIag32GKJI/DGzYoC8UALKUqHbexr3ZfXb6vVl1xcoqyG7JzrOUJLgAoIRkZ+l
+ra7aAI7AjSfxUTvMhU8m3rpl10Y1b8E4O2mdYDMcGv6qafDfAHPG89OKnvsC7ND
1jx1phlxAWR67MO3iqIP3pW0mhz4Jgjz/+mVdk88VYehApvX73PMrFBohjDkH1Yv
ymuk+XaNuzr4Ax/Gr17THuNVwzmgJWC/ZQZmjkpV2k8OVIn32LYiirZxwweajWev
zizTVnE/PoYkF61P+neC+wvqG4UvE6dCMCgs8WAYWT17wPH8YqXMNAwsa0c+YDqF
WpN30JZa8YLZ8i1qUEd77vtnENUwasxihxG52h2jAMK/Gvzsbgfdr7/g/YdCdAED
Teq0+wYNozLfifUxoo7ixw/7Wu4bucQ3CSQ5+4SQLvTNRSdfBW4eZKcM7PYSOvVx
GVnkn4G/e61qyEVzE7GPP4/bKw0KtxjrUv5Tj+MJvgyerY725D6C155nuQQLwBA2
RofEVr/qzk4SiTWJjYckJGl3Ml9AdwGy7ibDc3SdzTNXjLpTiST1u4HBMSlDnGyI
F/YT8LMG3QqvgGS/zgU/Nqps4z8I3y1wfilgGWc8I3bxJ7WkiG73hiEwKqA2W0G9
Dbv3O4RPzNLtGpSrxZ4FkHzlMfeCTLQkeS+lGc4asOeGM+/GU1b5Jj5h5DOq81TF
RJMTUhxmOg7U7yYS8T4vQbw7D9lJogBmQ1CngBqiyKvadpzrZMbpqny9pXPeEaKO
wGeYKUYpAIx5n2eiL3QYh7upBS/PvZtc2eqTtX6TYqLplq5mNoYpr4jlh9GX05gh
UWnrtt9Yo4KgxEK6G9nv5kXJZIdlNsZL+Jbv9pzE3kFMVYiBnCQEFi6SVbk2RcJ6
h5HY0FReF2/y4Ox9buFNxRTlwzQc3saVZO0PAESo4xwTZMDgVPjxEbLUr61bwMwd
kE2L412cNSCGCCxjgnNvbHpXw1LwVmUk4Dh6kk/K9l/bESFceYBLU5VVozyUsnk5
q7yyQn62G3JUwHbjji4r+b9Iv786st+rW6ad4OtwZgcFtxOT+fUZrxlwekIPUb4C
EJQUb10Z6I26cu9Cvdq1ZMeCb6KDkie2UHNoyX6frIjE0dI+LEXrS/0xLBcZFH0f
xeXDZ+/tMEJ2X9dMpYCGibfygZWoZTuvFDdJjrs0lS2F0VMsZX0rn+ENIHHOfv/N
7UfCergGEtREZdutQuxA7v1YQhgdA0xd/hrPF7/p/AZJeuQ2fo19cnuzOdgvrGmi
KqN39CDblfmVuiNXTN2GIE0qHc32VZmK75YtBpuzCefobypQ+xeQtA+ENM/Nksut
XOt4aGS3wDkh1CKXxKh7Mzcmn5OEBNzbqY8eO9YACaQp8/xKYF8iSiYvpfbm4Kz5
MBja4q8A7eMK9JHZ6jwrvEcs9TFvEo1rZRZp44o2nkg4hXMDCHn3bXWE6zv5Aor6
6HXZyjlr0qtGmdhpfKp2ZC9Sr4wRM6jehQvu55i/NdYN2t6JVxWZEC81pFLc5iq5
yDoWl4Lh6Akt+xUxcCSLzGsv/bFWJXhyu2Vs1uttNsXCW5YiRXfLhdyoyZqINCRH
/RGh3DZf+7bvRCUT4n/8xfps6sk4uL6H9ywlTx0kR+rYe746mGdA4J7E39fFVFBb
lfVv6CH3gC8UFMZ1msRRz4XXikrS1QsSPDgKKLoVVzCb19Vbn7Ovlkd4FUb2W6mm
zdQ65IP0BkwVrUoJZv1UdvNmYfje7xAohtiAkq+o/qwIinjuMSXgsfZ2VtIpEmN1
9buyzEFFtQcn23DeYbw2br2qYWOZigfmF2WIiKTanlCDGIWKvhdY8YpM8HZv23y/
mrTHQZlJisX2QXiugY433+Le5QfDP2PFqnoUGb8p3O15JrnREwOeWO4q0YgeP64q
ifo2uVIoaYE8Bnf8FrGP86NTx3cNSKz9rxJB9KGDBSVgeBMCBNeZ02FB95OxyHIo
J9m77ViihzLmsHWpujznVhRGnH0ATJ/7d7P04ftXfb1hBpPklHrlu2aIqSMx577v
Qat+7mmEwVNebUs0iHMrhWsBqVLpl270hZFj9CkToqxdXC/twFMnBKUEsABVmP/2
0ZNPfCfVmOS6jHZPawh8AlNEt8jbu8A8Oi/QSQRebFADNMblbC/EjYyvgm9JmsEk
QvJl9ppKfTYbcxz3LabNuAAROAgDvU3Ex94SGQ7nVXMl4HJj2HFhSNBOJrHpHDLa
kwy6gHVSTYy9/aVscCUvSOjoG90WzAGjPRU7Jyjxr+A4qLFDyTvJhImH0X7DfYlk
b5x/1hTcDvbypx0UBEn09pdQwF4lyB14naNpHUzbwzGQxQUOL4Ume2K856itbxay
5yPd+xYx4v7tmCiQtpmJfcGR2QDORlxZRbEHyvnqijWMGaLad6qX5gLhm/e0dhzM
2MY9Tk8cLVU3MQhoHtvrcVXPO0Z2cSnz5Aw36CLjkYV6E2M6dGh/0wQbC1y74ojp
aLtxF95kgw1ZVDINi02Lo3QcROnTkfNsMw1MjRmNKexmohYvv1rHpesL43dIgJuA
2C2EFTOU0DeaBmNxVLCzqZ4H8NjZptdpTzDt7iE93N93nQTplxCH8wHIiqYY4A/J
Osmae4lzu8VNq610i+WP3vRHuyAfyQIkTT0yuJzammGMDJpvMGbSkQZpH/l5a8Qx
vgCEvS9e51uW6cMuFRUd3nMvCTElxSu1e7uPhaqZ8VKNDqno7GmkiWm2BLHx9awr
m27nG74wb0jEMrkQFxkhK34lLlfplyX8Gr0GDRjxjd+8zvjzmYs/hJmYfUaUSi2/
7vwI+a75piMUXgj/E1u+GEMdKPn3fNYUOGrrO117D8TfpElt69DDYdWb7clwRY0T
VGl+Myg+78V/ZcprY7x2Y6xh1bCfWBNPrVu9xfh+Q7FoqPwhqAO0zJgQJ4/3FsZd
aq2LDq818Ea2Y/AdLsVYe+9YMc3bzc8eoJa2xjFJM/QUy4FsZCJRCkGg2BeN1q2N
tdJQNIsUK7xFD7EPv7t9ZYhWieSWIsIWGY3n/salSEtRgtI/hlPWVNpaPJqVsznD
Q5GvOSWafpCeMZhPCqyyWeBHksD8HIBC5sYjtlUk68uLuJv6RIezKYza05YhdBkU
wjZYKsLF7yoxvmIA15Gr4grxsCqA873pmSayLi5VHsfDjTqDx2iH9u1vu12/FmwH
O+XvITstegSaXrYUoK0up2G4Yv2RQSd73fTgD0Zoofi2kzuze5M63Cluq81jOaBu
pLvnfc5sQDrc85awUZxS9SWbNdk8zpKPi+9axVwfNQjjaeJzj1LhsvlSAiwClMBD
AENDkeZz24RoY59GFa1Gk+QOeaXsRKl7OkPhy+HplLaTD+N8dskjDm/L8GVXCU35
JHg+iLecn/TwtNMx6IuznMkgVPovW+IQe3pxyogEKKuAr75lFLPr2XpCCrrwfs+e
HK5lY6BhPmJwg+Rc8eThiRYrXluYjvHjHj2McvkJCOqH4qqjtrwm0FS5f6gJRSA3
U7kpSieddiaGqho5CFE242e05vFQBra1XKte7ZqDaheHlBO/Cv2dZji1Y7EmD43J
ARQK6j6ZG5sl6K0NxUlFhxwCkG43ureK1Kgbh0hLMtanvCvEMXXF/STYnGo0Q1bt
0PbhWSN8zjSRWJal59m0x9sQfm5p65lYH5RKrhY8Ack0aYu3aZp1TETcSDPoucox
Z00w55kUyb3MM3KcO7vZfjRSarlI4cu6Ohk+xOQucygJHWe56xMw5Fq7b911OQl2
F/RCSwHmtdxPTp9mrX41OT7xn9yR+shc92Yh8QskMpT/3f4m8tSg+3dnayKBps5n
Pq2qpmIMd6FR7YCRC5bGxf9Vq0naLNploGKOFeOpDQSIz+dO73GkPXbSwrTYYw/x
dgaEj0rrq9SIQHV7uMO3y/yDPm/GVZkfksZ99tceG+t/JVjrfNSNcRjm2jDo2+ef
p1pAz0raKLBcDjjWf7HCot14YYZ8302S4TBV/u5EY0eXIXBrc/dC9ouwomIkT5gN
0HWeAfMOVCKQ3sGebLWcA2UNWUrgLNgl1Ro06eBd1GpQ0hL42F/zg+tjie0XouPR
5JeWWG0elNKCWLyASozO56U/EgjRAanpLCYZ3YvkohGkpyxRTUc90zGXH3k68gP5
rCQZxNCjzocsspL6V71l0yVUlUu5ItA4fPEJ9L/ycZlWH0WCPas4XMRbWdJgrj5e
rK4jYkXB0BPJqwtSg955e5NNQwlaoDJSSrpcD5JMtsygE594OryBJMyOhsMthd0r
C+2Wl4uCP0ZKW+C4LJLu0NxPNtURr9MYO6lkniNooJCS9KQbKUfyIN9cuE9ZiRwm
W/tKozyCBsTyIdNtNjqCgDhX+s77EgZgkZdMt68ZF3RkTiuXmmYD4wG+Fbm8L7Ln
kx77k26Znqz9DpRLxov5vcAMug3TreL+4aNxFgZRaJtM5Qri4Eti7PxeSdn0ewkZ
tPgRTsSn8vFQNOJk1P0LmbAJFGFxeYvR5wWM437BPqCe7YQw7tPSVzkBIFbWjrAU
oPBXEL4igg6o8Dw6mi9avDrqQuBVGQZwIIWzQzx9xZYfhfgSv4y2Cxf64nr3XwUJ
Rys0+niTpeRii2WyMBGQSBQM6uf97SURiyc1yduDfPz9rv+jtc1z7Ol0HoM6N+qv
KaJchC8zlrSin1yb5KiJFECNMNbnBp5+htOS17hArgq5R4Jx8jr41d8O6NCU4hZe
UlbxzPmUOuVnGxleo5ZoCG2Rzz4PxeYyk4U1JI51tWsP1dY62VXR7B50SUxM07jB
DbhEzlIWcGZeG3/onaCRu1G8mS0EKhVhuwx7yNYTXGjwqMKsYrXx9zsYA6/c5hxO
F80sDBuYvV48+4h31ijA16OMmxMMvFOaWfT0s+l9uZqyuqmtiIIwHfimpBPJOTlF
z3BDI0J4BqkdrvK7nJG96ZUzCf7OFt098L2OnLHlZks1SWrS5lPTiNO5B0DC9+VW
TDLHTfpvyXzfmQjJ8HtXiMe+qN3UpiQHcNHsxrMQe0Qc8+31mhXmPo/H6QBzYDAh
GZ7Vb0aGHTdPMaQ9lFd8LIn9Ur+K5ud4O5PgV0xe/UqcSOTWjaYTqExla8q66ufN
L9nJJXC5tCQuS9oAFZHJmfmNqHxFLN/pOAAn2Cj8pjEju0CaMnvVl5dwiZGTQPVf
UssC4MIwyqjs9W/Gbn681eMltSXnP6cu1Itoc9PxNIluYQ+sFiokx0Jr85CTLjZl
ofJlaJ2USLE4GxCtu5MPpkvFtEWOk8J3JV1k2yfLCbzgA19XEiz8QrYqjTzgJyeS
tsTJaGykqg+DmYdBXzvY+QpzmTrGny9q+5FA8xnh4Up85DQRxtGqLxmq91Y1Mpw4
BQIrnZNipB/xnT6cFCndYKGeNWYb1osrxJTR2qzU9HZTG5/bqkRhWJ78ZdhQDnqc
fBAMge0bI48D8K+tab5pbdLivpQIl1EyYPsqXHZ2wrm1tUuTfyWtXFkLtfcAe3fd
8dgdIClyBClRodw3dYGBeRlRhCjPyyO2nB9N6y7VPe8fxHW4dyn7cXY/2SwDjBnG
wyAS11X4A2qNyoLEzqjHVPRp9ZqTM7ExCqKXHEItdE1iOJIeq15LXexnU7+UHWeY
HjsZCIxjFIkR9hCRIZuohca6lbtBmPm4Tp8QXmhE4aAtJJoT1dHjVrsBEnrfPxSz
bzvyZE4VROfbEI8w86uvuYA/pNSa5N6Qfru1XGKFqoizEp1CRoV6ZX9Bw4x2CZGj
fMNo7TOWb5+OdQi2i+0eibZzYIFaF6YAAVdjvQEUpsA+r0njhduj1aGpnPUG9KyS
Pdz3KX+GtlZc5rK4QnqzwGZY49HX8IiYrQzdfjOC+KeO8ewfshDyuRmXdR59NDAa
IoN/0MGv1d96tSiWFCt6vTA7Fmi+wH5+SxUHiRvW2Y+KxG3wnv3N5TkjOz8/dSO+
MnUGcAIDxSqnoAj8Nsaq+0F5FaVjhuM3IaU6dJnkXrLJBrQmK+8WLAA2zPmGdWG5
hubxB8yNEcNRCXBXjugQEaTJijhzyjpoAVI0IyDhbasOlJ9FbPxIrxbedFKQae0B
YbqP6ah4J/CN0/aetzyuCtXvsRrsiEybWuXQH2/cHl5TxKKuIpU2+huhh5N4qCjm
r6eFja/8fTb3pA5b0ytUNfR/BYy7syZJOzDAx90Jk59zUzzwTvGSDcZc29dk0AKw
vMs4s/VyVRsRijnRQD/T3hRg0VjIkn/jPz1vT3qZ6gvkEGKQw3RR/ciOBzuo0qNA
MrRFZlcbDFhlH1nLVu3WEzMaCscSXL/Itea4vTnPzOt4VvNPXex9+zeu0Y8GbwUj
0vznVgtRgaytzTEL8UgwbY8JfVRdu34WvNFar8yFgqaDV6jjv5sRNVbB86AUjSI7
mSxHv/zQk8Z7LQO7SPrgLzDwixUnSC/ErTWQKsj9VZDg4tlzHDklGQ3ZmhSjvsIK
GVbPJDGviiRgmBH88ww/7Fc8tQXhtKPXZj5g7gaVHtkTiIC1Z3oYQwfk1Mg3LF0Z
6CJLzrT6C0R/LKjkbR2uS8Qgtrm+H+7RNaS13UyHU4cqQi9CuA6GaYZW/6MyxaiC
zbZmimhTS9rup1o+tLS2k+38RpMkyaxHdN1aRT47KwV8B8W89iMocV5uNudNLU4o
n/cUwv7tXxQUwhKG6hmO9778jwmG0Hbz6T7Z20Jkf9HFpB5wfJd/KR8jv5NwJmpK
bTb4oIbi4vgb6xkNMAJ3pDFcAyBUI2lgp1phsBRkHkwPxlPqPVrCJKo878UYHhZC
PKYYo9Ch28JJbkDVm1kkY6WtCIZ5aytXlIPcXK5YsO5btqxhXN2hTxfQsf6AuDZZ
8+vHF9gGBzQljl7I4aNPgsi1n6E2/HntqbNV+hlcZJrlsEyMQQFRyReZ2EPQO1to
seuMNS45XShPaCrHRRdtUhUkmjDAqhDOHr/3d56OG8CipcHPcWwjoVhbTnAFzWbO
Mtysp8qeOBoUaaeJdMWVMLK0EOLksKC3Swmv+y2udI6Tb0G7+A61Vtp105wA+kGW
oUXUtP3Y4VSnFIlc6XHrGFyGhcAgpZXlvZn+sxT2PabHw7kgaCHwWWXYCSULrNdV
r+L0ciAhGuqw2nwYebKZ7OptbVdDQHWz25REZgLOxBN+L6EJKbM7FbGmDXWnCNGt
J4+1n0edDE+7Jzsfs3n3H7HGxMtgk6SYWN99C1N8yfIF3b/hzkC3IRDDdP2hV0Og
7q2zaXJRCktQvdMK4bGTPI+JX7rjCDoOQHAnuR218h0AISObEQMTAWzZ5kqKeBkX
6KtFkYcr9MUS1A1hKqGlQKomTqpYQOvXHJpKHGUTRTL9H0/roKG9Qxz+AaGq5Qa5
Ytr0OVV0drYEEZB01Etj+PVeJUx5uJI99bYt4fQ3mwe3ljPBO7cW0ZUUaxSPusgC
O4Y5ugDEqVRH7wNTBKhKxL1o2EzWa6dMGTfGnjomswfrbyQvBqT6eNeGuY1XFphN
yK3Af2emNSbJwXfGsrXcesEhdeOFS8SHV/iYPADpLXF3VPdjfx6uUPjg+0YCIyXz
x9PqwypRMqOnywoocRAA9J06QADf1abe8Fy5ByKNp3NubJxVk5cuZGyoKu/QsZel
l5hyqV0dty/CbQOXAQHdt4Lt5SR6IZl3uJD4K0PeOq7aL1vTKt2tZRmRmCKxZoxp
t5EFMssh4qKeNCmwz5llR1o1ua8PArxuI3D/rcKhhwRkd+zgpnnMYHAHEBOH3w1v
uNjhO41c9GVpuQJ77MoGeGYz8UA7KrUyK6lkDk3EvgO8KpJD95hCVYdV6vrx+GMo
12IPSfVEtMmSUoDLteW+uI19CSXG2jrumc/N1L+cg5aoHho/jH5wuy5W3FacvoyI
rv8T1cldO0n7M6CFTCrW7uY6laWv9N1kR5F0fYCmhs1CZWGIHnIPgTuYa66hbKsl
8Augu+4gT0MdgcOx8uIB/3hrbMM+I1zdRryymBD+GIUCBkUj5yJItiZUZ4nMbxhw
gLV6yHVXsNqnLmQperlYlgTWwjaHDmcdMts7S52OykboNMGdnfoMuDodm4E5uGru
3zXj4h2Gnm7jSPxMBn+N8gPVmfOIQ9Sql+X7MFoxah3vKhjRoY287uEfxD3xlip+
Gr5N+JRnE9XTkad05syuHGrPPGpL+U+9GFPxq2mkme5fnje9J06KtsWwrb5Mh1Ly
kEODIbopyjsMhhngMRqeKB0jkxr3UBL1htZLWeBoC8AlKs6vjNtH7UwnS5/cx1al
B+GXQvCMimL8lG0GI5w4fQxzkcpH31GEo7aBrCi25k6bvLJX5WE2iBTuIIwdUxcG
ibfPbk8o2y4Lq7hElE7HrcO+c2Z7gnBi63GyzA4hrGbuvpC1beMFe9DRe5+wEBhi
+BxbRB3f+FLbo/BKwPGrSyIxD+KY88+n4cAnaaP+B5ujDzNMxJYPwYuE9zrwH/jB
M7TZNQQl6wfE+0CnEqwfRff1DDHZvMOEoOQOSfb9CoGQUBjNruGlkovaXNj76TUH
2pjRg8qAefydzJ9Ygq4cWs0snmTMiARTR92HM3dFXeHES/Jjmvu+x1Is7p6UBgg1
V6+gvRmGhQYYCOoYMSTfpJ6lO9zMF6NPcwFzBEtBAC5m/RrcelTDPV8zU0Stcceb
51wPzgqJiDSJ8PMpkjcacE3XpoKcJWN/RQU1TDFYn2KyNy2J47ec6GjiYhuZHVph
0H/uo4Mey4jIUvRjbfm5CtVQ9fpMet+GvQon1Mk2JERepORZC/5I1AkBiRLvPbOr
y8NSkcUSOIB1VBawksfxb8XgNPllmzlYY08LcZQe2IYZUSf6BsBBW6bDzUFlozHu
a34RLZtY7vXtkrp6UGOylDCKrIA33GeHgzpRKTsssPR+aw7vY7yl07PzlvObxg4t
Z4ZaQsAorXhX1SQvReqQUtO3SjfNLIJsMeTuyOUP2ePvOYewvKfyYRpdDQpmaq2u
tSfz7YnAfUx0XphBRuBezDtdEEFnMv4ErQp6/JPrS1vQS+bFbkKRfukpCRbzpHr/
kQ7rg90fhrReUjJsyyimSs/sacN08mEVR6B9LJYR0qgsUfpySi7F20k+APVswCGt
hM2WR7GP8WsO2+1DyC3M0HkhqGXOm8WlgGDV5gakYRv0mrZw2J6eBu83uaVulbiS
jJk7uymFb2JGiS2qv06U6MVqFGP9br8wlWFmzO8h/+2xXCgpC7xCdkBvZ2NI5EgE
6fbB9OhBdjWZWQCkAcLfjpwSKrBRrS4jmPIo81kFvws9t+6xyUr3lNN0+CRUFU1k
YjqN6LE1Ykd2zi9GYLP9jrXVz4FU9JOS0Sstc70Jjs5S5lX7FONl5OE2Ea64o5Fy
OfO7DzR6crfZkA40GE0RLKbpUH4I58yDOOR6v2mbtARpbhsDeRfIvILMt0Va7YLC
5NQ7m+zO/2wVj1vA3BsakWFQJ+WE4NlFIvy+0CLTAWvvfhFRsYQBWMOOKqxk2Tav
l26SBROetkvrDbDCj85IR0nvBRpZRgTbFeOT0nTaLHKXYX93mdz7P7mV2l7KH+AT
LgjnayNffV8LjwP753aXKSw4a151VJOZa7S6Op+SClc4i5MrawQ8O772RvMZihRo
oSswCsgLWSEUQybNcXcCYPf6utv4Zix3w8M5U7LYAjZIupTMUsBMkRGg0t2V2awf
pAarYah7/GJvWoNVklH26XuV8BEbM4gAAqSJYAFLK7h5J84rcICSdaIRPglnESG8
T5CHjaPVf81N6d0PAyvyc2dTCZV4t6r+Utpax5x6bAY70maOYyXvKzX/j4PWEc7p
pNzk5g99IvzvUErfUBNpepfKPFscktxSifQlONRKADjLZ7qfvBw9UMhcelaQb0qN
GL3XZKXE6+dU2XyOIcGTGYVy+vhYYG16a0947Z9EBYW2gKndIpVZUFDnCwlrQXxt
OQc9bdo3WgKnrihkUViNF0xlehXXpMGpprFslY+5qjDvixB5G1sx8PhnnDDGaCXN
a5p1NepfPsXRP5Yyok5lvR+UsbaqF+cX0tGspJPXUq3J5FHQW1dNtHGTpoQ9ZOhu
GhZ+u4zDpVH9eyJVhpndY+lKunQEDe47BzOFdJodJUWYBSAix7DKSxPPmTu1VJeA
BtGl089N6GuH0zATzh7mqmX+EpEcxAlgMSPxTJ+Bhy0AcIT2TLOHZ/cc0DCTWFpA
X7pqghaRosEKFNtDvKSP1lbVVBWpes3h84yBNJMMi56e+BKchGdd13IlZ5YiVhPn
wTkdGI0TIwBckzbPe4gYrtNRphWc1yHxKUgWt7o9cXwb+ATKUgDQ8385QcQCng+B
VcmHUQ52U7hQe1lu9d+7z5FKqpoY4zPiEAQmnwwwH4Ymt4fBIUaQ+8StecVTEBrX
Xb0CS7Fult9q8ueSju7+4L6Gtcakub/gm20Vkl89xvX4LqD8cMGZdn+55wV/6QBb
oPU89o0n/Nraxl8GdMCMPi1wxdp1gT98oKLqlEqXvwxiWT/AcFvh4ilN2dknk22L
MtFN8tYmzSyyBv6X4TR6+peXTeg8RwdFXcsnRJ+KZj8RUSxnqicZtCKICqijd52E
4VAqVzzUtqQVsnt3Yanhm9kWKpexVajmBvK33PJ1YhlTojG2WU06miDUNgZKsxsy
a3t0kqbRM2+bnORwWbEcDD6dWKLMLTaijYjKlomjhAtuM9it4drzIukQsBLcK1MH
dRSHf5+7yn26XtOU9r8Fp1Sz9vxi59e1H7NUDK2SKiEG/LNZRTMvMZ/CRoA6tIVJ
dQ8aFzhxnD6wL4r+px+kSnNeQfcGfKtb/8d8ZYtz+keTmrxfwNMaDDmS3K099+u9
cRf4FuotCAFVbQFbwO5VHDa9Q8OcLXgMxG2MQX3/VBPsgpExJoHvgTaH70KMIPxD
//RV2nXqOL0FfD8Scq1wOVG87mf9AfwWJgWd62NHlv/Yue6dBv3ky3TOIvJKPnLz
Ow3w9CdDUZ1sqISexnxO7OohR/Iyl/ydStPMCWSARjLEEfRFBEFCESJialVyo14d
445bHw3FNVvO1o3aK0uSt3fnFzeRmqdivExRiSkp4bTJpwY/G/l06FfMJSx2iZBX
0kHa0nrOoQD8z6YPtLS5qyDslU7wwB0HC/5QyiKBVONkscwl2uYFPueEmR1MJQ9T
OvFSvgbKYWIhKu+Fmh1KHy8I2w1QQu4wnHgPCcIShRRdchBglHPkSVGLkem3YXcl
aFiO0W37PSmVjOcryb7mfeGSjS2cc2NEhSEt5nKNtNbeSzgy+4hQ3Nh1fxnkf8wp
bW/Kb/sUyiRV9fQOaroEGQQJNjtgP+WofdX71bdKb/KttswXXgMMUA5kEoCYndVb
zwp6K7xavJsxM8gPNFFrSnm9IUAueCK0utcvC9j9L/AsPS8kdKqBt2P8TQUyOw+g
d98wsyQlRH0FrPzT/eOYqHlpvgyKc87GE+Trba+vkWUU6v+6UsSBX0OWT+Woskv/
aKR0yW3LSIpST83Ch89pfoQxc6xiVbXQP44PEOVAZE73ct4R35k6YzEcgmkaWgGw
ci98RX816eeKaKMUkanA/aEpvP79DuMvuCw4wUl1MUghk6zWA5uhCwitPpxnvEi/
2XykFeuvyyVQyUjYfcm/AX+dP+nR0QGk4TRC1hpWfA4T5HoBIPTBONP3WCDeHxNk
aqZPwHYOofFMVQx093MZfw3pUYvgVHXLUNRQRG/3kuigfVLSVZmLJ8H5yipvZrSw
e2jjr9f9etKVvHtnUMCttOKl6WAS0Y8k7zD+s90XOMd4RHvKiUk/yd6bw05GzJr1
vxLLqRXa7F3mub/BfG2aCOmh2sv746J/zn6V0QDWFcMBNEXmwrBhXbNeLfJB4Cn/
KesPe9IMVXICRre9drsM6w8621ImOzTtaRJeEY8KntJjwkFG8cz5rZoBuvNKHXIc
2uGNYcA2Q0jdr4T4HLPJIYbETuoo+MOTRQC6DUhxePrLufkOt19UfgxZ8FZeT3fy
a994PlHxgb996656RZAL5HSI59zz0Oab35nSg3/oxM+Fk35wnkFoEAUrk1bOtHTQ
evZSc1HjRQsNnhL+fcM+AV7LA+WrjxWcz2ZdUhYnL+4gildE6vt+zH1CFpn9YR9g
I13309GaCxM2vB/XDwIz8ZRlw/RYkKeFeeYrhOeJYpiR9vujIz6nYaPtZCeIXcq2
WaSBm4rbSBEdRJHW7pOeO8lcwaqCWqSshVZdZHXQI7tq8z+eA5+mVDCShFTOVQRH
7tAJgX7YpZEw4pBlJiTWDIZXXu11tt8nC6siIHLftkiMAO3oHHJvIf6N/F9YR+u4
5lXqAutmrEpynferg2roJo7rnDCVaahfeS6vthvoQkteuVotBvl8WH9IKJe2m+/+
P0Az8P78ztrpEXQpVFraV5RD9xidI88wNAraI/lrQ+HDnkhYzaSIIfQKTNNNO5NY
kdCJCQ5/wKbQn67P5RnvWBDkRPmDWoh1f0uZZkkBAvkg/tdiqMuJG+URPcOCZQk1
m04jyhWac23yqkzQGzNGfG3GrzeELGnJ3hnmSCL4Ecc+7l19fZSNS2uj8mSD+JeU
HNBtKxJeYZcqkBvJopiVv4oIrQ4pIniTqpfN5SizFYYCm7B/Qv+x1XhMcS4Rgc4O
LU7YCkWyfpO5Vs1z9tjBUl66FP/9qfPFnf284cSFmzvf8Lu+ezlB/qdYgERsn9sy
6j4rjFxBrv3CPXHqG4LUeYCgRU2PuQa6li4Yf7ZSMmSt3Xpsire/pu3qWXwMI1o+
6H3sKu+5uMOAWk/xSdXY/a4XzDv9GzQjBqQGy626YBj6vzmB5Rk5rElAMkJKybC6
zSVrtFL+s+Bw2T7VgKjITF7u4Tj8fblWiNerqnKdHn/25xHf4k6Ftmc/BV4sdNSd
PfjI7/JtUQ3uSxo+EnXhaKqCgEU4P8tWx886XOzcrO9Ok30/W3KQI5bk/EAd+twu
616RdH+6wnYFaeyILb8AUAXmpSeSheVZD6qeoBkrxcLGUF50BVKiE0ut726Mvie3
+Sb0DH8oR73XFeYCnCgWLe/+IiPM8vFpsQ4JFgYQT9kagq5goC5KKlYFGqRvOd/9
fgNBIyLIo+rqly/PPgjnmr9Vb6R7F8ciN96913+I2H5BskF2hh+Go4xp3AGYo6Jp
H7dcwXwKOeV2811jF1byiJYHWxOZwargmDJEohl9lPrAxQQQhkMEA3sIGKPZ8jgn
1RulU8kjyreEODmXlUJwDdG7XlEU2BD+0Ds0GvlqBL5dY5SjqO0mrAE9kbXLA2Pd
/w1SmP3Bsy95JvMMXwYxwC7vc8yCU6vYGeLmmUn29NxgyR0XsnYHmo5CELIxGhk1
UnWUXXIJw9VZdgUE+BQl8FT8dlFPyI+8hcnzDXREzfiryLhwXRwt4xFvTqCajlYb
wQGmVAu+0vbNIfzwX3jltFH93ki0huqbhrW8pJnOdThhhonf4uzqByLflVFld0MT
kVtCN/xt7h7Nsnpd/m8hu8NiVdsI0dgY+ptHcqKFPVgbBWOVksFKcLM1Yb5FkaAw
GqDJcA8D7iNw7YCVRRUedE3FXOujktDv7myqQG+i1sPSCWhdyI7XZizNzYqydzoY
uAaEg1+tlFV6N6njzGx628DQRQ6Phi8U9iMY1XnJzc5a4hO/ubA9QW9BKi5tj9CX
pvAZFWNfsWTogDcGilWQ01FsTlEvyfqUZoUXMgLocDRt4c8fzeVCKv56Fj7F3K6/
jGG2meZgl0gBscXD9U9tBpzphjvuzUsIP35smgL+g7tBG0M+TAXA6SowS56B+JLT
r5ymFocn1HC4IAoZr/t3nutu8fxd2aacj1KlLIZhanZRnulKRRfb43olsNI6kpBC
BntYwykk/wvNZNXPijG0HEBU1TyWF1bXzdaouIeTPzF+UKmc2RhUNPJ7+uF717N4
ubM4N7u/FW+RDEKfawOXquyK1X8w/lrkMIgkmCKwHH51azYvpdlMzT7jbb6AmJS1
AkiZuP8VJcC3OsaSMNyOGf9A06J/ZstKF+OLlT976/6cFNIaUtr4NFqy36FjZdhz
ToCPHmtM1UaD1n5o5Cyi+t9yYEhY0PuS9JzcRtKDyP6TV2goZW1NMDYBk3+SsMEo
az6b4x2sjcAZS6vJ78y7+9sQKXPUsz3YpFtlYVq2w+f4zLCHwpE/Z2XXc3eNVZsR
mkXqxq3vnXGTPPjeyAKimmMCSuvJxjEM8Ki5eRYXmVHJkLwmRLLNp6+paX6Viz7W
Wcq5ka3YWQQu6LuQEw5VqJbNWlkzi3whDY0HYjs1kCIQADnGG1rVIQd8uiQdU6ts
5EkGp4Ssw0V/UUIR13pF9jwOnNZwDZwTeniZE0k2vSLMxmDFXyq05nz6jX5+Fh/B
ztUfMeeal2IMmiOPKRhS4c1Pvo31US91X+JZGjt+aHHeXk7GU1Zf2h9fooZ6zABS
BPuCnu42rQUo6cYmHcTA89DBPa3nK6SKXzXTpGbLpurnVGgK4TtvzcQr/JwK6j5v
tn5/Y9wa8KNxR3cgcSeVNak9C2J4xWg2xPAJmVWWgxWF6EaaRNtX0hgqsd8vaeXo
5m1ntSIphs4Fc98tZE47eRu3BLIcg6PmJbsBxuw0feF4u3M2YKmaHkrOI207iOJu
TGYgOLrYp/28XK86t/ten+z6XI1wPyYTSwBTeRCUVOvLhDtmt6e9Q435GZ8JhrTV
L57eaJBHNRpeGyoWTlxFL7DGSqcwaAhKMm1ciWv0fSOUbeSadqTpXDH1zAbo/8S9
L/2Ju4ayHcFL3BtneLeP9s9+vsmQc2F41ieCR1IbHUa1jgs6U2wJ1NUXqC7EVyRx
LKVWPEIqTZv8eCpgT5Lm+yrO940565KK4xJfuykVHLpHPkMrPCWJhIqqsGXssEzq
QNCKrc8Mxx04mrS9h1jm8OdIfir21dfKSMA6WCeA/JuVTuwIPQC4U+f2QS8cprW1
YhFzqCRR08W1iv9Lic5Gc9UTdoBs7SLg9twtrqtPZMQ0yQpADv3Fo1kx2yMhMKhS
njzZNnkNS4dBFz1i4jdBt/QsHjARi6Ofxf7xFeqHthldm4s0GqFEmqNCq+IlYR5t
PbHn4jj1uYkcPuO/vEuFYzGU0rnRDvZrm3zLFlDi9ys+qZifghBvDRSfLTbrY3S0
4W9LF33PQce0zKe4PUr9K6mfRK5wtCnoQ2MWJ9aHcerq3wWJn+39dOWe5Sh0UmaF
WuKQfLSTTsJhnpV0msq4/zC3kIfk3cG7iXmU4lJAYOGZRvzd2jBNs4nGvFqFsoaM
sVDhRXWVxM5ab0JkWOfy4cOCGd80B1hQqdFghjSlmNhUZGH8CxnwJ+8KxaJcP+AT
F79eDSCTWwseqdkqCoWAckZSBVVokASDjEmdky07xBfhJjhqB2JZ9fLlhutkgNPJ
FFvXHGAbyE/+29th+meAT2P6LKwGbyDCpJ4TolDyLO1+fEJ/nS1ttYsnXaKGGUo9
N/MpdL7MIEf6VzxKf6zRQWG1SottDJee9CwKbiIq9/Tzz/Ghk7U4vDwNXUI389zx
gnwwaaH8oMWtaP9pQTyA68YSgMWJ0CfGNNX5CHV1WRlOoRIUEDIqqsI4+z3wXZLt
ibURBm+XocC7hq5s40qd5FZyFWnHuktW77ECgk4xdq+Z3TlJ6FLBEJpZ9wYCApcl
U6Cv800SIHY2RGY79uVChzFc5M76wNDIyJ/3MokNvz1Ai1dsv42sZRr3uUelClGr
icNrR8qr7dG9vr5AhzHU61QvvfV5ePCkVl0pUqM2j89hAZHVvDOy+i/8I3uDOxMw
SAQkh3mjcbEPHG4gWv3PI9UapDWt3ienbvakNyJ0tWbI/wpA0Kirg7QV7k6ZWdWf
XPS5XMOEwgvFJXu0MoOwBlFbshkj5edpvlHN0k5pwM+QKHssXim3O1h3RnivwRzS
d4CymNbP+J+seXplOAI74ECPkqEVvva8pSD3LKeDt4eRN2T3TmMU1mZFG3erKGaa
2fAnBGPj0dlpKK5frqHmyAPxQX91b+c2qJ47TPaxxKpQrNK3xQjYfnZJqcftlQsQ
TWeXzK543VoiyELXCQZhjBPR3p0IUIKW7xZHi4o0wa9VtUkQIhmrJAHW25jpLZ2R
E2nHB0b/CtM16hSP1FsbBzU6jTxA/6DTwf53313b4/4uOrNIo8K492pPXdnA48gS
n0qwKCzSN+HlFtp+pxRPbbM6EXU9P5ZWudYO2uxF6lORcyrmV47+MvUDXCoEhCHL
bx5o8SAsieWsJ8hbXNgtKiyFuB+1uLRG8hlFnpk3eS29dWHuTWH+JsO7zhqMg5FJ
ARB9DYa1YhPQLMlAb9IWRObTb1urewyWdxSrYYFYuVruk4gCBSKIUhjLNQbXXvSB
5CBiW172sRQPwQbHSu5LkJUabjEXWnG0KinEIHWXteDjcLix/ARu2b84C/t56pUt
Vj0+5dHOtG+LoFivq0Ogt7SNBgdsY9bVdkMYUYg5zm3fHID9EQDiyfAe1cZNfhMr
m15IohQQA8BE9PRZAew8pjuCAM3uWwBjQp19vDjFgg9FODyUjiUowsj5vDDQp/Xj
2d3mamq+u7Fxs1KS3PMEjjxazHAx5ZvdP21ue7JcUE+XfcW5X9Rc6ud7hlqd3s1M
wT0sJ2obPLtUDKrlzerYDH8ghfDxsNCOjH8BF9RbTmgGdLSeinstBbyKgcGW8WV7
cncIDkDJi4R9A8SBj9ejC312nOe/Fkud+G7BuBzUaPx2FgosbAedTI7TTbxZliIX
xDyfHFvbtk97uaFqYUMCF27P/05fC8E+DBXr+bcDtAK3Juhljzpjw29PMb0r+KV1
2RRgsuvuOXhx+iYeKW7u0ymTbfVnsbOkNyOcwestVDJzDFSTBwpcScCH1ljlC+Vu
+93RI3rsA27umGdhplUa0RfVwrI2S4SLSdg7McqfUFR5mq0yttanHBNYh/GWFj4a
ayZVimsEcss8md4d8biiZDOp4EfzR8yApbNJJqVZCq55S6Mw1CEIHNkiz5Afb5WU
rmoXrJkmyCMi++EzfB1ANKjCOMOmzPMsxTza8T4qam6HjwBwI/bgJYRORkxVEruW
wEWSfrWJFVP1g8/mSVvbaSshat8oYfowuNei/J/GlP6mMMiqd+HSnVodFXzhpbYH
grfk8KnaxdSG4DygtCmNVN4IXheAm+Q7WhYydCl7Sv1f5vspUtHSoy7YKwbPHzrB
vPp9y/PZT9S1jk+q3s+guIbCJeZ4jLRkcNTod5tFEgY8GvTZrHaCzGGS2KjUHSsh
2RwVsy28AmaNkIs59uoCexATCDBIiOXTmdYZ3lRV4BADjXKR2UsB+eqW3TGCV/kA
cuNx5qFupC7eyOP+3UUvT/6CzmPA8+GMCsjhQYo3V02Yl7yd2jBxf56+vqQUZLTr
SyHZrcK7HYwB8D+MrdDh6yaICbKmautJVjofEdUkwo1F8TQh1U7WTZKxaWAfMste
WFDzZiaYu5vKQ3ZeQzOJzzlbR8xK4jBdgUeYqJKapQqqFjqr09vtGoRA9XDx8d6q
GDjSOZrcauY64TZKFenexd+zTdcxj5LR9gZRIzMJwJIl3O1glwF+7jFM4BNVkQf/
ZZ82OeV8bDEp6NX7Dxg6+N/osNtZpyx53imGBntYHX/emdoSoYwSbuCA3nLYfpWA
waQpavyP1M4jNyDqyerKmcqcPw+vP1HuujfXeA4wpy4uBzrLFPPkOlZuGgmKYXaU
rSEJuZt3oz8GT9KidHePzCGo+uF2sI8exMOR3k/PT9lQ+KshFOfot4iHWKfmFkk+
rZEVTCcIIUSzItmSgm/hQXCQwlIZom/e79mvNcL/bSXdBWl8mAlrdgA5Xa1EDfbK
gey/CGg+F4KOBqB/a9JaxBdQzbUlYXvpVZg3kWBljKB8aBPQb8PVfd0IHKs6cihl
rMFArgCcLRYALMYV+rcvSDrLrHsdHlImm015Bu2J+HbZnuSQ8/3B75vt9qwmy9Ko
oPJ79dax0rLzBihh5eTx1RNPSKNHrH9SHHPRgKA9fFq9lVpW8WKbmDjUJBPiHmT/
VAcZY9CEM6moZIhn38t/yMb2mC6M2HT+ZTbI2YkbKnch4hYrMVhKSGJpl7L1o1Xj
pcOVhR395wodmK0TGTnxBr3wxpuKDmxxBaf2jq6dNgDUuntLSWefR1FJQzw+52/n
ahNL+01OqOHwpNL1Z43O+OUzRBJa0UayAGBOTnRdvWj3j8mXL6n9K1wjf0Av1zkn
V4xO8wcm6UQxhtB4H/CwXP3KCKy5hPBe+Nb/u3yWuCjlfLM7T1iqVHwGuh4DOU1i
sg9SvdJTZ/2hQtCAimpchmeNbh7B9Ens1KhkkA3ckWWObmnL+uJanWjQCR+bjsc2
3oZ7I1Mc0rbXNFZi0oerlpsTdYdouEDsRCRh22rbC2SyG0dliz3KUoYVWL4LHM5J
jjwBk6JPIvdu5Vet5T6tdJKJavYZmdND4Gl73X7P/a1UIK7d5PgYHNmo85KPUVrP
OiXblvNoLPOas6GGVgcHRvBB8jWqwcnV6jushko2bLz6fK4X0QrYcUX84mfZK/w5
aPLosoNdXZj3erDff93dSNQHDuzhkX4VjBZkNXBQlSvPnbJamox9U0ukNXlwhTUJ
A7Wnren8eaR6/KMCdIabZGQLWVSVFaOCdDtIDI3WHNoMBmp6TEWywq0j5vUP8Bko
pNFfTxMlw+dLKJJVcd00+blzESOx37x66BWxiAmmrlo06nMKaLbxYYySWLIdTlHJ
N1HBUrMXWqT4Bl3QZV9EWDcdQ6Sv7FJcwDkazwOUjISZs6/i8jC5+siFKS6fYLCe
ylSlYoqGB52jjeKEOmr5X4vRSl2uAa3FiG7KWYqor43iN3dDcAYvHZbLEXw1CzaS
dGjTj7uSWGKCCrO+kx7z6ngOYT9/1eWUyxyiJ65y9hPPzL4emwRpzMsq4W1mCxD6
UqTQP7hQIIc5y0RncLQ9LFJEjGt09YCjQ94LqcRLGSKRxN8kJ1wU/hSbmDTrhrqB
2v+cNc67Dd/eIQO02ptbsWgHOeMB1hmPF3o4QyTpZKW5HhHUilZ36+hqaisJmZzh
PTWEIH4MlhYKsnjzDwmu650DkKoO/BaN8ht0/i/DAYBZHd7AMA/SlxoXKbokv6Pf
mJ6GGd9u1OLLgAWR9OSU+pxkKyIqNXlVbnHsYpxDnWWZGt7vGPH4vO8DBixrvdy2
OSIMIoQ906s6XrP/Ad1i1Rs3EBzuTeGVoyGa9rO/R0BIgsjVR9Cgq5swNnXIshQn
39UK7KnjNGD/c+03t+O9ODW4TouGyuTg3F9I/SHnWGy2t/zGj82NwXq+RU++Fzl9
KT5js2PFwsx5w0P0o4BIYAwrnv3lPkafDai7WaRAUkSsGIUA0/2YC9LrWtykuipj
w9/LY4kPI9JqruT7E83i/zJLxe7TTLpjjHh/VLnDwcS3WXn5msLNRIlLQBIxtw3o
8k+CtGO15Rw7dUFP2XR0MMljhTDhExOuO6arG1IVSvG/hzjpH9/YSCbboSp58B02
mJo0SMKXqUNWIwJLPC8U4Hhi32jfKGjIBlOB2rwlHwS5345VHDEphllnw0wtUEFQ
PvMgjDH9M4tPds15dU4n4l2WCXhdj1D4ojNB2sdqVBN4Yb3utX8AFoCAHGw7OZcQ
bFLxgI7TzTf3LwxAAgt3YqiGJle5E63hO1kgPV4hM3tiwUJMIXU9eoXW6sfY1VU/
kOaNZSdmFAMzgwT/+r10DZ6PwEoiqJP7E896BGv1sQQs22TCYuXxHKHuSoKKN4ge
NwrXvd1vaPzKWgQr1kpaatQgt2soRW8LOoRqAB/a1lt76jyDUp+LjeUNZzxmKQMD
xuu3NPmL0KeA/8G41nMPF5NQFc4aAdabNof1mRAUiGCQH30mDRTGRL95T+78zNo8
RmZok4uESj62rwQgR5R70eRO94x+UwBBSAEBrfTq5mhdiWx8MUT8zQM7gfUeQ3mS
r+C3oz4qfSiv2oxH6OiZv09phlXwl1eWvaBEdwps4F6AlH4Y256evZMUEElsN2Ed
kp1D7fxv4bKBdxvlyG/JOUEMXzHMfq7AoiFUt+dH/7PK8i0gIG3kAyw/GGL9CKhP
5ynHV5ic/O74At599tXd9h42+h9mX3YPiqQtW1ryfOLd2Dgc2qM3AXPybGejhOR1
aaVC7RK+XkWgM8GTp8RNosrzADuQo7LrrEOzk9eep/mlRyUphS/QyxZmd0q2qGaM
k8lxKHZQQ/kVvlCpgI0XbGC+1B7WGBvBFbplnGjNSAJJlQRJ8ZIxY5I0qDHOZ3OF
VV3QKRloyiPgMeNU4kq4nUlpvHOhA39v6nudF3G0K5zPRqEVWLkOgwAF1zJ13rza
/POLsYnlijgyMFkChvfhZc3ni3ksb+zdfJbnM8a2ImuFDb51tN/tP2zf64TLbLkq
2v28XUCEchWFvzo9fMjNAgK+pCPMKwH7op9wYmWVGIjdWvMGTgW3weckwRn3QXSw
SxbaWVaW1KVcd3/5CocznorLYOzIYeVaQoGxR3SL1WfFLa0En2Q3Kw/SIpIgHcAG
0DOfI49U2QoXJWQlqob9pqq9apNL7iGnHQ1WXyjdECpu1u+Y1Bd0fWxf8WdsIL7L
9+zP3J6coTJtBeoH1+yDr6Vla5IhN4BVjBtMEQpOBvUI6XFlJAl9T0y29BygM4He
jZcZP5aR08WrYp8g87S5yg99vVbuI9JvsVYDxukdDbdQyY7MKRDcfALfQAcJ2xAW
MZfn5oN9DixQwkwc8BNGH81/G9nzaEtRopR3KndNpoLyzWcz9VkP9xwrXIp2jexY
9/W2soDFUljolFDbQrrUaNa/NvywhaWAATCTcAsDLAZoC4mJiP2e2k81O/OE8nbQ
LVXm7ziCa06vwD7iERDOTdtPyvQ5fxv/DVm62JsQ/nRtNaD8zn6DF+rKXdgVm9HG
3ObW4CcP2RtUrK1HMSIfJ1EZgoXvTN2XhEVPF06Hn7Aa9CXdZTh0PDocECVV7u1m
EGHqaLDGDHaESKG4U1uG1JfCaZT+hYYsN+C45MmCvbZ/yKik7ALl+d/ba/2KORXk
OIRtCoJkoO5JK2J2I7dwtxIUwiDVer6NzHF5wR3IRtBY41GQYJU17skRAKebVyiQ
4gEAbfAWn2vTyNpLZknhlJRfBFHXH6ndDFheGSh/8vxPrECYAazwYDtvXscmjppM
DYD9J5db3VYKqOC33G/BImp5oxDZDUpHGKCWHPs045EykObHHdbXB/uZd3KfP5mW
qxPBmcO2GfL9EwSPu7XI+H+YrgLvc0i8r2Zq9nK877aHt9ngPR+rYUmcfDFMNuJ5
tXXS+240kmFJMloZP7T6nZrVzIlifsWURFuH6FH4eZBkHrBqg8OWI8NDLIwsJ6SK
34cE0tg0csIWdXNK9zmJmpWdF8eRErKsVPjwQ4lNNvHFC2QxE+GBUoclVsUQoU8u
ol1mOWJVVQPlAV0y/r3KLuni3rlMUkNx8cViGj5O3ZTmWEog9NxehFM0WWKy9hSp
Kwy/VDJbuvVOhS4CF3HxCF0ayIZfssJAJDzzcymIrz/L6Q7hBzUlbHJg3ROwHP2H
Lcj96OwkKPIgD4HUl5ko5F3z3qTi3fUUMsalopIy1OWFYNoauYkKM0O/uDjeB77L
nmEj7zC6TM8ftXCitnH7I+06aVCXdz8R4t+5M1q627uNLxRPF+10h/R7JcWvaDV1
Hslp6GM9JCYGO2RpoSApKfhqHNVnQSx+aCujSP/3CRf9qEvGqHzvejAqlM8BhDOO
X7Qbr8/AOowO39qxJPxuqwwGpvEgYu7eJ/NM+tDi+myhlRxWTI+5eJvnG0vZegzH
Os1wSJz7d615gf7wNvPc1Lzr0QkS/25Y2XskKJaiEWbP03iEZUNsQJr3j4zhP1vm
T5kyCrzdiJwWbZLelLTVRocLAQFZm1GPEFposGBGhSUFeu8McUzEAoSSSrkl25QX
aBZxq4qHIyIUwD72eKNyriEbC3suDentsvZFrd5+fm2XBsxIeGpuy5S3ZPHvILF6
ONTBOqRBjmbveMhwQgu4K2gwnVq2PhCljoLCH064LbNVOHooS7seT8A6BKY+KYp/
pcYifQJ+cznJ/INLoX3TFXkDedYVwmBhhFQulCtys0vRhe7Cfe5vpCUN42QJFNqL
IAeOmMCeY6sPar9YQTS98fNoUkGfkDvKETyFsNmL6jAWzxCuSnwr0tfOrYLJ30hM
/Np17YFEOAifFeyvVDNWc7ogTBbvj1lPa54Ob5XZtv1biGD93bsUegEbVrCOe8mn
aMOXk81AKZu8JPR6ePYCfO2zlnAIHF/M+sH2rhr+M2xxRMVoF5CT9nzN1Zp+GEsW
F1dVBBjg+QUjy6QHzzPnaF3+rv6n9B+mDiZ2ZWn+04BArKitPkQSFf8eE5Fanw63
4bmC/V+4hoegLKUuOoIznjplefXS+DVMPoLRh/B8gMLv9eApI85QPnFQfGzzTLWD
/X6Clfed7n2kAEVuf6sYle4Rwndx3oDgx0D0ovJVDiDKUpHrdum3+dft4tfeumxn
ktP4O1xjhH+RNq3U9z6SVkovFsdMgROZFHTlxfL5pqgkWJ9So2vqmTjGiJMwLmvz
MAspTSsPOFLYEh5M8A1RYe4SYuQPsItdCcSUYABiFNBDWAB9Uq4b6NY7YXfkMr1O
1gdz/AtkYG/s1Z8fqCCP/xNdFqCsB5o4amGDdz0C7PJECRBNSsKlKF1G33/+ewL7
Ysy7kt7by8SMP58fLhncXfs6FR/MhpnXckFMLKogT/uJPPfVEP00HsTyT7Z0iH8O
/R7Ap//4kvdGS45FQmUcBLa6NGXfOBV93txuiJVTA3RyqnWR85BlxhvtjxFWuzAV
UrxuqkbJ3hqqarXAcjP97AAU1wU3Cq2o4sha1KBCxn52IdqD4EHdMvsN+cJ9Nwvn
nzdaUAxYKzpoZoXxeFMd4NPmFi5EInfqSmAuAdB1XqO+DNf1vsWwIuxHGLQMN+km
1O/aY68nsZnEmNxB8HNgR07FkZ+bbJeq5UI4/JEroazVMjGQ9DqbThVlkAFnI6AB
Up5rVwj3csPM80vLR2w2a4s3R7GrY+4TLrUcGigAm6shlrZosaGcyI2g+qpzXrOf
0Js0ALxpk1C0o7rgehQuvoQn9AJqyFX49dT4Vbg8kbDlewgYFDOXUwFKB6RQsFJ/
OUBApXxhfyFa3ouRbqf4oS4liUFbFdYWCKJR+O2tGJx5oKYBMyoNqeUQ5zy4FhLL
cc276LL3MhhEQpT3bpA1baONzVwLAfb3somRMXeFJUIknLr8ap7vMfvZ6ICWOHIo
6XkKV7o4XDN/Z/TCNFeODSnjaBzkQe9MV9z27rZ1/R9Hggl3Ek1/+epS3xyCIDed
O1S1aULtlBwy+wWPeXphS8ooJTCiMi75jOOCzv+loZPAA5YywjZYjdQ0un9vCe5g
Q70eD1NurQpYmRvWxFVu0aGWF/xrQwUlePkQTbqRm1+dMhSO7Xx49MJ0E4ZT/zcC
bzSxc3uvAWFpv7IQFA+l3aBscKho9x9MBx7MyruyR1IoiGqx4XU6Rh7oStU1DLRS
MaPd9L3uYHv+Zx7MJVy51ukHh++CRlI+sDvulwBli9Q+NYxo2uPN9soSjuQ1Mg3t
gv9OYMHS12Vrk/O3k8q2eU3InQ+AKEkWzhn84MRIhe8sJjJxaAJvulfcDzyiOrh+
ViM8UjJJQ3gqAcViGQj9eSaTamNPxoLdjajl454h/mlu0c1iLiZHMWf8L2lJddAY
V768LiBirZH2keIr0XgUJHZwXxKCMyLQ3w3wmRqABVi249LmPxpbMYo/YW6X6Qa8
y/jcFQJlp595LaDrkoO/ClsuSdmkXAtRbbgJVp7g3uSICoY32JUa5xirPqKvxjzq
9rdrTWe3xPIOsXoom4mbhKkUQL5KBueo/8btz8fZkBEcxRZ6Dn2D0ztk/HlOa/7r
euZlmCg+IySdmI3NL1U9iezyQK0WK8mT0Gy4Y2Cb/zOagfKYq1t0eAejmAjVQWXT
Wrc//Mug2eYbSInmFByjk9ifQ3f7PbJftlYwzhiq3wbiAIXiq6MwxPzZAY2Y4hHk
bXV/cTSyR9P8TI5tiE+AQhkV/l1fWCddjNmgtOLN7tLy/+WK1hM2q2MHJY4/uEaB
I3TMBruf8UwA4Hc5G6CXFG8/8eYwxwHMBRy7iyZEBECIhSlR+uB+8wa8+kXMShUS
DQCaSXgC40e52qjg5h1kyPdfqosKDE5l6xpulV+65HO4/PkNe2LqGRWuEnyIkyXo
NwNJws7R5jRO3DTTQCd/KvzrPQ3PxXyNl0LivNG2WQp9EGv6aDMB6E0fQJi7Cx3v
khDdmoghu8bvfcTRJJ37oba+f38PXFOR/8e10lc/5cBjt9vTN/yprmiwdbJb24mk
WnqYPirvc48AMk6vqBQVvTBIVTNCeC3ktHArP2aVSBCQh55AbzydHddSmCv4WSpd
ROs31pSPZDwSbGXVJ3tlbRt5uxPF8N7kiGJ9j1EL1Sv+z/WuaMqE25KbT17RzzFX
yMk0viiMmitGww3LhNs0qxYgJF/rjyiakPMl8+RzjsKh0Tsrx9V53cYEo1VN6lSD
/Lob2e/yGVDWXdxAOR0/kLVAtfFse0lG0VusYOIthiySqxKZMmG2mwqAqDwWlmc9
8TByw4tGrau3jhc47llspTguRtGN8NsjtgBjMJN6OXJVh377fsXmbTUuUlaqALTP
y1GdX90bmLNrUebNwB2KaErVREKe+iapd+XIQtE7lMeoy2PlWdo7v2AeqngI2Qhs
76zV6TzWruUDqcyraV96sSLazBme6KYseLZ3MoCEdt6UkqBl0P2uUgcpQyoyedG9
psnb6ZxWygLWPDz2G8vHlmjT9HTSJi5Krhm1QCExzXjtahq2IbQ+1wHMLgrXCimw
XwlFagaItAAcCefmBQvB5P8h05Voso+jfzjqYOBHIj4rhhxeUkYLlA/u/ahab8LK
4s6x46/iyqfF65bb9n0H6DP7AwkoPJpWgP6rHYoCt1PF3NEB8TCLJyuBGRYZRY4W
IHqKk3kUd1yAPlbh2KAZBXEfEZ26sFBoTXTZnGevtl9Zqn9AgUGMKST0O7qxUDSO
DDu0cF1cGnnMQNZezmhBw2Pq5qSxZMr7ex+S5FQA+k8hla9AGteHV2T8+4zSyuQn
CUXRy5/kmtKpu8Niv+rdtVJB5pgHo9e3ViVCoLyylL5mrcQBR5VsXvacAD9AKAtk
kpBda3C9yTsLCl3tCCtJUuTMIgwp0YnPsmVWZNR4mZ0+ITJPNh+4bzPjv0RXtJYB
CPOHlcztlqYnooX/kny9IdLd4/xafqL33WNvi2vfoeW5tAwqcx5zJ9uWJYbg/2ci
GZwUuPplj0e1ka8shPQi/YnAx148z1yxbVXe8PS5jm0wAba3GFmqtOgKeq4wSFWx
CpvGksv/y36hJKW3SkzxfP07aGx4gyCAxz5wTNKKgy4jWbdhuzbCTQPnrGx80lvg
xuEBf8x3j0DGa6eQNNrb0YsCVWazPCRLaFAw0oxwTn2nhZQGPWBnSOBnKaGSC30A
G9WtrZILO7Q1QY9AtCiLR+VnaBxlWegTmzHSGc/T8eypFwmQg3EZDmAqOAYTolwS
q1v43T9a1uM1Euv9MpOmZqoOhoGAuvHaOeA7Vr71N/v7eOZbSoes8BJuv5SvNccA
efXnknESHoGd+cgBHvAiHx8TYlafPkrfHIv2wpN9BkOylQxQxjZjNQ04slT6ljU/
OzXTCda5GJtSE7TIWSSpqYPQ/k9t4IZnc9/KF3G2wOLYuIqNUFwyY7wS2ALLR5QR
D5aqRYEHNZySi3Yp9jaDN98qWHgICQ1PIwfO4ASNqOV4rXH06tUo+PYNCsLE85+i
sM89hXe5v4i5aZi8UtnAQkaOZiunjykuovXQ+K3r+Sq7CSulKt/8KlH4np1O/sMN
YuGAHns7r6wpiM/NIcgy6CJOReQJA7Cv2T2go+CeIpby4SkS2P0e9MAVfQKl9EMb
FmGArRZKtwi41Jg9HNkuTPKARL1Srpvjq0gmwcTYWDZhEwuigBo5RdnFfbhozrb1
U5D5NDWTWn6TrR1WJvU8Bw2x4QcL4cm0/Y1ORrhlT1I8Wy7Cx1eAcEkJD4kEczpj
R4fiPFI9P1A4vAcwZ+JIQi2EIH70bitXx+we26gBZ2VoPErseCYlyYbNH3RRwE6x
K3rdiMwCKBYAVAg11Z4nzOYMgrc4CNqt3LPHu8WxEjv03TAU1RzsR7y9qTkuMzGU
lkWCEt6uP2UhvqBYZWbiY+52BiTA9W6JJBwD1cQs0N8D6kGUhCe4A3ctMM4EQVtV
KeC43GxNLT0XuSALT4S/8QiEXJ/EGRq5NaQNfKh/kaike1iStWI5ie8KanDUsANj
JSSO90jPYfdfwmou958ml5hNLJ0//Tqd9q6v59MwJ/o58IxYqDS8nCPkgFT6gYoV
mpG6t1qH5fcnrwRBOQLQXfYvqsyo0d5snTWN8GhdxrpinmlIfNh5X1klxuJIqBH6
JZv5WrLiRcdhZR+Cm8R8VvCyJYBCbbC84lVih4N0R5GaOR8NXnPcbsIdfZJWycq+
FhtsxBgAJ2uGue3jEpJUSNZq8uwsmFYaCzAEsK/Gcgb/od8nSD/HdoqWJ/0jnGF5
7gRAMnlZGeTnNuxDAQJkt+ArN0/nUc7oNXF0E893mGAvcYj3WDmk6RzUhlYhd18M
BASnU8umuj2g+6YxImASISqkm6njNGQxH7CqQLvgVdSoA7rlW18yQOA1Z6+lxyNq
IVCHK8qBmgsa+ENbKMbWduNI0rQLatQrInuw6A2F8SS65+dsdkuCT1wGAyPoYQBD
tVlcRdKnMwXoQkfSjG7Rnv7UmwQjFysBxLz21xyIRJadDaodMApvo3KsEoBfoWC3
52do5l4WZq2oT+3q+pYG6KEyvQbfepUXCfdN/iq+TFCZDXwtSvXZSgC368KxhXK3
lG2W/tiaFXLTShGLgRYyMERz98poFaECmoGsVnGfk8nw4ohc/Phd715Rt5oX2Ep+
omexIHnsYszuOxJvJkQCVRdGTeTwV3RjH8pW1l05ykPGWxvH7Lxs/nBNQBGhiFP6
1y4wE8K/vrc+S6c6BcPlccSCz9ce+OlZpqh+5FUcmPsuKGEsupJ7hvlugA4Flcqg
uzRra5AFPFif5UPBmIM/SQaGE3f2NKbZvrRKWIwemd2MAfO86TG0cDKu4VwMaHGU
P3UD954M4xCiZYbIv6dVUKDhmpUBPPqZ1N05UE/+7gPM/Sxj6pPWDWWAqGCg6ZlW
jZgW7kpSVJLN+Q7tlwI8B4MxQ4Af9fMJ4smXqewoRxYVY35b6D4jZqdLjtxVu9ze
f3zW6RXq87MxRdjQrgaosUwz5Ay60TwuMpYQc7ilT1bwaCRV8Nq+a6qhwJ2w8sr2
ih+D2mYxyAOyoZIJfkWubljpOrjAAcwQisAT6YXtXCzse13qYnbpcnOYjTsSaKis
Jg8tkiRIBIx4BNrfjdclP8THKlpSk1okfJtuhLOirTZh5ZHpiaNKmyczIuOMsC3p
7EXAH4PANRx4pzpzU9AD/9Z+dhr+GW2+y2Wyd/6HCPX3VMV1auccQ2SDXjEha6of
OKupSznlD/mjYkcwc3Y4e9zR3ht7ZxNg7Y800xu/4npv8Mef7kmk4Ky3/cTOevl7
6mVrLdSEh6aL2e3PfT1zxbd4fv2338s63tsdDLLn7G2RxR0u6Dy+pdNerKkyZKRc
pCus58EO4EXZ/Aoi2ENZzwX+aCF3bYUPyX5afcO7E/f5Goi7C8ZiIdMrIa0J3y+J
urgeTfp/Rp7/GUY5HNuFpQhIvUXOnhh0Ty+a6UY+JeJQvIBo+Lqz6dkysu/nTj53
SMFz0yUk/ap9HRag49o/AhFkshwWn9afozyQWRa0VRGk0dkeJDNnUZOGVYVL5KlA
Yotq5IzqqG8aoReWv5iCpIbzlnhmmur19oqPXD1PwAHBwn9wxNnSnGMKMKhbpZYy
bmF+t4Db3LjN4Y/Z+OyhTkxgO8Xvk3t943ixcu52qsztjjzMKtbzKMecgNAWCR+V
qy2QQoDN1Kc8ZWbhWAxh8hbNVzQkFLrLY1cqfihPaDl4vAjUa2o6LVAyAaDHc1jK
o6bVz69v5nAjW6DMxNKgGoqnO0hpV8RqiYPcP1TOcPwGgdN7DNopXt7vFak8gb4I
U9SrCtXTw593BYmGMcEAAppeqk5Q0Phu+sKS0M9zYAX2qql9g3BLTaTL3MPx2j8W
pGGYJPb2dO3jEednFG1/YX9WBmlo3KfOB1SJWCuugksT6WAcBMCOByjPwVZ3dSH7
rRNHY4HvcWncNyzq/Ii1m3DvIJcukhHon4vyvCcJ311DADsHOBqHCuw8F2kkHpI8
LFZYvG2F4qnl5VCkBTz4esnHOXZHUzu9oNF1BZ5MqmlJ5DBDihAxhc/Hkdto8E0g
BrocAlvf8bLQY6Z/y5Q2AK0bZ/FLNoX4ev7WOc9Ogl5aA2Y2nwPNZo9LttS22wSi
Bkti7MYnboQd6ADgbB7QEgNlxmsYV/2MlhPHpMCF1fJjrUOjzL55CCc81BLRQ4Qf
8m6tzLe3xl04fAkqusqczk1RTDZN/C3AHBcyemB9xffmhYSj41WlnsZcufJ4QQ0i
GeBAWOVZtZnyXI1+Ux/21NRxEo3rbN1wrh1lZWk4s6fShatGAioGgOj0m+rjVVB7
ZEwdF69EYiivF0+QbSjvUWex/5BqUQw4NI6QWvgh8FrOob7Y+fHEqzypAtN1d0G2
AQoQgrLNzLQraAUUx56OQFzSWtj42uceOZozaw3Es7PY3qSVamsUThCUvGDtUqRv
E6AHZso7AFA3s2lMuBQnVv/qNKbbXd00rTaKHVLS1sqgHG2tOAWalFHGAfk2yB/r
vC2mlN3daCUA3ULZTaZoW5D0MJl1stjZZFaapb2JnCCb7yK/pD3x3aGQVoWTqzUE
RO5UWkNh3SckzTFhmPstGsO0yPEWAO5vpNcHAgjxyMI1+hcfzFnSRhLB3vEgQF+r
6LzHG0qMTDh2kRsvcrPN4CywDuDOoRiadM11I30EUlfy+GigL1dTTBxuA1v6uA5G
Ee4ovOPauBksB1ZCa3jwklR9JxjSoArz9Nn76+cM31coHjLROErD7talQQFpxtuZ
R/wyUw2vzU/BffkkylaihfpogCN/OfO2dtH7W3ut9RApug211k1cPpnEdmA7ae39
NwM7KjQsIQocFBoPEOLmsgta24V7/pV/yRRgrSysIBmCW/X0Tlg7R2C3BS1ewIDL
q39ySPiW3b9GZ4pGYCzwtAIog1fDgOhYXHLVHeYRHQXE0KbWlxExUvaS47TgaB+/
sKYpYcjFYpgZ5KmYKf2bm7HMq9goZdGVpzamFlg89lSCSjeojUZN1Gpi55Ya2vXx
HJl5kcJDGkK+YTNvXNyjQ+I6xSSFuZpv51YiUVvQ/blrg8pKU+1wDCv1VHuylptg
Xadml0kTuU9kkB3EHX8xYGgkeMM38DZICpVb2cwbbuVqITC3fKYrvfg2idEZiGE5
XPMYHerBOzzISvEDlwkoMmbg63iVwkxnP2nkA4ar/fdWkF14orPXPB+Jy8Knlxyg
uF7hyWWz82fcLPTvFH/rxork2PXY0N+MGVGnfbDwJwhJtg+4Etep3tR2kaW8QoEO
AyiHEYqPXmKb18JIU5a/XVcJh6KvIqKOH0K6Uk+GELOf7g7f68H2Yx6Dhpemaf12
Xa4Iy+e6vazDgKBFif3yUuvNDiFthwJC2HCIedfsYb4Nf6xHxWMhzOCy1zzehTCF
iHXNvMiBnyyEiKsmJEezb+4QFFI0Ni7mMMiZZPY0IhywwyX5QQ+du8rIQKSWf6P4
VRfndrBcQQZAQqZgv/aA26spJ0ga4r8ogwnUpfG0vUVI+FH5cL3a26zGJmf1k3Wz
DtX7XSR40dbXogPNyaSn16t7a5L8/MQG9vP5H5mQ0dc99YVB5FHRHvcTowHRSbR/
DdacU9TwTXsqkhb8rw2uHlW7YPfP8Cqfy0x4JCCnM+VyGy/aq+fjYtLXYYATyrvm
X7kXMnsbzCjFYKrfE4S1SVFqG72ILRbTRHNHZuINhuMxiM7+SohJrJipzf3mXa0K
ZKNAzezhErEtbfADPx4CZpBWWKgJ09cSae7kQ37/xolB6MhaatGUF2xN1BqtLmqq
cGSRW2TJOOvFCHoIQUw1ZevEsEZllDJTnfZj46Kk2/kgV05l+gX1fWUI/VnnfUWE
UG9RgiTU50Rg5sxkoiS8dyQAbpTIKvoQSW1gLQnyN1shIJzQ+eJiJobkIqQftqTt
oNxbMAcIIpxplGn85hxiEELbJmwb1sXQRs1vTYF0Z4IJNNrNqrYKaQwsKVn6+Swz
Xw+BXlu0fXNRkFhFPHFvyt6yS69kTbCuXI0m0LdNrqpNpQVGIpqWoaN2NpYS0ISi
0QTQEjgl1Vnsl+NWJULJ0pBLIiVoxJ/WQ5g83cU1AIrugLy44fDqK58YfsqEbyru
DEKCykhz4E08hgJ1eQPieYaZ8hQG7sce2JyJ6JgCNkRqb1CB1zd7QcKZ0BRqTAIn
nZ3CXq3WI16XnMn/yPsArsOdCzCJQCsCUW+q7RBVJjL1THny9qXCK4gn0RNLCNGY
rnhvzFLG+YMTAslWpmpjI89Kf0RDBMNxsPT3Y3JpwVacMLgFMPy+wSRj/ZPgn/CA
sdZp6br21qvxRvbTat4DNfYIODssLk2G2X3EDbn+paYrRrD3ULah3jKsimgSazjZ
A+93S6Qo6Tk83/NWBrQEhh5DUzrKZ3I/pwrdvkPjT0TypUIE/KRkxc9LmGRRjD8p
mmIJJgMnqo45h29SqL3wjA/DgatstWvbe6voJHgScpwwz12v2fg1bVLjQxG/xWSs
NYKRHS7xdqm3hbfUVJ2258FXPq7XXjtQn6VMh6y75PAPMBlWs7WOybHFzv3hc6D/
w6yaLPTjnUwNi/Q23Wb6x8bdTTqv5UA8BtQvsg5ujgWcC1b7AggY9BlQDFLyPPZ+
UmDR3ugZLfYITB0e/Cm2GNDPUwdPtP16UtQSfTzB2nHgcqU2xkfOwmxS+sfBL70A
7ROv+qelcsn2IiQrfSV7AveV+yjB8npvBboC6lhAEndlmW8amm6IU2UMpkDTdHG6
OKbhcNm58cZSs1jvMBjtFEW2zQL/53R95s7JMTSpqSkU+nUtq1FE8+zymQQJN1Ps
U2pu0vx5RRO37KsuurAIZA+fnNS9MBFr2AAJyTAu4R+O7gnfh6CxA7CAYuqYPoW2
bKqOa8vhdtvVr+PdX7Bi+dH8JTNsVkXQSE87r1jCuJrQG9iLyP6AvykhbT5jM/ka
010WV0xCzt0Ih9ALkSCyzlMx0dIGd2gvhetz9jEKSD71KWsqqMF8xmsYKOaxLXik
g5kfnOnN5WP8HSW6FOGbCLG/9h46gJcyPGl/v1RaYGvtOVko2jrEItjzzVls2Rs6
UK2ofABYo5SK9GxShbt6V3B+Z+gyrE0LfUZexsyLJwkomTK+Dg5ZtfIzNN1aGFIE
wdh+CF4N3tPpSs14GK3hxKLP+aKuvf6DcJ8m5dohjIL6d6Pfn1IL8Igcs8P6aj5q
jFTLiLKWvMDeWLSQE0ehKJnZ//s/vhusnXKV44U23vn26IOrI2VfFxTZZa4oSFGC
MetqXYmRE8YUDwQdsyFuER4CIqEJ8Fb1l0a+hVRilh4/Tnx76JKp3SmCJdLoPE3r
QefVeY4zKZ5lbK8uzlhJkN1OY/nm3nhHR6T5RaXldktu3vkfgjWpGljxzkFYrHBP
4dINDqUDsl1Dg5GHQDVdzT6rlkl4dWEmGDwWiM074n24Y9HRiIoxyXVstBuD49FA
fvIr3ArQNDJ6BGyOp7jThBZ2E2eN4Jk6uuWVNmmYyao0C3EhL4wYlqfO2zN9+HA1
mpzV7wXLipyO1FGvcAFy43EBnvVjdR39lpfVk5MDy4/Whq/MbuOkDha91aqrLT4v
vMFfCd6NYSVFFLgbm0TKpX1XgCgo4evv6XR4AUy+0OMkoWuL2pZ2AsZOKseos8gJ
Sc/iPuNMnwbatRwUVw2GhliWtIboSU75hXjSgalDZ9cRveSff5h5lXDu1XAuPdCk
nSrSOG8CpDvzQsnkYva9nALT/WcRM34TrMjpX6PHHjOu7T8+n5rEc7ZPnFfzMiIV
DzI/4gZ6tom/+WucWACocJOXH6/+IfRskhQeLkHvKfBtg9TKGPBKpASCFQJfZ6lz
ro/H0JCBST1dUItqXcrZDtjiaViLz0lSfGxLXnYC5KCpwGF4hyIEtiHSRkcTUir+
y0bSZJHUjpg1pSZdfdPLzEvdahxqA6TnAhIOQTKarOZhecOF2SyfJurtKjd+YkRb
LYHdVWc9pylIVkr4GZJLQL+T7PDADnzF8RewOnSMA0HT+s7urfLMz970+KmoomPy
OMTuDECJWsATo2k6HZAngilf8C3DaJDK+sDVe8/Y8goRNHPcezwUZ1fL1ak7Z6RM
BF5C/1hDWjgRZWQ9cku8ADLyfEMQXtoDOPamSO5jBnfIUK5B+rpC+tZKpL9OXsQ8
/hKazwtegLH1+v1yPdp2edFWrAma8OUvWXwrtgC1VVPfffZv6qlmXedFECd+b3hi
FRHPb0Z2f+SleJmvCLLiYEyay2wx4ZOdlc2wB4D5iPrHCaGC3iZ3ANMt/A/yR5L2
IqAM1kcdx96XBBWSVhLem+U98+wiktwgVSV+6dhu/gaql0dheq082cwF/ev5j8wI
DF2604ZEOu7OixuHPANjXNXr8qiK13SCffmtVNdrBk1XapRuBnk9rMg/Tr4ereR/
ipN6fBRb+ELNpSRjI33Q+6yXnYME7pn449ey3wh1hW3i5mEL04OIYK+BOAISOO98
aKa4p+vyFcj3rR9RcvrH4SKOGZZcNzRUHv5LjQNYv0Y5pavetgsBaFxk99KmfbZG
2H5VckMS82YnovZcGBS8bmbFba6e6VspsfnmLb4CMB1GTF44+CqWp/aaylOe6pJd
SgvWeU0/DQzKGoBcGiTFDGmSjvIQSsi9grZrLAT1bC5oBr5BGWWVmCEtnaO45Ci0
Aeluw4NxHfTP94omCcxLer6YFPGcRXlaTuPfyG3IZMWZx+jd2z6QbltFrN8OKH8s
yG+k8o52ETPe8K5aeIB265nlJQcpJ2plxvYKvbgC6miP9+iyz5e1/GH8kaM2tsJF
0wv8WloRBPLMq5cEQ3KGjKJ/KxB9H4DteaLNZfVIzfMnYTZ+tH89KHpwGxGuzxRl
q4jGOS34Gv4UpQ0e/U0PAICeiT1GuO1lQd10xqFChZmGjJ7j4bHDro9/8IJJWFrO
miwqe6N0al7ym3aWzanoj1UL0/Kb2U1I73vjffiT2RETvcTcPDj9NOMFEViBMav4
701yroI4MqTA7RWrwcUWy9OEGQ43ZgAlg8zrOZHDznBUUH7vY11MzqtCAybtvXWO
NnPeHt+rSgPiQxqED1NSA12TdmFwdLCdpRIhoLRl3upR1kSE1uaB8+0fHQ+dtwVD
Yd1colB8OkNF6JKwiaZD1qXxBNJDMHQZRvgqX8lfuStIK2U59QEVJrYFJKUdupp3
lEtLc4KYD6FdYGIYElMDHjH2n+tA9IDtN4yGHJ3XO47dXW5eUmG1o+VfADS1wxko
VFKY8h4j0g2uoAQj+3q9fbP2ybQWbFvnIDLQlaxaObAVEEuFUPLJLkXLBALqpjIc
JHrNMVyNq8HleghzDDGZlKV4dZmfxI/fTcu04RO0F55Q5d75vMLMut6AUMUQdOSX
W4MKP81w789TfXAoyV1FG5KIll+nsMhcs8HDbc/n/22pQ+niKmGC2Ss97J02X1eW
QZBVHCuzdfdWKhFSj73cn/0HIocyGJWhcHeP9GcwP2HBqO1fxWRic93JgqUFuv4x
Y750WuEm59Ml40fypIVO5+/+MflIZngU0QvG+KTqqZSviABt2FknS1h9Bf1T1a6X
mwbOUQ2gdooFI89TNDxX9wzxbBNsngm7l7RWjskRvS7KCvZ4STGPhwgAtslpBTxI
z8z7KnEEt2rY//+XD2hOWtDEoBFxlQH2sgxdPi+RXOSD7zCW0iHI0ScYz5s/TLRR
C8mFFYSF7nqTJ3Nf0ZGwBgOm/1/6vMKhHRXI/G+CPMUt2spt62UjnAfPqAemi/D1
plxsdNWFx7sCcNPO3RY93m18KT1rDdR0FiByjotNkqQBy2H9SMNxqaTDxpwjcVXR
idYpciqVFp7rQhtwohasevdUUllzBpMKoaPdeyRqoyApwL4J5R9peBbbuWsce//p
pJ1F7xY5oCVH1D55E9N9dTyOb7bax44m+3LRv6iOdEd4Xy1EexYjoSjX2wVgOkSu
ClgahIN0Uvdo1ol6wb+ccYnLyneL0v3vGSlO4NguXKqdC6zXBG2BtUyq2L7ePAS+
NddCiW+m4WfjAdwHE+WCFVlGl+A7DCqVsRDoMNpyr10I5OPbA+HNQoAB+u7eixsC
Z2CkRGFXNiuG5hluan/ZnwFSmfBUFsW0uvPPjqpCDCr4BPmUh9FIZSk98aeG7pZ9
TMa8bxbftM35nzV5azLw97LUA7APX7Cz2N+rq9L8erMKZXwWIPHFD62UC++ABNfu
P5MlqUeQ6gshkYBDUE4BfSPkc4Wavk73YQMCqKg6NE1y+1hqYsQsJJMcsbh/6n0J
FUL9Vs8qQFsvC/PiovR4ddCQYcF4iatBwsBuFl3ihNdJDFfJejo2TYthHwZ6XB63
D4p2lO+7m2tABRlMnWj/2hYqb1RiCMiyk4dSzIEbxCF5hH8ENWadf6IcACz464Vp
2k1iRu0I4pVz+SCzAt0nm5CdckNIWqzdW2tpd3Th+Lz+Dmt6kxQ9qyd73DlbqQFP
AF3jfOLI35Z9xvThGNY0nPIa8Y4P6Meg4JULsBU/GNlF6Cjscf6ws0kLdVcEtJji
Wa7+gB5VXjbOb5AzKkegNd6wN/XJMmJAeZX6eIP2hcta9RDP6/zKTjVySNeJPAGV
c/tTngcdAJxlVPT2mJX9M/3nv9O8OupjtlLU0XhmJ8atJ70wOb9rGHKviRYrwCMk
tnb6g83zpx2mR9Ke141JnYcFg5G6kwwWZhwhRmyuzUQyNAk5RzKp+sOoXaVGgGK5
2segOpyWtRO9LxWHZbViNbSjjsSUgSOMBfQIytkdA+dm7L5lIXRFAzA1mteav+Jf
I7qhg87UIRDOVNa4bG8DkeGp5suEEocOBuVjf6iZIZvMW5BKaY7jzYph8cMcKz54
b5Ju7njHWK6XMiKUC6552mHEjjOdVtbg5PKZ2nDZOXvGFuYG0Fec9uwhUvkL3/F1
ky30OINRs67fO74a+R2cC3x5H6lKKkFEx6h4BuWQX4i6WD3J59JZxf4kyc+YAYHT
QNr/prL5o6nAfEnDDBfInIVq/tnST9NL2PMT3JwdCkq/9vvzE6IGTY6RSfFXqkDR
rBJLrDuUQGoRWK/DYIr+G0Tvk3sF5w8TBrqJSWwjFApW+v1mlZ2DaYPw/BFd8TND
jgqus90Vrqz8xfmbpS5USeZwpkJVmd6Wi5shOZIJbbY4VKDOmPPBJ2+c+MHirRei
iA0uJqoB2CrG3jXEIrwvGZM5F9bNI/hf0NV/lehfS9AASv6FEFPJ6C03ridZsT/+
ao+9gTByp8UAryair0GG2CHjOZpSGgZ5Y49h1XJ/fJ5VMSc2KiRgU26fr0P+It8i
5ceSfwXhhE2WHHWRs8VvBoFWPfrAyBPtI4peCqGIwQnDeo1iIZrd6pwDnDWWrFa4
dpDUyr9MHyq+JnYu1BYMgwre9x2Mjjv9z2Z+2qj2/fgm+3ETIvAVHsp3YkOAX47W
1exixNcmu/9TfWLdbRJYPvmHXxYgTj/XW83xF/iATfXH4jSBYDA6EBCYDNMJtlmd
pthtIGbKiuUhANDHjq1WsXnRLLVwV5r3ODq8uvBy2oDk6GPKLKu/9MZrP/FQfh85
Cws1hejUJieOPXyQ+oN88xgLS6VaQdLK142sPRoFPB02KhOy/EmSS+aOWQDDUJHy
UyXKCNf1JrJUT9WkJr+fe4rNvNRTZZdPeNVQXIO0L0egh0CzIsQJb0OK4JQhGMA6
f7ccOwkRxxDoiGZMRmY6DMFOb9E0WdHvaeHrj2ISoPUZZCgDv29HyEXnJEXlsPLk
fv0MbtbM4fvkJeXI4kpKvMUpXs9ZeVwZDBgDHzSK6OJrsGFdhGkf5t0qyvamGmhp
p0PbU3zAqMcIaEeeao0RxxLYL4y830mhJtOyn3//3BFQr77ZYfDarznEGgZwQmYo
mI/U5yllCmSSWAjV8/J2IWAfucyUh9td9Mu/r6CsRpSPUwxm0lvFS+IKGqQN4ORI
duEPPPveAHSEUvG1ASAS5/0a1BNszTMftJ4YIG3zLFsFBi9MeMTvcUUNM/729CVo
jxITzAn6VUaYZwisZoiLTGe7wiWOu2s7P3ArGM6A+AxDk2FPoqeB6AFbns4KBPkR
EC9cI2f1SvC6le2wyevube+23YyWp7/pSWsNdKVHxNNYXEcQTL6Kc/eA6zGGhE53
soCiNUkUdgOVhfNo3oDNAmWS669vI6yls2oWeqikdZQDCzSh9bg90ze0IGVk7LLs
XClGZd+YvVzwwHtPvESGpTeEJlfrOJATf8d42REJMsotNAUrzsXohXzwGfMyBS1v
7cQe6+neN/uxXIh44A3gYq1hD9+znkWyFBNHjEVyMNSqx8Apz/NJu8OyzuO8MqdJ
hUBAnXDTPHNuJco+LJ8E1w4QgXAK5vZ8D38NBDyf6Kc9uguN4TINCrzBkEF52/o4
bHK7cpwdAAoCn/f4s6315GYBWKbTa/8lFWdeMDM2+uezsvvzWCG7b5AUBNhvfHKa
qQfdKcUBN0sk8vonb+wYMpYJY7jcRVBDvnY0Hj+M8guLw6fMr815uW/MGRMkPwro
P6h2/1RcrewE662pCq5Z+gvT9NCnn/lYUM7pIuH31gZeCXFZUikXpdO3w2T5idvd
kM7VZpEuRTHxZaxLnOmiPzknf5XjXwSqO96gHuygs1pWLsW7pmANP+iy8V3MBuwx
kVzieLSk6uBiyapYnfxNAoOoZtARvXqGFX9wAcq8qjAnXmoTA+tJt+pxRzD1RWJ9
jCZJegYeAhKrh1QWSzG8GM19YL2/XAQaGhulB6w3iPQULHhIwVEG9r4Ra6iAMN3s
yyx+KkCV1FC7ubftsf8H4c5ZG5CLVc90W4PXdRruFTLt0LFDkjZsAIL3/cPRv2Kj
JEsrJwGEd/MIXnu1DwFb17814Al610Rt6L3RnW7pvS15fMNmF2nEXuclrofvUYVY
0+0QHNag8KRtCi8IJgtxvpspnCED8JiJwvLh0ErkuwS58EN4Xe8ZxSWJ9K49bLhH
VgAj9cElkWLkty8lK2bpIkakSIsjTP4bOgApCN94AxEZJh4GGifXxvbad1DtuA6A
0NHal3bibWQE0bBqux/b/NPc1M2uh7DqInQwNqxmfRixIWy8pOJDaJZ83vB9bQ/Z
Bav5GzNlp5A/exsqkM+VQ6ca7FvXDPYraQrh2A/5yjA3xJz748i0KETdpZ71fnNE
GK9O76YIa+dM+g5SkOZ7LVkfCcDlki7YdROAqCFU27qGLHHfQTxV4ohRVIK7dCX+
2Jrp8x8yXFF8LlTe9/kyV6o0iqZNu0LlzVL1cAArFTylTdnyuZcWKmy+oBO5g0LH
M5YURUiKflBjLysK0l8COQfJGyPCKzMLq4R5lFXvMZqV+VyQX4mjwO9n5+Z80qLq
+2R53gPWoeJ9/WsTc95ycWUDdYw006Q8Pm6ttn2NZCZv+lqN5k6Qs0iVrAJgFC+A
XcNk6s7sn/g6EgndBIXJqE20jsUAuBF7VEdVXHZCks+y2VLVZCjSFGXDbSqbp90L
KQDGvPFPebEuTRenQ67PGwP4qNC92Zl5bdbi/XG780t+w4RQkVu0ya6ayrYoVyqO
iJE/QV54fl2N0alYtwKYuqDCyvTw+6LUpgYS1ZJBjI3lIAUp0LvxhHnmzcqxIaBb
zSR2YxQzk9Q/zcHCqYop6jgM5uoWI4Scj0R1FBHlm6MOuKwIdPL2m/8LHCI2ZCW3
Z2462xHdZg/OtbfAIgA3EU6GkFNwV0Gczik8QD9cy8qqM0NuVEZ4mXouh9sp3Xof
EZShmvKGtuSUK/Rd1p+2vU8xKsKBIJcCN1+hb4o76FV2+xn3D4oTvxglVSKaVwU7
Lu+I9gtoiEqVDRrwGdkv3h/tcHfNFxq/fbNT8GZURiLqK3olJ28OOTNUKhKYq4YZ
oEoclaQkePdsUngdkZQs9k53zwx2RYzbc1pm83F0A4yAZ6PnYkOMfEWMaPvw+acv
YzvuGXPlOaY5fndka5xj6f2LBpmBQk7y2QxbevOeZ/76R5tcyTy8x42gjRPXrDPb
nWkMbhjk0wXcWM1YJCiNUDqYjWoYlTj+UqD/hkogTNHlcFeyqAFqw9jyP8ZEYFSy
SYE26myq8W6/lw/eAT+TMXEsuXIIzMyEWNf4Yz5p1JhMNQahgJFa0ouIw+JwoVFi
v15KCCavaCnTWOvxxero+TqBgWxngwt6nyZ3lkXUU+m716srwK2Z5wIRulXsrK8H
hleM/1WEuI41rFhB1+X2whcpXU9/ASQ2CQFNWaWKoNUlbxa9WmvysXoX0YrDjhEb
KwWu6ZT6G/B+/2uTUs8H1vp+pEAr4onDdxn7zDav890HoS7NB13TFI/m4TAzqfnV
Y7T9V28EXYmNulBFE2DAgD4aIhROgMer/0akS7PRm0mlKLb2WBa+KS0FZvA3TviE
jb5xWzJ6Y5YxM23448sSgaRIJ54VJnWmBkrl1Ws0qeTuFRnqik5gPX0nwdmCcugd
R30IkuUUJqWpScTg3xwFJEUmsFxiwQmV5c+vI6ZWlUFbuRIrDixB0M3msfbVipn1
f2WaH9LZj9K2RXouapg0KzlVNvtyHM6L0iRuVKbk1kMd2GGAj/MoQvVmwaTzPdGi
Bn5PLGPhfOF/bsz9D3zPONQiwqQ0HHxwCUzISoFrhoffezveoU1xWejeakpeIvWs
wowMuMCLLzzBt82U6YlyCTeT4GSEsZGcUrV/LkUzalXapsmFmYnnJYytpYAYddCA
jL1rREAFVmtn2vtDQGmQA0zROI9BMlwmZzzVPRQNMihnazLke9HOzs9pwINigg4W
JQj2W+YKu2qF4/PC73oPb7z70gXUXescIqVpyn8iIK7hDamZXP3SafJpanD4MwpO
tH4hQQG6mm4Mv90unlR+ezj592jGxqsjIHHkxXVKTr471mTGZWPdxOxb/Ss5L03/
XIiZXR66zpJTB95znKRdSobQCo0+J7vVtv+houbdRZRLpWEmeTZd8wJZOMTE49ha
xPXmq+NIi0EaRUYVxs0hlVsmaBU9Kl9eZbP57Riyd+uO71o7J+Bhs5WrQ+bocGJb
PI1aewtqWAFKdIWmbZVwyC9hfrBuhmgQnbNOISLU07v2wK9sOp9r3Z05AUKNwRv6
gGC1D+stBavWp4Qk8QMHeSwb9ta04wVa6BuUjnglE+26nVthuYt32toQzt933IvO
V2q2DZPc5VIzrqk5mqrgfhgaa1SiylcMYVRHg/nzjGfEbPxusRfmc8qhAJLVEyIM
RMvsqcZWbRKEZRszuSWvVm8VYoujHn1aIdMghH88iQxdJfd7TIhOXqMB8vx8e3nR
KutHZjaKNqmM/cJurEwexmCj+GseDTDIXiRmPZAnzA5kd2uSzfmOCyMaKwZn7asp
oBEoBs8x5e2UhHqqxuz5lPZ8DNJf0KhnDEntlCu+RZWmPRfadchp1eV+pOcr/I1n
Tb48Q2a6RzBogYgF9+Bv909G6SziM3hAgD8bRj+1H0kVBFqyVEax/009xGGBxTqy
c6Gw43EIPbmLlpWs6t6bQrMLr3uM0OU1CkqpW3aBRT/MDYPDufrWKfUEDT+4l6OR
DWlL4yjqe6YLiWkqne0NLhoJ+d+8W8b4JjLINzXV75we96SZmbkQM0x4VQ+wa6e9
PjILIsMMVCj89FNutaAC06JWWOZStlONW77g9oIJ1tRS78hIAiy67vcv57GEKfly
+gy2mF0iEvtHF3EpPgXXfulpqi+xt34H1GF0oAVF0XQ3dIUOVHugLi7mrVPLT5mb
eFMwCIyt+zgJl7JhZ78fzs6xtLagfvr64zWMWgWxlkBuIayjOQC0WpRsqHEyR65u
vD2DV4mI23bOVyJ7jX0wkS2tgj/eNq7k+s7aBhPKlWOvTCu3dOI8FLX+5P9BnBGB
KfbmWpoQ23zNhpSOxuPCR4nABm+F+bvEvx38q5RrK7sLJfaIL6JAcw5m8J4gd2xr
5BYN0n6aHhQeOGnzwBeeXMAxbdNxRp5c519LFBpH9kxeP3FDnLb+KNax+xyJmA7H
rIimh4okZgcoJsxPxv+vcyOxaZTsSaXMSHfKsgK0bIyHqCiZMoH0ckfKNc7AKHHK
pZhjSn0NiW7mNYDdCCbQVOHJuXugMOrf9aERNc0Wpch0K+ibKZSf1cYoVxldqhwk
DjT0DvNfD2rrJuetR/XPUY78JTmaBvNdl1XUyZ7YJB5tuURF/Y7cAjdrSEhhGQDQ
dCvIkwxvxs/2kYTKYbxAZSoDXrkn/83QSB24R7z06Q4WnjUeS879f9qki1BPhSS+
AnPKxQZ5JL/g2dGqa2W+OWvsslvFnjcBE/V8hceZC4JMfsiU+DDdf7L3fbvz41O7
nTt7Dn0scBpr7nUXoXudGM+2iOFvt3Vji4tFP/zn8RiGJzoehqOgUwDAdpMcZgg8
zojPJHcncWDzsUyH9eJyFp9a6hpjxxKrdR7KiuL78lTljEFRG5o6jdGDR6M9j7eI
PaCTb3bH+zRAjQQEoi1Lp/zSFhYve7z5lS7BLUv75a9WuyzCulEuZZKaYOqPB33a
x7fKw7Q7UNC/7YK/qvcDvQKVxFMWRr8U3bzpt67olLCATeU78bjVyq+7Lz1XnzKD
ndUtovUf+iCszZCPIBSzMgpb6Il4NkHFTNxlA/ESRfxUCga90W7AXu6VNakjekQU
/hMDeq2pFAz9PQ/mZBO2WMHln8bVzLNBQl07qHNyPMA/EI+yIStnfi494xF17OGr
nHcGQLf3Ku5LKO42GrQ1QWx3LntXUOogRe/NACl5KlYZfdbX4VDK5WzXfkfSLEfh
1Kjj4X54OZYnXvWtSNxhCVLXrkLFWzqtXzUrzHEN9zLKIf9IRDa+dPY29/WzIFiW
ArB9jIiVFlyrL2zqfEWRBiuCyXI3JU8NVQQ04b6XcHUWs8s4HVRDLiRGK8WFzooz
t/Pe2Z/INiqzkumJ7vgUM1RrW5+bDMg1PPzWuWSHsZUXH6K5ThdODBxASIB3UPI/
CSw56p0lmx9XGkHlXjhR8P6JrhqhuWYO1S3kFcHpgwD9K+iDlM0sPVfxE02N90r2
7sWZv57FgOLPYD6nLInIQQUxogyB5rg6SLcCnEt5naxODGPoyX0nEDOOnNXACVyB
Z1X1dm4/cSYmc10qwNe8d1gq24N88Bl0IyEc2lY0vwd8da6kPccnklHFnBRrHrmM
RW9yJHdVyicxdQX5YwCkbjL13S5VpKIGzKq0TlddB504MMpUMGTljwL2wDuBQdPf
F97BVFzkWRj1hTEwu9Sq8YQNccHsLgV46CQMSfF976d6VjbH76NmeCPuVCOKLZ7d
BsPqoizC0wjDEJgNjy71PJ07Zf/GIMVhEjNVwC7Nf47dBimYgGx36abXa9XT2Vii
77QOkOaji6+NTTP2p18P3aOtv7mBKWazaxeoCORJ3yvE5E9H0Xb0443ztpkoSBfH
HAWor26M5nzlbv0Uqh3koTFJCmzZwUoleZGXfxFlF7iz7rAyKsM9BhqFk5XnpIHd
sKHJSQil2YaRu5piNWpUyHqCu7IKKEzocJqdI+o2rgBlbHaIAnr9OFHPL8+qGlt3
YVWHrh4u4fm9Q0zyOgCJMFLc1xkFMUT6S/s5OVxNysGXN3hXVJ4hnWyF29+j+oCy
U0BQI4OOS+VAp79EDRTQ48xsDehIcd0TlyEc2AzSzFBg+joargjVbRYG1xQZXoPh
U9x0l+HCsOIWeGRkcU/izqoy+tBQ2NAAwMj+hVR0gtKRNj/O6FzNhrDQ+zkwswnQ
323O0BcLCeh9ycnorzEEqY/v1GOa0uC650RXNzJfTssYwqo8YeRXN2/SWNoerfUh
RhOBn6IurUiWkxwG27+8BKGIe3y71snAqETyIYctgeK2gsaJ5aaiQVVWwPez09PW
HFT/y2jN5bLRdm5dBPHsU3KwFUBEyG8miwB7w8wFFroAv6cn5Qw3nCCuwPJh6JXr
o7swbDgRvsEVmY2F5KLbiyWXNOXw9WU0lYhxrB08xNNuoJxy1bYZlR4WHwqozKrL
ju3/tRwh7ycQCaivZlaZG5bh1UOYvFTtXyZ9zu8z9fw8dZ6CJTtuS23tYAA7zl38
9OjE5qCLoT4Tb+hjYpyxgJBCymfyr4I3QR9jKTwjCI7/uEzMJEuUnNwdh3Wf5bMh
DFHMMhKgYa3zRLVi4P0rTRw4oTi27exJs+VFgUOWoESJc3fXv11W2BbhslVIgKM5
/3EsBGQxaH5h6j18XdyRQxSVmZvX8RiONKFvaNJuXVedr5QeZ1y7yzBfOOR4j26o
3Ua1XwUSyf0W6nUpZ5NWQyDYWmjJLBy4sKBqCDkTtj4QH7fziG0xNLNXwsamw67S
5gZXI9TZx8RbMcmIa1Y5zZADHRz1nPVftUR/8GqODFZ3UmA98dmOiGpgrfJZ2bXs
75yW4FwwhGEOfd1XhXjLA4CciJ8HxWgDyUFDsxiciYnYzMUo4yXECEYy6mjiRKSC
BL2zgD8vQG62C6aDGA8ubrEEQJj9OaWWBfZ5G8TGkPHjuSTL0pvad+QBawhoQa4b
8JE46Lr6rR9kecDJ4V8yd9uvqMmLWVepgPaHKHwUkAH2qGFOIHVu9Lq5baJm5SfX
Vtz4EWJ4Fr00nOWUava499xmmziASL4VEJBjx8Go5GtAGzH1U/4m7m0/UAjLH5co
vbHmH39ksa1sSzYC3SBgG6OUwvjz/SCXnrvKpwQi0WuXTw1Fix5gtKTz1cstxoYw
5CTXXA8TQtgJSK2gR0+UBDkST7bY03viajmUHKLO0i6imeiPPzMONORCbz2PriJo
tJ6loi9esVidT5ztYb/PhvYwiylTCycADlJXBZNgDp1Jc8wLQemUgmJ51FtdtNc4
+abXkEDxsswHhT8TlBoA5kF4jkX/XFiWqKHZzU3mTwi+akVJZlBgGBfxXI8Quyur
G0tCUO+KCRo/w3FUMhkzLVewHwfVx//T74xc1Q6UASATsq8l4Mpowlaz5LPMDe6W
uaSgouiSy2iOgr1VNp5zD7euYMhBmjScFxrpCGa5KAxVXkCZRru/Py1bvoOobf9b
JIvPzRI3EKTuoSxAWJ0aXHLZqUQ8mobM7HrgC1c/5BFkxLGAxtM1U80GeOpJSSI5
Momp4e2fNP7caCZQaq+Ry4jyQsu3VgiPugjvOU3L7hJYnd7clkUGMCLoiAb+KQ5A
jdgRAM5RAPmrsrmL+VkAq8qGtCcICSiZKjWbYqIsyEiQErXi8Sx6xVBKvK7xws8f
QJpL85oiK05wR1l74uinjal3zQjph7/3J1J6fYlJlyXG1Kqdi5KvwPTaU6woUgW5
aTYnFu+nM1WZqXtkn0JdbfC1gHIpGlRjzvStVE5M7PQePPbM1EhWa2OvB3J+4SeU
bGqPe7f7bfAoq9jqdC4fp/TcZfAaFLM3gf9vL6bOEH11QG3CD/xZIt3ir49tP0Rv
k1to1ryUxiDbQ8s0kUa68T1pBYO7T700IxIHIW/KJV/hMJIUTxRMISEYsIPnbSPv
mS2jT4oEd2qBwFkUPN3FXtgOwjbdFIMKd7wkMUSQLaRm1SoFGQieMgn0ceKsJ5PM
l2EoYeM7OPIgrF2MTPTA0+Gl/iiLdjnC0SYjFHivNDkMKCIL1IwURdBMCZFZbj5q
iGCLwn4xbjK3OxOObZl2U9PhzY/9h9VadG11e3D+2GtPhlGs0HbYUXDa71XhDglR
5p4qHZ4fI1B/btxQVfNjAqzvVy2zhdq9yVZNwofnrCSVxgoqylNnags8iqyJmxcV
zAGgMQzZUkHuNehx53CapWa0QGQ+CioNHE5gkogZiV86WDTK3OjfkYN2A0TgRRPd
IusG+CAwGCJYrpBn4mN7VowHFkpG6C74kxNF+WGvCt/LMJc3Iu+8pnTwrBabZVJQ
U2W2nHl+pz/Ii2yYHYrH8GWmZu4e8LE7V/tRMczX4fgKEKHQTOJc95zk//5dPQon
UgAhXlty1wHQr3iXzSRecd1fpf2865ixxXmW3MrfPJBUq9Im1YDv3kp/aI3E/k7V
m7Om8pOCqgqvd1/1yDKt2QLPgli2AZvWXDo1I14ds3xgSSv0mdf59bm21UaAdUGw
fQm05XraCS2WJX2HK1ZJJ/gkPaJZvMh+wsld5Ro19cNVZrEIsMUJ1iFXn3w+Vj63
lxFp+uNgEeJx5TeRHaGOjZ4WImEQItq+zypbgQ6uoZ8K2kh+GSNWrmQFH7TRo7rU
DfRNdR8NdZVVXsf1h6MeM0MaRNr8918yr1UPgpMK0ePiueexz1kljMCokndAIcgM
9R+YbYQ9PADV3EwAvFvO5y44OBqABS8YvM7/WxYIU2GJh9tXiUZL07lJ0fEjBEaV
xODjpz+IGRdt/B2RcDP6iPMcfgTQXqdk5BxSkc/EwbvptvrGOPcWD3CWZx971kkr
NR37tgrCTdlI+qLklVcwVHwc1fIp/O6MOTF4kZt/W6tRyj9aUDfijbcLNr0qmuNn
BqrGHy2UBug1Q8Zw2xMyE8+aUp/DOT7PnIapTX+ZEssqEnfc5iGqA0/Sbctht9YX
NuA0OiS0oZ5vGGKFVrbcKSyFkAID10pOoCBMri7Ng2RzF5/5fmPDyiOCorF1tn5F
dZrY1oXJB5N4NfJmIqCwaSub/eWmGhCt5DipkBfzecpA2rcT4WFTJHdxUHlglWBI
FjgtjNYNVUjju8iXxTRoRna5sLmYtOqUjcjn1SuyyHaUYepTAxozmmrLogS87Vpz
rawyPK9zGJE8wTxs3wl1ldF+CueCYRmxGm8gMEKtQqZtz9XCCPYTeUvumFrtzFml
bpkI2jt+7shEsyKDP9VRu/RvCDBfjdewFYqmS4vzS+gB6ZHcff8Hgo3rEmU6bqfK
CJXm5CRpcyd3MCj4CR0X+qpbdxJGw8IKOMSPCeexNvQN4NTgCALlEsy4zxWAUxLB
8t+fBVKArOGqiUWY6Mmwq+p/RMQ+w/tDtkpn/Pr9yuFxXPNyeXxPJ2AaNJDlHmWe
MAY6LSFE2T34oeNQ7SsQmpLKw3BQz9d0nSpaGEwcMMm8lMfOQ+Jcm/QNizgJm1Aj
OIV1w1CFwan9r/ZTkh8XhgY2E8ORYdni/yhW4K9gt/83Jxb61VmY+pF3/FV4oCSV
TuLNTLaWbbFMqD2dk3eBcS2CMQPNSDcQENW1APX2Usck4OjvXxluB7UkNmA14xXK
QhpKpJuQqt74T9VY9UKqIlPX+7ZWV9juIt2DGPpXWilub+BdMr0OAbbx5P0OasoQ
mZ7hbH7lOKUyiL8mjZu23UBGIXR8dC1R0xFi13Fj2fHz3LP/TCJ7o1kcwlWOWnIL
l8D+jcEHnCWduDT4Y2lyvrDiVatjRWtvWqiFtC03DdnPc1VLA7D/rGmG6z6DeEIi
2LARw2zqe1IndwB60p7d2WLg+xbX/Pl87UavZHQb9I2Z1tb4xOLBG5HI2+Ce0MMd
UF1Pri9/sqroyBCuSrbHx4+Sw4jstTL+OHbIoC19IrnHz4Zjyp4PksLx25JTSGEe
AGaqRk8jG3ZNPhRfxtDJnoe4e3uyU6EQBNoP86lA/zxnwW2IUJAaSpaqQClj+0yW
4gGNvXoLGChfC1g2NDl6OzMeBTm0GwEM+jPAsyIGvzCBk1v5ydpcKJTpXyhfO4il
LrZ87D/vhqX2+Sz9DlaA1r659cg9xacXu27s/R823nD9OTy/sP9FBg2k+Ojgyz7H
pHGzdYHVGrCmXb8kcjBR0iXYW4I2rIqipziPhPCAzLBDEprTEM++kGzXLre+9Uvs
vz+aeucU1jZmK5Z8KXd/oCSU6vC7rwxPrwj56MEYJK4IQ0Rs1hwIklh0kqw/mkQZ
RPTEKmmCdF6tn+aLw5XQ9m4t7eUxQWav/iC88jbpfxO8aZmgUWpwHiZVVXWXP3C8
V7Wae2AglgRarsjQlLE4Jzh8TpQ7xlvHq0LXw3yKdFy4C60B58y7n+C7ZtHQVx1q
Fi18UET1zH02eJpWk1uT7TN/M14RmIdrKgJig2m4xvNyy/l6zqajfnBSkgLAg48A
rmis5/Z9o99lihmAcep2usOnxPy7flxW2yYcH6r8RVpMTM6xivSA2wqBpb3E/4Ey
Efby83yCZfUnWXEJBzzJFmEUFU/4S26CN+pzhygrNcpbhlCqkpl+ajbUTU/L+joU
jN1AzTvzejBbu+Cj2fDvCpVJPijg3lWyYOE46PrLrfuDQvneOBZavXUxXQiy3HDm
usWHM3RnAZJYYqKEUyLSi3+/5E2Gxi67sYeNQb8ixDJvY+yh+T92rN0PO2F1PuCJ
hqd4L0Kgg473PaSbcRvhx5x3EhAyFW2hlyAv8ueqC82MuZMsEtWYRph3gbOLZxfS
sA0oK/j8zareHx98gw5xcQq1TZtdkrmPCXQ8fTrmAV+TaOElANiq81abGR5wj6gT
uzqjAA/BRINfUH5GJn46zISN1EDgrPAiJfjvbEiFe5NBRR3q/OqYJj/zq3KqyaHG
8JS2mc/xG7jPClfStIuOwYVsa0sRmHvvETM2dQU01OWvJpNllGxX+QLL32rKROmD
H+RpWVKpb5wys599aAc5D1S8gw1/VDlNpdeT6RCk6bmDT8tC3oJE9pKtK8bJLAZm
Pcfn1nBjVNXxUpYHeHd5MurYxqb17iCkH1xqxt6JTVXVPt9ILite0PE6nkQ+4a4a
gcWXVJR1YUreBkgXXFmQs5AGqNDo6+gipBLi9gWP4WEw5hw6Sge9T8Cnbp+2G4Bz
cHE0Wd4TjZC/Tcg1pMtLJpu3M0erYzazSp4rsx+PA9x3nneIlOvkQ2W3Rs40Osh5
fIQ5p65Llv4uVgAdoBzWg90p1RavjwV3D8fAw+K7gRfx5u3A5ZSmCaddYSOz9/7h
7ai/EXo1IPX6admWGtYJ15tFSeRkrE0Ez6P25F0mSl/nrNVJ+3Zy6Wke9z8Uj/yg
AioKoQ735IeZfNqt/iTdOvVRvgr8TVtOnXNZKGEGbnzY635hg7gxUyT9YtbwIgYx
DtEaLRIXfubNexixFuk2XccpMiuCR9LNs3+AAnR1k0kxsxFTM2qfziiqfMKZHPq4
OXr6afm2GA6iNRGBXMVakXN3Ehie/lQSa1lHRN2ItXeOiU76NhRKZgb5yWCXWzQB
/NAwJPCP3ayQFlaoVTI0Hi571jg5FYfc2EocQpURZU/1mjc1fLXzx+UEHNfMhXfz
Axmm4bexiMK1GGNWbtCTR4PpvILoWwBklEckWa6cE8+Teq6cEFmAToxv0T46DQ71
DuGBc+432eH4g5sUmhAtUJDBqqQknrGeDEDL1mkKo6UlRDBzhxFtva0RwzjXVAdl
dvDwdelwlWtTFLII0IgKcOxVI2Qaxv572aJMTdx3MLp78mNmAvuNPeoiNyf5MjRC
8Pfl3ENWb331t/NrShYrP9wmp8zldhswocVUEOBKVYwsePdr9v5I5s8FdfZ2uNOq
eFzDf+GDsKZux06irWCIU+XytTEy5JeOaT7KyLbQTP0Sci6SUQL0IN1fEDL/3Lai
zo/TEX5Nvh9/oeVlZGvjuAeBqL8jWFW0DfB6gHVPrj38yUc0ZpGkkDAtCrxjsOJ7
5tKw9nS/Wzm5Yp0mFEBqNXLkrv5Q6IqaNzIJRWj2d67g0Hjr6uNKyg+RF599BWFK
uGL3wuU+doaFrHtFIEaAL1JSb5Dw6pA+ozpDKFMRrOvS8zZNCyHQxYbeTSvAmS5m
ymu5VJkPRzVHOcaB0RMSlNAidLd6t7rSWSnKNTLKA/RjiflUeIFQAfD2dkDzOjia
yIOdNqWR80fZoZrP1PTVWctrwxJYe8kowgkhZ7TX0Ph/BSKwTuCeEwRdl5G81DVe
pOgAKRe8b+UHjraRgp6eFOzODlckywEgLNcllpBBVVFS420ZrAPs9TqjURvwHpoM
f+DSFvNAq90TzUg3wPT3HQtUIleCTiR0erfdCIUH/MLSAsSmN1cASGf1A0jnpA4M
iX/X1HO675c8uURhV7I/JlHTw8iJ4/Moz0JEgDxVbNv5mhKlogHHxmlDAIelsSth
NJIC6y56xEZoufPylQOcviirwzLlKmaTgODlw17UO5AS8dKEYUaVra8mKPeg0ZB6
U4hi50qNLd0J7ZLvpFSbv+JZU6oEsayGyjHCBksU5CyeEEVswcKLVBpG+VESnzh2
JJIyaGqnUwNNXPqLvIUvOA3Go5zJgw3srHZjVjCS8A8m1OIK8e5RcsB5tO2X5bYO
Ge6laSAr7o6roWTmZLiK0ZRdpXxedy9yMrjdt1uUhSKPDHC5Xwz38I/4GCf01khm
z5gUyHpY/vedpZP0rb+UcZiKFDuLtdXo/Kh5aL/6+dzRhmUSGcQcgj4BPSzxZ39m
8VgMmh+768VduFAw3j60KW0Qv6s7vrJZGJI4ESe1ZpfO40PSPgk0U4GTCLERI5ol
iZAxeKz+Ybl5ilKANr17MSfeOQlb9X5W8RXh9ggbNn5RknAB7NUm8HjaMHuunRHL
lvkrxrbmrz2nlUl+b14WB+sW3Lnk66IeuuyrhOtua3xovpm0+R8mdNgO8W1Muk1p
RQcKO8TFxpwsMAYv9vKEuHJwGUj6105t6tPQucMjmDapIKyRLAW2zCi0m4cPN+8a
HImL6ZRBydofU6mVh3k9J/qZrMyPHc07wO81/KOJi8tldgw+Sadz32k+EJJ4gLE8
VonPaLkGo0Nm63v4TGFmQCJWMDpNMmcTmZitGK5R8Kw5is/oBnZ5mdrjQVjE/Vns
+nVU+i3w4iF2+tPid69uUzjrpNnHVPFlOqbzdl2Klx+h4AcbFzQms3viDDEF1HOp
fjpPHttlwpZHXSyPLs0FLXrnuiEzCSOlOYG6ELfypxW1jJqZgFHY+MCCn1L/0ZYW
tAZ0w3SVXLwX3MsxJNlQXINUKwGkHQ8fTMqvOpSHVxc4KOMK5j2UbEJo71I3OoWh
aXBMHruM7YTWs21hQBqdyROHTTBwnorKP7USsktSL2MIZSeDKGg8HARMqP1OJtUr
XZqvHxZN3BlMYbBOjWXILb+BbERpz8HwcrTeU/eBK+iDjpEezI15jLB5DuQYfb1u
Vc9MkEVfB5hrWDeVtCk3pdxZwnZu04kvBNE9JtSFfU98C9np93xnJ3l52XzriilL
3AbBolR2zYPlSYkLkTRKnNkq/PtnyQpnVsKczd0eIoUjn2O895P1Sn9D3ZW8ZDjw
Kou7YD2lsEPOMqqr9KUuFr7+nRZVC61iwAYLJISO9LD/y51iC674NJEA/fAT09Oa
L2xdflMCScBZBT2dCydulBLeTo3duq+iHeYe7qnjT6PQUbWALb5RoTyGpEDEcNz0
/Klw72XRAwUKIpOaY76nneXAH/REMro4s0AtebUDgzOG4zmPrATqKx4YhHUK+HHG
Y+vDOFMT3zcHKIr2uLF2a0YSaIpbuLv1xPlx9bpbbpG1OLr2JastSqJ4N+i56niW
XZ67c2hw6wUQfd2GZrZcADy7dfT4fe4foVPVNQ4adnBvkwIVmdbaBxI/LkG9anTP
5yJyvtsavZLtSAVEf29UNX/hM6oe7ky7tu0X3b8AmCaRcrGc67ApR4fNbQ/4sXIH
GcCDCQ7Mk7N+HLEO1elhgppGvxMSaCPryjF5a1eYj4rSfq+pkawY6Q1IxYHU+MYo
6/WEqc2z6QqmuSxJa7BOwDgOQSQr+8k6sgVGru7YrQsGtrqn/rKy3BPjL6NP8BlR
XnHjvvXzS9YFCLniWrQK5EF2sgPz/fZlsI/bIVbiejig+gdABhRN7q8B+aliqXvl
T/d087x++wRze7+2BZQrNY/VYQYBPMwCDk2IO3sTFAyeCuTC9ZT08uQUo3lz/1qM
GHShKM6dk4FcAOK8ZvSYtzobs5YFaj+Cl2aaL0/4YC9SdHiCptrATGagWxqXHrN1
MmsHlu49vCP7HBrMdLQ2SDDaL9SuJ60+zgQL9A1nTR7/xBkhZdfO2752CF8aPnyP
hCkIoQCQzrn4mX0ey88ocDkLCVTs29gruJARoj21++ihxk5pzCEPYUJ3VEWlhQks
zfkX9oRNpH09x19BD0k2zE1pGfuJ5SQoQX8otwpW7lo3Kv5QpjRv/9UJDn2pSBJR
s3RmBSdOF8uuGX6L3eKu0rx6g7nr+KcgTNJvdd+YIKWcaSOhKOjE74mmuVn4PGpI
vdJoPq/oh/w9YMF8S0+jJbHI0PjSmIWZ6Rj/KYu1EjtE48+6clHlpRtDYABkPy6X
7TD+WMVRuT/Rn478oGoUpU1NQxJZPHDsdY2ySD7gqTISS6jrhCLAmfub/Wme2Gjh
Oo0QTT2tAZdL2mFEb19oMoSQWxE2tddyExlQvu/ZNE8Cf1LEVyGCPxd5TdOC0sTc
NB4BNttlD4rvQgRQQv7jS6fOqhqYqMX2tSLsAFiTc6jIXhKzKdWW4kZJIuyR3iDn
S8vezqiifSh3WHj3NEXRTJF5qLB8wpfZZfcCpuHMFsIRywrieica4B5rcuwug+l8
E3hc3gSibF12cOHIq+BPVkBSTnT2yoq9zA7c5E0ugTRtQUpCnHrLEBgv0cfv9hxC
9dPJqNNJdX/jai6kXcHXvwQ0aUiwnc9G4v4EZ2KvXHq3n63oY7p5vLto4GTQCkbK
epRSNbaL7X1Ye5sLUoXiJkMFMtNYEcBtYhYh2pSBB3ENaIpYQe7IR/hy2oxlEfVd
/pWtstA/Lt6vycMx48N5g6hl3dtsDPWbQdCyX8ySIayhoZg6MmiJBnqF27tYYvkh
DTw5dw3LhZJeQhQm3Co0FYgF1baNtSGzLnFA42phXAuH+8CWZ1SjKT4vGaA9k8AL
tskRBfTNL+4WeSDPtQM8C3naT/S5c3DHdOB2pILTRQULX8Jk1xVY5Aiq3E374rtN
DNHG1qulNfKbwzh5/1cH49bGyO+dvwK34HdqYZ9esyt8pZ/xdnEPnltCBNyjRf9D
JFUdjCwOz+tJkX5oMno8K+bD4xo8qXsIgJzBR5UBYoyDgzK8JIQj17NBwN083jkO
tEIsIC0m35XXSvDoGhcIhICZYCQJatXo1EbJemMw3FIj0y+ppOi3bTeTaImaRF1P
Hw8wsD9zIZpN9TPBjbw4bAiIp59Sr6N5rfnrlC2H56rgYJ62V4A9b0xIIjcobe9W
AsBbk6iDCHtGyLt3j4wXQS+eNkuWTV7mZKouShr/cWmFbcShN1apNUvz4X7LNd3a
Zq/+zCaRrmDMljrUv5AwXnwqltBcT9KEQR/n7mhNCXPuR09pGG7P6wW1AcKuzWVS
hY/CrdphJdFgw6Hr5aV+Gjd+0kbFnOYF40jBYpvSM9DVoXvEpWzt173NzV5fueqi
K4HquXSTH6VvuHS+eUagWq98ywj4sY+QkoLt2XQzPYJHTSRdXAyp3IhaGOPGG1Gp
OUIqbfVr8cTKr+5eYq3t5FsDiI38846jlg/z7Hf5nPASrjiwiBUH/yLbDII8WomX
Nd5q9vw/lwFOLMUayeir+wAmRbctKGEW8JuswmVi7za7tDqL2HInhZeTGGu0AZo5
gC9MdtqxPL5czWfuKzAkszcjtJ5yyqOLZnI2+L2P7qTjLRL3rS9JGJ0zvUeiIqNv
FJUUwLRxZ3poWAr1qt/2sPdZGaZQvlnIQQCgpmMmuFwg0yODYl3ed1Q06sD/bAUR
uRchCjaCGrpoiWY7lNGzSH3wsHAJxSNGYntdPaQeKY6i4+5dxVe+82HebKVrfoz+
UbAFmezKF7IqUms5UftPAMHaw7ceqBsfe88DioJlZ6ad4M0oEjkQ29Bc//ocxXWY
yotoR7QA7D6w1YM3wxknTr5ioDSAwIszmuJJgIK7uvqD69CSATOYDEOHjsESQL/c
j3KbAGrLoIilf45ZUOQKvke1r8W1YUvHF/VXcJV8nwuP2ieMe63r6EKLZlZ/wrS0
TX4aBg5YNRTl6vkGRvSL0kOkyx8U6S9MXgGND2rrJcO4gvuMIjaSlZf1V/iXYOae
Dd1QpBqzcf14hnO2Y5nr7UkzsWr/9493GqR+Ec02FR2jumjidqQqHcpS1y5z/8hN
UMcQlvZSFCOs4pEYrsFSV5xABfH52369JM8ajm3aeypgAFaHM8phO71OmDqUIJhV
iD82XzItHwrtxhQuwfVUGon07azXdiNKISupfbVfLvbCTJLQLnV+dyVntIxXVQxQ
komu1D3+zVDDMLZedhJxX73wc47epMszBbhdIfi6mzygQKwedsfHIFSaYaHIE9y6
ZeOQtZSpJKlPHlqnG9wCDKpR96/KdwS5v8sxCslpl1cvpyHdWJ8k3ClMRR27SCxY
4Zra+z6dinnyJ3NJKgX2z+h/Y/cuwYzkk1rr39hfYo7WXVQZUP+g6RCJ55U0XgUh
zpIJRh5dCb4qD301GDV2YOqxpcUWXuyTSL2vov/A2jO2VdINxn/Q9c+3VUz5FODz
wy+pxYuNHUvBRXDOJ1qaJyBboVrMFQPq1YlrEYnOSxa+4dwKFpFn/v+HNQwOfwU3
gIwaUtgRzBngEPAL3weSA6ZOC++cLDgGFfhgGr5ccb0kT2Aisjh8Z5IvvEkGkll0
8JY9003ylrkahTSwqlB9/87NGr7rU7ap/Br0IJ5xVYmb53lZkpiSrSdZ0zxW2gvR
rig68PR+6/o3Xw4yVLSZnulCCdyI+Dtdq+YcSHYaio7yi5w2RVokq4j0y/8X/2nl
f0Ukn7Lkb5vDjdTXHDqcQd2dH2mhbuSYXcy/IN0kUla1VjaM/fl/wrfj9tlZuK+j
a5+Tkc2L6+lDxEbfG7ahK2kASSfiDSnnzIIc9nTAOojlENJ8BqX5ykp26rv75KV0
Svi7FFcE+Uv6ZgT8xsjN4NtR9XYWsWAWBHlT95rlfbS90zxF6KM3W4ST/MDb7TGg
N5QOUObAN+KuynmJ+TznfJjXDBQw9TKptZ9vwp0xgOW0Ba59qDgoJ5Cyrn9LQVP9
xItq6PIdxwxvcs638hvy/tgzlnaBjMZ76F0jtw0JrmqGwwjQw9vRE6w8oGpZoIy0
731qSWBHPpTDDeqM2PPow1eXL4Np5CRBjCFw48829QmzWuBSaYzA9C7HVfgTFd51
WIfkaDUl4Daw9XxNFKtThGX+sFzhaWnKyvezrvMkwhUdHvWn6LTILEOgBsCsX7OG
b4a4n9WBBtD6jHSSugayas0UwsJXGUWDsxToZSyeDFv6kyKBP7h3K43dQYPDI2g1
rJ+p/TrfabZonjbhqezpmEbkgc6MHpKYXbYTciq7D1Md3tE9I1G9Lx6Xp8wcxK6n
7399o86hAaT1mKbGnD/91lVz1OYo5kRRXS8ZK8fywA0oALMBWCSBXEFMB/+yHcgJ
3gq2PdvMPwe+xWwCX+A+OXS4ml2zIjhMzI7X+R6w5elR8ny6o0jl6CrbvAv4JqJI
bD5Vz5R/75b1vWXWU22d6ITpDZYz86UZsPC1KKOWHAoZ3reJQMJxL5vGy2ZNhFkY
Kk4BtM2OVuokrpSm/yJ7VwFIJZ5p2Hpg9BWWeq7C0fvOJpVrnrJh9dbXD9wO1Gif
9Hoh/XkQnY40lz4XxJZtEeaNwe3SmCL2zHCwzuFlxGdMf+2yEzCgVyHEPt3VPCYX
2fgh9C1GC0x2J1+t+Dhr1Ypboq5pmukeWeiaXVH4LMr9IvHkA5r9uOo+BT2kILsH
r1egetMk1AccYR/x/Mvo4MGjUiDTpNmL935cV7GKo85AyTbKPi2H4ipP+OznCGmB
jhVGPxf2aqQIEqYFaPLojIHHNl0ZsoeAWEt9kSrSZ0kgkp+iwmvhUjY5PHxR/Yno
Yw4sPB131o26QnEd4wEExbUnsMufNTN4OCLc4tCzIZS72Gn4p0z4O/h0y7kWrW1D
F+WwhFi52+fYuPmvYW/gwYurk2dC8uRcOry9No27Biy4v7bT5vgUSPxex9GBmNGt
BxX5gJOVC0U+canwK4f3QSVMiKJOxj4tzPGdJWt7azv4asYit996dozb9SBhuNPg
NsGHwvlq4FDG1+50d92WqBaBQFsc3ja4ONAe88moD+pLB650nF8+CZf7fQrCa7zt
Mx8HOoVoKkdSGlqlm7i4JfB8nbTaw2rDKx1EWoJp3FlnG5WS3or8ufF8cIbGWYW1
YnBfDTYlXT/7HBNrE0/MZYxzvoKTcYCT+57knmoRmW69oX9gZh97uAdEO2IJm/Nb
Lh8P2LY7H+RdR94Hr+OToZgP1pw+c/XGxOMJ9E+d0R0ww82TNC5HoxTbOW2WZqTH
GBBdHGkJ7YhMe6fuAzhRL9BVWtewfJRWxwskoPXRLTygul295wTJ0XFnzO6guutZ
ihibEvNHKj+qdr742+/V3x1QKgU3R5wpqmVZN9YunyQX+58DKI6WmhCLn3e6cL8S
6znUWkPokYiMI2JV/B3RvqlgpBTimzvwGNjZFyv4/q0ytxtRIR3UiFvKlLh2IGiF
ATuHl9GPft4Cby8sPBhIKBjQfKpO6roXGNvydL4xJDpPZ96kP1OPEt6hRyM2gFBU
zNSRHfvA9gwBYN+B9QJy2/CvbkycYEIrdHpZCt8hCiF23eXD3rOHTxTk7/oO1Qka
TxI7PZ9HZE3RTnStm32T4Xuik7kUpLsfB4/mTy83qDulA/I/P6omqpOKAY/mzBDb
+yI3eLBITALtLJT9hLU5aC00O75dbQqriNscdPAFSdzptbN3pGGd9ldqJi1ItydM
C2e1kWLB3auHqggOYNp/GRmGEEotR5bYUsGKxXKx5EKF5AuDdVZFcKuCDIV67PXl
TM+nI7X5yZL/0n1rk77TsDAGant/XGyoHQ92+FaBbh0RdZqjTZElk1zVxT6OolDy
mCI5tZFXBnx2jWGKd0vjbXsOZMT9GX8P26Kv459tm/gyttGRxMk+UzpUa0dnswZu
Q3Jkz0R/Ekw5QXjvt0iDW7mfDqCpBjOj0WujEkd3FllVfgAjGNY1nh7NcNtr9l9g
2op/1npYMo7qer8Ayg/kU35bS01CBmgx9Ya2s4edWZds1vai6dZtug9RE+9Z4rjK
21+sMXNxAYaQMpf2lH402zmMznNPp3ISPZayLMxHJoqiplY1tH2z1mje8mqJD+e7
7HdmUXN7yJN+8XPcQabkqvTN+d/G0NaCe9MwATw64PgVMEVNTxpm81nWYCLrUW1N
c94Sl45fnjqvMB8/Nmg1yDlVIZ6fUkUSBhlFjPNas+n7kqaNZDHz3+fMMxvk7PEP
nnJr0w5g6Ziu9di4VHjS98Ovtbf/qrC6SQlRFZQ9DDEWw1t1WLRhFD3/6tpVriZ/
t+uwlwizupx0B4fTESZ7rOMp5d07gH3BDGTaNI6hFkOz1sT7n7BGAhGsDnJ9LNzr
MG6miKdHaMaHnfcoxXPV1kkZ9/5pTjZ0oYawuQu5e4l6LgcdEEFw0SW33kuDxQ4p
tk/lSmZ4KOxpB9KZ+KTC1tAoejDA0WsHS8+GOWY6Z9nNQ7IQZqA/vgTeoLvAVvOz
t1iWiWWOPRKy4xLB/1TeYmVn4E1nkiKlaPGRtxdwM3cfci+6UzFRwnjXaaj+Omid
dnlTDRIMn/r8ZcjayzCOx4qnI8Gy6BoVZBqhGo8q3iFx750yDts8pBjiRK1BxUb0
0fuqjK8IhpZYN1idlbvNvVrenQFjOQrSG1PeE8N6uhei4MGz8kGeX9mM5tq4DaP8
nKKxCWDhvU7a4HlEKOvjhFEwPXcuGcZM7g8H9TPElsVv4Y5WI3aBftwFcLnTb/xd
vQS0LkaVNhdYpfHKOdXJ/Bj8NYUTowPUN75fxqTEEcup0Ymqo5YPm+HMh9X7IptA
bmSIt36dxdx7yaE++sFPFAsk0H2DXJ+fcnh+EwEILUVMMPQhGvttaS1+72uV+Dd7
g2pBpAkihXday7FgAla5VtnnFXP+al6WMrG5FOekMUJ5GA3ftsP7AgzVJfLT+Hss
d1z98bTZb9F4dehlyTk/Lq8n/pkMaPoeoDAwILuxY/RUS+Z0AT0y6pwuC0MrXyhd
nDkrMrtjE1EQJg5zHA3uFQjpNvvrS+iVtupuZCWqVIGqYEBPxSKQiXgvyCbDxrC8
f7cnXqkFIZl6qxAiy6c3jN+jNhyQdAkljEXv2XNMcxAMIR5qW03r40lkNNvpxIRe
/uIh7Fl4eM7Yyq4BOgGL2rWooht4x2FdU4uysaWdPCN7yxzwygw8sQ0uYW6xlhQB
pN7YHsbkfqk2ipS9sUiTle8xNvudg09YlZEPDkfuHialXLpFjLZldrUgoWx6a+I/
GeTxfYL8/JKMM5osbM4Dg3+3ABypsOc4Qugoe7kIsy6ngFSlRJTYInvzboDIQMTd
1Le1+lAeQTaUeY/yb/6jK0sQvd9O6UkRo2NH7+BNbQLhz8LfO9OglkfIXZ1Kr6XJ
O4VnYLflhj1MjfSFDxYURbNPaWfF5TMJXY8rwzL4QdK2MuqjGU9WxlhlzWw50lAi
51RJ3UNavyF5QjPp5bxCttov9JfpG1phkoLUJ4MCnWBDi+APld3ap9rUE2O5MBT2
q/9RXC5n1v//jK8blnF9r0jUxdN49N8tGcUfclAvQXNpuMyl2bhQ95+IFnSRrKNi
+3UPFBGsIQxKbHMVyANtIIXe/VkwlkOxfQwsd/JXi5JJxVMkZpIOJHClg4mW6tri
Fanl3WTEHvDIZHkQMMpJhA8F21Ua2gSnlnV+CRSaB4UIXqdFN4ElFJC18LRhH4Og
AzQiP42ok1NNrYUBMxRLtPfhbzVkpcSiSzAkdRym7NuQf+AnKPxB9TQvh27E5xxJ
Os0R59hidExIQh8R89PHhl0TIZkyFk4nmpNbQnYqVbJ5FkxZU1F5dIvQUrUFLTA9
e506knBm3qRLTMH2ifswJJMdt9+wV6ojsoeHRmEYSGkPPgKdmroZTzh4DveCmO+A
Gc+BoNkTe+nVoOp+CY/wl9tjUP7zZNgTZQWNwTdrghylqPcUNNzReNLZAn+Zx6BG
ehLg0UWzvdX13KVkRuI6D5HpQmSKHvXZTseuWp6l41dWULeCNWJek3mfPZpqNJIp
cOnlmZjcmqdTrfiTBZ4KjMlYYJhMq9d/1w6Vfp7yp81m9eOcIE97zDxnZZdbxz8G
FTgLC+RgbYSmE9DM//FX0MoiUb6HXugu6JcOs3Ep3t2wbBx//7SO+YSFXz1Rq/Gu
meHIPDSWzFXd0OYPzEnKsBg1kvTsjnl1ATDw0Xq286yDys1AFh5LDO//L/jfvyKa
7w3TSSdZ7es79yKlG9VA4sosV0LOERe/BpNwHPe7yALqmWglvtCZnnD3YTgymEz+
aCuMZ2vOC+kFruIfEknVrw23WG6sSIHmu9n4LSCuH0d2pw2l/+/Cjs6pGRYTMEAF
J2aXNbjISHBkujw206yGaF1mNvRYooAyTsVlIknONp6Vs4LwnVoqMc5hZhNk0zmy
gUjh8/0MegPx7ujGF/EArDo7zyKyemxKyPd6yWQyMVaB0hP5VlQBtR9iF8EQtCSA
ZS5P7AMuqmDhC5o+aGoPS7MWOqR0HL2WulZQhrDlkXsTvwKTSgFR3rk5klnVt3N4
KRYGYWiMMyLhlhyF6xnKW4Bv8uE2CjqW5UELw1Gn9Hq4brmnBK0cPdKGD+5c1OiW
ZTGzFer4PRMhg+XLtIvpNSBgdIh1MUM22L+HnVYL2bTmsr4ih1V42BrfEHP3uFpZ
HTRaem8Sczw/2WgqcSvfJEhhi7XmR9j7HiENErD8LqCVrdc2IMeTFRI8xNFJtWLs
MRDYkDRLaCduZsID2v23irsK3V3zV6yjXeMbsdRbVGNj/U3eF21npXVWYOEbuK3Q
VgIs8YhWp/nAg673RDjlyZysaoRbQRpEQKeMmi9z0QUhoLyORvftnvCcicYJr9H3
gcCdl5bBFY1h3tzr+04l9n0y/Va9/pcpb924BwmV3LCS0reY6PIbWiCrid7yvVPx
/IUDuzs5J/hKoY4yYXCD3oXlpVimDKjIPmBPmq1nMouDn8pewQIIM29HpEmXV6l4
ZZKS4T1xWukWT98+guqtP3GGWcwja9yyE7QduchF6Y6BVN8qOtnEOmgCZVBSNTfw
oRnL1p1ynQJm8jKV17Ud40m3FmF+TnD8kJ7/LGcFb2GZAlGY9lxG6IIEe+meK1rQ
9Isg9k775RyofBs1iMbS+r7yH98tIvKqw3iiUK13oMrgSwrMuv2z7n4ruvBlw5aa
M2fuMhOAiEuSiYy3W9LTbgO94j5prfN2j2J/m6+P+aYkDp2jUuOI/vK/ZIHRzT8d
/+Z5S/jGIrJB7wgTamy14p7+OEuED5yN+bMtBOg6MQX9WKAOQjsxy1r88mQER5of
1C2MRcJDQTx+yFQzvs89wB8lv+liUl9ot+Q2kDg1VwF32eCwTSgj2z+7WUSvA93S
XqvlGm4/TwwqSlWpQXLjaSvGdjr+uBlaf9uVDj9TbhKNHEwpeThtAHXEqPSdXm+u
IMM62TRn3ZOWG2Wsbh65b6aYLW1d9mFys9n17Qr943YBknWSAQuyF6o7nc5R3K/t
o+gIWIsb11j6UpZ8rxMf7KXr21q1xdvntN6u2bMWGTYwFTLMiKtChA2TOmy9YENT
ZsI33S/oONwOQMxE8pW1ZASU2Dx5Dsj7YzAtwb9QR0XCToqbs3enjqkDT5B2VSgM
BKE+YKsFUlktQ966ECB102RISkOaXhlh/WjY+mFtYlL3E8lrsN3yLxjPD/MgeTW2
nPULpINSO8smqKIC5wasLnSHDQPj3/M6B2rmLeIKX8i0L4H7EM9rYr+GtOrZb4U5
JCvr7SGhEpaTzlGVayV7dVV9M0LA/KHbMu3zIcwwtC/F3cKRM0eQdYMr2RX0tb1v
Ox5jr08O5BaGbogfPuphqA8StXzFC1dtlXNQYq565vN8ER8MbrzA3KnvfWFCBTiE
vkBmOf7cmw7lYt11UbMyrmn/Mb/884hO+3evMANP9LIm9xhCY0v+GTU04asTOoxd
h+sQYxDAPCXqaZFsSnO5ZNFHvrBeyKnFv9xtBTHow++2IzFLIKnqOAUIv/DqYwzl
hJN1EuYWrmq/dlHJeuWf/lQFksA3QGHLpEDrqZb4qXCv4LCVgdFP1hstJesdoW1O
0LEdhDP4yAH3NBpCqUOuVe5AKVa2QQon8uxdvLak64thnyzOag/Yf4QtrYgw88R0
FfMwm/JEmE+L5WFdnpSkAuP/bblQL8S+IWM2cYBQyp1QvZzvfym0IViIijjR7bzd
O/FEXs0GmkQKLtz8HK42gCzWt/8onkuloPVsOAi4UbgyNLyoA+o9EjQx46WT0Ynp
hPLSmcnrKhRmwD/UPGebln1rIimwU0Tq1n55Gm3klYb7lRnEgmY/pP0r7GDen7SE
6uiRFkD09k5QwOb1bDZdxaZDK83YLImnxU/L8o7s1JveoSZDGg5lae9tuz23gUTy
G3Y7KqtsfWKa5dT1S8NRZw/kLEUwrlgbcsWq7I5KbeIXwH6m7WyiXgetXc6i5HJ9
iRsT3uI6p8jwi+dGMv9Odjep5w5BCNwpItqa+KDFF3H9w9Uzdjx06ETuyL7v56UH
WWDgg+UouRJvptZ+mej8LB/UXqaiUKJXucgaJhM5Cl37s4TXH0bejzmbY6px8TBy
6okkF7Q87IkdfVI43rb0U1eIB/2RHe/Oj5Tc692KtPNoGZlURODb280t0Q+cu3n+
osoeoPY5t5kieRLwg3VTrzgWoAo4jSLN08UtY/nU4LM8WwpkBs4brv/5BewdMoQR
YwJDY0kHS5w+zyLyntD3UJkqZhbsL3M8Fy4DqUmi6lrwwjoO+vNTVP5dnh5JHO4T
CF0ZQaLD5jrsdlHxoesCp2jSehlicqho+2cbrcwqjRDpQqgstItxZVV2MZSHEiH0
KXeAhGOhoB0EGykJypoVEPinAMKqqsUpiB6pTMBDxT6crFuUs7St2AaXvUQY9IBt
vUHoZy/qEBbabLZVV4ZaEnFyNw5VXKMQLUyjcf6mUwN7s91zjtcxqBdH/N7O2kFI
bINnWXvBzar3DE8FivHM3wGVr62GgqJuejVCRypfOtPqLu6HQmaAArxvJuAp9Sis
z6OloYwSIRAnY6URuEUwYdGGndqL8sbLh9EFe04Qy17xSVwmW2IpJZ6aE5jKkomc
nhgUXkebKobu1ElBjyaV8WH6cj09ogwD16ctEG6mGm3AnMAuS5thKPeDwy8ao7jf
B00zjPMkQUUcR/2eX41Pezut1OVNivwxDts38OEcXXyI13gwnxdkrRAkefq/P+5B
NtiwvO4F+9LyGiUo8ZY9qHoD4TI2OBcoJDf2Br3VSICxNUCKjCqUjAWBmnnbsd2J
maR5jLkYuVLbqhyffwTCZjSQ8QCvCJMg45MetZDiAVNZR/SHpbAqRyhFUdpheWtd
ubs3MCEdT16xwDryPaLgMRVMPt0/W4/6GS/JYMoEw9Hvm9W89xAlCrm0B9m2GzwG
ZdUfgDOiY713GlEWGJxWdAqTXC+vkUTr6afN2n5QGt7JkD4wVg1KmMgW1AWYbBIT
YJ9Vc+Cy2gZKLgqfuyh+BcUsZ33SotT67ttA0k/X+pWdujxYPJrZJvfzyVZK6WI9
8/U/vUSEZwHo8grVkl4jSarYQQj75TF3a/2y4KMz8m0Z1FbfCPZB8OmVAr+V3sOe
+FaFt8rN0bAeceagR27qdoJlr6t5mcLSDfk5bjJtH7dHrdw+ipjhDToMS+ziVmMo
CG7i1LMXY+A62gOkYX2+/MPJrQ+OFAsuqVtPDyFEasqq822vAV7RIA096KO9XEGF
kR4eLY2w9hGywEpxT+78RDsqbJg33tTwmEz8r4YfHzF57evQ/4a2ZOw1DFs9OT1t
NGnQCKN6qfGKBlJEPJFTSjxmsa12LqLpTDx9HkzEDM98s9uN0Mmg6kN1VLIR+qvE
IwavstA4yXlq38ObJkwYyvYpGZsgkXw0udVKiG5DNzOKoxTyznxTTq2l0ZHA8tX4
iYWC3BSaZ/SAZcgZGgVpbEYOJ6jUui+F53yr7ipa+oUHDATgyM9A1HK5yOOexh3c
t3Ko+d6mf5uJh4a2y7/5jeVMbWoHeRmlyiA/CtI9U5LMD2xOzslPfVJpLGU6o8Lj
SqJkViODferGCjtt3beL6PqdLrFhbVtNJA7EYBY/H65gPA50d7q5D9fFqVKmbCY0
IljSVvJuB8YIoLT3Zp8r4hJePbzZ8HcM72k2THU6YGCQ0UtWRdRfjjITbGBGvjBq
lLMFXHUZa6P/tJN0BLus+BT5+0H7bGLtJoUR0/uCjbe5rRu+ePO6cIfSNjgtBUZu
GPnhDbVBe/aOIM/h3mcMK2RGBpgIGZNxLiKRSjUkMVJv0kueMn0R3ZaxQS+igsfA
dH/DWH/H6FCr5QFonS3NGRjGZUnFPajUA2O2TM4/YJwsCVHtACMts3ohwRyikH4u
ztT2sI/biCdAgAwSMJmnO6DCMNNvUHd1HlCA5wwqH9eFOeZ4h3vTS+REv2QaougR
Wtvz2po8grVMXyAd0GbB/GbFKwRi4CP77qBKLoXzv5lx56wJCV55jY/MZcDjU5o/
t+hxpMaxxywJVPvjV8MPdGACDTuCOhQF1q7fI80wnvjo00uDM+bPPU0dF8QcFyOw
OtpHhUb92ZFLgOFdNK14TjLfaN21bcTualV0LPKskvCu+l8CyX96CxfZRl2M7Csl
YPWpA6Brohz4VrnSImx8p6XpdAwn4RUWmp65u5N97YC1SiytUfdD1C9SVEv07TfX
FpDl4RPqEpBL/m0VXL8ETomLQEMetiWRp48G8kn4zxBmryoM8VD3+b1eWGbx6IhM
h1mFggarIjnuXjGLMLZj9Q31GFs0pHziCa0DCZXfrk4c+HMf+wH5AbF7ASI60He5
a9HhbX82jLPkVhIPdnxjc8Z5ZLD9a4PUG2SyE9py0mDKBCvxzM/XOaK7jfrRrsrp
T2qaqUQ8Nth5jMD5StY/RSpNiS1iidQsP/m5xc5xAiKbjgnWKY2SbJQjddYNtk/o
HG2B1+mZo0d6UGvpv9U/Eg7brdPsLg7gftcDDEgT8kNsbs5cYI9BoVmw4kheUs9X
TZ/XKpImdeETZ3jsZFoZ83fgoYzSl8cR5v6SBTTYTXCMFp1ONnLKpNrOrO8z6NTw
6x5KyOjykpavcFvgvdwitAApAn4tl4dOZVJXGwrLZQ7dRCs7g9Nca/7v6m4bx0lI
qscyBizMzPqRErlJUO+bdRUNziTS2xbHWhvzRAAdsDuPBuTAUYqwn0mUOL2M87Cl
oDpcZaoebP/FAA02ygl57sb6F6qDCtokRhvNK7enpU5DBfxl92z4IuNaD24jmdgd
ptl/a/To5TuNFGxeIG78diOEgbNFHY3nPqSI4OKqS6TenhHaoUUttq/99pkgdSnR
mee5fIrmZJO1iVzV1tWahbSXy/3K/sPacxQ5u7oi7Mhk7EIJp2x+tZRlEOvpqnLE
E1kpSDJ6mwdyClB1dNkI5qXodudwM3TnR0nFKUN8jC93NyQgU1Kae93+pTqHY4SA
WK0sRUzPBU/xRHtnDESEtdJMMypEeeva+kgZ7SaidwJnJJyJ7t4Hj309hD3JRGMT
IrsFYYt4O4gJSZTz7Pi9lu8x3pM0dW/tixYYKGuhqlvYTVKjXXhGap/b7OVw+uCg
K/kYbRBkRz8JW5dWpqOIsej0jNHzh+nik+z8jOkNOgq/MpLS+XRkLmF/sGCoNdSZ
mLZERFBV7raqDd+W3FPqoz3yeMw6cS4ep7GesiXa8ccI+fLcUKFiOzpuUwFbRwxj
MEJD1Qf1hR6bxSUMBSF4oGhyxt86CyLgDfELXiSQcz2rrxEdJiat97yRUOS7hBul
3iZGQGW2ikUKoiazxZGx5PYGiXaN7gg3bukDWvr9AnSOH/NkC+BTP935gCK3jfbi
K7MSQksl6NjtNI1TCgu+cq9o4SJA7WYxfCitpO4GXRR5cm+uAjR60++OkfdiRQ7p
XW2P6Q3lY/BSpUq48GAokjmSIv9NxKVOR1TUxcPZB92Ayd3XyIgQ9yQOj0xIrJyT
0eJKQR8D4FF+uUZr+yevybzajKYjhk5My2UT1ET+xmIxyFVLb5rLDiBzBcDqIoKG
dUq7zw67Q0PGp9vqbIfK5Eb9+tdZOSOGtQ9I9me4Tn0TBRNjkAwPyPw0sxLMB2Ps
Gbb6j/87DjluhCsh9rCdgBhepr1ixRfpchRKTnNxXVTZtSi/1wfYvdZAdPt6p1JD
YeYtavQrHYYl8DnojStAdTicWh7i4E8pQgnEiJ97ufxjYdzsMq1JEVcPqxcVAzvF
84LYtKY0jTWytXeDgdTetMHmz9/FLs9rkPY+ja8mZkts8ATdgjhSa7C7M1Wcnte4
k/mtLA6jm3u5nw3ES4GqjmZrD0FRHbDSfQDIo04kZYMrphN/yLlfBhva3vwgCOxD
+9niTGIDCS4S+g195O04xkEkfGEQO3uirLDxx8ljl5iYqzYwQVioTHIwUA3RwxZ2
sn7LP1wKr28L+T1MQw7iUBLmh+FHqgWYsNcWo1niquJcv1Kf8k4bUPj8Dzyt59xr
fF8cBocU1PgtyD351P6CQAq2DyneD5mTnBWUVdlICzp8xm0lftw0SNcO++S0xyA0
CZ+dD2jdgi+R4Txw3JwFXw6NQ6WsPHtsoE+hFnP/U1cRI7dMexSjFVgZNuGhPpS8
K9w5GSHS80qCWqzn6F5xH0neZ3xLtyOU5Z0KXiBEXRTF1+RKq86FPlG9npNK58Wi
6dWgOQ8qyRo9530mjkhKxDXE6W+8trJkHX3ShuEoN+D0tijqHIVJ5Nh1DCwma3gF
rnse5ehPE3oOmlMHPJvkHkWVEMmjx01ZGMD13l/Oq5k68IbZ8paT4s5p8LdC63Ia
D60AUIe6QowwMrbn5/k+bjC4yD/kUtCM8NGxai91haPIhtLzmLcWn6nYsf40+9QN
JG/9z1v8csy0Q7IuUZU0PLrBPEyGV1p34lsBWMOu08FIdhM1q8qrJ2bK6gMwJVNO
6VqOum7v/ACvQ7uO0hZuqO8x1blddddHecgGrGNkJzDa9SfCGyN8Nk9VpSkuOarb
gzPLQzHQP05GYgkzd9LpquGbP9LDTnxoTN6M+OhaNoMfJbIEeN6zsDCgHsQsQW5w
oUI7kSiOBhrDhPlddvK9AJm8NNcvJAS3isYQp0Zg1rqfmnaTmhvNg+sUpWDoKm9W
a+7Be9rxSWn4tzKlIIBwFpSLaHUDtwlr6nYIHKCtDFSPnZ6I8GrWPa+Y0LW2Okqm
8lnNi/I7bdH/1qb+oa7fnOziD4h6OY2j9Fb/BCCfp7TSThhB5lfGE183pIIFeuU4
APQxIlut2LuWR5uEHklHAHJZp1jbQew+Z19N+xTmf2GGmwY4cu94z1EwnsVoSa4G
ayeoZbFa61OH8l0RWs9SoZC9vmCASI/8hgDgtmVF7YEWHOPd0OEVQPgNSfAnPIvd
enFsteqspm6FRzJYs0ZuFgkD1StgagYhvCp+tl2y4xdJXQHxT2wUKRINQbYrqgks
5dsQeeNz9aheWWf179HqM+4iNn+8qwYe5zBsEmWSGFY+5/6K1g7LA7QYvxKJtewn
I93+6/xhxBIb453MlV9q/fiFhj2SRDjfau4dsZ9q+c9prvhOJ+xIQI/JcbICwjYD
iN3OY7L+7J/jr1EKHeFIXW84Z/B+HpnzKjxvx1xvvl6b+m64WXrrWZEp2guTsWnY
N/NjiwezxkUZ0Hrr53ZbpKdru3y9S+gKfto832YAjyMMZ+X2d0HmLsYnJXLiPGGj
l+bUvwkwto3NAPhLIf/G5WWmN9ZOxZNizKA5aICXr/eiI84s9WFDT1+0vPkNYNpO
ncgLezBMw0xyva2FmIG0fkdFTObxBM/DegJVvAndx49B1HKa+26dK+V/jJ6uhcxh
HXtf4BUDGdu02vuOiVnx7yQ7Xyzuxcil47fWUxLEsHr4XD5DMtZYKAfosUJff1Br
s9AC95Ao98ppYOP8pdDGZx0baSWfL/OOlR9yFwCQUO8rJrEzk3MtZ9e/S+oA8hza
BfqmZV3ySReG2iyN4RygIvN+MWOXGF/MRIZ+TwDMN+WOxY4TrIn5sSg3tvc3LorZ
sFytSH9QjjBaDsl+QsIc/kqLWsusI+KjqVLQR2mIp4JFrjYXwFO3wCx0FHBL8W5T
OZtA/HdQpizSz4osBvoYiM0u4EpL+zwKSQTsW35adAy1FSf/asspgZPIbb4czR7N
7M+piuX5CA8g0lrIxvffcNnnX5XrjmC1yiLMfE5hGGmMwLjibD5QhVU0wiA3o/nh
vrdNSbfvaMm3kETvoyx7xQNzUmrAks0dWCslhrw6nN46LE1Mrw+JJ5sWUtc3s/94
voYQQl9cMlSf7YifZ0pgbFxLuUMriBPawglUZa6hU1mXU/+gev/DGe83dk3iMTiJ
A08Zcbc6W9k+NdrlUFSM9ULX1ND1NlmUtDXRXqH8DW2PaK3HQflngYiV65acqgYX
OGKMnrDufFNDXo/Q6OOiJq4Me9PexcDYHc2dab5iKpU95+gu5O6mN7TsuTYpxytW
5kqYz3UpUTLL0+m6/iyUz1MDwh75CwutYbreOQ+vdm4tizQELcoJa8YsymtYZ2pu
U4rB+d4e9Pom7mAQytovLLLKW8IFEM742QiogB4wZzTXbN4vmHVeZLDBysD5drXo
VACnfCEyZL2czMyC5OLLDQVWjXGFAYfqodZG9mVqPq/zw29CBfIGN4XDRz1a5JCU
KwvroIt2YcL+XoFb25plJCVSK/dqBdODR5vFNVjzpB2ZBUa8uS65E3QgES0ZoTc8
9rE2deBBckpDaRKpcRNElsNYpaGysjaGaqvnWXcEdrCVwvHAoZoqeoSu1CYemoe+
xfI87Hx7JVd460reN8VFxWBtCUjWOZUogqD8h1H225XRGsYT5wypl2lvkSb/I5Hf
RUD9hAmLOLb7WpkYHB7px/8i6PnUbXR8vA1jXZasXLzZC7mG3Y1KPEV+mB3PPm+k
N/SRW9JPWZGJG87b7Oh1knerfZrc7bZvWmuDh/nuIpi/HTeBCZZUVrB5UMChfSKO
jYUyRvSUIFt0N9sWdYWt7Uztt6va3YqSFgMFSTF5a1wctjQwhn9uQVecVfqJ8bvf
CVaoQ8JsTp6qnvrgDRqejxFZ7DJIy+9HqaX8mhJsVGUejjB4dMCQZKrsCHLa/u7q
an1b4i9OK7i57Lpsnm46vfYPuw0ojpy+/a1LEG1wBdThKumZiQMDMAwhcheQxiMf
8Z+68bA94pKbYLb/4epVRiMCVvszxaDv1GWrLhTHPmb6DwThSMnVzX9AGVezch0k
9r7nO456F34H1JNQqVA5F74N8nXrkVYXvTf/oalj/hA67LvqBjkhzkMxNLKppHTK
jIiGHKUIuwsh+Keltdhzp6l4QqaIlp45GUVqH4fJ3KUCNZvWcmJHC5X34PcaO8QF
270wgOgVxEyXm3ZBw8uQVXABVBEsu3VSKoDk0Szud5HALY9r5fNnbEjaGS6cyK4P
HIo/RBTJwmUN88984fTCSuSqVGlaji7NZgUb9RxJ176CL5S67/otus2ETOhWbw79
r6ir22ne/KYtClvcQ8DPQnxVpCHo09QOVBqAuZerhKH1A0/GRlfcDl6nez5ZJG0y
V70zjnYvXhC7TKuYn/IPLSxkqJK4IUsEwMFkznA/bTTBzHk28cO9nV3YaENW4SFV
zj/0DUMIRsaytqsfmZiFSc0GGVqnDIwQS6vYybabT2Mjr9NTPldoz8YDpRYOhkBh
uDh/NWs3V2c2y5nsuO7uteuI1GplxqUw3Y7qyHAi7pnKv6qgwl+Fa+jinW8PXjkc
gUbEJxWgRy0pO4SRBidAkUW2sBQw+R23A5IJ1gjfVIzPLNqMsoQHar63GarR4BDv
wJEle8prtfkcbyAnwo8j5vtzd3ZB1bktem/F/H09fNCexTkJXORVlV+1zK4cc+dl
VK5K7+MfhgmDy3dFCPR+Etu+U0FJDcdT9C1j+OnYepCX68LKra6DVU4/qv0LkZd7
i2Hu2nsypOdt4hbTciibNNgayNQGGrPnl4/uqd2EteSezcTh8OZXlAb3/ffQ2YRi
cj3A83NBJIrcvqCI5hiFKdn0yeyORFRbl7v7VZ/xmPrntjIDbXMbzPJaeMSSwrR0
/r9HHWPfnJOTVJSGJz21umxxo6wpGgr4adbD1h+OyVRoZXWzO0RL/h8igX7q8Cmu
zYqzM0uW10UtAPm8mnWRkowtlye0GI7X6iARHcH0d/R3qqGZKjM4aVF15S2pEe8+
VKBOUXS3Y+sQHY4nPadSgZZxr8ZZaRCvgEKm803fkwv2eUxynB1h1a1whBYu89zk
9TCjRBP9rDZyLfq1X0VqJaPHi3fYGLDRmNdMaHc5Zd/5uzDZjQpe3QjCvxbHGcIU
QoK3jNImorbHdruI2LlNZVS8gkv/ZtATSYWFokXjPYvIfG0LqFAC0SUBRBkJsa4+
LJH2pqH95DbYgVQzH5CzD03vOJe+OGNz4PotY/kSzmIcqJznBBv4MY5yOvPpOy2n
FiNKwEsh6FvqhDEOe3I70SOrBhaNdzFKfAcPY85Xez4y2n6rTH24V2wEhQzm/+RR
hDyc5Ip9crGb90i0TeoYjmHwh5d42uSQocydoQRNmin1+bbRkAaDeEq/ArUqRBmb
Oo433oG55jjiPbqlbVEe7CgHhLKABPtceKBwGZvmFrby5eVwNpeGb8Jul4B17jDm
xcn3UfM5kMxUVKzB6t5WcrseSbBKRNuOFi6I3Qs1HhRm1leskCUVBZno6gn+Ywry
ki/650SpgVJRzy9IQmhuj39UqonbKJeXYi5A/3vpOhcbIXQy/u89r1UwAlj7v9c/
p0vso4dY5kq2Gj2Pm0mkcTWlB6uh+z5mM7SZiX7Al6CvG4PiZ7RzmZYNB5ppBoD6
6ztE5Jr0+NtN4RWeL07vABSJCJ1vf1Kx3mCcEZ/L2QrqtoMoDz2eJXSnvHvoiT0e
48YcvtJY+etiosfmm/zjI5//6Vfa64jbDRWKHiO0y61IyfueX7VeKywfPcG3qShL
HueTQSlKeYNxd4cjqueFkzhTOXdlYTYeTyNON+qofS6WFw+sbhuSLwDGMYklT47H
M8OY+e3CJPO2Xo/c/TbMECfeLjM4vvhxHpla436Jjxzqt/tjenO46O+RsZHoxPB1
a/TofJDRKaNHxJE4A7FV3gaEFEpm7OjSz7iUDdkFtn93O2BK5VDGDmqw277rwIMD
NlYyqFJKs47mtPsl4HSKlqxvZjiuIE/LQOI4NTq9n2zxnUd5NhCNbNzzG/WfVIeq
dDGqcU22y8RP4tDHBHkEZ7X7bpKpt+DCbutTCgDcTB+iecj1AUqmdskyaDJoRpOD
Irn6NMYrogpCbYvTcqiR9rEBUOE5WhAAOsw8IPymEsI4GL2uI0UQg0brsnsjezNZ
ovCnccyfjG0n/BcY3tRO8j/9cstLoYLSiN5OVZtnPlDnt3c2UR59OS1touU3akBF
zBsUw59vgHlZgq72ke2BAMVMd8OHc4WdxAj+R6njrFMNDhTNZiT06Fk+V9NBEtWE
rQBxQVbiXqAv4KMJeh7LNqWLiIp//fl347jbEf3UheLYYyiu4QuVPhz00SV+XEzu
VtlHVlZlzbGsqvHMCSu1RdoTGTHq+eBspfxW16NJNrlBSVG1d5JnPQ9PEJMlq91D
KiqWDXvmOQ0QhEUeO0Y8GazrqkGNZcLegyo1N/xJZxl0I8nUhRvpFdh3dNIK8HNm
f/BzviY4b1nU8KngqDG7sGDuNYppFiTen/elAI3EhqEnCZuidkCQmXy4g2ylHJPM
KDXfmwwI73Dda6aUdyESGFAm1u1sJHfOMlh6Mzje9slZ8UvbYwlCcmKe/MsFE1A/
Q1Gvn2WwZhZWh4DN1Z+cM+4/ZjXHEy8X9s7sheMOua8tI1A6J5eOm5uAevs5Oy6t
RMbd0OpscKkyY7H00ID8rSDpCg1hLhl0qqS3m4z7qdaKvv71mexskefs/Buit70r
lZa7t8hyTWL6vKRK1wSH1BToeg2uz3Y0n/oEJvI5doZrhuK/UGAz29+6m8TET46U
8E7z7RvBbbDKWylqMp8zlVADM7ZzXBKdziiMYpWsdCOV2SDO2Yic35imzR7KeWvN
oREH1Q0M92WiPjlh5lNZzcOXQ1VjElwDomjtXE3q2PD2HPMBevzfGMInHb6/q0Gc
Xmk0s850nj6I/7fy0nFKywAJ9oRnfqODtByEH3ylHv5vTQH6jbh2R/XbXgT1Ykiw
kj6dwdbd6M6kkLmTnnSUqIB7T48dlCnZ0PGOYCMBL1ilI0Q/Ndl0tzSKjgSNi7CW
fHhTcsdfq3JYwywNeJTutjF2Y6ysHG1EzSnuk10uTkeP0I0bVEyTNUfvMNGuUqoF
zPi56F6Tkqw/ZB8AcX0og4vU8ROURK0J/mYmWEDrx+ZzqVmCbfjqL2uN44R29nMN
va6TkhBS8E1ZC3u14x52mVXGoeYv2cuL1GGh5lDbU1CjhOnnN16ypowcUpLWSCAk
rA1qhR144msoIy4kdFqW1rNOAmlnUoVVsESBoIjj76pwOfmkVENrr8LY+meXmDAn
tOzhOQOUieMsBESCHvDDjSbo40w4gsNF0IhHiRwzSRrMdkawXHZiSlRYgR+SABjx
sZw1hw2/2x+L4tojKYsAhap2Fx/HNSaSY3gOfGvO+010JK3ldWMXs7t21yUGGGeJ
cw8imzeV+DXzF8vweeAVOpg6TgxfE7GLd0hdTX9dsRWuM1Vmm09PC3ekybK4MO1V
v7m98Rp7VQEX9I2uR4VBiIyQVkqv/NRwITE3HenyRzP7HRfXp8k0eMvBg48e6kGi
wxmTmacSO/iiVG7yIRBRnUdle4+7rdXFELWakwRC8/ykGDaiifqUOgHISwyM/Fzn
r6X1sKnnifrh6IpLOVWjgi/c9HD6RvcmvpyUjRF7VAlc85r2XRL2TAqJ768USONa
71eXh6Svgxh6rk3meX3FhhMeFcNqwIxvVN+x19rzwLu/yi2DsXEr7sPpjWLaylZf
N/OXksojc7ejucOruEMhva3NIpgyyB1bNdTFmBFRSHrC1qiUrzGg22N/c0kHnS4p
L81a0NANNQ3gYIB3R3zu2Z7mDf1k1CscA6vp//B3t57KQPAQZ2+irE5AbWnvhIf9
BcoFvoIJbBHURFqwGolnhU/lIOzChQuJoIAQtAwTaz5aMNjQjAUtV1DtCaFs9i6E
mlwyzzXzDQKsz2MrkE5g9KkbBHM3RRtDyCIMC5GUfAdK1BE2ivFYBzuDGS8tVLZX
OOg6v693A98MlkVFBVmh/ufWaFU9nWAcGACXAyLvq9fyScCGRHI+IlmwbqwNfbBN
VqcnI+9Q67mUEZvOm7AjDKfoJZs4JuwXZNWsSO2ZSrlDR/IW+OfNsPdNLGsTQmG2
Qpukd087drFUYERKbjmFYJtavJpZiQQ5p1VQu2efht/HeALXXYW6twzNgbGV/VMT
ySrYFJR/uH79wFkOgQDtqaavvOOb5PNaGdNaslquC0SBeX+njtOVWh625gGf+ywW
jnctKiwgkvKGS7xWVeULAbeRHqr/5thsjpe948kdO9Os9QHQhtofx2XJxG/ywE35
zqHq1Sa+jMELTYqX5CHqnqruJAUxWqNkLii/lTV7pGfebtlsKuu7/yWtk3h/XmZ1
U5R4Y9SIZci61fuQ4jq22t/Q9OSEJlUR37EUHwHJy6lWUSBccIaghbUEKPYoPyRT
6dPkSHzkQv9gnq4/z24W9+ebHeNUjTDkwT/rn7l+2Gg/5hr8ytHG+xKiGyfcVFx9
yvd6ythn8AgbyY5AH1GgZwrqzFaIbyuY9wckgIU05LNIO/TMMM2LQHkpISIrk2Bn
kZZs2hfom+n4xxeHpm99ogrcpH0sTc11R2NPg52b5+t7j6GUtIxEojuwI9KIw7uB
WTEfs9LpG85nw652ZtAyexDuNdul0NB2IwEj0Zir/G9OLV9MR19LN78BB/ydL6tE
aFcxTJi/H+3VVfC7ghe7Ijc1IyeGtz8AWV7cFPndqGhoDAodfN4bg++/01IoPExJ
p84DX63bohdBWZvMWICt+yStrSV6HPf3gnHR2+P5wrV2kkvddylf1PLk9vVjLGvY
jdR5ln79Lfmj2sg0ptBGqRaKjGg+6BtTF3gPmZYSIDxj0Y9zW5ROvcZs/SKw7tqM
yu60YAqoHP9S3e0sMq37279mQcKrCv+nVPACg/1FRcVrTOxVwwu9jNedwYOFKuWw
ehPxduasy5QzokvZxjgKd0H2zBQQwWdDubYL7QLAtvWs9XAyRWqm9LcQ14KxLMTB
7Mj54qXKlsqFB0/K/1OpfCyNREsTn5DAprKqP9gS1fMw4ix/WaA2Jtn8WpoD0F3Q
LWU7I94uCWGUMDw8GnC8ZyKvk2XOLNLMoOJCsTUoWBWXL0D+upBQci3Z1Ljy2zzA
8JgsSpncy5GbYgbmJuuKapkPFi/xlyQi4Esvc1D61DXSPXJ6kgqn1WL+grS7jIAR
mb6zN94Yn/8Y8H45RHC2K8793RToUZ1JW+PTBp6Vkz80X/2NmH+X/+wofHH3D9gO
ZFQPtF4Vm7Cbp7XS+HqZJe3XsbakcmJWnYa1Gks964VX2qpZxxrZiqOQhsZcGebV
M696zYaYw2mxhEE7p9AdW8f7dhiCjy+rNDTpULHKwWhzmVoC5PZ8YE77fWVby2Oa
s+x0bh2vtz4XA0Ih45HP+8WEMWENT/7z5WaCDXTo6wMXlghyeNcqlCA5JfJfhOXE
MjNcdXpXuJGdgQhBXROV+oSAhJE+mcg9JMyBlpaObJToJ03HttJIor3TWF7aZM/v
wcBmE+2mOYMk/jxaorDftj9wFFgX+6r/yNSnzuif70/wzUb1XyxccQSAeyVLmAui
f0UpeVDdVbAM0VZMcYOtcDGk9kJRBELT3uwL1DEx5vD6bdbhiVGnP33kC8/CLzr9
VVwzJA/HAJMpMPvLoAPNOxw/mMNYhdm9pmCmfH9q+vAw3KFJuCa9jFDba9rIz76j
Mk0qRpH1rXPY60HhG+sAbiW46GYDVJ5jIEEC8kgrhQW6B18pa+v+F5q0ybNPwUE5
BPILp8tuaXrECRvKv80ooI2e3jReMTwH2xwhC3UcuAd1M1Wgcbbr8e6g2Nry98Yy
+FTFHdFe/pl2DQtSSJ5ZOGv5eV6bNQrdQn7mClj/ULzGPwrR/o1/ULmDDcBO3mCx
X408CNLWp6Mvk2wsehd7HRKT96wtipzV/vOCC7Fl8K7UWtCfOKBsthzYWjO0o/Ie
Pm5khztLtON3etT7vPgza75Wjeh/xBaKXLK6RNmJjnDgvN1q39sW7BaD8pdppFie
LeK9zTxRp90Eo8y/Imk9DDrJGtwq4Hs+vH+999caro9DhRj63sto+NfeSAIC/shC
1WCmo+diB5VjJxK86lvIS6gKGBpICrvur+RqiBQsKuA0IY9sk+hRWrFx8MmOU4VI
hs5rTyQaC5gTbMyGmrqp0KTEu0NSUX1NLDEFMhVUT15h1fPcuIve/nPqcZCB+thb
y7ea5I5yBNUTpJQtsyqfr6DFUBnyiNKuT2OwIGMAAhKSli/5pgV182BoKPW/+sjH
v+K14tie4AHp67lYTato0U/lTJUKzPD2sT+UE/7nC232xS/KWSyFDa223JLocUwI
9iZ4PQn2talxzFqYgw2Z6VUsEIuraeJy7W3fL8YU+Rk84wSG6gZkc2DLDtj6w3eo
StWsRupareFUsPjfcMKpFRmyVxSCjKS8qIO1g202jCmEyYR2AdmAhEI5JJmc1VGe
NRtbFCUuzW93cug4T3uA8ocVYRcA23WILdJnvDFFTCmzF40vHHoz5EuZWVChdcWZ
fYzd9P4cr7JJlUQ2FEvHefb5yaugPxhgs44MrO1pJAI2GH+JcTBXd1+Prtstr0Dr
kEn92YLFwJUHZTIYWnkjELkCFGHcUoLPdZc7ID6RerNDJYyuJoxVM+k/nrl0DAJZ
huVjwS2hjODJdvyh3r2BATyX6vS4ExBimPsFd6oH4Gwk2bAkyhZmvX/qqY5Ayoo8
BwFeF/zS/zBbT+kTybW6XPtQNQG4l7ptW4TL9sC9inltSYJ2qFIbJkd0iCfgg9eB
CXna9dNZ+OtHsYnRXVldMagaglY6TTNkafGd0Ihun4e5LNBOmCBvTOUgEnf7AaA0
gVFeov/m+rNva08E5FoOWx2TeuaM+yh5MltXTnpZS+zkTcPXk1vU5u7HhPykp39K
iCUDaJFgx4vSEqn4aed+0IWNXT+GPgOpAu0Vk/zSYzBUAMrvDWrTl+rINnnjHGzN
omYUWrtuWwjowgdZqMsi7QC99fwkN4ngWHXMbrAKKH44shq3soa6CJPDr24dnEME
NaUBbZHV9gN57Y0rOeUDjui6fT952wJG+zoBDpwGhFdvTxPQh8u8jb8OWz38pUeI
muZnxpl6tpzu4Qg8Cwc6ds+j9Yp+8Y1fiCSVqdlgSxI415sXDbrw9Tcdrub+FC4z
aL4nC2j51kfNPKQUDZxEgHjLjWgUVhwMtQH7bVOwQbHTqOB+bST2+Ga3/3NHaqsq
MoRaAQiCQVRjP++BwbBhEOq0mGzdHBzUbQlSmbE1ohLIzu2Jws4Y5OWsvmu6Zkws
tncdzUAP1392/QSl+fSXoJ+PttTQ76K75g1iFot0JhQf55D3pffoV3R6vovtT+JP
hRNbp+tCZxlZIPYKyG44T3sf0sF8faX128voQKOU8h0p5zZbgx5rEt4oazXpuIFm
UbqLueUIGObfj6qBvNXeABDApvDqih5ubS85pHDHu4F5SWDpuMQ0wxF9G1TPeCb1
rv/BI3vLbFlZO5gVuRtvAyoKxHpr52OqSmuaxdWbIOOtjaTO2A2/vgxIgY5SIokf
Wb1i+yGwLSmLT9g+ZPz+ntEUFR69M54IuiKNjXlYhdZT5UUpVXSQWjdUJ3NFZfip
VoEs1x3jaH8xfcigrAbau/6PN3MJsfCavUITxa1QGVEXApuApNzqoumKnatL2S6d
1/vVLTmokzC/VDto+75kW2djohUbCZfAOfqQR92Kw4yN8VeR4Cm6zzMk361QUMLS
Zfa0kj4fUCEe1eaPoLSAjfRwQzAxKBdWTM+6+dEgiNGzAfnByh92nTSa3cv+4BxG
xair0wlxSJqRBPFawrTWI87GQUm6MM9h87gCsG3fZCAAK22iVs1m+EkG8HGAOV2V
4k3QW6gFRQmSVGYVZItpuNwCh/qxxO6mqcfkH//FrLaB/jtxDn0Y0IBY5k4qg96n
31/ViGv+SBTTrcMDHrMIMaC7vIjq/okwVj39dBioWbI0AwT/jzlpmljbpGA1Jsu+
C3LwC5ouvHGXpr1L4OspVLb7yQrJ0xGNjyaaIIx/1DVy7uJdWcuf3/YFnHgzEYcS
udBm3ECG6ga6TyRE6TZswl62es+P30LfIKa8l3L2prXp2k4K5WtK2itsW5k+A+dF
AQpS+NM/aj9cC6Zb3dHVuPGywhUEbQyK6ex5CzwLieBWiQJDU9SxldEcMv2R+yhx
2qYiI9Nton++I+8CaungLfliHUIlUok0D02uUZPJsCt4ytBGT3vLjSBrPyaL3jVF
Zb80EG7unqWoquUKWc1+9rkaNaPPx0meOoFGeykQjfqqjV/5YD9aeWTduYUlZTQa
SeJzNU1fmBd4b2qZxOtZggKZcvhOZLBYuxDQ86QP+b53Ma44fJWedk6T0c4PdKtL
Y7KlY4E5cKyFxs/HZYS2F6n0zgquFNw4yRl0FzJCuOBwunYOZ9ohDbTGnfbEGGpm
lUq2zkb7ntPpHHpNGIoipXTv1AomvPwAx+bl9i56CH43JigMrbQtwnqbYaOIMVYZ
Sgg9Uk0KXvWObqBiBPf+MKiXD3PIDpLCh/Dfktc6gO62ANh1Tbw26B0B+boQlmIX
6EXoIvQLsi5cexoLqgPoSOGBD7wG8gwxlUfLuhci50n3IQ2nYZfhWFLRfuZSMJwi
o0dXx9morxl5+vB5YV7d+r+WsJoSBEWDmtX91/LtgBGpgNn3kZGsuDpH8IZdBRfv
Gmj61YnXd49pFd4z9jvU8klmF2V+ketqB2J/3KyzjLkKHKNYBO9uin2gZ+GMULn+
MqvJ7IgfqOM3arh96gGxfFgdVRl7ci7t+WdBYsOwXoE8dUqGRNFfTigY3wq2wmFW
roRHToJsQNPxHov6SF9mvhP1HHaDp37SyTSMgdcKv7rwNZJaIAVB1x3tVLy3F4R4
xr2i8pF4rem9TxKj5FY+IvTvZHjN+oJ8v6doYFGyiHIOShx1SYBAXisEaCPCOSiH
yyHTjU/VBurmw58HXbYk2PlzTMWMO/GbWMArJk6slq6F1USyLIyLqyQGErirA0pT
aF86S8T85CD09PP/mc+HItvPODUrekjZyV3ILoUrBMniOYeveGkIRVwM0uP4PuPG
unl4KMaGSIzELVEAfF0XcvCE/wEO4qpJNZ0nx0ebkeQCqTTanUr42fX4AErvbQTf
Ce2dkDjDk9xD/9GuqwJbMO8rIZoyRFPGGhpwo0u626zFcUTwFogoR123R73Z1ZQA
uqN3LS9RmJplvPBliIWCRytP3SnP31g9isu806MeUfRv6G8KsF1qEps9aiAyoTou
VpgHOPQAtNbFigPAbvY64N/kM0E015hEekB5qlitGjIfuA3JP4RAFOdaGH5l1ugR
ya3anaPcOdxjNhwAkBD4DPSafzz2oTlmV78Y1fDBSwN+JQdhc0nCrvk11ak1CQ+G
qHdGQxFinOXOQfWKDDHgK48vKMYmtU6Xlue4x5Tu+Hq1U7VdM40YDrS5hxplp9An
vVSheGzgC1Z60wulGC8JHL8ITw4N2yDwKb77sZx5Fm22D19evJN6hVwVbg/t+kM8
Mx9sdVXwA78X8aLKa4T9CFG2DgFJ9qh0l2NweAI/Tv6nBse7Mnntaf8JPtGNPaWe
ThVLtQC7at8BdnMpeD8appD/5eZVjgeXoa5IZ1jh8R1rV8YoZ5LZ6pBG7m4Qrpfd
KyLp9mxOcaTMLvi4RWH66cPuBCaaia+R/brmqaFdqAa+pi6MWU7Wx444THjL2XlB
/A2GKWbHyTLY3WN3xixbGHPCFFyFai6u1q0Xd5eckMdgCNQH8jOTe1XTb5rGWS7E
XclZsTbDhRdAjEulxBUxGn3bJH9OlmXY/pUgbth+tVurMGmqX2WpggmPwX3yfSNu
yxHeCxP/vlDlYdtbZGB5Pt/YVo59FgKp8jmFSJb+ADGEE6UFySg7JDPfcYjrIgKi
9N8F+6nkPU+2QlwGWXL+V2jLKutBjx1uthf81t8v61SoGc3MnkMblc8V+FzMGMID
2B64E1e1zJ3AvwWQPairlJx7OeAoDRX5fojGMTkE/BcUcrhixoDcfJ6rYUPD2iOr
sPjWJSVDcetbKgqF4huNyNGo04vNRBK34xlsVPs+RRON9iFBExTUrlvcFh4jk9x4
8PfQCHg/JgUhPb8nc8ComlM88ZVKSvB0vn2vBXgVFweCDZ6tK+7Ot5QnDuH2v7vh
wAHT9SqSIutjo6zbumBW7y18G7atq92xO88uouOf7Zvpwt0ibe3Uh/CtbOJBuqvC
66/ap4bKhDl/66p4RAf4Ty+OU7EHWcrKrQdYewbWnK6eyZmPdXlld86RxMuqzUn2
nsYzjiZjBXX0QRnlmPbUbQTrHk+YNOKzV3+KSUqG2BnzSxAX5YARUOqDHrtCukkv
gkFu3OWyKFTVvSKW5JLLKqt/M9S93FrgKwOEqipcIlLjdKgbHnfq5fZODN1l6LZ6
IiVmmKT1OH+HXUQebIov6YUevYjuKDpo6QFWlUp93CWxTG7WiJx2XeUudxUzsjCa
oP2TMPmTOt6wz6w6MGs0acs3oMfgk8BIm4mIPDVBCzMMmVQ9TD7XjwCNPmZ5U1++
ttlHslY6YoEn2lzON3CT4mNMPFsUyOAqRz7/p9PD2btckqi9kF4K9XN9YfY3AJFN
YCgYrh4dOrS4h4v/hZk1nhx+HeZatAzDYOYHNdnPVKN+GIWG14hZEKRLJTKPdsqo
m0X8ld6GqHKqiwJkNQXCoO+MfgZPVg6CfLhJuwWbhInrdGWmllnlDnU8n3oY6b67
jf6cJevJ4MpPkaZGuECkKDIzkTjeBiE6iMR7th3BZ7xGXrccXuWYL4mWzsFdBZbL
z10yC/HXOtPGMRn0P+4AWlu8j0OKgjSNbfh11JccftxKnkGE++710jLm1MXEBZlf
UWEd4rY9jVWHhHuNITwbeWOUsXPzM9RHM4dQe5YvyfnY8dNZRQifOAcHyzEflynZ
K1XrcCPQjZUm3o8PdchTmkiMExlkd/Nu3ke0Dt/8PtxyQf3GtmrREWilimdyQei3
BFUyYy10YafectB8rYrrsrHSCNKs5caXeXYNfD+f2ZYiIm0LfYCzX6WtVTM/fQUL
hrn8t0m5zOW+iICB4Tmm37PLeFEjizCN9FioB2zq0BStVLBnZFx0DS71IGnI0XcU
vir1Ir2WuiF10eLFeXGj4yvHFcipMYlHerOTG5jhYQrCFUHDVK/R5JejVI8XZGha
BLo3wYuq3us15Gw1ZMFSElv47KRs02sdlEN7+ynKdChZjl2ei96KWlwMu8BHaR3q
qtpFh9GJqBunfro3l4Hju2vQOp8mWcapbTLBzMzDwMAo+dbUj8oODZztFOSKljEF
8c/O6ehKfMBV5NuIYovwuVRHVI23S0PihwIVKZm37uH85KG3e9mB6OmLKbdzUZy4
N8ZFy76/8G4UBDy7Nn2jAAm1x1uqPGapOaicvjxnOEa5YMVXbsyGLRPJ2hEo05Gw
6WSKisjbC9mt1qSMe9lnM12ZD4ePp2HtfDQ/xP8pqHzZ2nhoJfcDReFACwYmBTZo
8+LfO/v+gp2cAZgZMC95rly9Rlgf9WHXl2h1ntapYnWrnCQkqh/4tgmTla/EJ+nn
3zCspEmhI6hCAnxngBs4fmGP/ZlVGxKsEXL5aYSfZP1aIawt+cgqvpFsKk8JnW1V
fs2cJHm2DkDB2C7/sZHuiqlhfnP5MFwtTY6vQEIyfhVxd4LqOduR3QD+kPIph3qC
qHGk+2yS9khqLwh8CXSPNIBObzcx/NkoZeKVUaU2DQ9fhES/Z/aPpnvwOXz7FcAk
xPpaxcpIFYkr4ZUGtYutqc1aM6TzDwyxu6PGAWa/CpL4HZSYBTPtBSBt9zwCIwMy
M/tzSa4U/a7aecBO83vc55FwSItdrPrsaCWFkc9kJ6CXqTyGswi2/H030SZ4Gloj
cgZBcmedz7W+p9TM/VV6QufaYduv1FcssG2HUurcWXd4ZUgJpSaHmTJEcBDXVFA/
N4WtB938neq5k5felit4GSeB0kjgYHdoCqfapK05L0GuznbOru2H/ENWWAxY1lkQ
DjjJDU3FMh26bU3EutTkHP2O8a2i9epzyzEvfxYMZ/1e4//q72sTr9C/+7XnVonN
bIca9S82sqNs3sQY+uASM1Udk8dBIJYQbqmbyda1z1+sqIxbiocENflGsBk7vMIV
ADkQIdnZs4udOhRlWbMoKOR9aGAwL1KbloABef4TTXp7A7b5VuMJyMzTsxiAiNOn
1tDG7DROPkcybs8ckVv0UU3Wjh+CGoQQegScmImzMGxZAYsZhmSz8ECZnigFWprP
GZpd00rGKArarn+To9u0xqEqPYbU4NfpFA+2yIXpJ+DW+AbeRsh9Mdx1bZ6CuQ3v
pu9VCNt5WFTwnycZwe6/yW93mKdNpzadrZtc+OPWYE+/Wwsv64xoJ8PJUjrOEpn7
SJ29n/d7FaEcwhXcNkSJlUR44E11Af4CEG7HDUhMF2mvelxoBGWSiKt9S0kHGXHF
Jp8NRItlzMVfOzYmksG4FbHH56N150eXuaTvZDPNGIYdeXnYKxFPMFnACkniCcsK
4iktLYREtKwXsp+FSAzuD781hjbVMq7OofYjn8zf43wBnA0MVvGMvtfijCBan572
705w92G+919TgxmUWtBpKnMs/WSRwSSS1Wa/7DhIlNyWxvKpLFT3rUDi+GqTOLFi
WKSqEPF0Fv2Zux/bfU9wOek+VZg+TEm538PwYsd86tG2D+vBSwLFksb3R3aD7B6f
piOBkFy9iqv1fcxRFNAIVWgNPmrBm1VRfWkdpZu95UqrXxZoJfh2atncX7F1A+sy
FDdIK48nyQGMXLvXtUfGAvKnLlZJHxZyVNDq5o6t8JsDuPGL0bqYQFAm31248BmB
tLgTpCx7LFIcvnjEOdAmh1jf3is8g9CBVB9YD3IPau1G++rmyEMHjSwrrEzZlexd
MZ7XYsi4SjG9V2S0xdSUvHBcK5Tv2MzeSDI9cDa01WkNu27NPh7GaWDwrM0Vxfr7
POapFHDDlyWt7OhamxU6EvLBn377y54Vp4DagfaARNIi4AChp3nUDovwXByYmISp
NMdu/eGJBIHJHVjCJCzcNWrpLnkGWTdl1eyDYmvYs8Rf4Mn0Uo9mPlQ/b73Trzwe
77LnqZeCib3aJ/eGzH/S2HvtBz0M3LCF9IcwbeO1JyD6YHoVMRLm3PquBK1er7ah
JDcD5XqvKOfNBw4qoLjEWlG1c5wtzNFnmSVD6QHMDQjZ1kVHT++IZHWSfOLpHtms
3RB++ozFpAqIhrwLMdA/4nm5Ktym6KogQBLFDOM8Wsf33/iVNLOL1Vz0QTSZOWCB
KTX7eVdm8iVVFe0TinywHpWYaWdzt6u4CtosUx1VFIy3Xvt8TIHjQ5yXqCxmIGVD
wdysMYYvNMFXBGZPq9PUL1Dpj0PXy47QoNZEZatnRNPkoiNrDiLr1w2SbXNxxrWP
Zdddpw9j+x/0SsAN3/yxifbPjhdS4F+WCN5widERkR73eE4EDs/MpKljFRdAirW3
O9GZuEvXB7eoTRjTH4e4eUHm6Xy/YYl2DbqkBJn3hld45eF2jffWMP/ygjiPPYkF
4CIi6IkhkHabtxoDOUKpFX0grFYVAo6/riZfSooXLNqczAA5eNWoH1Y22c8LzNRR
M8Fjzu1F1n5ACFLQfcdrzO5Pi/ueeDEjBZpdezESb9ZQIFFsOHf569FyOuWHPn2H
fvsmKY0Htl4gqJYOzhNY+NBzr56v6M/VBV1MBeJj+M5GFt9UWOYShHLql7Qh+cAV
eknsRYCt8kYNTNMN+PiKnazb+sGFJkIbgT0bz72szEwB+6B4Jh+EayT8BZYMAGbY
4PlmGL+HzcJxmKT6nMNj5P1hiBwIcVHVk2DrlopApDQsuHJEuRlR8jPXzwpCZdbx
XpcJm33oLkx+68BulTCF94ur7/0UM9Rh5nILk7wVNBn4SnDK0IQnSe5VAhFOiYxg
A+RYMdsiZLDZZ/zlcHaP23K3tORFmefVxXpBtMVe/eue9eOM1mFmd2bRL6qL367E
gYSo1kDsJ80zaFgjN1LxJ+Wu1Z79MuHu09zdcAmgzhYStOZ4Gk6zBQcaplBFJim+
cjwc0nPF7crr+qQNJ/W/iazaBXrl4DF2XHA4YsWeAdCnEWqbHbPeEnn7mMydX1u/
1bHAQPmo/4uv2KfjPhRNsff1/1mnkdXJyUzVxHxou3Ua5eP41hxxFUDpD2a8WZmM
kKskTD6SHslD0Qo2SA0dzS7V1msIU/uDsfFRWc054qsD+iABQFvOF8k1tEi5Oxj2
cBTql8tCqVCvseA3CA9vOGdvNwjpxdmjnXUT85bBXyfumxRRg7ADVFrmr+rDPsdQ
+5TKF9YsF3aOCxQrLFd4iUfzbwzudy3kUcXh++bGNuUiKXoGyiP8LiAM1tvVu7W3
9ByRoXLVKyvd0fEda0SmP61+fuBu+ojWGQlxb0Zj1Xj/6KC0xI3943XkzQtf0SeH
cY2J/nHPodNZ1+XQUj4sG4d9Zis0vCN3QFgDJsFU/n/q6OC3DDi26LxWfC5ygEZ6
ruoQJ7USvW/UgoL/okkfX1K9TGskww/dSX1ML8hk40S+dHHkeqAWwiQb3g6HdnGx
zlwvOKPhUq8ECtSmUCP2jgAip5loq2HrrtwkZQKHYRFihX2ggOKcr+HN4rkfVHIF
UN3vHSYQP7lvzeaKMeeNKAVdCCOEDcFZAneM1NuxqdyoYEH2J+VmB6Ac+G6vDYYQ
IrOP84dWOUIjRI1R6sNzBDgRoqMiW+6CdO3J5mg5GxIZWdtCatT77NQsVjUmIhPb
2mBHxFTDHUKO7obAOmv/1WkEpK/lslKaXah9dh7BLY4nHbZEJ5PxUdMgC+lj25UY
YHUGj8mS5yv6hggf1ZYvi13bPH9IlOesvLzOepcSVzYvhxjoD9rnI72t8KLEjTUZ
G5xMMKIqqG4UD79BDaf2TzKqVBF0OYUsTeradtxOinYKjT2CuGAhbZvP/hIlNhWF
g4fM4Wo/R0cZbc7oEdy0yQxYk4R0Kedyh7CN43yaOXzSmj9MunEulG3vrFPoEWah
vfo1LzhM385IZ2+UPrk/HtQ8n3H1SvxcZixEJMeNAI396ZZXO7sjMDaxlyMTFEMe
RmlNlZiHHpu3kElGl1/D01d3Pkj30XgQOhhu3zhoxxixolqJMxsKlLmBXOgX9aY8
dAiglYqRnHgx0JnIt5YhKVWLECHbq807Y9zLzHxJPlila20SZ/Y73CvsMQa4DkeC
0S5VnOgUl05W7DN6IvOK5QYP5q4K0X9JNr7+DK6KCijfgECxQmOgIb9/lS4yw0d4
CeRJ8WG5RHIZd7CfxprrveaZ2e3iMs7IlJywph5X0GWCDqCFaD1VNsxk3/ijZFJ3
Lr7LHs5HqJOCHg/oRPGuRJ2MXN0oTTK/gCJ2QAT+EeT3gF9rZ/cjgpxFgclXCAqs
mzFxUl2P0PYPZX4i6DbsEuzJBtVw+6mOjIFO3NTWsRQmiz1F4N0PGmmrgxdVvOB+
uspd2jYDqM2oibjloSvMEi+N15CtxxOuGcAynBw7iQO273+24OsD2lAV5+zI6hjY
C5rD/Xd10SAFsJKO1Z6psarEVptyFqaPGYsBZO7RrhqQ1Y7HAgrNq0om8DCy/IN4
GUkJkTq5jnB9X+baaGpGtkUcGvfhSkp7343m+1UZoEC7kRYs2z9tOV5jXONdGRfL
Jdj/rA/T2G/MJMP0e3oUCFvjpnHQ79upbv8pRr35zxfT63yKpYS7OlPj3GDQ5fRR
VMxtpyPoZ+G8iEV2mIMlBW/2Z7x4AUHQGSsn+cZiwYBz6lKV8MoKVttAaaPwY6gn
WrALzcyDwSJKQJMCJQos2gEsU9jsIK8P83nQdxQ/T168iEG0yIb/MLL7j4V8WERa
7yqGeNWdb3k0nQkxRhbdlv7il4Okcr7lNh3LOdkQ3NGRTMU6qoRBSbQXxFvnR+OU
isdxZYF4m75rQyPDWBs26k6sWaSz6BHGOrHAHNV1+vyxap4208zh3BSg1xCQRGLg
uG7vqncpWUOd1AmV3LPWnCPKau6IyIvfNo9x/e8HE9EPh8/4CtoeZdGVN+i/7iI3
04i8rqmjFpC5MT8UflOD/x85ojRSjRoU8gmKwWeWo7EdJHQTjc8XMk9sgMYfe9OP
8Z5SNhsK1m+gPMVD9xRqFZBcFJvOW3vuzsD8dyEmcsMu51H5Ta6qi6u7QdZ4IWCP
EQgE7n3sxGjmoR3MGkT8mOoTuK2sNl1KgjmupGVycKWnHReok2ia2pESuHF8A51a
mza5SLYnfZ026+N8BzjYHGzmOspujGCsvOnHGB6VuNXb9EE+FXXnR3nZSXGcgWaJ
nGsS7CayD88eyvCqUqrTonazEa9MTvVfjPLLHFg94/YwpLien/3m9YLv/Hc4e3c1
N9j3ef2+O/lEwOmvLtqCZhAxnBI+oGv2uyj2lfIlEouW+q6W3QzqlapgOtw5HldD
u9jh8pfhiiIw7gdguooargzxbGp3xprvJ6mDakk9U9K7sMyWZxJ6vdjFQpx2NJnP
672iBwTEokE1FmNNsjLWgmnFsY72ZDAiyTajFOIZAqPyligInmPbLf1xq1LLmuTc
J3GR+vicZyTOXrAqsUEWL7OkaNtsEtLMGH2RJpLT/dpDS1MG3ZPbRDZJKOTxXWq7
mfUDPa637fu+2CeiyUQt95G9AkPi9zMFP8bMygEQsi1TdlbCJR1dHtgqi81BEGFT
qrvWsdi/gdpTUY9DB69hMMkGHq7ccMxgBK1N5RUxiDNe0Zf9JdccEUNLjx0R9qe2
UdPWqU16YDPKCYcuPZW5XWt9gm3sNsoPP+nn1SZyPL3HHqZq95MrkDIr+z9dpLvR
S3Y3w+53XRGivqfqjOjOXQYWRkFfdziBc/I2/PtHY6EfbXPfK6sqEBr/uDXPxl3J
7WJmGM5JP4qmBPNch9HFGmwa7TK0hoQOZ2OArdeuOsUTJ1IW1yGLG6TVoTkwvMvC
EWrWM/oAv8uyaKBqr95xc1nI2dEb0FjnsSZ7GYLlI9gyX2rqcoISEkXEm8NG1oWy
RKlSCNwA0LsapZi+Q7pOy/1N5C6idJBDhy7jnXKzewBi7ZlYIUDuHYurDu+Rpwsm
HT/pX2Zj3ZO/4vK54wNbA9ZBbLrO0GOfLhKxaAa1eayxfD1mcLxstR701bXlp0/f
PowS7JVLWb94co42gTAM99Xz82yYbiSQq1mbPoH12GzZH7oznggj7xXeIYgvk3Mq
Nuxcmt9s8Ym34d6V1UxpbHvke5+6emtg+jHCfS8PhJG5zfwiIoO6ioKQyrlhCSNf
U1LrYNqlH+VTE4/gBZvhtYiYPG3vWqJ5aPXGv30pF1MZSrLHbe15n/tItkUv23iQ
qNAt5c7l5CDhVzZgV3+9FmXOwcf6Ai6fqWdWhZYBvn3BC2zO5HXHXd7A3QHCpaYG
vRrbdzQ8gKR+wEY1GQGbSzIuCFdPGFhQM4ukCSyynWkMRWnGh2gXh6HBXFy8Uwae
WWE3jYPcnfeXqaiMbtAp9RQrOqrFVjAE1JMi7nVs/lE5FbMaEhSQp1D2BBHFIti5
bGhSs1E3hhWozlrdEeWQkJpGGMmlqx6WhuDUOj7nDcYyJx1XoSdWZEazmR5DVWXf
RV3e2wK/mPuhQKlraaMDsLgoEt5Bx124TgrmjwgNRQMK6usdMcZ1hb6xyvnSG3ZL
Qe5A1il5yrCYwrxPuBae0By/mMNvS0sycUHnU1LND7vjSVjyo+HAaYI5/IeFM5mE
H0XrlTUhbmIDonYI0J+1IzP/Vll58lmo5h5GAPUYqjB0OvZetr+mRbNx+PBOE+vK
2FtyjLqj7fMvOCzFeLji2g7EcSCUzHoGCgDg1wMyFeLEIpd3NJRv0M3ROC9CIkpx
1WBKTOudfEh+HfRZEbsnbyjmQL2YsOHviYQn1MIeGmImZVhHlUMlbQBXYGeX5PlP
VY8rupyIHPMbi1RUJv5i5Vk+5AqtI7tntAxUIiSnPzrkpfsoj/MM+1mgddkxXuXf
x6++PCRUWu+KgTJUDcg2pwwuwDAthm3Jbzeerh8BkE102eNR52a8r6TMM4Qz8wjY
fvLR3bmB+g7et2BZQ1rZ+Y3cuP+tCAp7OPEz2e8OZud1kGaqjsuoNL1MKzSximST
zCeUspfZtB6IW7YPW6RUFn4IX1YzbdRpWqgjnI0arIR93F34EATvjz6f1zkzGX4/
DSinDXdIsg9FcEVD4/cVIp7h/GvWYRAGw4igO7x0OoNWOb4NQReVKGpWWcLOAN6x
CZRJSZgFhPUrqmjCH0380hwiLz7FIhPvfzjqT+iIVvw/4C0H2NpfmlQ/WS1z6iqn
o5KKZmSrKDXK8qf3vqxPYYHsxcx7uYc8tBIK5A2ObJ807QdRtQyjiZCAcBdUv+Bg
50iuw91y/TJnzd+kLFuT3gewdhgUKZcNzwAeOpnvldfe9xT0dH5KFRogRM7AaU3O
cCJllEmn1fdfqgP8UVYG3bWK4zFpkHYh+l25rMQR2i8lQcaMxEl4Q48grPlm71fq
+NehzQQ7xWViKik3P16F2maKSnLHuWgTOG1kUbzbvy/pDU0XyvafOasmQmlKpNE5
2JvA5SXHakZjbwl56lGt9j9cqSfNTPFGn3DBNCmG5Qj+JbHtPxnjy2P1pN2avRUt
OQcZCiUeJr/6pMC3N/HUE9JFru1Fri1zuHZmJ5Oi8pn5NNKYwAHrciQDEHMgWJ7t
PI/SLth06Ss0jO5ISfhPB5p81aSmgHJjUsgeKXjV3VlfV9XJ4dpDw/mDQ2+UyzrK
IVKjG7IFN91Og2UWEmzONQfeHevq5y9z6P5U/LFotPqBuIuRuLNjfPdSbUkQtXCn
P9VxTcc6eqYzbyKkGpT8KIkCOtlBSKqNFIZqcXZTFIxSzqhhJOqZu4fVndAShvI3
BaFiJoh5BPNFH3FzSoLNDrY0wK3e3mStdbS/mZ927CWtvGYL4Q9I02mixthRH2Yf
vgBbuZkXI7QwkyIho5FeS8JkpY2LNVNbrP8KTUXtIlbj/090FAgCDAyX1n6iwtfE
vf/wrfc760Bxnh4UySQhcbsvhTpKHGSavSlD78KaGpES8zzwHIzp9gRQVMAjSXM2
BE9+S7chf8eQHjFk75V176oSmYMbeL9FyumNV1gEOkNFUqtJ8KVDVJ8FM6NH7nXi
9LlDJNRoXwREdbuyvAuiTy6b/ZsNSqsPd43pdACvivY7qA84GXFRHhqqXAVUTX1H
2f/6rU7KNOkEoxdXUT1xprkpJrJEKMUBHObW2g697myvOCahkNx5CleVWyEjOErG
1O2KSY0mlSehy3ZM7RdYdspODWbQ+UnC7QmI4BjmoUZFNBp2jOVDBVYWimERNe4M
pDmnsmraoQRa1+QmwGPOYKg9DTlQYQ6I4lKccDIxPq1lQYUCujsyhrWOlR1w4EYt
5eHiIZ7RyY4bLEF9LfIQQvwPRa+y/cWuJ6z33S/1CYoSeOZwWTn/UKco2Nuo4OZ9
HTsjruVaSwcVbcZGzZCMJ7hVJ+jRPfqsYIbbro4KZSfCQL8v+8G/UihOb5llhexr
0zpFy4YklUVaHLokYOVXcNp+pxuFfUmRjt15iFCDHd6QVvtUlCXFYoBTMec2NEhY
TYkk8l4q9KmXpj2/hOFxaqMva+pfAFLpp1a0tqUOx7X+NTRacVrz60a1yhzg0glm
wVpofmSxKgRyGTdVHaoxYLxRM/nzcRsxTlO2GHbN1JYijULpWtv4Q2u1Fpkq5Sr5
0ooCymUw/FYg7gx+2KAoM8qIdRxUqNr6mBzYhDGoqP7B8uHj+ONKYRVd398uBq3R
9ciNd2qpoS7FNpzMP1Yb9DwrHcuI5ibApEkUBYhQS1uVXlaCnvwLwNqHZL8+DtRQ
2Pqk7u9VU1Ihjn6folZ1rVQyBej+jLIuZWaH5XKltDNzPEX0pEod8DSPo+6pgn1X
rZrl9FQl/eZrb66u98PCQwiKr4rixbKY3j32k7HwIPwdEJqxFkWrnxMJQyrNYHBt
vo9osY44JR59QS1GPx2JBUC6fJ9TGKYS4V2fgCYOTZbb83UZc6O6Wfr070NP6ajy
mXnWkZOEXq9IArCBm7UEegmCRq/MoNnBTkT6rt8gu3GCUCu8JPhmG+fgV0c7ZFmK
LMs3ZZY9Qyqa+UyiKSEt+g7t5RFVDIXcdVOVQ6bv5hXq6zZyBqgh15HE+j6OqBaV
cymd2pGlgHu9HXF+Zck0Em9S6IOI2ysjAm4a4hevPb/X+cYIO2sXFmgR7/ul5Ibf
mVlwrB69R4vJmPmg4sJ/Xu8PLImIqPH8XG63pweX+Y2bsWaxCG6N3klowCXWYyWc
tbUvqoIUR8ps2U8/dZBIR/cot9Opl8BPx1zE5mWn8WVINxxv4Hq6/DTRlJ7t50eo
9IfNQfW/xYmh2mCBVAC+FlHCxZiX0DVyUmUxYflVEcPTuBuaBFVgbZgIm5xB8T1v
6pan0b9vAXGt221tgaoh9V1cESYN7nseD5pZEHCs08HQ/AsvMCaLhzwB0Mfii3Rg
71r3Bw0NGjh8sxk/UhyC+QvWxcxatbr9nHwfDG4HCsrcbGhqKpjxIDHI/7iAmCK2
x7EmYeFIBqb1BHhdo/KVkFWYq0tVB5X8XdornF8XFxcdjHEseCWaYpVAMvZ6XQ+r
xrX+5HjSEPc7MbqXfAxGOWWcN7vKGFLfZT4V7xW9rEoPcWbggVXguhCtyoKVrm/O
yWDVZ8GeWKbvedun9PEDPGlPueTqUTn83uUuTkOR59k9+ZxHeUdmsM/0JmtAiA1i
gQFgAjIGh5N2ACZupWWNRbFUIrKdKZfREiZvklSlRZCaTdZE7UrjTOd36C5dMEIe
1EVwdfO5mPSEUCKLigHusorfkaHMypiFk499lxHlXvcvlGIXVjtMP9yLJgIGgVQr
mqtfPVlwetzWLnHNVGLvnl2tW6+0nnTNd4qbvOSEvhTf56iN4t89Eh5CGx5ahYnR
RrjIIfjxeCLnYmunHI3+/a/MvKESkiis5AqjsKoln8lohUZr/kVd7pqrfJuAPwFf
FhywXnfH3bFTQQGgLo5SPfwMvp+B/rT02yXZKQirjbutZADzmoZYq18TTcdKmiKY
KGGwjq9MpSAH90CiVEebqPH20Lgm5NxMMhKBZVXwMsT0YsuLZ3/DwHeP48F5dMwZ
076DUi3MXD4CLjkF/tDvHf9UnP96+9sOgqryBMfD77lHZaMKu7zQ0dD1l/PIJXJp
MyHrl/qio3HBV2BWOHWhiPkD/i8nYbL9Zv65RnlG3ht0F/iqcWDZSzZg2BkQ3RQL
RcprQs2nMC6vwFoq978pU69orxk9TJgMW+rIHmD09OACPyA80h9CxLUY5OFff1f4
S1MZYDFO8Sbm86U8kawCk9v3PZKyCUY12lVNRRuBvIsCvjsex+adlN2fCuJ6dDSX
sE0eD2i1tz11TAlPuW04fUpsztdn3XI9cWAfBA0P0yQF0JDjbn7c2QtsIs4AEzUl
BHyPsdfYbDl3QzJVkMTxgAo4O9G/50L+kNmLt0z+8sBfkioiX13rt5lxcwmmI3bP
4J+FHRLwXVEsigKRRLmQMKlb9+xCveX3zE8r4mUxEPr/ZLSeoZ6HwPYd7BJx+X6X
USbkGsYaJyFve62C07L9VEtSWzg2qdEwQhJkhKAT5c29kiNxw3/HfZiDyiKLJup8
c1QZWWQYz7YRAniHMV//p+7l18m8tuiRzyrtIkYMne5uNSFkm8ynNG7gRd+7b7xc
oDWm0K9cSy2GUs3AFpOJ14Ta6oo6YNqeOHD4ZmlwfoI90vx3qYfqw3mcliTZZBNL
B+nQO5i5OP4AWA3WEKA2Py3fMUDiE2+Wmu4lmcgS3R3cMV4qwSvVEBlbNqkKwSMW
/1m0Wcv+CPxl4WsyFhzwRJgePOIkxS+VbJ6aMNn3u+ypmEaBuLf8NAMeKubESnsh
Pw73pdhhbF/COIQ2yrEt788zs9JW1cLIgPYiF1xDAkm4SzuWFO8VFIpAngPc8G8G
+7OYme5v50EXESww00MWWVTu6QZWeWo2U8Dw1MhYrGLBALk8QBB5KE61fxzYPcIQ
bfWjHfKxpbNejriJiQ5cNU9V+ke3pQggAM3/egrbb7RjkT7wMzxSxMLfxNmi9Mz3
wtHD4NWt0kYejJg1vFxWFC4m3Vsu2lZn2j0e5wdUODaMqs/L5gSWQDdXcPsxk64k
EqonLlj6F493ECYyxxGnDF6dvJOzK7CzoaA0Fm6l7l+ospkxPdhheyUyvlgIpDvJ
RYvyEtvTM2NCevDel+Fpdptkp5rz4mvsHwiEEFNIsvXBL1y3kB81dbUpv3HU31Qx
jCBB/fFJ/P5pgA2yB+Ohx++/++bYhLOlumN2kV/45Lg8mK8g6jMrT4pbIZOKqHqc
JSJJSIY/ITJ/7CdxZyz7tdm6NSepcr3xhjLcRy9XW489OMGC+VPYYy22wLLkfqwA
ReUGYtBm1z00GLPOfEuko1rFSxYbAXyuXsE0im2z3gCXJMYa6y1ztMM/k8wTJkvr
BImI18hFzmJudamcMGn+aaVz1ntFSfNnp/X6Nhj6UpfaoDxoxCpJ9TH4gUhDSTnL
N0sb0lHvUmpmgOP8pls+0anuF6w2cA4m7WiUQmP7K3q+DyuUXBS+xZDr+QpeDsIc
GzCwC9Ae7zuB8hqN/BioNK8B1C0l285Ibgv9S1rQp8+CsuScKUtdwD62PYxwd02H
BoOuWbRM1HLdKxhSYZyQ+dTO6J5wpmueG1ewPwzs4b1oeBQJWqBKZDFARl6t8E5l
bh2flpKT1SUfyHQePli+klmtcmTp4PhO9gp6Gj8+fPwZlJew6X0Ce/cApf0mAFme
IAtxGgSbJTZIvSlf0g0ABL5Lt6Iwh7p+WNN6tGGqWvrB4yKKcZ3N+abWmqBzeW5o
ScDrJ9tv8yloGXkDv4iU8IRnbwqr26Aq8N0utfp4tvZp41vtiUys1zDPo7DQnQ3a
dwDPWdJMjdbDIFtzxN26GOad1i/rTK+ER7jsCFNTX7YrY0Z+G08AItFzehZ/6TRx
+GEplUGpdiJ/+Wb7ATbwNZlOL2cW6VX7hgUorqjSiwaA08ytGBjCUHWrDgzEWuT1
JuG5IUoPY6E9iWqFMS3HW07XYyiZnFETyOJyFa4s2JPhHPOMcy/UT2/Bah8xshDX
3BadYtitcfaYVxA/aZ8gPlEV2fBjxpPl48iv7qnsDKxH6J9BHQVmnyXUr4wbeBMU
iBzeH8JqrXuS/XS16PeZcPrZFupBfQLgg26tRdFxZ0xxTj+Qh46nz03ZXKUQLZqP
Tz4HMuDjIEwDjRK1bc5xFTODk4bkixOS09AjVSyc1K9Wo2iQ4Ljjo1s0k0/HDRuE
wO5uCAxR2NO9wqWAtOgBp3xSI+dUwBjb/N+gAY4l76uKGXIull7B/M5Ttt0M7/X/
T50CRIOAiG1wKENl5HchNmBerZvxdka1IqXcbZ3VjF3TIZvDo7K5gkFnPB2Eli0V
q+LJAlZuBN1jOt20BHHSUMG26QWavjuamcc6BOyoFJFd1V6s2BrRI+7nZi+LQFSp
UBxJKmU0Brd0aR/WQpPIvJ6/weNCdIG+Gz8r+llAt/OOlrOpjHjcvV7F5u3g1RqS
8lsNEFICkmk1lcB7vzAyWSwQtnfs9qPjPJPchFNZhPps4yhbR2HgeL64tBfiQkRv
5lADwj33PVD2d1TnqD8DSZNMRVeBTptIySt+YFqOcD8MPwx64QIA7dMRHGcfL0RA
EWQzhcl0wTTYkK4zG6xMkpRWa8hAj2+hrmXMMwaO4uap2tVL3v43tE9BfRqNd6Cx
LosDQ4JnwmoFTHrzi/9RJXO9Ipr79W0rsXZ1GqJAsXLN7XzuUGeVFUBJuPT2J/MG
h3WDXXmTcAJsf/8yZgL8q/DjKmKYY9GwRXQbRcSTsFeb14xIfra4S2hpSDrXtRV/
nKKXffPoJVfCRg7t73h9AFW7O2upe2TjTvESPtWMXi4EwvJpcMGK/tFQjECkGUWG
OTKex9Z2UYXD5hdWk8crMK6JlYETxDL3sKonDPuAZPEBNWZq/WULMTy7rdeHeQsD
/ZdHOdTVI5i4jXzaB93KnXgGZnsUlAZmUC3D0o3OvPVAqnylHtCj0xT5XhPtPsb3
azFMCmJkuXiTv5NOzj1q4tb7GmPMDzztxm305lgYwkliyxRTZ0C4MXA5NnHCks6x
oKlOWHKarXwgP3uZxvB30C7Hzhbh1K0d9LfvdWXBidYLzAz99SvvoohF0C0pHZG8
5EI3dRUNcOaehx1co2WU4t83T0TKcMwcdq6uvC+wY3yIX1Z7n0usInYagO4ycIPi
pMLu2kMyL8r0VJUJHmYBdj4NZNls4ZdyxicUPWQ4QgfRL5xYJJ0EoAxbI2XzIgma
eTykLH3Q9VDU14e6WCeKOA8rFRw6DEQd9g4TvV+9/8pTF3FMbmwyTDUeBHhGdGtH
ppB4u7zsEwXTFn+0vbaRymbf2KEZqoRdz1NuuFSLSlmT+5zM4BFrQDP84xaQLnZw
3YoPTlxKHps/VKSCeX+PaGslIhBGUuH0x6tU5jmAuSQ3eJ3kekfRQAsiAzwlSH4Z
Mt7p6fA42/tbkgGdhMh4m07hDDL/w0XE3P318/+Gi5HsHC2Op8ymy2LmgRX0dsly
k94jKXksEXJCdzuSt6HHcK7zsClYBvFIuFfRm5fDPl/yJ32rOVptipiozuqehc1I
kOcD3WC/JmYlN0H+eCwNs3HDR/tN5sWhXc09YlZwfJuSSsix4fWd+rqNSPt2Ry4w
tDyctt6o1AWCTclJlGMSIJMHC1tvyPOL+/SS8Z4PHCGSPoCeUnngluM9YlN1MH5U
31dmpGlN3vb+AiVPHA1W5DH7mIoTVCnrKnAkr/q0EE5Rwkj9M6CKk7+AawdRYQAT
FkaF/h5nyjD4mP53Jj8nyqmPzcn/aA02C+cEyuafcG7xACbQp8/N0nz38RbbL2WG
Ac4Bgp+usB4R+vyxClMrO6lfkfTowniFgDKErAKmVMTXxHwpotME6Z35cPZjNBHF
UmfSunj5g1SqDTcrCHpNjR/wJg+2tRSiy1lW5QNkbJwVHsyigx88DGy2Hk2DH0oW
FaTvgwelbA9qSGtLKY7bypHNIVEhaKx1U6mBf0kXnmtuDxcqgevUKLIWM5rAp+H7
PhLs3xHJfX0AM9nELyQWhyO2Eozczj3FUViLVd6sdAp/uTIz0bsLHlGTz9E8Czz1
+yLqOMrvEIGYdrHNlUywyLMrAp6A9LcZsqlQVD07H/MtKldstndvngJJ5ZS279cB
+SJnqT/c1tfO2Ft4vnyvcrsvY1VZPBiCfSI8Egl6xshahMU9Iu/OknjvuTn7cM5B
r8CMZJlG9/nW7Aj3jD6mz4UL5oz38pCjSgxgC6JYPX7q/uPSq9Qu+twUPll3LJJS
rt6IYJo5OP7N0ru60s7jY3fGAjTvLOIaAdGVhbqPVI4C5S9YFy99DTaRq3B6zfNO
X0M24ZjhWdpEAtOJjRUM7Glw6uGHWEe9zo0x/fzYHUM4hCVtIlYtITLqAKxFaC6+
FaW66BHfH3s59dVlt/GdlbXH3V9sYG959j3qgKbhRqfYQSE9luDbRxVj0aUR02LW
aWV/2P4JHYmL12TIWO9/ZXwaLm/i/1hX5aTEanux4NJd5J2VRDOiCxkdozxrNVNj
WWC6whTjTxZswF6wr6lr8zOuIfGRIp7pEp0bYegsdKrZvpoj9MN7MMW02Yvzbulo
J4y9VcgH6N+rNPyuZjaa4erOVZjxDUWB/41biZ0dl2eQ0aNMJJgGWWMkUTPOc8Tz
tCPP6qdzibp7RUffM7PniUBY2ak98nuk/+fDkReU5QAUQ2yptznltrXVRPBctrUh
ZyO+dY/ey8fTcR+9wYVPAM5CsDfQshjONyMyg0/AYNPQwBEy8pfNPdnd/u9lvaCK
WNpYC/+X6W9qMSMaOGEt3tmK9hH61eIa+M9B/3g7f3ueTSkFszA7eYCQlngucN+4
Jv/zX1PtZVxAlZc0DoJeSaAucpWvYg+O+5kD9y/hZgMuLTUpgzqpj7cu1VCtY5S3
j00auHw80x1CKRTm0ltfgSKIX8kO+/+zdsBsYe6l/Erg9BmVN791dS1F6gndfq6M
lHNrNo8BB/FwbmgnyrLwEGyldDSlxPF0DfZkNFTTqbf85b5Crr7WDDE23s/DRi24
JD/pnqPRN6YojxeMv+ElRYUWaDVsWsZ2NAwTJevbln2rkOQ+s3UX5zjcWoCie/9w
nxKkJ0tHRAQjS+Vbo2IBmYFKWLlGaP1nydu2lIVRYYxPdNYEVst66XP4N+rFaMHz
4wB2SoV9zrbd0paOVcSksrZsVVTWQoGCbuv1lJmDhTOoZyJHR4UXGYJrsoyJmtqa
xspyaqQAuwQjwqDXFsRlrbxEJyMuxFDEUNDOwE0C+jG5QafGwr0PVNOpTHZFHI8g
roGpp8j6i7X14zA8QSuGAYCV5gZmPVFhh8+ytGSUOwTJgVbOmKJcALBQQzpM6SBR
ge2RnWRH1Rmho5P0EK4rn/jgbYiMeIp2/QqQWdajj0H3ztJzGh1yvHTg4Ox3C9ZJ
Arxo6kCvoo9wfxr4khgWOllQ1avto1OHiPDr9O3TIP08h/O2elMheUTWeOKpOOLz
YSEim6JZkCCOKa16g9rHDUZx3QXPwGu4b+jMlg+ZsxWZXvD1yZKyp3hUzNbOCUo4
hrGKnTylpiI14TCHEVnXU0JwjDk5VwM1qh9IQ/an4w5GIwhuQyug6dE9GHoSx29Q
qBOPmJSv8RBOPDGnuIR5WRS1lD7khIaAh+Mg5FYgF0lHknGYsdMZ96QRYQDkQGDc
h48dVGid+bXSuCUb9i/LiOzQWFgbZQcWibkzpZq/jaeZW8c+ky3iKd8S9qXpe1W5
A2XpC5H8U/Rs8G5KTGhOtNZZXPWqUJEFNLyq9caPa8i3pib4gvhMILZ9WpmqYH7y
l43eNt8XXP6sB8Has+0apjX+W9lkmg5qmh3A75r/FWnyIJH2TsCMei4K7LRcgFig
Ek3aV66TM0gG8m6naqMeohuKmWJ3ilpltJquiDC70jZRd04qmDZ6TsdQKUurYgGt
dEBMVcCgqHjN+szLS9gqobJM87C1PfyHx/fr9zH+9/VIUcetSVhqOB8kmf/N2dl9
SSXN1s/Hp7vAW1MDmVcPGZTkO5sKgo2qaxz6CRaRJb9+uHNu3t3UizYTzwls8LkP
inpubkhBJiqq5YJMAW4uPc5+KNqaY2JshO8lS7hzWEt/LKAqGLUd9j5nOQIhm4JH
kWzeP0hDvzFg6dkYQbdo8q4YG09Jd81MMEFpNs/mxL0bQoQQ4JWsTKVchj4ojQo/
Zw+5m4XCiF6dKYyfeM/R1qbxXTCYzfJ38B+Jozp88mueOcWsrWAvtYo4HAHlQADq
chVcXrfQ9UFdWnC6qsrssM1+xfGdC6ZoEWcAdmM9vjrecIM15FQNr03NociivzKs
7aqUfgtJCCN7Cw9119A2pavozx59dFOCY8PitFwb8Sc0cS9ltizOEFI4FOqVW58C
x4r5PPRu8YaYVDt3Jye6/4nTiYVHEqYyuNW/yXgKqF8vi51BHE/mmaFSuT+MWWsg
IKLUQlDglZ2iiGLpL08h6y0O9lZ+IMo9nxRb9QMO7NfYiBQct1FHfh5ifdk52mXs
qrWefGTgbscgKfSPyvmGyJ8Aw11fSj6eDtL99dXWJVG8X3c81RR3f4J1GiPZ6Q6s
X1Z4El5gCbeTvSgx/eTHdgdgqi2jn8wX9lG5Uwb9m/EJdHyrc+Rn3KHVF9QR/Crw
/lRgpIQKRkswLF1JCX/ub+OBtXrwXjwGbo5ryGek6CqRTApZOYWagTZVfQNA7KYg
mgUi6865+mqf/4xU4DDE2jMCUYykm2UDVvygWKD6BoKxwl/wDEqrodjanQFjIaxl
zr2g4crHbsqxDGyFYv+J9ejbKRV2kcfyxQy8SI3KciXzsJnO0SNyM1QxqeCFjmRI
u32BNL9FY0O3f0O4sKaub7ZCso0+EBs4jXt12soHtkS2TJVtl+zN4E9bARaprqJY
Lz6EbQmVMc0pnvFYYAEZdHoOFbdm1pSJ6Jou3lZWEDA+ePYVQ2u/3vZh1HG4Qd9y
wEogpgpSChiBOg3gtNjkUx7wuF+mJNdRXJHyYYI3zZZFLJ0wiIJSaeD+rAcBPnV+
25cT3bAqmjel/TC63iRfMfUUgYQeisfggtbUG0p4tsrHNbu8tTsU0S5UmSqImhv2
owy768gR7Wc7wiGaMLRnf4flMv72sW8X11zay5u88FEBXcxd71106L4OTKcUzXq7
cwl5WUMzNsrZIiIc4wQeMsQiOAXi+scnzHATmXCpz0pbKyBzhPIse7wKpAgZmmem
d1BGIcBrg2nNvQsedCANK9EX2CUuH2JJXDIQ+s58qklCW87VsIJfheZOMtPTTNB1
LxBVK3otUEYBHOHXnjC7wbw/1B5QIcxF71c3IrCci+jpbJkPxoEoKA+eBolkKPAo
4Y6KyxkyC7MaXernd5V4J2pXmHN66uZcScmHaxcQDgQ2UC9kOPrCOUVU0wZZQ7Sn
2VrIcktXtHAAakjJQALv9UjnmLi0zPTcPihgq416Ix29uE/el2g1qtjZgpz4htUJ
T3hZUy1wOunSJ2JJ5Q4Bm8jtGlllOBCULOjV8GzRxB5GaEcia0H/Q7HBqh1JZOHA
XV7bCAiISpdQK6oAt1bbG8LjbssfDaGDvDzhqs/hlJrNJSFcbzP3dozsGmArNOpJ
tdgtavL0uzdVtNT4wfBxkvBgt8HFoVlbfbKZYw4gLrQA8gMAQem27c9D0LozmbpW
MZPzCl2tjPJPeRZpJdoNKrhCPFfGIXd1lLrXRVG7EjSHYdCeiOSkvfxNcpciDwE3
I/I9qh72qWly7Cfs887w5IU/+Aaylv8S8j1EJstzPSu2xFyTrt3uhf4r0aWkhMMc
aNhS7fd3rhejwzW66h2DsAfggRyh4zxiCw0wNSpEPg1UoEW83U7aH67NEdh8KDVz
Cb1Gxt1zmI8d+50MKN2j0TakvTw9UO3hII/ZRv6/0IGEoei0JXNl5jgH+XzMTqC/
I9zxaChRgodMESdnNWaANJIJLlXxGbmH0HY5m1Ol3PjP4BVDIq/oEw96w7xtn41h
tc8DC4LSFyyCSD4pk5wsbBBy42hE3nIzUrs8Q91V0a0ayCrJj1k1VwBvrhqRiw5x
++du4g1aLVMOhPpoANjVL2Ec5wT8TBOsNF2wLr6aKHyK8lutg+tuhUyFy92fT5WG
u7P2RQb22vUSNvnbXTbLUHYftweKZCcU68DdZtnaJteOuMZnu4x/D9T7Sg9l+QLD
CoTBSvdpYefYbYRXFp+9cIPPtiafQcja2+p/VVPxLAxwqFFcEOCinnRSu2DFLQ5+
icqSaHax1tuTJ6Cy6WF0omy177rxbABAMsP6XZg0naEUXA9ssQKc4xSsp/CGzSXs
iQu3ctqx9s10cll/VMDAOp14xF3PJJaVNLPkgrV3XqtF8Fs23fe/qq3mMStqMj+A
vM4GAkjB1HjOTezuYtUzvhC+92Vhx8loj4YaD7V7viFwdWDphExnyLCY8H1/OwuB
jdcSyDRdU6fVFMcHo0HZCuxm/kdNGS0DjzbBEAQiIfkQbHtYMUHAOwfUI7D1csak
AMEyQ7V7ud0Xm2nX7QbgVkmaeMnCMskjLZlZDOgsVoWC3jOf3A9a8lT5VlXEIm4a
zdv7exBSlwLWVbZJvr+LShgbrfHlNjGEmuh7SjGR0nLqzww+tJAK8/CWN5Y2LegS
9DXDySl7CZcKtJuv2BYSyQbmLM53ubueQentU0QfxSkqjMw/7gEaKoUIVO8fgT6f
nB50bvSir6lSFAD3UAJoUuJY91170VCJQQ4ZqlkxFvTB7FkawOHRtXXUliJqrhg0
g9nqjnTErXxhytwb7kkyf0LjH6fJAmCaB68qfI2huTwsd7Xa8tSSHYMxZ6gwQE+G
kBfVRSBZnAzpVOF2HmsLMisCYtLCwCsEUDRlYeVjqzRXdZlewUH1UALUq53lreTL
l8bYVQOhHxTMyvMWP7sbMxZAb7JnZLjsFW17Lp7cAR2CL5g7DizevSElb4pw42iY
wVAz2+hS5JOXmJ9lQHVFZSqal/ynisfiKGC9+7qezfiV13MCSv5+V5pwX+RArvZU
q3/D1WAGcRVgSQ4ilPsypX7RJQxzGoDDHDb38QLnSdQn0pwfU4/bX0gb3FoNTbz8
6XsLZ3/w29+W+cv+THzWRN6qMW/UTNZCrB37DHRm+wrJLlSd/GAF3f6bZpcoKJX2
KWhU8hDKV97HWdRZX1/+NnTDJD/xT7uWopYEUhW9ZJprEY/7P8RnaJmg0NiO+WKF
80wiDYC5GDYksHNo/qa8Xd2JELmDuMdO1yDHAfKgpQvMxh03IZPTkcv7o3lWQpg0
4avAeK4e6NELp6B2RT4RWr3i3R1DZn88RMjpm+8Gnj8AhaHzbijZcJVsCjELWOiU
ZZ5eISwdwVBW0Hjuptox5aJfzARwdV3HaNTJHGQoXq3J4QZr0Sxu7pMKT0XM/nli
S3z4PycLNaB3HzBeH/6SgJ9EGou2E9bFwsO0rRpiZ0SCbi1K6yw23pgBq4RlZ+RY
UayZYp6JmisdBfdQXBOyWmu77Xk+4UkkW2/PAFYgB/FqoLS/MbCPOIsH85RphdQa
jPgqa7C6NJY1DShYDB2TGd3o/FLN9aoMfpMxH8CG5JtihShB2P2FEcGFOZfKj6lv
d+RNnd8UbQkiJsk8E3xFpxUuhDZVpswa9dz8BjhbUzxGQdYL4511/vHwtEEUauUP
m5v/3LBrPVoXJg9TmnjDJik4sGOTVPlb+uNrmQRc/4hrFHLJyMONh96t1nCke3fq
1jENRqxlumuqon1evYRpP2IwcNpUSoq8+phGQW48HzEajvOVlKbTHYCc7anGq3q0
cMsgV2LxaAO54PEd2uyd6fZDv+UtL5QgucldAZ0I8OEK5IMM+VHPIjxcouYJwpcL
PNlGADQlmiyDemNkTOa5AXfcpwD6JBYQFp09OKCbUmwuMZb/PT8q6M3lIHcjTPQb
bWxMHZRXlL0Zwis3ox8IlxCbou4NR8D/myI/3f6Dl+SRoGTB8veLp6BQ5McTm+wv
V6sh6YbsuG6rr1s0yKj+dfBWUOUmQ/+vXNO5XVDAvPYIAFv04Kcrssp22zupYBAJ
WHk3IdA79ZNqJTQJe1o3eOx8GJEX51n3u9kx0BFhTA1vAcvZ30fp/a+qRpZ38Dsj
+lophK4RSYVlrcM3KEongzDiXm1ZJyn+Q7SCSv8gyZuvzTdMbkvPoTpbNpODPpc9
bmVDU4rScKBEWK4GxTJFZU6vAae1Z8pMLgoqcwDiBwHl01Li8nHBhtbi5lq74sIa
THin82jEmLgxo3kagmCC5HX8ql12rp1/RGj+bDaoVVO24dB4DNE3rx45UV4grOf5
llYcAA1p7+Mn91xW3Se2lbFgg8B7PbIISoy8HAZXVR4w7+D6ky0U/6WUTVBZUWNG
MMVwVOYP7czwdDZTqDvAqua3AqsnCflhAFJvfn6zbSC122XuEqnjS3fl4SvscuqU
806+4JllsnZ+XGUdbq203r34eEYhYSLZTrncv72W6p1Na16LV4Xgk5s+06YNWVgo
2A+FcSRdfq+o5TUbqqoD3grkFG4tAjEXbrtLuLXuZLAwaCz/e/peHZzkuz45d8Cd
lqBLKA8dl0hQPxlxSO7fSpryQq0DksG53iFk3FBlByjg/zFoT3Ueo6HMhg4gm604
EuC1zOcUZSZbgbX2ok3pFQybhGc3A46LLhJFKo5ziA7yC44VV7vjlfJssYbvr/KF
6DLw+VDp6sBStneZwIckkwfcCbx/tF+OV0OYAWFC+trMHIsqp120Lp/BkDbzohBk
voG/DjGNOtJ6OOT7b/Aprow5ocBFdeUz8M1TSTtOYV3SdYyJaYdaCQio4bJJ/tKY
E+EA/UQCYtufN8Qv6ZB29sqLdv8EDEYJnjvemnfeI+zd32FUkozomKJbeIr5agHu
6f3kNoc3cGRFjtk9AXaRNsNf65HaAGoZdl4pot3K9mUH2xr0v+Opn4MHsv2R8rLR
kkXVWZfUipe5WYddPk27j6T3ZWTshUjChKAPNy5bBLfUijujEYJu2OnjbaXvoEvR
Tgjg/refvVPbwxjXo8h7UDMXf6yFljQ8PbKA/Rm9fHI1vIacMhcXZF5DjPdWv5Cy
sB/Thk+Ge7saCiZUd/eYHxDD2fnQNnkNyZh36QGKPzYEQHU4y4qwTmktzWf1YgTt
xoZ+AhCAgGJx3Pk2VJ3hl9+bXBHZC6IqpJ6NABt3lBBoOOxZLw8EV7Sw/mQoWYh2
NGcLMtYVt9gWC0d7/Lt2Q6Yd794vA56SGKicp/0nQRD5P5vO9UQzN180sVVOdpxd
SsdVWLOhoZMQXMpXxVr9KqVmsgxeL7GIRXtE+Cj5lDP8XpqQmG9o4+QR62dnz63b
LNUEZ9HKrBD7rKSrgEfDgy7FhOdVPhbNVx3xiZUxhZK9J3RZ4ECOgvKoBPTBupmm
ZH7f3BSufjRVcCGMepR9wUsRRJj6jj8Nd+SOqr+II/CMwYxb/zujFddYrFDF9fru
zDc1P22P/7do8CJ9puRKEzTNi8ijlhoovQQKpEuPZGSgYLbuuGP1PVKX6LojVzfK
HklH724QQqw+DuRGSU8bZWScDqYZmsght/3HSb99Uo6ScwUdb9xWlmXnibcyOc2e
yH5gTc+IOO+ct5YMAhwRAzBu45/AgE+IXaV/DxurI0C1ICCfEwVkPmyckLG7pInG
UxBLaR2fbVZ0MXpVaJOmX4d9cGnMwnFDH+WTkXbT5XuWfz2/FllK9tgza6zSZheJ
Z1zpqUIutEE6kTymgEb2MpqaxuvSd5nf5wXJANgQJHR/OpaxX53TloSLxtkUptAY
NVCXW2MBEHdn3+6Ea7FGBcC6iX9GvnHa+FPpQcp4pHZ4PXTIanhk9vGI+EoLRCs7
DCEgYaDBtNO1Az7JiR9+iGMfUTdNuvnFtiq1i0H+gC4jjJqrlTSUqoeWKVxpCv9t
MplzKJAM4MQ2yEHVIDH3DAbzYnsyD5E3PrKWSKeH+x7iuS1T4DwQfKI1U/tjlavY
JhcnRp5J7y2yUnch72J9V81J+s8DoUSYbp/50TbgA7ERSDyqjHKRryruxGpCGqSs
PSqUSivGEoJ5zgKfYTVI7364FJFLO1EXgPOoDBmVdvFuR26b1ffoiZvnBH9X1g7D
5GXfsZd0rQZkH1qwM3+Orj8lw42+yLE+Kq1UItUuK8cGVuk/TtA2PP0xrDSzEhOZ
tvcx8d68xn8TbUp/G+EcwiLKE6AsBZ1/uDmR2vds2IDNx61yi2Z7pqW1hobM8OyE
ocdultbW/YZJ0DNFbmxSC6UiClF+OeR4z8+hJCTpTcaNj0KAJahGRdNdFaNUciqg
68t93Xy/5G6h6RNc9UGYWKswEEvHLmaIDKjVTjQDvYJ1eG/xSPNfzk8F7X0zxgmt
BoJV1hY6MlVk5X59U3unjPwKPXobdz/ckAtz8/TPmwUDOrhCXgWwO5YvtU2NWfRB
VWlEVz+AEZ6ain8KFnaWyPrEINQXF2aU/b8ubqWa3OMTTsn490FCYK3f4Q5rMqZy
pjXANnlmxPaw0WDg9NUVvU3Ht5uNjAVWLAbN1Ktnbt0qkIFl/NzR02BrfvsGTPzN
BYGLprcSuM74sPFAA+kTDNbwxuqNki1JfuUjqxmMOJv+NvOPhECkdI7OuWgvCYSb
xtx/n8wLqp6416goi06PeuXiZzRaI3RHWzcyIT0ONygfptUjFPb2lDUNdDSBuxjl
VpqXiDb0i7/0luKgcPYEYtl4Ggnvi7TMvSgd0AKvpaAUj1j5k0h9VEWiVcrp1gHM
UvROGCVMKLHw7HrPQeSpUkA9ErwNR5wk+20tNKMmgnzg2QKigTKeSoyYgEPYMFG3
wlqDRWE8+/Baefp+ik48fQUcaGtdH683egLD7VgMymWiojzLQfVf6prsLtsGqjrz
rhDsIIVvYMai7py79hx7YL08JRpQG1LX97WElguFESfkC2IkqgCN5oZRg0LCFW8f
W+/DFsDIwnEar6zEJOKwIOCoS76vmMakhLWko5wtWffj46vzBxpXLyLgLRXPduaC
njgrk+54p75E2kC3Fc8K0upmCikBQ9qQKBhy58OtPR9I+HAk3u4D3VQz9pJjLpLl
QbH3dWYCRt0+QIBPFAnpKBVZH9Ge1Kb2IEupx9V9EoL3NDl+PNY0yjU6zF5fi4Be
tH07RmtxZXT8+h5o9mtfWW/KXq/6enc16GhKY73qOWZZhZuzpteLy1p0yOPZY2wd
+xej+kxWW3wCQq+eecf3/sIqvY1AqeoLiLP1N4RYVSucMxc5icB0/0zd5eM5EPYH
HesIeixotiIBr9fgJaa4BAVVGG2unFzcTyqx9+8rpFHjWTe0DUZnj8B2QLqPET0V
K4ub7i7TmUSnA9FBi+qjOgDCj8o/waKckz7TIWD8bCj2XvJE08T7Yu89/N9zAD20
zZFTtIBDWRaOYu7I/Vzsem3z8VRLHRychRxTkzIh0T8Y3Nb+IhYZkLmyIUE5K4Fm
QW/z/1ujpRh9JTIM4QbmDBB/e9/r6/Jtc/SrkWWKoWfmFpfqDlRWv8Z9+ZZ3jja8
qerIlZDaaBfNPCHeP5zTfKBjxUtqgFxx8il9+ngzrFjFAUVGmRVR2tKEHh6bRKnJ
90HsfQQj4fN9p46e6OJ6cWDqcmXk5u4jvc7Q1QP443KOLHDMe3nmnPff//VYOprv
oxhA+WhDLwwacaeBQSWqVyXbUo+WeWv4s3fDs/WJWUblV9FZedvjgQ5e+foWK6xg
cQcF0q2bFW+M4c7suEHSMKGTuuNI9GicTP9TW2w/KmQOB8wmU4wbYUX/ZMPqwhyz
G7CVeCt0UEMIZVbe9AUEDaCusu2R32mXYYEiOzasiXglcqA0Jo0/Qd0CMCdbRs1W
I9/cXY8GeLZ1dkCMedMnanhvnzf/PTPelalJEzRD0bXptj2Bd4syQXkkpdwcv2Ec
Ytf9mx5lbmjbN7S/jQB3PwTLAnGrqdmNR6eSiygapQWe4Lkl1ZJKClnaF208Xmev
NfB5ZlvBtImnrefYYwyZtV+v9E4giPZO3rI0+rA8lR/zUs4cd0+mASicqyIKW4R2
wAY9J7gHJxSdkF3IY3NZK3HC5KGwMWLYcmOKXqIhth2uNjNGe+oNqV1vh8Oe5KFb
fLeDcGrTnm4ZJPlU06K4rAjQy16y0nSvpZHiQT3SL7C3IPpTGkypZZTUJF/XK9rG
i3Ern8a2fKo1119gGAE0t822cf7gqk2Duhl1Ujk1KblpUDqquSzdw9YCPAlLnmmT
hGlalypJJ+GEBENwRsynvqN98jdfN4A9/W8TP+DzUdQtwxeCaX5KhTawoPrmU7Ok
+g9vi0e8F84IF8rZnlrUxuHEAjEK5ZaFhbpsioAAWjhg02zEu7WQR1HdMdBL1Qao
fIP1l/dvw5ZKsaeYKjkEAW5GUDriU/4cq9PNzm5x2mNIRRYfSAcymngycXXo8Zfh
MCy3cdXa/ca4PLOnyj33NSzzBCTTxUnj+rr3mXF9wYdM7nWj45ujmyIEKQoXjQ6k
5MpVotnDez4yCJ7L4IPOL1Vt2HahiYLFC1l1YFeDCLVlB3OvrfgM0XhsqmeJ8F4g
MWvDw4eaGC8vCi8djgR9D2g9X4iZZFyZoA5ziKwsGoDWoA0ZZ/IbV9oOERLBdzxR
sifNphEadK3SdIYSRomPKcsdO/W76L7L7Ze68eGQRCJG11+WiE4A2wthyMYp/JvH
wv3zp657N0Hi2CLA3SDTOX7TEeNv49WOgaSF2bfiQUFfuA20v4Px7bG1wmy43IKO
IN/k5LzfVogpBmm9i5S1kxhp05DiWMlJJJZnw6pCbcs0BaianqedHCr3+ZIVx5bI
wbYlYshaoKpuFXqXGOe3a3y8lFi+eI6lqAR3GYd5x1fpx6NIAbIrE5p3dO8nIM5c
4Nbw4QpReqY4fRpIBGzu3L9jRpmYSw5zdXPMysx3TjLyMFYnkGFavbFyzUTKWaPz
gjbOOMEDLB0UKtlN1UkkBbvzKemyRZfaNVFOK3PblQBLO9b0v1OujEgTv/Ew61Tj
PllQqrtRt1By/VJVOrQPebX4VK39oakDB+1fpYtCTs0iMMWrbY4NSevyzbX9Lmej
T81XbQPf8CDfe4YsE5paAG37cFmSrlH8pHY9TzOK2TRTN9EMbhC76ENHHoj3Vh9X
kTsdD182WkAemWwQYBbtrwtp2GaiXF0jUZZGbRTtdj40fLLA0iEK57seva0wDNhh
yCYJfEwlI/pHqMosIPAfxfG19KQhc+RrHAFuXtorAkAXI47vEBlt1P2UjF/f6rcK
ExfleJRE7oj/xKp09x73ECW32C8KS5sM5C+JIskyDkwwETb4YPBHgcMLixWSho7b
O1imNlC5YKkRw2JDmDs7XbMmnMHcZ64ex/psUH3Akwooc74RJtlBV0d4F1dOJnLm
lghqonuA5IKFjKDTJt7a4xolJGYmAHzBH1z2cQxxk1TAsrnEqIuNqtfO0tuhwf74
BbkhmJvopSb9Cg151xJDvsoSyZU6RP9w89kgqAQq/31IRNE0B1qQjIXX15mMCcFa
pGi7fTdEEYywRH2QxSMjjv4no/PuDXtsM1vha41kQNUP6oUaleLSIk/iz04xKsj7
jmdALC0ZeeXWdHCBu/aRE8vdOUNv8E6wzUJ7sH1X0FCHNmZQ7/auCoIUdGkufoY7
2AGz/D6gopNi+hb+tFFiH2Bx8dh29be5lx7ld7kP1ghClpL+g/L6azMrWkNe41Bo
h5qaojwV6jUutmnoD022hudjBAIlMY5OFSDQCd5/mc1h+pFNU0088XtSvrwSJITx
nPbKyVX9BNlvfIdiMZkd+Id6GonvYHicRd+fq1O6SrtTn5gmSj8iDm5MAAKhHAwi
z63N8LQnZ9cSZ/cgxYIL5NF2BD0o+33GmFl9ZXVLOl6V/rCgXefomHj/xTvVKIGL
+JY2nFAE+vWSyZ1oevXCzZDylRn2++LQLlOE30sh6pMBksywaEZqby49uHJ3zEgp
26bAmpWY20ZEc5McKaiw2Aoo0raqMm6CNsVA0pdzvn2udgR4uBpd0zmvZH7BxYNX
c6QveF/soTTAI7Y5bYJ/4U8flaOdCdqCJMeBtUqunS40pEqWjixXEkhcol/lr5/j
ihvOC7L6l/xYSauEVztTjrccu2MsWQrt6rOK7CUr/+nCfIdlMGcLwhByPvsgXcTD
JXvgCcLme1VHnCI0rKXCFDCW9B6SzqYlZsEAATr+LK0T1TEGLpwb3brFzDTzsSq0
M+gmX1jExs06lE87cEIXYSkaTjHcVzu4S2dlfRAt/6/jDVJPqFn+JpAPqPEWeDyd
RLyqPXQqU1JbA9mzShXPNAPKlmPoan98g+vBBM+mqW3o93kLVXZGHyh+msb5Jorf
4GyenrM4aNHJLblsW+Wt4H7/Nw3wahyLYBMFqWawUiNm7qjLPPNDKMj1OlZwG2CC
PzJweo+/wkdstgw57Ep4KxttBj3ktdwFy+ChDq0hRXhLqtpvUdQsmjVESJegsM93
TpLBocI1sQ8W4iqnW5addqIDARY6NEND2EPZ/Jm7ZzYdsMpF8ebEc8aHFH3ZV2uP
nK0NdYIBZpe5q3wj77cQVkROTv6M+op3jR/SsBGdhj06ZdOSMDOzSn0wZjd4r9x9
DwXwd9Eula/ICoZZt53AaSn65L/X2LYwf/7XaF9KZbZdslYwQDHicnzov6KK2oYj
1jzIPd2xpBYreIUhRXLnHQaOr24w+cBs31t6lmVvNVvGFu6urCbLjKGMeFgjBbxB
jEM/fLhH7GlnssntNjZXIplkjaivyW7FL9zCwoxqfArxdchFurSCqhYn453IF5yh
VPHgmZmNnkT+V3nzogUnF/1e11KkPWcchzBN1XivAN1XYfzMoC5SBl20SAL6yPzr
C8PIYJ9bdxBGwQ2IXe1DrVeyetcksZL7doTgqvfQlpUG/Sw/KXmEZyDB9aDJqYWi
FwylyWMl3OE90Jp5sxMNqwDYgN6yxKVIhbl+HAgO1AbaE8yVdeCqYHEXXxXE2YcY
Kmhz9fo4/Qbezbg4tGw4+jKXWXSchy3pez+ViqM5pma9HYtPa3/jlnB/GrQq5j4A
gMAkhbwgKcFl4JUu0NGRoPU5YUDWD0QbgM8m7PzlJ1RVYCEV1cWNCwALtm442L+0
KlI6LTm8PvlQgp+ZiPbiIfIgnjoERFu/1KKz+NRG4DRSlw/80agdO4mq97DMVk/b
L0Vj2+eLiBj4wmJmQ41Mg+OnvgecqYj+wyhyf1VdRGW27XRg6aJMRbX+0xJCMulO
jAj+QRYE9iHm2bqY0V6I20+0/ZPAW1QNQkfYlDadIGmjXLICJFd3EPuqORYTAi47
8zSm3hrp91WGCvh0ESc75PGGfkY955EfGS03jVnErAYA9MEFio5ZsCJh+Np2NcAF
9iYXn8m9O/VU5LNTxakSxpjq6svKns3cujO9Bzqx03TwTyLpZjTbe3Vdwfg4LOXO
QeUIlM8XjGhO7rGunXw54QeLw8uYyyRD/JTLsUE2uRRXoRpn69/wNtVFd++dAg5a
zn5elD/CkBhpo9AcN93te2H0sPzJ+tSZwjjbPFwBv05771C2XnR5u9WOyUsNyXzc
Xyvu+d3hXdYxqrp7fs9FQU5M9R9D/4L+BfwWpJE3Z6sr/sYvsywPc4grSgdTzcdR
TfU6JJuDkjqPlSWjKXNrpSkf1NrGSCr3W3G1r0+Id6iW9IAGbyvh7erdKX7lLXjt
xB95DRPEfSH3WjG4Lj1PKBsvUcAvC0BdVdX1sNepQNnLGz3xmbItb886AemykvtA
MMx8RA/Q+nbmL68FzHPWZPZipgY7mXYwdJletkL4w9RA0UnHpxnBUdLy+uzAZdb6
1X10ZGK8hfFzKicvoO8hqFxbOJflufZlw5fwfhZ9qBEYXXG6HW1BaaYk3lYK4hVP
YUKoZHTgHIcnFBfnyzvp/cKXM/9dwqVit0kcH3wqUi0yC30pHbdMOvb9oq0jWVdd
WsnnzZr+lDvwPqTylponrQsnwKLRyA2eBr+JZedSEV35twgn2uXXpVutnENBKpC4
10PNpuAnRWjSSwT7oFKfm+0fN3LBi8BDPkGIaMkeZMW4EvcQEJkT5+nqiTq33VXG
kcw+Ck9LjEW+Y4lg8X7hebY58aVH/bTx64PfXMbx2Ku8WO96AK7JKYZmX6PzFm1d
71E/TVjyJEg1SSmXG0QSbpC4l0C1HgGYpOaX1pHfEXQh0lITIXyeJ5X1CeFqQQS9
3YJ+7pE5lv+jjZnN1/xUuK4cLHnKkJE7XUtiL7mhYm+pcax38afxMaiPoBBmNTT6
6LioqCKP4aE0H+g7r0KGb90dlq9z3W4XkZBNqpky9+I/ci8IHqoYxxvP/J9eZrpA
hNzLyqhlA1YoYK6r9HeltL+iufT55Byo3P2/z+VVDKa40NgK0kJJ5qPpyuCkjoBu
dzQpw9+vz/FG+ajmDICVSmhqDsKLBWXRSLvQDBZcwlH9MpeBpi1l/Jh3s1HgjhVF
IzFSijOrKY2/dQxUvKaAQ/od8pcb6SoC7Z0CVsBDH5Aa2QYhyEOKyZobBysr2Cj2
x3SMTqrywo7BXhaxAi7q5HudMZsVQZJKwhCCZer/Sx41L7WxoxvRsLC5q9UtcB+A
wY9JxhAD7tz+Y8cqtk+XCGTfE0Ur5f8YDOX4PqcXT+qtdsHs0oFMnbFXcNL29r87
5Nl7sq61zyANnfvtUxO5jw0YuvkLpCkwa4RPpL//cyx6l/LgFT/07UfMfpMVX4JL
KDIMaOq/6Mth6oAQGs9PcvXt0w+tQntvPldxzyqsF5t8AXHmORZ5TgjxUQVbiZe4
75zE6y19uko1pzNiolOtR3RtKXMNvUPkCqT4VbZThtNrrr7+x7oXU+zskTBFJGH8
EvNZ0GM0uFucfTTYq+jrlQGwV2cID+hlLtr1dRR1d4e6L7RlvMuitjpsntT3qNES
ud43C4Mc/Q4RJLF+btAiHvtOW3AxRJbwRddXghvUsCq5mnIJ54o+oHEIqem2yYTQ
ioVFtPSrjD5/26I0PibVujsgRbyw6IH6pzbo1s4oGUec45CloswHsc8Y3H4XME18
+LIOOugWamHAggzbjRHr+YP4kFKK86OkkQFU14FcNYETrqwca17bclV/Fp4xKM2w
gBG/zvFTnuNyzEn3d4PP/fpMKO+SSXnIszWUP5QEv7f8JQ2vxz/JkzoxHvvkB8SE
mz/CMbP/cCnv6Qa9y7Ox6iSkazqs85PLaUCt29mnb330e/VvyjNdlU5gyZspEDEc
XEmdPgGN+uyj0rOr1fMM+674xvcB41vMwh/NUn8BtPU8xAkg40VzOlvA4/ZyP/z9
p9HitKbv33PLL8JTvmLcqcWOYtHqtmqslj7QxsSmARB2hQWGLgUTy1GxYU3/Z6zM
89Tqzt0ZkqF5JglQFhkvZYanWf/SfmnrXc4mTlXoXk8SfCIvzFOALvhI1j0mS2ol
dLpOkTy6Ik/I/hM2LLsg4IqXQ1ynY88BWCJ2Mng0jEfvL7mahV4tn8MB6qshn9IW
TQppleyIFoktZJBovOqtpzPI554wq00LSQItiFc4Ryb364zJy1Tk7+ZYmttr4zM2
8zo4rs3OXuLNabifzrBIjCAILGppK1VyZKWyDPLlUTSklKDTUxo4irjIUrR1fPe9
ykG9B56sW5iNhpUh8vcNJ7cGu1p4bK7hYDqamHAGLi0rnjbaLCzuH2HWf1Vrp1ee
VIe73Lw+kAAOlBpKXD19nQtcyzkTDnqktGLSpFW40jEDphnlkvf9oWEv/Jt2J34Y
030EPCCuPrK8/0dHSFE6lzqQqiBobA7RiqSjwbNiTLIs9QHzVkzVlB2EpCAohaaI
AKfndRq0KZUvOtq+TdXw3VqbzrnFdsQ4NjcicIUgWL17BCrxy3jWZFXabAV79V7v
Agyvcfv+y8+usnMtS3C/OnyyUpdzJk+KPXcOOymmVG7gwPLVP52irdACeqfryfu9
JRFYJtokQ5KAyjXG1D3ekTqEva9cQjXYpSccDoixi5/cGHJv4rD48UVaS0VLZPeE
3kHMaaqJEKpK2RcLzOXwg77oPmMNqLlAEEk7DNfL1nFcE6MHAJ8DLa4Zuln6QSO2
AGhoTLbk/FokdBYFEFSz1UCM2NJAGAOPub63gh4N37flTL/uiZ1CJ3MXZI22TV9P
ptKGoPzsS60UVGGwSIpdpV8tIvQH42NFmqd681zvDndSJ5TJzEjcPDhhlFd/7/Q9
lldrR34/Et2TZcdcQbCOHSJvB4PIXGwqJj3PDpMA8BB4B6PQIyu09h/jaiiRCj3p
AUEil46kjSpbhXVJZgnvcuXCk1aAPGbA81CXh57p/EyJ0ED2AhW3irawjkvd60+m
XyP4wiwDFuv7WGvWWVvqSSU/x+A8kaPk07teJlQRQHMqrpGndmFm38yiNWpUU7eD
CQImFxs6TBH+4PmDpGSgxxAI79CBc12CtFQHqO0mwN0sXNmEz/dPrYpxXTAK0wsM
lcETwOU1omacd3aXwrb936Y7NhW1Srit4CvSi8CPd+zkP8D6Fpo2p1jdO6ukEXuS
JyDuL1gcXF74MJaZPdOgxDHmypUIKnsV7zZCjlexc1y/FGljFy59uc5k4kv9YK6n
zNKrZOpQSC2zNeEX6+2ItYrjG5eGDGLZRImPSBWHCwzy+PrVX47b0w+Ztd0D09Mz
Q4YwghhSs7n4yz/JulwpdBdqOzzTe1vmK0AfOoLqW2DweDmJhlvPTJKqi3dkzT7L
a8zNb6gsS7HBgJiUE3in6N5DRKzZ2slywuI42VlwelIGO6r8nc9lwQ35VLQmfQTf
RCJHHy42CkB9chz6NwLlR/0Y0yUgxgD2KuXvJW4vxqJ6ziOz81scH+OpCPcJLD/G
TZsgJlyB+gsimtWoOGH2RGPogpNWaCQFw5MsE/lDRLybFBfnm39JZHfNY26QYiAo
SJ1ZZExxuCEjmw9VBOFwDH06UmQeZQ/Ij9/Sf1/vsqJIB5W/x50jZgyEDQtha/5c
EjpO7T/89FOosNm3nRdvU0XWni1xguGm4R6nF2RttxgMIAepJcTxUN+KLPEcqLSm
Dz1Xez+ho4h0fwdQ6+iFsckGTl4nhro69LCC57PEUAZPoh89LEneZ6S14LUDK2/m
XVavp9zDi0efAXQa8DCNmsTq1UAC2yvyWHgaWTCxtd36eoKAtf82q6hT0zNAzWp4
u28RWgydrZ2ZpuR3NYkh9Jb8NRTrp6z1fPJpGALAx9JOs659UqHVpit9BgPsH44W
BrudI1ef78QBsKFZJHyytTH9ZF8SPQFr7zRavkFZuIEYPM0p3WPijCATF/4xSNLt
gbPjTF4UVXLcxn53yzqi2GGhdAnVmDg2yOX6i4M0BFBpDf8TZTqd8lkhBn+yj2ZY
IHBCxp8VCSz1b9y+gPDApip4yKMAKqxJgkiK4vAfa3hapPIQnihUaeE0SKPe72mu
rMVP5TMSMMCHLQXeuG+4CrBKhy6aEjSfC/q2RiVG9XM760HKMaQ37506msF1In70
VUNUR0Ypobni/YwXIfKTZ8ldLhsVkI8CHkrKFMrlPdSauOjFjMidK9VC6ls2kc/V
r9Ls6mGOZUIOKEiCtdMGUbs5cei7nHEwfzILqmGXZaUmD6/HWwsPrLAbN65U38R9
0XEpdlJW35x7ZEJ0FvC+7CGTsokBjTmjBEqqAiz1e60UXwIIDP7bhYjcj/Bqv9mU
VIJjjY3JZxuG5CpzCehk5wDEu2U8pkA3Fw6h6aN+RoB7wT7gda5nNFWFSBPoW/oR
k5V3+B8pyJ4+k5eHueursuVaIDJ22CyeXXVk+Sr9ZCyMFArQ0Jlt+2PCVn1N8ycU
Pan3CzqgKR6412zsYK/PPziK5i3ACOtpJyPLJpRjqpR2xoK8j6mxDS49OKhaCKcn
xh68jqnjGNqDl7DuSg6PK9LCnLNdgqUaaJ698/54KjhrKsQOXNO9XokR1tC6O2c2
HGlpK2Ppw3VyS6AroDrmmUEd2aqiZyt7gXUiFVgdmkZaxGSkpmq1W6cV92gReFBp
WaFBZ6sQJ3CM6hpRnRhjxGNXDQgRtBoqla+W+FKpGe0pMNnQPp8RL/VaDFfF89z3
ieUpzYHNNJIaKRhiU8ziZ28lZNevd53LzQ3hGl5f86p/7nghslIiHQsr0bnp1a2C
4uHmJon+mi5s9wGnFV8Upss6jeLJGPBLpzj9XovGII4fVoH0DlwJv0i14ZYxM4Bf
mcHEmie17oexryDonC0gIwJV60tuSzqVqCRs7OWCgD5OwTMiQEr+DpQ7Y4Iai45B
Go+p/W2sidgFuFKZtkedjfo77f03h6ZDVuVJKcKxvLTDwuJqHr/SYCM8ih4Ecoky
LDdf6Jq+cH662fPnc1w3KbbBf+uRgjxGI3nwvGHXfEQMuBCBRpbE6Peu2LuidxiF
lMPikchtSoL9exu5yPLzpply1mg8gmmQWu5xq/WMGMBRkYShPqkWD93B34Ac+wp2
3kKE1OOHSohrMFVQ6J3fKavth0QobqYkGHtYf0rOIFfrYin/0PTFOPt8yEnnxrny
kso8YLdVsIolE1VJtnBg8P5ZPGLpPwE6YoB9e+YNoRk0P0xCqv5GPTnDAXsU18T4
lvBweryeZFfKSaxbRmGIPd2INu5y1oBotIbXts3nmaTk3Bb9EvXSUGzFPTV0da3s
CDvLGTdROepCxjI19dWWVvY5iloX6UP9ZLnIQG3GoxTWklAxjC1WTVDpRKTqiAsQ
a9Ee3xTfx0sEe5KkgNFv0r+SQHIBlTdGC/44nlgR3iKBWliLt3ms9RPq31ssESfv
Wl1DmYFWbuQPqDPc9Orw6uno8UNRjKuOUHXU9Z2Z7G5GEP/g31prCafrGwBM67zN
wzKPstNZzgtXnfVQu6htwx2MmXe0ZcLpqn1dJOlvJC71hp8vnU4BLCZS1L+NrC9f
ZvsqdtKTuPvLPvqah/s79v54k+OgdTASNY3o+AjG33SV27GKKOSggMxlt7mFWUQ1
8oFu0WTpJuKGDGQ2AcNXEfLvZAnU/usr+aO+LckZKIV8trnpuAB0SNa3DPpjV0g/
2h/e1An2UukzCz9nLk+VqHR2FxcEWGUL7VOnhDOY5vUzmt9tDlLgq2YCtaQDtbRF
x3BXSS12OjNuTP0em7UiHw98fWvZeSo+WkUUIOB7/8eQCsl2mQPOYNgS/QQx4IUb
glOy7B2kjnGP3jonJootPq9S7YNbZjcraaJ6NwCUrxAeoZ9ru19FlUgC4YK+A0vV
w3F/74cWswkwgH/P6gkJz6AxpoZVT9fAvbR3NqLQusUe0dQxm+uG0W0zKfHHaQQt
uga+y2pc30L/bXD96KFMF5xh61g5OSATQn2/y8BltXiCoFYr9WgADSoa7dylvNbJ
onPb/3KLoPqIY2GuQcneIOLl8WdatRzGbZZdpKWVj7VCMex8QyF6UjjuVktMkgtg
eESY5XfjbZ7ixLdX3eZ5shain/BjX4xJoM7uYK3mPCD1Bk9YSebqMfbBbuZh2mLe
rk5sm6o9FfFTy5/4wbHFV2X2DCxmJNXoSyMQpoayaxUA5mXYxSXDmLav2SQNwpS+
nOiqUxkDH7oZCx6CPz1nOIiAQeh+SAaJIduxOIm82UnxNhy6Via9v737GCzsO2N9
MrnItqBvSl0fcEiZjQHG962aqpiFyDxwZBriudEhx6YBGVN9xeeudhP0SA1mZQZ0
7UlQmUjGUHLc4rJuGgm8+UDRwUVqRmod3ppLzuHVIs8ineVHHRF2Oh2mNGFdG3aJ
LyjQa4plsixKvpk76QILIBRk8gyGFoeSJFMj3to30VbIgMIEFZ9pb1MlFJYqHpuo
ndfunpm6fNj0I8KI7v7ELu/+e+bvw5cWZn+5z79DTWcUF+0vIq7Sfnlw8xpXEI52
HnWA/ieAlq5whTvAl9Qgptd2MFSPgx5RSlT7rTmDlA+hXOz52OF/WOZopmVy10Vo
ybS9vNQuAPuFrIok0xTXY7pS9GUrrIrfZxGgUSO5oTnG/3lnQROCdTTX8ecWG+6K
vIVowqVOu+IT6++uhrnTEfhjApMXY+GXWdwAiPwJa/wnVRg1SiavyogMKZki4o5e
wFp5bUid6I/tJDRP+JMSq3daiZEtYXdPRAWxb5KZHovAVshZEtTQnbIu3D4xCEs4
8O7jfF7Bk2pzqOcYNw7lEcqssDq06boyt5Y+L9NFI2Fn6kiXZqRvefiSxFluncgz
Lod27UCu88f2/u76SsZdvh7TioUzFXM1/4KGJEG1B5wFhkmjobjHVLRTc/PofZ6Z
9hfMQzP9Rl50MQmppuJNvJWVYghpOYDacr3/3kbRqe+dU/bA9g1hhwXgP+a3zmMc
vBWH28AK5jyD2GtzK3xV93K/euBQHZwqCLLS+bHVwkI8dM9XZcl7q85JEseLRa36
dxb0DljAvc3I5+zfBihWj6iIOA46OBYI27Sb16kMRy/Wz0KovJ+3Arvlm5X8+z8h
r/UAJCACXqhaAFIyI4lTh71fMZMMkfBai0/llBZhPr4Bb1szI9txo5OhsZ0ISAMt
OwvDgsd7GyceCXdb3zkpaHyfd9r0hafR5odd/BhwVQ+cxcrilQLDX6MknJUydGNM
RDr+ecxE/LdnLOXVttAY8fA0XLuGoBxbuETVYMPGXEH8A9QaI2KtW6hIPERafbl4
C1EYCfpS08D6koEVzqyUDuk2O9bcZkAcAVY/u6Ra87Ns7cHaP5mkzozEQ8j578mo
YGZwO80It3VAmeeCvM+MlEe+UD6PIuGVHFvOiJazsKiiLZWPobzOauLiOu/QtFoy
RtUm27lnCr5uIWgW0ux+/+ae8OJgQWWuJsXDOPkwjpXGzzLAIbwJPfMDq7ix1u0n
b7EmZwnf9fWCudyQMMBguTxPmmfzkE7YeC4MQ5OrCkJ+QE2SY3MFAOQyXWBiPdKy
k1eCfx0gt1PE+UAETyjZPZSe8gdYtj0xeXxct7Iuh89jrv53ajXzi3M+tbYQ4rbC
zNORQk7Vskr9GYE0ZrUE1pqc9FO0YwNoswvZ1Nmwlyub/+1sKVNbKyC2Bzh5bzjP
8k6JtTeQ1tLO76T+8pFkCoxpeKO7M4+TeBKZwcDD0a/AEWmi+DcpuFR1p3PfTslR
lAjKwNk6KsJgmayRDhwURDOM23nQrtx18GrcDc8Bsmdeb+sUvVUdOFPYUI/QyC06
CuOu590nvFg4zyldigASajWqBNHauzY9UowsifyUDadJ+Ur5/RRGdxLbv8N2L6bW
Kf/tV/HaUwS+Fd5NrJh+2sGK3oIlgZs5lEoYww1o1Mgvs/0MA6eEn+rASFuLMxcc
N6e4J95CdtsNvVm1Ytw3Ci2PKvWUyZdkTWGzV+m2kGTiMh8wr0DvxMFrHlCIuk9a
J1IQ8rwTRUlCbU+w5F63ObhQW/6FEVoiMWw1tqfQkJNKSod0DZ2OHIWurREqjPaP
SzVDa1LaVQC8NMbl7mMFbEv4ZE3mYyU4g+bveveHsywRdpsQzsqHjMrdwp9kLArL
Py6kXNBPSU8+UAVt4UftIfOPNzdUhS2TeXcRD+k6znBhnOdRuTvUSt/XOG4fpmT/
7P3djPKCoTSYk3Sy9Tcsu4cix302aVA82nxamrVBGR2wJbB4FOMrSrUn2ZOdddfU
nW5gPMO9klVRqGPm23ZDZgmDC/77zxsnKblRjMmL2Z1IoO8RLOJHp2s67GTWsssZ
0dyIaXplprqcUoJ1o23u15MvsASlge5wIfaev2chGUPkeIlWrdeVxg1l4BGrFlph
X+GxqywWWx2x0yXogc/NrjGXJScyLEudswJMKZ5Iwu8nK6JjuCV40EQp0iBtYCME
XhzPrsO3IU8a1KeskwEfkgJ64SLkcG9YNRBDhQGSQ3OkJPM6gpgrxiRBuuTOCBu2
Bg3g87Cvf6pjIZ2bdth9+RACkLnG2xrddILkXyayeFofhQd2lW4u3pkrCdIlfrQx
bHg3v1BgxdQX+aH4fQWTkV50H4EDC2HLHLqPJBsW2GdLXasGhLHdfU5QokBMqbWp
sfd2aG2ll5Rlz7Iy3/d4zUGFhhkxTnWNJzUdFm9UAQ4tXSCi3HQDZrxLEF1eG9Gx
GOFAet4wquGELzm2gjujJiVsl1CMvLBrWWIuv/fFeM0pX/PYP15JVze+PpPqLciN
gvIzwGU4CcyAMRgnvEwU8KilCLAZOpKV0zg6TFfnO+n7CBua8PDCO0RBn5ug6dzm
db+3Gm3ot5YXFTXqvBVUC1CN7mAHj95Pw94l5MYGbsELi1SzAvg9fyE3Y5RYuGLJ
nP1lej3HKye/h4Xwvtuve9FrKuBPpR9kiHQfQQK4Nxo1aJs3hDS/EgQwdUITMKRk
4BHIOtSP80mHEuW/MQ2XGWthko1FwVKQ80XgCqaYfvfZvVmUcCJCDrW7gFfaqA+6
3XykTofr+F6BOWbcBMLSG3rhj/8JqwWI9Avi2tHiQFGNLnX7pKie5tUQgZtSBbmC
od+5151QCrE3jsffuEwykNp+BHaFF0hvC4JrTlmA0RLMroj0hDbBTTqVXNRh7dqG
onrY5cVn1wZzuGZdag0nS9LE9cbV9Zl292ybah6PUlh5rhQIkrQifCPqjKTPZbS1
DMdTzjsppSo38OD7CWNWVuBWTwDJBy43zcbFoZT9qORKorgegMzoi2UX4hGYjGsX
As4xvLakQ7wNOpJqo6Y0AURuGx/dBJBWa8QovJZYwIFNBNToo2xdQygnfVwfzkpo
t2cjufYyk7B2FbLDpULZd1iQOW0Ox4hFmZz6Mb4+8/eD+vC+F9RExY3YvtwoasWr
EeQ2Kg0XOY7JEXJS0p4XZ6Brzh1tL5zPSgKGN6jEn10efQ8hKAqqUjrv9nLPYfpn
YajhBH6d/veNgPLQoMVotbVEMVdtLksVu/cftDp+/zJwhyQKZmWYMJdVF090HGFb
7dx/biwizIaO8Tdw7jCGDMv7/famZmqXPrs6hPkBNSft/EcHcDWccs4Fvz9kzsuT
hyezRJagUUB5daWVn9ehswvhTXPxmzND+lTMaJIFn04ey4m3EKu7PazRHhOLcj74
esTrbQGRHIkcRVjlp/f2sFF2nbd40jJG44iTt2DEKb6M3YzDhp5F0mv4lszU8bOf
FclRPl2mtsfsav2Usx58ikl2IDm4vKbMfMS4AglCHE/VR8YSuzsfI0SXlImvSiRL
XqUMBsB5yjo3ykvtK/0pJibl6FWgpCvfPQVdUvNrqad6hARkMTnKNV1NJrKTGObN
8UzpOUw2VgrxmvDyo5L93nFudZQK81Xj6Z5yEDrQ37ZFx+IKDG8HiaQh8o1TaL2m
qMWFS2bRiN4+Irhz7B8bZw+pJEn9mzFqUVQPF+AZnOG8AAGHK1RgSJB1zi2U6n9Y
3rjdtG32PPWebpCMQwVupjClnF62UgCyVQikzyR6cd8F77xu8q64Gl6ieBsSEALw
Bp9wKgfqJtVGQH+4JM4bhxF+9chZJX7Q55vurThdVcFPfaq2PH13WAcGId3kkNgQ
GuECSILUP5ewxXUjBJEHWiP5Lu47xXytPF4dO8mp54xr9av/FZcbdnBOEI+euj2R
tC+BgGgNbrU1KcGLBbuMBaN3aO0IZroWHjtf9CKvrrf8r/eC/wekueo1tU7bUHCi
qFDVrJ81wQAnouR+ttPWQzYWukfaNkLGC38fbtvBcz32DEalyg1EWI559HTVn59N
LAY6MIG43cNe5aHqVIt0xNQgV2Skwt26vEmcuCTzzbmwtzgbNIvff/GmOFDtICiN
flib1ep1Q4llIjo8HYilhmVJEI1EUOAtMfHiPr6TIxT3zCrEOoyzMFmcokb5tVAi
jw0+Qe+WzETSVClPdix7FFrtuGUHGYx0GQxMGCbQu6X2tnoPiCfjGu1A6piKBHWr
KgK2hGVlfSzmK72Sg/EC99xKIKGUisRXeBSHtsJ+6IfagfJ3OSF0tU4xB4bS+dKq
NkOJju03aiUcj3EQ+Ae8m59rS0ji6k5UZx2cZSOnGUQZEgFgfGvQPVm99j05gC27
LbTydDvGanMUdWfNtuhY2ou7RGHj7Y6wLRYkTXofcsQQ43gViv3P+Xn8JR+zkYVj
D5KvQGem+CSke8iLM6rXQhIowNEICAkc5cVDS5nNRYlJ6KcJVNEN7h3x1gqQItc9
eVGcMNlbsvMq5kdtbaLYaplg0vvRR5sLBJCeREXitvmsYDey+NKPDwY2wSIlwZHU
V9TKqRi6V7QyCGGHQXE4xCkIF4V/fvLxXY3VCjlnAejH+EtFAMmFfeEe/sb3HYzg
EtsA7/+chxlYBOa1TpgCZMyH/LafKLBXtYQM+iATJDw0JkntCU0Lf6Ll/jNT0IwQ
iZULWnhprNxxwIehmyKd3IK+zD/SdvIQkJ+L0IyU+nII9sYL7lxwRl/r83qYfzTm
FUtM5bmEQUrvbSEqhw2a0Kzo0EcNuNlsVivm0nW9ZLwLF01NMg9T/cWhNmrQuqpC
F9P7m4xW946+x26PZv3EVvPq6tMU1yosA+6bC3mNXxDg/DCZr6mtVn+Vzt7+ETvc
pga/aAPYucvOxCFIkOgf3gYAwPeHWrrwOMDFCDJZJWh+1HoRDXk6ZSmEZ6jtYJJE
fVk1xLwYdgjiIU9pfol17O44XpNph+XaJdYqNSsRfJy73fAb9lLmeExIu/gABlLN
FqJlzo0sq6UOJGvZgJ4SgVTQDbjvgimyTc7f3S7Se2OOxwdYdGanZruLgtafOhlh
IdSkIpIkUh/9wra45h9lP8mA9bn6/XmiI+CSoRTVO/3ki06LS6SOPzGETOhjta45
EnXwXY/c+pGHkQIVQNtnOytjYKo+Us2x7qn8EOAVuDkmXLuKr1AbKmz1K4Ch3vBq
eENzh8YuZE1k0u9gzJ45OJ8zpn0t3ObrLVFzIUvndXmgEn+aovrUE6d8ymVqufUs
w20FTvbeyLNxft49EJctPyw1dJTyLVnzP9rB9DhR5zHBYszDRrCe7+qk9sXENbLn
LtE0S7wEukA2q3RQQuJCpYe6vGZ20/qixANNNONLgOydtM+VZrgSPSsQQOs4AsyE
8N+PohcFFthjOlTZLgo2SccvxfldSbtrNcQV4OCS6feckE5tJ1ff1l2tFe3L9tWt
snBpJbl0cC41zNCe2rIwSeYeonsT+JMm9GCjurBuv8kjA4zR80lHMKbuWUj4W/U8
F/IAq1NV+OxeMyGtz4QkJTX52iHKdorOQN0QMZKcJ5rbuRI+w2xi1Yckm59kWbXW
ufkjW5wPUguHBnBNqdzMpm7VNEc3rmTaYdnUm+SWcTW8D7hKduahpZmZNfhdiU82
8kRDMwiDMK0gm1V1+YB0WzizGocCDR6iIfIovgcWqewA/H6Ex9RQ28a966bnMOTy
yFckSMOBUU2OMgaTar6KTqzrueHcfZcdE8JdTR9SHTw+zSu5+LImvvlMMBa7B6GI
TZm+Fm1JVpgR1qRhVrNl3mNNQ60bDpuIhOTYWHQvKOJCGLMEtuIHtiyto8Q/Uy5x
Fdjt427XYHgXN6CJozzupSY9wX4rKnrcaEo0HTiNipzshyR/T4R48yVGAPnYtbB2
BxXbIcXkahOaQQ+0EB1oy0a42KMk9tQXRwson93ON1V4Zk/I7+UQbc2cituL9Gjq
OrA2Dy56cMQVBZpk/tfZ6arnKb06HDWoeqr8atVngRyVjKLBvyRd1189DRRy4MOY
tCr3rM5esRHbwPenwEiqvAFmQ6evSAM0IwRewMfSfj5+Go7OUSD0xhkZTqi4hfmW
8GPZVqIgSbNPnO5pCZg8BlF+IDO6IMtSEJ947ayQlKAO/0lMHAdy2XNXvcP1jLfg
AyXYZDYwqnh3zIAv6ZMY/nGKkjdPMHTKNIlF1ZRerhf3PLYv3jYC3eoAaktlrDmn
C0rLTvpXmOFbY52zLJYkWvH2Y+i0J/0amnAWp6cngByc2U087nzCznzU9npJHeem
VFcr/NAkR+JtsEchSO052duUMBrEGs/vtzUXJ38k0ejW2Wu6oIVs2yjCHNU2uN8D
XveuGV+1cWbgDL1HCoJtA9jOvuBCXK7mONwNadLoP562mrmsZScIt/sQNCF46tVv
z/RibGDiGBC+j+5hbTnDSRqJXROPszk746sIxwLUvHUA+lhFPbPxaATlw8NXQHja
SeM/YS0GuTEk7trbbcdjvovaaBIo11knNs4A/QgP+JrR9hMxe08v6dy5knajpgYa
QdiYuOCBjqucqEplGhzTyLd/mM6QtqvqYIuhPzd/tuuKki2txzJqWrzjI9o+ixpO
zB21Lp3nj/ZKLOWyn71H/HO+/1rE75FI9M1/lt3GBe2EPOBAJtwW6KQlaefj+5At
ufPH23+X+zm0Es373Q7RF5l2MsB1E/R5Xtim7SFawYF/ssUnwuncQ5/Ny/UV6+sR
ar3CdZTVwTxiGCy+UcArg7y0GKJAxHIc8PiMxWMJLwZB+2IiKy+WSIK7AfN/1Uhf
snLIrQZGsijhyDmH+AcrTQY8JbfgaQjWXrDEUAAdv9gvXwlpuHHoFQtkFXrrAjw/
JVM1kS4bw5GO0MorZHqiJyJMTnfUk4oK6A3q3G+dPtw12ZtJvVhbFawZ92q8G2Mo
Wb/8Fm/42l8nUMglb4aRiqQ3L2w8hKjYDftCCjVS0PMsmVMgsEPEfrlfiTOL1WNI
e8EKu6dDxkPWQg7MV4IgFmClHWZMz9gIB+Z9fimOfiljqzbljaJD2yXl1sZgtEul
Jy77RTAFnfpjAusJygt+cMMLcLPokcZEUj8PYQUQzf8oLyr6XBqFUXsfgYxJZLzw
lU3VnTMXDZ1JorReRAbgskJfovyJ4yztBLwIbOm+11+Rs/zN77oSTsmwPYVgJ8M1
WGOQGQCk7AiDdXF1abUqk5jSPgebjaqMS8mMCmz4QYXXqGatbI2Uu4QhNQBmvzV+
m5aZtWOZ41nvPseWw7AY5eaPrLLMx8P8tA0grQxy2Ku6HjF4mA+uM9Qmzdoh5Kxu
4j2y/TsGMxZa4u8PqujJ1nbMsK8JEZBQxhz/qzNjTXbD4zfx/EzbRMIdPH8Zvno7
6u7o0LtuwXfQxPXwfrAardfqUYEQW6tl5qgwOGCwo1Vyno7q+ggPOdoFVwE3u3Ee
jojtibdYZacYfrU7QIFXQ4IT7I8i7kPzWt/GWd7wO50rR76jZyuv0eQf38jZFWrA
RP6g9KTFTdVPuY8OG/7NQ2cKfhV2Nuxe3y2NKqkyNf7YIPrspGKO8s1Up9fGXVIZ
axNGLG5SxRqDHmLWAYLjel+ATANUI6uxdEr8eQOYcsSSRXyiswGqy0zBGymHT/AF
MgQOKAD80vyeq5l8r/RmlP2cVKzHq0VRwku6CTwCeLt40FuTTgzxynOUqM1BdJYP
AvtVvIjvjyv/DKB8gQTvXWNLq+H1zVc1J1uyE5+aGFD/ww8as9/soNiwVbuTLOw9
n+KFmhDbHVqeBBPdfaxzPCbMqsg31SBR8p1XtaM3XZxQh6X91++RvSyePTRjkx8X
U07fBW4xArBFv4LZVVjQIs+9xr/1mI9hM8dP25YuO7vRNokp0JfuNnSJum757SZu
V+cP5IwcUsxvAzxxJ/IHdAe+o5vTGRz8Z4F+g8e96m0bg+o0SfeLN4RmsNO6eHgd
5UWkiIRrwIoJe+UB2xIVpKLpt5Aujsfz4oCWI6WRdThwNVWaESC3D0sW0VeWiBFx
3cart8dDQ3UnVZ0iWdhFVbyP03vIVN/lkY5W/LvBLN6+mQ1/4q7OnZsnM0sXFmpA
L/uCwaCeCZ0thkvGD/i/6C3o3q8TrPhqTmEj3D3to5srZ5Zo02EUdjrThJZPY/cP
t8LkFMKwzYaFWFHegCsIEA+W9DqDVtKeX0xGYvYc1hPVPGtsnhsouh1ypUld2WkF
HPqRWOQhAZ5LIGqLFezlcweW8pzGT2RRCPqW671N8p8hLX6nlJKz3MramuFOYhXr
BBdPnZHhkhOG+gsFkZkvgLlRo1iGQcMs+5gcWRzBspXfncGLecnlp4czgV3f6Jub
xnmMlyGiRRiIBBdbHz1FQtTKxmezOoAMpoBzBYe9WDDMKxVKONNbhojeuleX9i5z
QYNSsykkfMESPYWWZ5ymq44PMln9vdZ6f6rh+/fPQ9Eu4b4O/cXKQiCHAUJrRjZd
PAhRa+TnX0cFrSpZMLPa2SUQ+kUNUUGQh9T8xBeWtd+8YXsiqZXUSSVmpE2qbDz/
KPPlO3mjaXdRe+2s4QisbrzvNfwHyIqPNO3+JO6WUJsP9oM/bWKyTxcDOfJpfOLK
mb2nU4/f2+Ko602uo5K1JHbAEAAMKd1tUCIK2rTg7t2GSFqf3oG2UWokwPSi4GIV
MW3uPpYKOBM7vAXuqTPT4WietiQHZ4B7VSpc50ZWCgNRn7OULHUUPUTYoplwaRrJ
PH2ysh6ETKjKn/4fkYoCxrYFXNeDY/ve57CTJ7sGfzB2MRKbCo1hPr63aSG3Mf5m
p/Qi/Hets1mBDE2K71AVjToM1fk21ViwaBUEHAzzIxG2htZiE5UgLpm51myk2lAz
kt7Mi3zfh80nKpPLeabFVjC2u0vyCdbah4NpE+oYqnCpIa19bTJOUh088kA4X1yA
SRR9gIIG3Uhx10cxuAORHBEMxwgtnAfcfKr82LNpybTJwF4X96XYMi5oX/2dg3xE
po+4h8KSZvqOPYYPfwFVNI3exalmjD6/vvK+6djjXqamDaW2pilvTNma4QG+qSgG
BqxLgQ5WB4NaRG26iK4MgiPWSSpTYEyJl1Ng5NdebpmHVdI9cBiwSRGgupETD9e5
ZBmykgZfb2VmcRluYV+F/QP5joocrucUPIor2Q+eUjmcYEwWsc1CQCoG9b4G5QDK
VWqB6Z+O7GCdyk6vjYFzQ49eHambikSpvs9diViIRTsypK+gNerOfvc/sfU8vyrj
SdshobOUddZFPomCeLK312ju9XIAVBudD7Y8GxoTaQ152BXuK1CHasYXIUkXrFKK
8P9Q/JSLar7KzbXCMs8zckWNJ/KAjZD//O8fUH5UTNmPa1KSJ27uRjT1TvNaKHGH
33lWRVrg6BABXlsM98j0ZwyKknjKt0C/AQpuBMN8H+MCZnaCzOovOSxyN8BSlhW+
0NWgKCUF1mYt6Bd64y9+5z4S9MNuJ1p2hkOH32XgLaphjgHKuu/igNpbL780ljlu
KVykQOzr+iFF/PDw/Qcn00quPrZxKExuTr+md1vobToXACm0udGu+sRHAvXlm3Lu
mtGvevseH37dL70ki0TsjrtTjyWuz29WrORk6Dqi8os3UZJ8C+W7lUm0zBOOkcGE
04iE+sUKcfUvhxit3j7Z20yu7SNAymmD0PAdyYW8baFF7vlXHL7VU2z+6CtUYZdr
+8ruQbSRST0SRz3amaf75L4RqDxFSX6TimMrJJ2v5pTZvLNLmgJUGX9wU4XWHm1q
L6tGZW0xFNGQc/UWPO9VfKNKoCeVAh9ZJZDdABoYA1tu1sK5LQiPTgZHdUVmIOZp
mHeHHkL/oJWrFZVX/SW9dx2HQmz7344KJbVgt6hrd0Yno+/waPwVEr+D5mo5QVqE
utI2TE1Yjnf2zsAr7oNDH4rCq0XIx0iLVcnCdwoqCABSwIKIi1VN/3j1D4A1O6gC
z4bGeSgW0v4r5emikQSUWV5PgH3vzoGEvnyXtx7WLyBRysQtJMJk/rQ9uQ3BWGbK
3b4C+iNY+QomhEA1vkCX8b3Fyd9M+/7ak5L06g2TmeMTRcAhDd/9ckxr2FVDbNHF
AdSnr/nzJF1KB2fCCYY3B7N809+Yu35HjOBhQauwhqr0GZDMVfyWcu27Sbj3lP4d
y8H4Jv4TanRGPwezG0H+OTGo3dZBQ2NRDhLWhxVCVWrcGouQd391gLf4B005AFkM
05yizPFZvK4dD+iD/+lNA7xSjVwFVgW8J/MWRzI0AGQsTA9X9H9OfVqk7sLlqruV
E5uaLcTlX8mBNlwFABr9aHXB8tkV/qjMBhmiDzjLLLoIoMBfifvM/QYYULvq0Xc2
fFppm+QR+1433KWWAK4mPsWkrbLfxgq2MY7Q4kcPAnd3HMB0tP9gwkZEdh4ogHzM
pImAv/d6vYs5nnc5mf8/42dYxbXAltaMl0LTLE2O8s8L+d8/1k0nbFzP1kRFhvQF
LqvX5esetxUQ99lzTDoqL2e3aZJSwugGPl8YT64uB+UxJOTKFnFbV9nuvsNNzHzL
dt7+Q8fAI1dd/F0LNOYJ8ySQjkNmhpD7kiDoWaE6jCg4pfGyU8F3LNziyFAubS6W
NOhU6AreVBffA/4yjCzhkCGCbVBUHQeEcJ3fdpdZA25SvzCLJByKjdhQSnHdFMw6
WLn4YjV+5wE5f0TGcAZB+oNfwSVcb5Lp5koE92+ED+9WKhNGfMzkI4eC6dc0Ld4Q
nn0zSntodyVaJ2izKR/5g7wum96kDOj2/Kz1+V2+OJ9G61mwHhKXTPqpD9I9zvXo
WzHNZsjWsI6ZISfXnwcbr7OyD5zp6+rWMsn3rKYneXt+DWyA9JTad3Vxwg0AeZPm
y0vpTaZWummy3+O4unWABVbvObuoguIYTQ2Sq7Ce3tXxcznIJsGkxyq6sc9pYH+T
hzojZGBHW14grLtlR5pUu4jpZpFcEvcEE7BImi5vqPiHDI0ZHVItb9waGEXIDh7A
mreENUP041tJkn1S0rdwDiOxrPUBIO9wIx63AuiMqw8hhlH5kxsVamje8Mxcao1D
cwmu/P2dkj5Oz4vD6f9GhAgCn2hqisSl7lQ08Uhb2u+N6vrE4qQ5mR79IMIhiC24
5hdApfi+4Q7SNo1BvpSDPEQEp479x1ujYnnCEQ3t1H9IusqqgLvpxj1b4Y8aQKN4
ydavtO/U0qztHv7A9rrqfrnI0BdFmhGKJ+gGdwdXxsAIfqUWw2iHriAHoT5N1vUr
lKjR/oc+k+K4VHTZR3QauZOcaJ8uIDaoNc5LNyLMDYbkB9tQ1Ca64vyRxrrJE8Ln
PIepd0DN7hI+I73KuvFk8AQI79U1kZQ7eJjoutMBIEw+NPf8L0wM07aYc2fwOlXc
Jpnm3imp4QZKZ0RwVt/RnUZDXbMqj16NsOUtoYdmcPBhuuhcUiBF0zbmRthomcUn
1diYWbsmIHWRGDgeauVblvfZsKqJ7IC4czzsZxOd7Avpn0lTGQ0pDb1WfwkTyZjP
XjE18urZ2y+RZesRIdV8ndfp8ogIVQu172+F5U2e6koQXPNihyuRbSBwPJ5z1XXJ
acUHCj24wfZPZEeN3y1LroJYEUx7u04ztCcLoRxZ2EFlaOu0no/+Of2q5VWLHibs
uoW7RWFh2wRIMO1QCaIYTKNZQREkRYAZGZu8XB8+SVEKGjpCLoQ6+fbDeyyZRwkr
0g6GIQ6Md4f8qcZIK7rLGE1JzufQb0WG/equHtDwaC//xep6qBKoGCPFV5nMGHDT
RjmlDVpz2UsC6pXjyTXbX3YsnTMrj9i1XLwiDzPLNRKFTn1LDrEBAlM1+bHa0iJj
rk2hGDH+gUEmVXMIk/ICAmJnSLPA071wE9YsE6riKbYA12g2oOKZv2Fiy89yk+KE
whT+5qdgJ8xkLbeTeLgvNNe97xBDvPswNySDMlM1CNtBDPtkz3JPp3qCzyJ/+PGi
97bwrw6ElbWejQYcNsczw+9Vtf64jx2zEw1SG1pDbl99f6bSvce6Eud6QUps4SCd
os7p+W2tGZTsQdgxPqH6pSki6RZ+qh8OHPWqrHrEckN4W9cMZ/elkC9Kro+XnIrq
11FlM7n8cO/xFoxI6U1KSFzpsaANVe8JWtmbJxPTE6SHiXuUjtI4RQQ+n0NKCygO
+xtrhFgfsdK6+UAc7SAG+eWb9gIYUbhj3bJSOyABf8XQ1+QIYdEw/DD5UJ+9KRDM
TKHngcnriANBJ3ZO0kEeLlHAD0ZbomEhc9ShxjvXyynZYQSPEwazL7MkMzxuzMGK
rmKzjxOs6gDo404oCFaV0FU1W93Y23vPa1hA+z3/+Te7gvmsiWDfIlilKB5lK4b1
sLn3fRZahvvjpmBusvkFInm+Y8H3afmIihC/fqoAFXbKauj0yPyNOP8GrHmWk/B3
pUY9BmuF+6RZymvVJvwWFhWlcfc1J0+N1KZuO30+qDonLEATpG1HHxjM9uXqpPug
MsOgNbKMY7YwzPQAjUZTgXP/1Oj31h6K48Xb4eueTjtFoGbBNFLU1xlJ6/hZBxfI
LVYFjOxlKmni+SEJmRyf8SehJfJMsSMUrtbniOQ4+HQDTj+YUNPMh8kpSjGjLk/3
Xx41PKmdoRb75EcnBdejx3rLgiYTVnmfkRXP6SV4jwAksSsCFd7DryabML9s1BAv
JHQCHPl3eeJX/aj1vu3JR8nmmv0McMqT4lSx+XWK+7fGyXcgHmD218oyoXRC5uLP
9pbMDp8jEOH0GbmfmRbGnCe6b8/mY1LX+62K6KldzJm3w0XV6j1B+TGd8JVJUfa9
ozrf0skizDZ3bQKUhkroYJN8/VTEl8Ey/2jj9pGBvNs/29RAOy/QnZZYnijfK9Eq
z2yXb7pbMiZhfneRe37q7Toy+DOAwv3VrEbV5eLexrrHBZ0gDTGaVWPp3Hn0B2NR
IcrBvETgGKukS0sfcgYUf/mXeK75mh5nTvoy39Eaksm8WMDhHxXRDL+RF4nCvYjJ
MSG7I+UNnLa/fm9NZ+wWvAB8KcLYlSwlb6Qy2mJ9mPOcSihyrXnR/wrEpQ4SOAwD
KkXYW22nhZrdWw85otI6q6iP50UM9BU8xvh7XDZEFPJdVYw5iDelGRYDN+5bV43I
NxLyHgyRqfbFhncP4hpZThj4/i/5tzX8NzXSuyNkO+ePtwa+HvUKjjCpRG3OfpR6
p4ZfXp5WzYsdfJ4v8whaRlmddSeC4jOdA+8ih41JYiANZ5QS9kDS0WrFEt27ehGN
BKZNFzQ4eRJAnvB4R5iAs1ebdJ4I+8bTsmbLgUgDXA/vbEeRIaxbm8l6bDKfKkTA
wg6+1JuWa+yXeeMkqWvpOxxPj0u7xyUTMcJOoQBG+X+Lcaklee811LSrB3C+5xVQ
MaDkatNxUQv7Vl6M08dPioaFy84lqfNKxzOhs6qXL0TUQmJsC48nmPpY/4e3B4XG
4sTs920TX/0afA9IZveinXjYuyw4x7UDDLROjd3LAZf6K5MxusScF89fVlw6XLHH
WJxkyD77ryRpokom5f1UxhvooB/sFhCl+1yGyZNCUMbScFsbX+QZoNwYDcdEIU+c
qgHLjSamGvS8OgSXNaZ47DMioniajXKqskfi1IlvcE1hYtEtCjenVRit+lkD+fHA
Y6YAvU8ESe/S8H5W/PfO1ZuvhxoRBiBDVdmgN6EJb+03gSYdodQYbWLuY6uXjLJl
2qu/te+4bLOEOEvhiYjat2Ur/+I7t1rq7XkY433Lvp431LN4NVGM4d/pQrVZm2np
ZfUa2js90V749tfiYaIxvySrlrULgoJowjc8WAkNyRypt7qACI5zwpFE/yAdSChe
mw6TLFJs1kuEYKW5icCNOik/gWsxu4Y7GY1Z26Y+BfC+10wGEBv4ghNq2y+arvqI
ufe8031oYtqnp7U0fRM7cuAv4bD1PH9MwGTkbjcsM5uTX/pGW4FKicChvjyf55qb
vCade+WGsGmXVzZU3VAJnFz3k/b5+oDU6KhWHAxjwdZW46WWhXwc1zH2lI6BkiqN
cuGxhne60uaQoHOEmunh7TwWaMA1QQ8Wo2DaSBhYLmhRwu5ZM6zitWsVoA81vH48
0wEe230DXkpHhYIsgO8ZkU6ch7bwz0AiucNQP76NM7it4oVFhoggYwkdp6Lmrop9
2EXEmdSCaIKiwUhUs0SSaM9AxEpfJkuZGLjuXpqzP+HC0zjp5mHIDHxAapssE95L
u3YYIPAoJpWmr3n2SojrPgGpq+Ln4wRAb2Q0xKBK+YNcToePnEV6QsPhJIHSiqmu
Y62J0+oNyd5ybtQpYYe+Hm+UHt4G6dO6UvrWdDL50maTAXgM17HtPhpnLNVbsp+P
z9uXaQPcrHmLAm115kHSCk2hqQ+atxgIsQuU2uspORxVu3MJ/uRDCR8LSiItYk6D
6RL7wOhWnMoHaYvAb6+Xq5N1uZ1A25v911k/GzDDRg+ZIWr4tS1sAlG9F3v/sbm5
EhzQM0hrpXLKik4oeGinvGXczWrS2htlgXxHvb8ePqVqIHJSBTmqikjD1r1mAZKa
2r2J3HcI6TmWulQeeNyIISu0Cy9uFOJdtcbD5yCVB2KL/O9iSvqqc0/50iLkmvXE
G0vH4SyuBDK5OIlwslZ/5FNgEcL4Xxm//bt366TqvbCBd1D9eSvLqRNA7NX3vNtT
YLpCZ9u3+vh596Hl0ed8Y1y3toI1yLK2aybcMPCI5S1zNKWg8Ar9LxH739W0VtQb
xcnmP+Co3Eu5Tt7hm7v28brf4dGMUdSER7kDwVBqmZ67HQBhlJ/2m2NjVHPl3WUE
jhZITx+Emf4s1vfWre4QiWypSpwJ/2fDWhID4m1wsaQT1ygjTa7v4cuSn9g/xGUb
UPD6ddOw8M2QlDzETXgmy6x2LqjTW99hOZXg2vbQakaZny705p2p4sFBvSdzVQZK
NY5ndoX11Cre2tYW3GH5Zci+ry1nbaR8q4jkAfuU6PeGbgX4SC7g4MF+0HAc/5DE
BqrazcjyygnqcOycrd4ZEEJKNPiNVXO3iYGpJG7/i2jm+K21dSRkXBttwHka6EDK
x2n0LZsJ2kdDmvkHW2VXJbtFvNqY1VM4kdiNTfbWEHcc2Xr0fVDVRMQ19FEeIDrO
jxrClhIfLBMlxWsCA0+Co37Wq9MrbzcRlE9YE/v6zMPWy36g/YIuhpKVKWDFa0iY
g29Btt7ARDdXwCYplP+TBK5VJ21kpafQ3aiE6b+XNWSFZra7Kfo4Z/qFbe6Zx9bX
otyyiPOi8Go3PHSdExIU3ctlJN4W++R0Jc3bwb166/jwYeZMxGRL/z/OO5iBEjuM
4mZ3/klzKGM4zsV5kK58tYS0KEa/prjleZxz6stJC3xynGpSIQ/kURV0LG4CJ4zq
oW30c6vGCqyyUToNEnNAxO1Lg8OiI+aHdm7VR0yITecJ8UpfFSWMR0n4LDVQHSG5
gPp05fwvWy6ZxPp47SHlAWEfvmExs4ZLBitlhpC2r76FWg2m5vSl4UD0A3ukOls6
`protect END_PROTECTED