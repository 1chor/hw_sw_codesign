-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
T882tBYIMtvMSydiqVOMyOlJMix6PlI77kaDESAToo6pbz9ht+zNGy/E/s5zARnQ22mRGaFwFNiR
TsTR3bLzJQli8fnM7eHXsWkcK8VD32wEmV5r+c6aS0DFhwtVOLVF2y4z2ZMwsFH7atohxD2bY+Lz
FBur/zvgbtGHoFyrTNY0zbMWLSUDrf4U+nu6K4dzPSNXX//qO7vxd5RSsrZygb4tenD/2MteFZRH
jx+niHb5aMJUtXmyimZatExTccFj2+nYd9clgJoESzkT2HafEjf/06rLnmA4hoGLjrtSsF0kYxna
dcfwnXhnoH6XKJ4wmqaOC7SeaB6ru5vBNrCfyQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12544)
`protect data_block
ELgG/IQ3Lvi2d2XCeEt0LHRyHmqPHdBtW6nccpih0wC7FchPp1lkmM56/r4FMvqk/1EI8wZziwOC
FJ1JYbNg+2lWzZsj5q7CvVAcATUG6OG64DNGK793ZCd9eKPcVB3yJVMndVobtFLFG4cZC98cXU33
xoFmjDagQwbnR53q9fmfTaLQPzUkPgt4nwbwi+cvwpNArZ1oKeYHEfOqdlPy/4OUFiKt5hZ8FAKN
ucpZlRzkXnd+HQwIT5cGUE0bY7cSlAFbsDEAL/YlJ+Q29hf5F5o+LKleQU9f0i9kkJtq3GCxKtAK
fAGyoHROvaO5xlEpynvgC/pm9ibb3pK7NxydF3Gdu+wuGN7Rj1I/ELC8yKp+/f5q9UPX6+/FfFrE
ulB24C4DEuRYPkxoUTig8E2BL5VJcUV1HWyKKjQUjMhgRapr5mPEVUlZ2eRybTOu9JiKMCa+C62n
nzR5nzachluIbxtcY7Ttrqn01CqkcxL/nygQVnfn6EHLoEsjcYvhFcWWAqVWYloiFRKsIm8EdFYF
jQi3d3HN+3vQGFZ2VBnnYxPXLg3Wdb8T2d8v4bdrKo3F2GlHQCnYkvPCxxmJufrtBdXVQ3pQloaI
qlIUMd3IwhjIMWIv/Li5CBDG3+NWXnY6iAT1VdQOdvIaSz0MXuGlcPZxUFcZhI+TNhEcXNGgnn5L
lYTHEtJs2G+9ZFn25HzYs30sU8KLScl+GPIV/XckEQHp2PmXbCO1x3rz9JwgvPJZuGLaKtMVsQFD
rY8vov9q2CZ6ZPrb6QqtGvaZtxXMvVSDTmHL8BWsQRCJtoBs+byP3Oxg5Yzu4u1YeAzuYHUvBjUr
6rVkjGzqc1jfWTQ1Ea6rRY0WMGwSSD56oZhrmMFjy7YfIcnFwYNmxDLEEqO9CMsT9yUn54FGt5t9
anSFxaJOvTnYju9kNUVWcKBwLtNsxW4b4AdnKsTsaQDctCywfnP+4yzC2uWQz0nBZNkIzDdAVkqT
Q0LsmjEz4uutEPrzs3w/98o01lfUU8w5CZ/pB09K8uYS0Sn/W50Jx6Ew3GsAzNmiUpw2F9a4g6UC
wV7fToOOv8eJgMLSlPZ8jNxrTi6jqeAdlMawT96ozfKOn6RGGR1Wxa2UUCLq1m09CoSDG148DpW6
NS7co7684httFzQNO9BRdlClu8QzUC0604jhk1PzzRm9rmtFKT+UTnQyFXvA5Bn/rCjyVFhli0Rz
G5Uc125WBxQgY05aE3ulE3NoiKWRKYn7WPwRuSCMRvmwHEhcHLrV6icefT4wlthHdtU4IQ72EmYC
AM2Q5d7pHBUjdNXmuWk6DtMTBHgMBHzsgIU2iz0k7hCWiYeMp2nzXqniAdPz42IHSUiGpWZ4HFY4
a1OeSejP37DKZIESA8S2d2S0o1NiECzUKzJLBiKquVQ1hlrHXDhU4WhDEK7gaJ9y9hzfFY4MHbKX
D1u/0Kzp+qpFbu6gvZelWeP8w46p9mInFgxMpgX8N29+ozmeuZrzGknMYxYrhpgOlWlQHPk7rMK8
kwcA03f5MV+KSU4MSllMv9TPQSNliZq+WCPtqKhT6STQBY9OIWhb4KfU9oeFQLJ5bVMuHoSRwSMr
IU9moDJu9cnPEpy/rvk1SPfeapa2Ctkjg3IrP92+hi4lVoW8jHfYqMY9mCUmCfXhawpdU6V3zTIi
VJP6KmM5+JCXvh8VXsdisi2Jhx/3ci9f9GaK2FELFJTAdJhP6S7WOgK23sunyyStvnDK4MyjUErT
JXo8a5hl1a+Z5dwSRAhDclZMbxkqInsFhKAuxAfkHu+ZZ4lgLJvtoluuP0OrDiem0ZoGgLN3pEO2
UCFLSfrrVPBW1a8fjLVo8xdUQqpThXPfiIg5f9EOKHL/vGV95rX/k7vA8u84QzL5aMbJH7px95p2
XgStIxBG39GrBJRT/C9+/bmCNo8952iBrM5tRZ5e+pvO0aBh4Zv76IdUtpQLjpS0Eh/g8NzBeKhz
wDbg/CO+W2F7B0b52sqoKkaiOe0W0L8y1Q7vZURUngxQxKSyIQkbV4puvu0ODkOWRoxYIAR1OTCp
Pm/i01XuO8tXH36VR3SwFD4KmVUD4bcoN54ATXIz3iweuzSEIG8E8lcgzt7ka6RZg9fyKG77ejFC
kEv7foG+W/8Ij2pehQpjDe2uQUHxM8EL/8uWyCaybhh0F67Rhf6rPHOANxPy7KadWO1qNx1W/0Tx
R+GSszjnTBvIEiwuDIssgy67mXqw+4/yZ26tqFOtDW48xvtKD+CT6QLr2y6vV9R/4KAPnyiSXv1g
OLnaKUqqw7tb9qnNdTRqHckHZMEkGdFf770B8x5vuHR46HlcbF3D8CYbiU86FTDSkTQMegysj1C0
7O5w7uDKilB4Vv0bTdmu6g2N/8cqUy4OE6HR6jeVYQMrrUA+pBeZDagvZIerxoCSlzjZD4cuEFFa
pLOg9PKw3myly4CLbOswK0LnEDR0gMGH+KCmS8YJUUL7XP1GTX2tJMcIKRmX0+emINsAE7vGG1LI
xC2uPMyV4vUQWqbshoDDyP8zewGtVtCu8MvFoeQWQJyKpMrV3T9cfGd5jFFUOsBeJuOI9NgG1jmQ
azkrtEVqQ7Prb6GHHgQCxzZJZan57QXG6uclRMxsRSSZdGdZR8b0PMpDxNP1wnDYIElmNHdyP9pf
7XxrvCnm2P8rl0gu9W/K1BmyZFdjKJtgno5OfNmP9/3rgwcpx4baZuUXylPro0PV9Ovq1gZfWt44
MGp4FIiVafdif5Opn/U1JcSHh0F3ood3LrFFjIFPbaUyNEozPgWathZbMIws7ZaEQ2q77Ppialei
IETKGFqTIKDiXYIiyQZBsCWXd7u6XwLDbJ6VlpNbwh84TU33zIhGpY/QA5xLIEj/1dEOHf82Vsu5
CcIMBhCGq6k+k/IuL7N/G1MdIJHOTqHN/8ln4S8QNWiGJD6/xjWQ5v8ZwPXnA+PMKi/fi/O2HBYL
pt9TvBCIIhjjZmoaTZVyUDrohSlGK/ChoYemgW9QOg8LDVwrGd7xnrN5PzCrCux9PqVQeUcphUSS
JAwvqdHN2B1Q+05IBRlEgpB23PO3IuZeYVrBwUXZNY3QIeBUB5v95sfBlmnMrj5JmQYgwucGoRl/
MsPaHUd/GegIamAymghNlaU1JDFYU1LsBKrE5fyB3/ru5XxmZrbjcSsEbkjH3+fJENaoItQfz57k
n2ztGqhNyT2oLcxIlbaSIdzLJyOrl8TZeK70aGyZYcOgNKoi+d6ggNkyp53ymMNdTA3EUU/rS+0/
BOFl0r4KGLJcIFhkx28vMVDxOxbMnuyfdVVK1DwWFWx4CZ6hntqbR1rJcFp0zZZnj3s40lrXEC1j
Xn3TD9by+f5lgyHXcdAE5wR5il/LCTyITvtUzgBGM2cODi23/xdxXtXQSIfZTw21d5cH3M/zub4F
WGUpPGAXU+Pozbok57rzCpxc6E/z4izJNcJVFYe5aI3sPQuzUAP3rYaouU3p06CyYDQEaw8vK/Bq
AtG6gFINfi+1m5MXQFVEFUKe6e0FEujlYI/xzGCWyKWTZGp0Tk/eiCk4R9Qm+ySp6Cf+eB7Y0IKW
BHjAxQNe1tqHQ8eX56Q1zG02DWhBafTv3Alr5U+yrW9TcRp5zN3ZVH38VyJATXDjRw+/hd1vVRgR
WuJdbgRJiYUXaT/PE6TR5jKs+rF/NNXRyJSL0WYBvTeUZTBu2rGOgLHxDgvgJL8J2WQnXBpexS3M
uUOpEtJ/T7d0I9vNBWlsqdDcdy0WG0df8ZTmMTwTL4Z0VCXfZEqI0/kcn76fINfOl9GBTQ39u9w3
AnGHKNfMtQx1uZxLZLwUkuijTXxSRw60k3pAp9Ms/8WfrxV6GjNPHNIXnFb60fvB+C5l4jjvIYQv
d+EgsnvF/qsow1gbZcjkYh0c0y5IoOmLPJUKCpeWr1LKZPA9Nw563TmDea9lUSR1ytyWWq3+Wyod
7GfqyzEtaCR5rC8Rp0OpBbVoBZEQ1dcrhnlnE2yvdsveQrlj6p+NC922hy15XHYh6gr/PUJ0Q+gM
I+YoPXNt0zGxhdVGCBBCv5G1yJXbBoX6N5yv5dc47y91FRy63yPkxtWjl4RSjfA+5ae/nX+T1hHL
bR9DojXJtG/rKYl0VUHSiTZ9N2Iy7/qFPJdgHkGO4BpMktHQoOHDhB5vZWxjCMuw9efx34uHJK2L
GP6YIdcXvipmd5HcX0iPmGBeZXhyEcBy5dtqLZRiKfmyfloQtQDbAeI5YRMaxryw6Z0sIYzDY1pD
8BHKPjT+FN/08D52lPg/dYcpcGyXC81a2mAAgE2BOmW6KB/fE0HkMPCT8/Ctc3E0ix676f0ei28U
e/SLtBa7B6zypQt3lmY2+r4wDwL9CCYngqiIhjB9gRREvyW6CltB5aQGAXKgx/3iKYvlyysTDbm6
Qn4aoWMILp2G6PwX37cnaDNxNIbOUY5DOSVdSIDEIhYh1SNv5nT2I6EU3SAmJfCbOPGpak/AlMjf
7xNDsLhpa2ord9IHyM4QF2s75hCPbJLeCJdmiF4+vEzJ/7bdHLV61AwpKgu57QT1Td8hyZqhFTTO
+eogmEHbb4FCTDhx98NVuzaJWNNyRJ1IoEJyicZRO3SSzlEWvDAfgFYbMbV/qNbVhWUqQCCbd4Lo
iKR3lWDjk2PvE5opRLtTRXgXGM4RLA1Ukv4PrMAdbuf5NF9diiTpE20dpICUbKrz3ta44g+t+2EP
iFgeR346I3lkHhKw6ghtVm2qNn7dUVl5yvJmaBfbLF8abJfI/nPP+UR3YkcKVWQ6rGhfDWuDC04I
14QI74PKRNkLmbNLZN7356DrIVPVAsYeqsExm0h2KtX2Hdw7h+QKUYg6mwGGTaBmb3OjZOJKkAwQ
StXYLU+WF1qHbUuHbTqr+tzsW2LVifST3tYAzq6ke7/9rYfzX+wMS0MuH+XQTNMStdTWdDQswcvl
0W2UopvOEi+jj21+WOXMhXDccsKJvqwiqjG/UuIp/euFfhXMszWs5lkGJIY+8kY1duCnv0lL4hp6
Xo073UBLOvA3P96I9doLSxpUYHo2TVsIkvsraQGLn83sZESkUpYVQ38ePH3CQNxsVz942KTn9Xti
g8keJjKTrONdru3hyX+cBsvvAtpnDdaO7awQl113VOwPnBWiUqp6lKpp3wP7zShOV/LzPlpDKabe
qI1qrHCg07DaPMGxeKjefduSDA1Yu7yN+mbP+kA45kBiZ5A55qv3OMcdudqiD/2bxS95LsnYvpUX
9ba5mNUatmjHsjAFd0YQUBUqb+Nkhl6f+2T12LjIVN6a52U7uTHo2soWmhks9xNfScT+WZqsRVIe
DY65qlfg0Ig15RdjARJbUO3c/1CJakfY8IaLvgTaX8XuXUfTuOtQT989Kq9/MMftmuTdQc3X/5lA
7rDGAIpt+WTCAGlNxMcfpw/xIXWLV3alhYfHY+bx3FUtaqhgQ75qz4w1c71itb92BgBrkF6pa2lC
8uWvH2AqGAxuu4wOAmTT7duoiDn2PFvp6Idv/OXZzlPDwswnNjPnw2e+K2daFvSbGo4lys96OpuV
UUZmL7+dfr2LStzsT8BWrIbiZ+60f4O9UMZTld1WY/SuGcOaNvIqxsc/EkMsuNGO3UgH+Aggr4Ik
fuw747IKmaHHpx9BF9lA3r0lLRRLYwermGV1D0a4T99vmm2zyeTEFeVmwm+Fe2RziHubfNNv7vpl
tR/oHZkpoL/njkdfMJ3PptNFF8BDfu8uInjhko67LckGTyJSZot/MHIIbT2BGKymvCfoqRSS0Qw7
1usxI1zHaMB8Wt3sLFwQ3hXj12yI6U7jtiA/MAwrpK9hb9y5uM+COE3pCA8u0C60TCFK9gMxWEk5
lnGxDeM0OYe0iPSGHuduFREH0JWBmCU9SLb/CfTHDWJm/KJ2JFcYLGcwKD89Apt8s4zTE0BGUDpE
p1gV1GztBNRyBigYVKwEW5tM17oSLcpgWk2fHZROe3ryzeaMMNqEtLKABaleojD4jWI2KhFO5toD
lM4JgNs5hq1/56afE2Pv7s/Mn7DhOVTSWudSENRT7D35+UHtpPpbsUfYoW40xXVWUjje0h+tf+Ng
i7zA4GQzhnmyG+IcgZ3t4LS5Csgibd3b0tfXNO2F238ZLQKaQkET2fhQkfVPJRMuPRCIHJkHh+jE
3Xz4ibGMLlze/zmIhNhid9gn0H+9nct/+DfZZ6neCX5nr70SOP3UEAgOPHR0vud/2ihUf+a28Izq
0BWhhCI5/yspmLFXXN2GeR4L2z9dsTd9+GJTZ0QBylrzkbU78KQOzSPj87bgwhsljdlLLQIgynb7
tYbWzCtc46yjwg1a6uPczLPE1FiYXKpciELz4wOFMv6j+9CtU7Gb2aLZPaSMWs5wjfGbupPqwYUa
qaAwgVPq6ZiouKpZxl1n7qZmIRM2xH07WFVqJ7gXDbB6gHnewL+l45+ZvWHU8sfK7II+hDmuy/pI
k35DVaxbwnBB33KLTzqSOJ9cK5KiZ0CbahUtzC4VFj9FOXFXmA9WFIY73BDEc69/32WmrE2CJ+Lw
aBpgvsbGlKk3oTnRzISmHk4xVupxhmOmSss7ulzow/hJeDaRahLMcghEW+dpTL1J8ryNanUT5d9v
4xn/eg3PI45ufdpB2ADqL1aBUHi+KKzb/HyLGW/5XNNH3J05j7w3CQ7nL+jOu+ADXEdlT2T29Y4B
M0/Bms9cPuZ3F/yvBoPokSCMhZD1cO7H25B4/9PuvtHdQT7AfjQU2s5GuihR3tORtHmRrnkakyV7
/re7/loGRhD7hfjCxO7plUM4c1USa64RTys4KYCcOktH0l20QLGWQSF0YDAeW7FrETcdDVKiUope
fSOr/qe0LMIjLYeZWD4IVyLsHXs5Qm+AuC5S99a6U2G2yjY5ryYDLJD8UnR60uQ9umoUeLA3sBjM
CBpS8Ut2Pp1SSJo/+Cs15dvZB1RX8w9A5BjhmKU5NJ/f9hrZ/zCLBaRukiZSaCSn1d/5OSoqLm+H
jIBc5cXXljGTcJ7krhsKWp27plOw8UYZgr9LNIu9ag1CHtuC5mM2muWXoCA65bfMwd30rOBS1sct
EAip/eigezGST5foyG12DRp8B4jOEB8aehdh3tjZQFadEi6SaNN9W4OKekZcIOtKfl3RjEuscCAf
fp8H0cgoyK6diIxSifa8QyrAWa+fFUhU6qvs+aSgj4f0J+bvcI0bzRBKW2uUWQrCPh3jpMyLF9/V
l7jLw17zaCAup72nln0wYLBM8gpO8U1QsFXnwu2yeeVlSt00/EY/g7/vuLAFrIbwIQ9oca+Wj2+m
2us/kRdRZTt6SoC3lFquE1xAQ/hrygkmfOb/MpGesIi+kR5/ShBYOyGLYfnpR2VvY564P1K7gzeR
c+kPhVh+KyogtwGm6KGfOvW8NQP6pUnU3xC8hF1ZI+B835lfQ3n4KTD2ZoumIT9UFVIFK73dCFwa
Fca11z3fk1c/pZmo5hHpwVgCh97HcZL2daqQXVFTjzfCTXVF3MEtcN0n1R+xG8GRvS5jr4coZtrV
gEkvSVjycuG8ucTBy1FVGBUMDuHIoRjyEi92991cXsuYjcfYA4ssYGseRGk/9stgAhY9nKYR744F
mjlyFvYNhecjqj8IZOe91qYTXtUfidtPtgAAmd8pN6hriJxQc3ObMnV8Y5PNkTXAKpaRyZo8gcWj
2ccE0XlIGLcRAZTbpxchYbuy65oYwBcnQaQXgbvVqaLPLMBdCgJSDSO5SJRlNnfIBNak8jYMyjKv
ORqJRIM9KbEn2MwZotMwpk637A0BBCLzcZJ3k8Ri8UdQd03PClr4xcNW04EIylkiuiIHZQBDMMA7
pYUumvoQ+Vs5MkEn2+4N0zFbHcZ570TntnRo8Vpj3m7rqalYa+PunTTiM3fOQZQj8kY7J7gcYKkN
2K9zl5JYt+iR4YZApDunUAEUlRQVJOXM7uIA0ztXQFNIjc5wPud1DEQcfPs9oEqEJPl+lKSBLwwP
76GtVRWqQzd0J1EPPQb7bk38CXE0P6pwjC44dXFXMUcU36CIPytAUkuu/sE812Rp5ako4k/sX/jN
k+vAURdUOpRItcxzOC8Ua0Lpql5TowsBzUBuhIq5NKx/ZFUPo0lArfDNLzcCUInt36vr4gaXIxWz
tFcn13aCnRLgwietj8VuI6TZq+67SmdDUCrgnjcfZbcGNcAlsl5eWf46aOfxP9zqBmlAmpSr2fXf
+ymhQwa9ewRWkI/8gInlOXGx6nrHZ8V3oM41WsH5iON5ai6hG568+hRVHpo/iS2bmB0bLtpSBg2D
+3560KAiV18nZhIWEnrO7oa8Fm5ps2K6AlJ0B9e1IqwYbIQXU2Q+AcgwnI7pVbAVI0f9BejB7w6o
45NJld1quTN7DaKsZDJc1yc3Jl9TksdesRaWhseYh2QxULYfnynXltto26kpmtbZr9O/E+9FKMk+
F15AHcTfvNYmeZj+0lSVYkcbUqRILwlk4scwMrdQyt1WYIrqSlLw1QbddhkZvwKk0jC2JHxWNjks
iUa4fQV8GSqALUW63ezlfvDiI1E+ODHx4YDoXVpuxEAzf9TSjYZP0sp0ICzxkcQalNZP+CGJmjPc
xvOPGuBsE9zSYO/NnsSal+xssfO1TG2I694vIeFkj7v1jz8g7wjRxu8KlXDq2vfD6kxm/uMpIqLD
NMJJ0CqeZIgTt6fvZ5FCKvuE/WCoYcdeDUaOjlzITB3882T+cD9Y0KLI0g3CJX07W0fyxPAZg8RH
BBXINtiUY2+yUbO2KOVFIbSKmLi0ansHkjY6jveDsx/AHExmUyfQwNnyCNclOF+eaRe5t2ykntot
otzBV/V4kZaP9KzaaEhnhL0RbC6EEtv34xLbEnou/QJZ9byN/kz7LihrdqWq8CcRA5K++VeuOUAy
JfZ+5Ph91O/rQvFc/7Z1p3DwF2MfULIfdoTeP1GZkjTQ/IwdizK3yGyCxWc22LWC/nPjzdB/zY0m
GBTNT3rQNHWmaumHnrD8jg6vtyuvlUeJ0TiqISDOx4hyZ7CPW9zCwEHEAJW7BgROXuFCPLk8cGzK
IUompxTRfvue9hO9j3b/WRoULg5OJiQMXEfLlSMy/95wm6BqSKrXmXdnmtdolK2pGhPjY3rLlrD7
+zwJ+BaXj0kP7ej6tPcB8HqlkKqWbu45cFHbEsxnj8bRg/8VchSdmozcFZ6gu/hRo/2Gl/2abz4p
epOVJ2IiexNv6PH7LJOvL3lXwtg4kjXRY77u2dtQopjSdl3irYDEe7f5W3OgFqm0I21ZIqA2mCu+
27PODagRlNKWJlWMHOCsZtDe2UBRqh9/q2Rc4roLd6svBBGzioQ97/B7Z9yNT3u8pLYYp72UEuM/
ML3OkinEtIPEWU4ibjGB4fzKUr6ZE5O1SU4FwFibVpMOlWIllQ1pZAfhQPsKKQnYCW7wR2i2KslG
ojT+dC6a0wnJj4wh44xTq/yGj1vPD0+3R6esr8mZC030gx/nHONORBlOMYG6Za6w1OhUJHPUJ8uf
KHAQ6t1UnzgFzA1pNvCDXiDzS147w0rG4/FJ0n0YYrMP2iI9fRFjfllBzAoPuCpggm8CwHGrkuZ6
MC1CtNWfxzk3bQGtO70+9Y5s5sYVP7Q3ZtrB5n1q48/W9J4Gf57ZfwY/UcYeUYxBH/p4gZmnDou5
1saoGjfo9miHF1obiRJyUa2wS5Kvr3dCHeBo+tB8hWPN2hE2QyNrP4HnUMRnaRSh3rESKM5mPcRi
bFRhAGZRsKWNIjk4s8Rc336YBBOSVvaqYB5nnKRSoEUhRyyMLfkpkEO0G/QXwv7TCkSVnBzW09d3
QPSd4xEOs2UsBP9VK/iXcnahSRZiWwdhgasyCcf5N3Ge5AcfuUz9bl0cKs8OFjzIRYc+4VdLjZNH
J+f9rAxGSJSFxY2smkqnyTZQHtOGvtXalucJhdX4cUMNEaL2OdGTET887GYVycfaQBkJ3JDvJTLn
/aqFFGHPxRkHw6tVfiTO6kru0jDtIdrr70fgnvoOcvt80qv1chZMzm38mRB6sQQfUPWhmsDH8RIE
/ODrksc+tGepmJosO/32Z/6euVhPvE1MQl+PVFhZDAuMEokJdl5oiqOEJpAIVa5qTltgel4d1DPZ
1xD5Z0WgzW79W/xdEtiCxt6gWOo1rcBKtnDeiTmrFdxD53Yi0ShWq8mOgqPUeSAZnLhNkHXmRfq5
A+/Bsc2TglwGxrTzby8maTnWQ2aTngFc/4KKAMSdbYAGFDxMYK5+ea/5g9f7qpG1Anr61vg0qkCl
b2hh1W4HcYdMO0J+9Sdc7Xq/8pXPSW+PnI9LedGY8KA6pk8QpkFpruecfqM7XLoEYfK0pUnOqDyi
gg89buK9yKe4SXNzrbmqqkx4kXD4ljow6yEV0u4eJZ4UrsE2/a4gGVj6xxZ397nt4hVJGJim2Uu2
cPKqFwWgjoea3+4nnv62XK29L7AlHzRJGvvu4LMRzjJDxHWHUU9RMEHGsa+mDN8wqoDygsSgItSW
M6zRy7EewUU/fbk9zXP/4p2SS4jS0JWTdmZk7SUI8g+G2q2/YSI83jFvmcQAr7oGip58ph8jXn6g
J4s90y4zgaEdrsCMBN6GSd2+PaZPXk/Xl8xd/YwQ283qgAelvL6k3GBF5FHnyYrelv5SjSHkZlfC
yI1hoUQcOq6cQc2YL5pw0SiRB0AqketG1IQO6DcY9lrXZnVXnVPzKdoPDAkxJj5NC45eyWUQVpXo
6e+98s4zP6IPVVWC97SVi3uOgWDroJyYAcxP9gQwhaG7Ih1rkcEEmUgED+jwWCg/T5dAztSfASzh
8Od6vd76rvSvpUaq5+1DjbPhyckQ5+sEkxoqgMtVY+odHwgz+kE4Yb/zZFDx9SzGlKHHLDqbE6dE
7cPYuJATEqW1Nh3ZiEKZqbIXlUrhfBiFivZ+GpsIM+DQEhffXJCkrqQWLrcXoFiPam7s6YS8+nmt
2JSjRrHPNcSp25ECW5ZJvVlalJ3na7i4h7gpm4068QqfEdhghmIOXF5MHGvbEkcnITIF5zlbGy+e
fx67mS6HnZZoa2iYqWD7xG0RDC7DdeenxVDISTjHA/sc7yrQcaHyqDvgIFHrfyzF87Ny8cBIfFGo
ugFl6OXxZAgN9GNtSuWrezQa+YZollVAJhWNuXOl4zWyMbFd736u+8XSg/EMWDZZtQB1A0betz2I
vswcQJb/gw9gbWNqKD9Yl4+DNpoig2OFJ/HssxKm8foC/Z8UBfOX5x3zHOW1vimABMXo47c8OGim
xrCRfhqIbGupJKC0rzJoWjsOb8bXJUvvTrMDoE2HjHjURp/SqofsyLbR/a6bNsVUnWfWyG2eAWMh
v+nE0qLxsLuypTx25QoIgiC+aW+aL3hgCk1Nk58ErvML3MVoar6YkMNHZoSQ03MZVgo8rtgkq+yF
wx4/5rAOY6zepjidEO6b8qssjZ2m1un7tcDlvDqqB/7IcnE8EARAA0o7OZ1Pakc53nVl25wrHQZx
AGIjVGpAEBoyf0wwHuhByzoPJ00CJFhbvC+Yw+hd7HS2ehAbT7HwA/XwgiL6YDg8HoaA9XqfAIrB
aZit1WHB9w4T41oS/vkwN0wLSRElo/v3D1vj3pNpUC1wXutOZRzAQDgVl3E6nsoPhY2mDjEhzgbB
/dzW1VWAMy9U3HnShAZaLZLylEBmKAxGlge9xGTLMy7vE5eeBR/rrd8cLtZOt+dE06JTZrHYximw
cmaZDeFum7eGRe+pGHl7Erwkvr3SSjM9z7SR+QHKNKKVVACAveumbXikGgjbQw23wXo+3ysdqHtg
84sqmyb4o+TwPxrox4LnuIMn2jiQ+KO7Y4hGIQm887s8SqBdDRKJVrlV0xsOhtoJVDZvg4hoJcP9
4hBZqHXu/ZY/duvLWt9vcvdvsrMtqgVErTXIQRlMlRKXHzNX5Ybn0YFQLIKTA7dchSIDa5tdO7Uw
Tn5o67Of4pyzLJi4lkfwMbPR20ieLf0b5jbFhB+Enb6GGhexrfQpeqexh+d2AbJFbv/XOo8DAb+Y
UekdwmoSnQbVTdTF7YVXHqXUgPpnEncPRW83ZBCZyXXgZEzJGkZwBCnsg/GKwxNd1xXvWTtbShMI
LaIWupSq4U926sPZymr8lJGg/kGQSnoBsghYEd0tJlAvK8lfZnQy467PNftKdnrS4677abnzNaNe
goa0oYr4EflzC/FZPRnAs8qux2P+ap+r//n7Fn4VzZ6yxk3x0mrReOniUow39fp5RZxB37kXlWGa
DU+7cX48T0M6+o3dt6f8oTVBYMnff3GtCrGkn4TDbcXQKrSgUPWEkDKcIQIpLnTAcawmuIqlt7/1
j42xOT52vSZc2USmySO0C80C93wpcOFHoVhcvRoBc/aycpUOuPTCZUciNeH6QEHVJw/xavlUmhzB
WOQz00s6oAgRN3UTwOH5PiZaHUikAs0izhmi2B9p2b1SnsVTWfk2gJIt24Q/cjFPV33dc8u959w4
8FMDXJZGU4r1Ia5mNW+m2yj4YmKqPtHCLnvE7nhrUjZpbPgKAfgivEHujHaF1kaQI56s6I81Pqzp
3wHP2wxoTCIcBH5PrI0nqrdMqf4W/Xa4SX9iiF3OeQtDJ9hsRpf/0Q6m0fWGD7O4cuSxLpQUoiuZ
dIJegwvFxT+wVawCtGR3l0dSZ1f0QNwTlFhfZV9vC7daf2js4IgtkBS/LrDzF12Z7QCNhKTib5R/
Rn1YvtUGbX8YQw2+5f4FGrQ3vWmhrffUKhqC7tcfJLAUWex8PE0fZ+ZqnsD5yYF+8ev//KDkapuF
yr7jphVVrvjA3V8IfycIPVExcDL1YKX3ULuhvHCBaKuriijWK0csTl8TfrzSuHKVeltwnOZ2Sb2N
cPfS6ujCpgCRY8ZnIVbm4QyzZ3Gmi+Ycd2VrfMF4P7uIR947pTEyHVx1euXUL/m4hedugrzo4W+l
kUsSQp7UmvC2xh04To9QbExhxy+tJ30yQi60yhRIfRhn0jB/9o1V7MK6kER58Z3syp7u+0N0U7D7
7hjD7BelggytFasw+J+Eg294p5qPFNtj6is8JG5rJRAK2kM93LGwbyEi9fFlRf9CDF4DLS9mms90
xAxEF984GuIVSPrV7rjj6g+nJNw3Xc6NvoySHLXhmjOZ5o92x4h9DxRtM7pOnSSCMEwNi4Gp8cz1
hA6Xs95e4d57XoGlPy1CI5i6d/OAfacevuLsrE+BjhiMOxNl25i29Rg+Tatxxf3H5sUtC+juNeQD
4kbRl9Jl3i65DK5HnaTqVpNhf39jvDDBVxAK8j2Z+g8eklgh+ff+Qec8+68xjMvJ5EU1XmMjdkFB
htDOyZ4Bxl6zlJHBnAtZ+FNsx5icrQT7N98dWMm6sa6q2JS+VclwjkqvJfXhRQRbOqyY6KPFtaBb
LrBPyrN3wh2mcMzV5eSAa2Lxrt2cE9a+xvbYSKa2DpvjgNflvEKYBds0xwnuv4hUgJx2DZ3QqrNf
RNsudHF5+mdpm6ZiYLKaK94tHIWU4i1+iWYokvFTcRo+0aqU0GMO6vvji4wgybKaV57gpmVFpan+
8ouEbqBIsZHo0f0slWwZlhYBVa0r8cSiJUlr0llk73tqvzIoA1E4LC81mJ8b8bvOdrApt3TSzdCj
OpbV/otjsUsKeKvGWvfrQFgCKN8HPOaJ6ebpg0P4VgjhvXlOluSOGvCNTaj3zvrmvgymf8aPycQU
0oU6H155STcMrhiImD4uBG8EQWpPzb7wMpZPvGVSFf16ZLDHGNg/xzro7VERv99++l3h0JmEe6BO
TBXD2fA+nECtmQhwxk4U6UOXiF5ihPHeNWeplRl/stVF+avP7GOE87S3zLctQYPHttCohA5C2bH+
R9HpqXrO9NbB+dbta/+L5fNtgQjjZhZuc/J/i7+QmuxSFOqXhxBH0M/y8Y+n8XIJvsM5pQ4X3YA7
AXlHWl0XC31Hdx1KQ4uJ4Wv/4xPk5Brte5zIObuPMDzCqiVir0Dv87UkW+16FDAL14XgFXQJJMft
fvutgwi2srOkqc7Yye0or/ivmBCuMkyyIgy7wZwyg7Ny9KPyHtDoWUVgj9fAmQbRsA19t+HJa6Kd
wto/LsSIDEZpslUpVJwG3mmYI0b5pqw9/0KEcdJSlpKR1rPkZw0EYdM2gnXmwrhe4UBBNWyJ9uBv
giVf6E7gRkqTrg/qvbHa/usig9Oj7BwGrZxGACDk1wfimDj38/xiSyvl+50d97Qfva7/1mDb21/S
Khir2MyBKY/6TDTXSP7t8rC5VMsSjkELGHb3TfHXT2Jn63sbBtluFaLbhjjjI+kh2v/Srfi1feVo
XfBjQYh3QVMGcskyKNBbzDy4y5p5FrJeU9lmQXX74jegEz8Vz3tHBDB8EeOQ/+PQdVNlB+4j0Mqp
i3LlSvZj063pw2/4fKrwXMr0nNkaG7LQt9kgMc9kx2QFMevdrzwVtHfthBsjtp6qrmazbni/+HLE
1rUUQfWZoheQ9mbnTGNhBfZdkZcUW+NXoDCwKV3UQsrQI1d4sqap/rsPkhEEa/JE4ccEI1Vr/1ZK
+wOR1F1DpBYoavR/06ke/aZ7AT1vRhjgIa/iCFpJ4iOzkb/+1aVnNlfvkjD4L5ISWQPh+jiEkko2
0o0fC6ILl/U7EhgjpVG7KwGWCd8x34ZUuh8DPOitnC9ijpmNU56I1SdLy5xCQRvsgK3fNih/Ja/K
zqkccuzF0nWnnZ1tSPxalpmwm4coeRXgscj/sHxH9+lyzw6af+oFkDRHg9cke1mAwwB8wm6V+bHB
XlRWbDQma9uJbzKYTMxFiVUTKR9BuSiz+Ke2zF5t1rEdd5FHow+WkYDzApTl64g5IAhA8NapdP3n
A9ode2Sr0QlT3/2WiMPzZo/WAtiOqFWQG9MjIbVfyA5zJMyVObj6EJGRxYwMdOL7n0tfyV8lY4YR
SRBb3EAjUAxPVzcYyjwzTQuCaRjLcOtBusu4Jr9mI/R86/vg5OJf511r+KCYvcCoKVjFS1Y8SquO
2A0wJMZAisoaH0tRUJhmfvK1oejRUDI/lN+zt1BU0tuKZxTp57v3NQM6rhkKJPLpgiOKanH9Weed
LXVSz/Y3Nki/PvFsAfL1H3wZftoI2cUPhwPLFJwaCmZvvy/yN/Vpbz5CM5GMTGIIl1lHFuUPvlTY
FejSIPFzxLIfgHrottlTxBzFuYWTywkgbve9g5p+NCBSF5fU7XKGCN9GJeJvQqsAIvG2lyizWQq+
ZJrC78n90HxNf8R023aTTMqM9gZnOst5q5YZO3eXm2NiopUlksLhVPCAYZ7EYepCwiUP2LL7TKwU
Emh3Q11sCuxWVf19kbUlhooaxmSTY8RmmBw01FW6EPSzIdFwS5wcTqGJqA1J+0yDDQ/bMULFkyc8
LMLGMNPukK5r3khKHELiBxmiISgIFXQI9vp90gGnb7Dbx3pUhU3kPIKK31rnDsr1gl9O0TQR2waF
s9QLauExIdmmnJ47TqfwQxBFTjfJ+d1RWrkMNmZNEn+RtW91mO8HCl5JrIyNs7eyAHlPtIbh4YfT
uUvwqSXBfySWm0gB+OScrUnfBU3BDc6AwETB21fY2fnHIu/MmjJEyGipBnBLEUJLlQp/HyBB0Dgh
FeZoxLfZDCSRS+ftughE95UWKCN3GaHn63MTNJUMQC9UvFje+KzGM4hyP+ksnj4sOHFsTTAQ5C0M
03PK2VWwHw6J6CNSVStPs+UrK+gt/qI1PghiFmmReVHG9N2t4vpvaZxgWqfMkwQac52Qt6ZITz3l
poeEa2LZ+77YhesYPY+z2M6Q6hoD3PUHDOJvw3ilpamow/uHlTdrTwUjtp/1VIdivdb0xEKpDNe+
DSoDdFTEj/3QnXp5qGxxJ5rKLsEco93EcvQt+Bh+t8LwMGzmZOOO7Oz1ZgyXFIScyPieJYPAQTuy
ghirIQfFvdM6xxEMPa5S4Qzok9QrroSNa2wG4u39+FixNnOvIWnxc9koG4oBLOno4GK/JpqVbDtE
Uv0o0AI0XVqQWu0RFngo4YfgQLY4K54dLHKPPd/9ooFcu0Cr3PlrEUQHK5jIRpTZ9SeZJXkOpF+w
UsKa7/4p6D9os75TxVHfkGHlRc6XGKnFY1mGWp1V9G2HkdAm/nuQd5RFDZxiUjzmglgQtnlt68G4
dvlNaw1VeUV6hH75cpcPmJHwdEbM9gROEkq8SdvJzL2SpIcb4oRliiOC57NL17tsRuQdjGSyc6TQ
YZLpDBUOl7DWG6ODfZLMCKAxarA3k1u6NVK3ytQ+HWVnsvhJorOlENMVqTBVg/QqyajLjVOJymVI
Vfar7A8DCqe+EPYfpXajor+6vPvAPBcXwQ7Oqzx69SfFmEBSxgjkIT3inVz8x/QNNHbRYAliTYLF
P/bcLwjbi7t0phWo1KIPY0+aTUwAIXYBlDYek3/CB9TlntQ6ToJ1uhb0p7RjTDmn6RuesUiBElSq
f6CNDu1jc14uLRqkCvYtnksjw54tT2zqZro9CKxJtKEqENPDhJqzsUvAoLIHP2mDUdTnYv0jucy0
LO5vEbAYCGXhbKEgLHWrxRNNsDPfiMMkErTcKz5LxH3ruAqg3LwSsToD8BSf+9j0KR8FOWIKafA5
CUe63reZG7pFBUs7LwzVaeKS/ZALJ+NHpKRmhzQYLD1/dsQmBe80AUhMthMK4/7fBl4TWYwxmDtT
M0+otvbk/oLwQRwUJlxVm2MBUvqkNex/e0YMkW2x+b6hW6gsxRTzUNqnf9NYAs1d4+Q7e+4rbwmz
uklP7Q==
`protect end_protected
