-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
vEkH6doe5yRkJDvV1U02zX9fUOiSiQtAPGgE9Lw4Lo4TP3kwa3WKSclOR6S6cZmh
rmNWp+n5Tj0RSgo7hueRvySiBsskyuKZcKxpzUqE6GNsVc6NuVMTZJzrXAdswE3V
Mwx8EYOjLJTF04TVKPiGYWdqDccR0EwlWa2ogOhYgXY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 111968)
`protect data_block
ME1080NG01N+BGjhSyESnHmSBue2D5vCfU5695iBa2aCOEKQKaOy5c6uWmLX8NxC
V3szx8MyROv7G6B2lJg23SqrQ3CsXrNH/yLPOSqn3Pmjk25EceUIbsN8E21qN+Gf
bNhdChPjYlkpUO4i3LixB7S/N6bj3YTtTdRDTLhwvU1QT+e34ulvsof5jhVXAdRW
ucg226f2fFZuJgHUZu8jPYEZ9VPdwbybuOSUNuu1lynJl6JWw1OFT4gw5ehzhKrn
Uvz0AkQPNKwS7k7oR+bSyxBSme0Pv51c2qyLZrYq7a5jJysg63/ecK+zq0iOPQdn
g5KPTWOu5vWLI0IWICTr6cCFSugpoIhmQMq+X6cebQygUFS8amvrcNvdZPNe4qgS
gk/Cb7OwieghNMJneYmQfYov1Nou+QP/66NhgbOmFmxIkgFiaovsgBMmH9RshL4X
nCQVoHJ9HhVeww2ut5EA1wZHA4lvIP1If7Q3oWJsQ35hpUKMw8xvYAgI9AydexzR
gMbIN9Cu7PddzzLcFzFdSgHQmePaT+Z68aqlY4Ccay9cyff6Z01v3Rf8ZiyN1iqK
gtZ4xp5Rnm9R/vBXCgTLiIQkdk1+zsFnXoDgDnQhXpQ5HbJiqNX0HxEwWns77GR2
j+hM6C7cC2854HKEBXvx4SkLPSQY5UvWb8jbMB5XAVBAX6GqyqpR8BqtULu5wke5
XG75QVpUSOtFY4AWTN64zgmUsfHhYadtZpxQ+qaSlv05MvtYQydsOyka4/e1eLwn
xzYydvj5usMatjt0zsvPOJKS0bIKgXY9wwXk/gBze0NeN3GL7Pg4Z0yaRrNGU0Vj
WH+DpP8LYZ1TTeatTQMUv6taZEeXk2XuqSV/q0Npb1QPGB+zR456u3lk0WPi07ll
U21TuaTYlednBSc1aRfr8/wWzAYA7SejGntABGJu7G208Kpd5LGy/twI9YC+a7Yo
/i4lLdqhox6DFu8VSlTjsiCNGgoom9z2Nydy1BxNAYG9U1yziJY79gyT9raOPuOP
4J7zGPao//ltTEMfWtX/ZKHaR9AyM1fYj6tU+vN6SefzawvmcSQ95Jn/o9gL0nuK
s3Yeb2pLTUulYnIWW2YXxd5CvPlXDZzUarEbmtNgDefDHmfa7z/QGxW1kGt79CNr
tjv3xfv3KiKSwXVrdZXvRFcO6pxs0KaC6BiCHkAo5fSm6IscoPON9Rmt4gz6HTPX
6D8xiae6ow3ZlDIeoT7BziJG9fjuT6xC2r7lACYgujS7YgkjL/EioBxxeyfxQQpg
A3RcYbGC3uO/IH3rJLPvmWiLTR4yLadxNijLyIt4cpeWLx61He1xYcCi/Xc6WJd1
j0yZhsjabHdvfgyZlCF0PMB16O/aHqyHhaArF8pMtzthf+U9wBMR3dut5rUPPHvU
g2n8HqbBlvAgJL0EpuINR7k5IaIEEveaHS3kfLqWOMSfGNejqUp3nARAOSiXUa8/
zAlq1SfN/xPTEPkGnxWu7QIkreu+ZdPwb8C0QNSXU9LxfOu4HHT+z5QS6bsDXLAz
GGTsyHlfCQl6BC6ITnrSX3EWlc1ywfwvMjeoUt+QflfDXNOZW6LosMh+1nj7wFqO
InRvB132TS3mSVbLiEovDCGD4e+6ARF2KV8vevBLBeKSvPm1wQXEyV0Sv3W284vE
5E6Wn0w6mTv1Eo9iZw58WqpV9ji+jrSzcz88Akak7ktWnue/Yi7CrNMKhJ/cqGMQ
uVhWzBDt8dQEmpWhXyY9jDDMFH4z1ARVh0NSW4RAY4+jHGxex2oAx9ZZ8JzPAcfo
x9jQmweTDQ4eYOfI318W6y3vZhJQiaBu2VvxCCHPF1b7YUzcm6Rf3eHM4Jw2SWqb
qFp/B036IKPZgXCobGwOmW3eL1n2URjqk2A//yFL2LzWF3xRwJVCvghBe6KJvXqw
CMEcN9dbGnaI5mCyBkLul9zjjguOheX6xR6EGQg+jaAxBNexLxn3IUcEFy64Bjq1
7MyC8f8ZoRju4PXvXEe7v2UYiY6rA62clSdPwys0u9uy8g4AGm4QSp87nwYZVv4x
9EZjKXsLMgIw7PGPAWaI4+jHpDV7BWmRORrMr2q3/wOhWsv7osLk30MMZd22J0qs
aVa6JFt7/vXrRI2+CVi8TzBnfDf8h7R3iwaEBe5t14OA8lDjzjo2y3uEOv/CBPZf
1ROdcc8E6jcym6B8HjdQFqgTBTlqxkRoxzlijsr+SbkqepX8sNyrmYdwGLMYKNUr
EexWAai1X3DA+tix51YWN8Zwl+ovd8E58UPi2AoWHZMDRfX/DHAKV40Ty4B5pI+d
GiqiyGYQNvBiIq0D+DbFxoEWtnOMzSgUlXHfRu76vQURFUzbbl7pyRtr0CzxHQqD
HQudTlpPUo9LkVhG9jxMrMF3wGnmXvAg1p7IWcVorP7wS2clVJALv/NiHpHA2Bzz
rKzG+kGOyfQvo4kWFgo7AufJaJgwHEuXrSphfqII0ChGR1rw0cpZohjvyrHQw6TO
ODl8iEIeEDRCVmBzC7k4jJT4HSnG3qSvgL8gzD2BLmQz+0/CQoiRjxd2YujbPbtW
v7p5eQtgsN0vthPwGKdSYq5mmA22GEGp2ZpNPngO7t2++gaNDtMwvt0HfZpaqhxv
G5DEmLUiHkb2YQZXHSnZbCMqbxKv8Ck4rVLi4gnvYQ7MgWycPcNEWXtMG2yB1qDi
isDRkY08HU3gDEvh5PBEkzemCun7N8gxYhCchY8OO+bnt3hkBRhK4AhWfpOWcm48
OW77KgxDXk0OOlx0/h3Te+yW32SNodwkANM9SkIK9qfO/Bw6S6ICtRDnRTbEsBoK
EOJYMAkCoj4zX2DSBqDC+TyPEzLnCQmOsK7Fw8WGNkifHsH4peByslOCLORrmj+W
OvYQN9Ptb9/pVuDS3cptx/+acMXparOVSX3fyKnWqiKbLJMboYHBETpfXrelB78U
i4TCYIdD0iZGB0E0s1dOjjnH8Yu3RxMEPn3SKR+8zO47WMtOAT0qej+gn1RdAS2Q
C42sN4iVkaovzbfZSk53Ry/CekyQdM4co8kg09zpnklLc2vwlygwmUlNTtCOjiwg
krHif6lNa7dNEzyNh0sc5nx4YcrfoZNW9OApRlHMvHzs1DGgVhtHgAVQ9glea02E
3DJ5Y2E7yUWCJQnas1tt//3VJHrF3w0hCBe+qFgETUqwLJvlLcTtNbZa+E5P8Li1
i9aGUyZ8EiMtBD5rXMTpQsV5qSpkfw7vmUuJUSLnJf7aCX9JHgxb8gnxnok6pknN
Bol43P02vkahmJU5iA3i9RsMF1h1SbxaWGVuAb3Tbgdj8Q9oqYMe4ge/Ic/LSu4X
cEneIZyPQF76ztPzJWaxrzQ/Z2HnNtQ3npRaZlIOo5dgnGM5r6k++NqpnG7zZixd
SYX5NCqCR0JldiSsYKMgtN9exRm4WLuFcjbde0TinOgyy1pxRivbVw1trsTiRzTu
Lhs98b3YYfwEOUvR2x7fL74eriFEzVoN5FuReKUB70ygQFrWGk1mVxTlZAKliWhL
vK+Y7igdEzGtEKX6jZrF+MkRxKsxCjePJZoH0d+LuysidJRl9robwbMIcfSqFwxR
osDzvXYunYwywnjBU2sAP597aG7bhT3pYM8VqMsMRdTIi6jicRrp/ZOhjBxU160g
NM5fM5lC4LJQbInsHBPiPjhwgjVl4TmtMGLu1XS2gjfPackw/MTZ0HhfFUIwT4s1
VrokpUQhEd9AHvv5cVTK22Cn/UG6pd8GawawsSXTVXEw66AQJXY16lfgbHVM/roK
5f7R1IT6aze0KIxuBBGuIvE5F1EGGCT3TCxmPjiJjDzKVcKk7cUPLRmboz2jiE5I
gfrK21s+rLpAr7oEOUlmU7yK13hfkMHES4wMo0HBMBdh/HNk7IYz8OznnXQwi2Id
uIocZnG+zbd+PxM29cg3h4TdTC6/qIhW7seINvRZRw9w//KiixUhV+R2QyhE7vRT
sa3l0lUj//kiV0qRTcIXUA5dMkv/CoduBsMhTeZWOnh/u12aIn/FlMWUyTjUmoF3
JC1eR/UWbCmZqqCKIMKoYyAld7j14emm9l3GatAk+R89XBAG9NgxalVOBl07V+zK
2bFiEWI+KLbirttpJoBjKOZhQl2eJxS5sdvZKLeA9K4OJH9J1puqaZARwbQwG6KY
3RJElvJ5fZV6gkmQXyNbqWD5DjeqqIHY+cDq1w4LUyEd9/RTz3z299g8UVTGfAA5
JSmBzHXqXnBg93JnaLhOWkhdpzVzDVycTrbwqFMehMzTueKSG4akn8Typ4oJE2gi
vKnjjotIySErn5rOvbuDLaNCkwXrZ3ooQfi1AYDINT89Jeb+gelIJzp2FgBdRnzx
SxiKSl1mmLpez6t9j/tUJpniG32duOmWPlUVLUXGKSQX5hI3iUgjYQO3XjMv0mU/
c+Tfq8Xy0HFHn9q7WLIwd/JrAZxJriojcDEteLrZosDoO/devbNPtRwmCBmhRkpa
T9TLgGv9ykUsa8QBXHWktyZ2J6AzXuO+R78HoYzJdYI3ryRB7ZCWJ4543ZElh0wt
ZwbO0iznaf8umvRtKPgk0Aocn7K1y2TWxcFJoDIgisndwsVVHh+9Uu0zGFmpWqsT
gVars1gvbL2LUlEKxb0r5Q+GeqzteIRI5ILK5bVS5oiqOtaonSEcLry0yWv40lCp
pGbECf18ya4RwVgIzohqPuQmRTBhvnB0PpY+N+9BS20P+8lvOl2md1lkguY9xlyM
VlxCvfBKxXdFCSo+mmK5DNHT0Yj5f0rxDcRFaiFoM0m1gAJ6iV1MpIOsviKscoxq
gECmbMl7KBd4WZcizPCLimA0CEz6r+uqbktnbu45z2Wk4q8mah2qABsQz+Ri1FNx
C1u8w/5prOauJCzcUkeSlaiyJIz8yA7n6C353BZvyZypCBvD42pgScXx4ctaIZoh
zcSXguKKTF1UimSYjhcF73/bkFY79W3g+6E4C+NV5FOlramdGYTu9GIXH1mlbyeS
FtNv6W3K0Kpslle6Uc5uFPvUEGicrkctQChuYJnYWLAuXqWBx7nFneiaKHNBJZmQ
mx400qbp9lmHjZysAjraMeABBZzyI90AQMqQdOTJrLZqLMwDds3mmAbFn5cVjgwj
436USLWeU+uessPSEYj2b5eIP7XZOjNftYa/TI37hj5DeYF2v/t2TfojOtTp1PEr
PuSa0MFRrxS6T3SSrQCpkYfoUgN4Sq00wB6mDxwiS7rA5UW3DNGCXc1wlPoOfhos
mxy39LzwLts/21oIVTLTKYFI3scoitxEh5OAhxC6yg+wD5RmKisYLgSMO306q15L
BvmrvzhRsPJ+RquP8daX4dCCvPo+HhdJZrcAOyRbj4A/hP/3Mvg1Y43EqcI0trux
J+99qHsQIDH5nEEV7KMcfdhJzo6f+7b1r7EM9oejZezEVhLFyI+42d7xhTVz1wzI
TEdj7n0clEVgRkBmRq00PpKYWsF8YPumxwnaP6of+0zGuD2/o0kvimY5z2/Y+rw8
0JOXQL7o9K/GpN2H8vYj0w/22AsIkQ3se+BdHTxlwtDMBHxPW1D1053/VbprtoRP
1Pk7MoBZTa4wcclIC9RmdepoSLKb0Qj99ihj90dV44VKS9wizdasifn3+ZO8/lHX
obsfi0qVkhNpLfY0Ue7hOOoh5nq2YZ2IfDP1m6Yi74ZNVl3UzQrKQy9riCi7q2Vv
eZ56adktTG6ZC19jhynHBHHrd18eAGshFCBpsM9IqljpIbj0NWLZiK9jVBpM0cEa
dcFQGgkxp+OVAu6qalDXW7yV4lZGjstoCc7ZyMCDiadvaNfyvgxQ8qyecvLw+jWa
fk11YeXux8DE8XJC2lI6r3rRAnpLcNVy97zdgF3EIfEFYl9QWFwr/gRkvIHRv2Nb
edc1cXqPvWp2RninT3Tcj88ZfV3E40djh928RJ4uNEw2Ihs+oTDSZfSWxTHEq9Hw
0a17pKUtL0a/FJRkhWxVXy3/Y03N4HW2IICuLGYlm/9LSuw9Z+Al1/GRGOFlT2Cb
LL9NMQQgz6SPmv/LKglMwL29nELtmtI+vYU1ueASjSRw96tpRuaAoBqAOFAQD2ac
JP3Apbx+I1JPSPHCmdnaOrxg6NlfTlm8vdeMMOhGXMBGE/JHYTYyZjIFeif6ujCL
dMTnCztF11TWFav2VTNnNo5XgDaXBcg3D6/AR6BCAxmILvBrW+osebuJZs4mp0q9
wZQFuZlTErKdQu+TBCHVriYXNtOBeoOZZpLWV/rDHE7V0ElmLDr6wGk/rQNx42tZ
t6L1ecrnEacGycSh8ABCh/0bFmgB7DTEUm9Bn6FqitulUAd0CSL3CGC+UsszuMSf
yzyDliCVIihAQFg+zCM+eatpI3o8kRl74W2G/4AqWaUpRm64ziU4sPTpFxEEOqun
ucegOfQ0pzJgQj2pMqljkxKIhnVHI0MXYVsYu+QRCWhKoa0AnDyXFj6dNkm6CR8t
O3CRaDFtDb+WEgCTVXdlSulWzb8jNlcGdCamGcCTCLXkaj/pIigV+KGaiostfZG1
Kae1LwfvZF54G6NRAfMcU+E2xUKyf75ztmDf5brAPP6MpHhgQ7Ca898HJ50GkeMG
Vhux5R3Wpi0v9ztLmlenQJx3dRaCaHP69GnWDOFyjKbM4+i9F7uT6mnigj3/nDmE
oGzXLKiSkGAnEnK58g368lSs7fEZSZdJuh+LcmYHF+CSQgWYWNjkh4oyBkdHoQJE
IEGeNwvjS2yjLzMfUrAsoGE15W84hVOh+50/rDNDDP856IXH3E+QDi2lOvAUK1D9
yjEzWJamcn+qS3/MlIj24EmGVWLgGPfYrNqvgYcNgSb5sRSwKtVfAAFyTEVlXQpC
+BS0W8Y1ILuZNXSSDRhJFC3drhYHBGy+B9ks2rTuZ1Xd+JefAD12wBD7BkQyWYZY
LOYokuUX/D5Hz5SL+mpF5yDoR2iUsZdKC5pAOjxTjFtyNt9COgU5NffE3dg0mb9n
xyRHRI+nwH9uFM9ifjUKbJ01ybP/ICY/RlGrpZK5jy7yCo6tme9vCw1N4eJDSO6w
38Gv+vEMA3UVYvoh9tmGQ3fb//OEpETY5r23Swmh/fM9t6PVJGuWk1+ZCqJsiF8q
NitMcaOGRShTe3YxSRMqdNec6Wp0Wz2+p+ToEjYK+nEkmvpAg/3HCFdGHWZwCE/n
uc6rE3YdwJS/6veaUOTe7xHb3OrVdCg1S4w5nRUr6O3RYNK+YNYcK55FV8voxpmM
eXzfSH/B5baWnKst2u3G25+TLV8mlGN5tSd6mRGbeiagm9ktjDbpzeBEJ4qN+tj0
NEpibkEIDe6LLFvgkH6mqf7hHohyTpJZhZrCKuntO6P8ALSjpk1NS3Q6GwS8vBX5
NaSM93DnQRiffIAwkrALDpAcEkCv4qUFTxfS2ct7+FKPUHCydarBH2AIFrdcQ2WG
8sBizM4xCAf4ABkuSI3oE7GF4Nj2wP61jQ2PMYfNl+pwhhigz8yJ9QCHkAFJ7cJC
16odT+ru/o3Dao+Y+c1qqleE8Hj7J7HKCHZrPpJPy5sbqKxdgOhhb8F/7pEtYSHZ
/OyfXfgBFhN9Fi6Een32laM4Ohs6wvnayGiJbCQvd5IeSPftJ9IFXDwrTR3gXzV8
x57dd1FgIjXh+fMlQU/5PbjE9TTyFNDJLT0mJQmz5zh7LPZEEH8AXDggJkea7T1W
30zgUO3ja+WjzMJCRxRDF+3kTMORQCO55pCR0diY23Gr/gpyRRX8uMSSoo2BC5Mw
mvyaS4YaXZ1OuP43508VDf0oFL8uw+Xt/B5T7DSg1YQwUWU6xZREKtNmo8d+ySma
jtgAPeIVqKzpHqq/UOjfnpXhh/O0HKClzk8pjpZeeXJDqFZQssoQfnIQpxbjUCWW
xu+ZTiXeLcX/CR2Tl6sjJzzginX6eHqbcl/ZnO9odwOoze2CbpmVE6HlbiS5rnk4
gh37/yIlGYiaDXwuoHrEZBEDLgcpk3D2xjbjOqIZXlSZZjMvNxItqZ/UYPwnhhCi
bFW5bf1IIcqf9by4ckTUurPc4FKylIn0wRIRZxTocK1D1hQJ0qYVVPhWG8mlkkhW
quvcncowobjdMUp2e601+0gGcyA0U2mdNeJ4Q78r0lFyhaV3bwjK8xE4TxA8NrMa
8JTkhpVHRmqM7v24CLmKN+Nh0IjgNl7hzBZSKCbrLZEgFm56CS4wRZr0AtPaWPdl
8sEH0cDJty1a4WkunR/zy+Z0wDdSxWb7A15gdT7mH5k0WfLIUkFt2yvvvFu+mJQK
WtwNg9qnK5HiKoqPmUmZ3IC8A30jmTFIbKLPqvoITWppG8Cj7V4vs1U7UGiMWwnf
CNXpNPyZ9V4dSKIcoAX+29BG/dcCblC8MXNHJ4dUUtn+evIU/sc078rQFXpbALxi
m0ExOG6yGrL1FBhYtj8RMrTS14KEPoXg0USu0deryzilCKpLPVEtabpm3+DBk6oy
uxJECeV1nKheG+5AAO12E1phIElsBBtylBPfjKztlh8EvxQjXpqZfmkxuRE2KiuU
Ud3atbHoxYTGZ7Fl+YHbWqLkh40rWw+suKIG5vBKpRKSNi6D0Jex2VIUf8zVLoID
Sn7VN1DYLft4JJBm+yOepUCW8o8mokLp54GsCLVORpT/nwEW+CBSUL29p2/QneoB
OUj9/QzddrZtILsCPs0fw0bgJQSwM7Gbmsy2ciDrJdQgc54LIxV1Yy2+YwloshUt
Y1p9DuUaVw2KqbXX+QWDH1dJZencr1amNR69178ewk2QlN7Se4ke0ow7hGvTaXKP
CoCi+GFfQy5dbQlF5R+NRD4/oXZCsF8fvazvOjLk3yHtm8mswjXk+cjjFdtVTnZB
lPY22axc3Fq0jpsY/ZMDM4oI6CBr7rMif4OiVqckqLgKv+l9aXtYAaFqj8YS6f1c
EqOtGX7ffYolLPaHl43DdnAl0USgpQCLIwcedjXP8S8GqpfTNU3TZGaZSe0QD2nL
6cY7HIffbiKdrYhJaFNJsZCIWA7QeLmSgXnroykKUuhuKZ7XlsVXF9gv6qkFz8AJ
lmyKf8tkpZf57F03CZ1yqDWfw8Rnd7D9pwIEc4eXFkybfi2pil5GxtH8NdHh7dR2
ypRKVTh+mUwLhFrUu55+lITfluPJrIEIgXEXQ4jRO2T/NIckSslnErpgEPEaviMl
tRkKKFJM4aMQdVHnOd3Lr8vaQyxrvuXp81/0O4HlPzpIOUZWKJKjeT6qNsYslxDl
V5R7dD0LnoR3LwNeXwhS757+N+mPdywCtdhthSPtmmHGEPR4ZJ6nwa5ZIBJN3d8y
uslAiiEhPvyh99PHyHUmazvvxcitD8sBeQynBdVnwvRhYxzcd+ILGOYk71AebEMt
bw7YYasFzPNu0QFDvsh19HimSaEyYa3sk97p7wvkblDihwS4T3Cv9KR5ijVEOTol
Wfr1jp3Pu2tC7ghuReYHF34gMNSJb19fTzOWf1KjUwcnVHo7/CGxOH7XlJq40TxU
pD4dzQbhcq6Mm/i6fyzCwMNV279+gqKWMb5Js5ScyK/ZJpcceFxdr7JA8Rku7+ow
alUbobXNkm5T68AXMW6BfBrAnwXoAdoJMxEwDHSwUZUEGl75aYrh7rMulkdlsRTQ
Mv+Tc/A6UtS4xcNnZPNU8y75Gt/ceSONJJ5xTNMvgFq/NOWMwP8ULEBXQkT5keYu
+tfokpFHOajHoaEzYXuP286xctY0kcM21AGZlzCezRpxReGA7/y8Mnq1dc18+u9F
5hzf0v+zEP0TC5x+18oIQvXlBxcsdEq/bB8QyVVaDFtM6TymwmQ9A61vspBzsBv7
x8lTP2lA3k+vtp/p/RtNZ00QgJobLVNHufAxmA6M/ktR7tj8a/y4n+JclYWdo6Gp
lL1Mh35KMI4ChqEUOFRZbFOXJxtqvl5/tLLAUKutkig+bTTv28S7XV/ULDtpeSjZ
i1cMk8TdSbDzgLbYhlh7UOPXObKB/3o78N6rRsFhz9ZmT+k12rydcX/9ajnJgvK1
3UJm9WporKit6nanPr0Ss9zT+H0K+Oq2ytplufzzwosyegoX4G1FT1ZdBTk/PjJx
GUR3N4hHe/riGmkxehW/xPhZ9uNz5FgXyk04A+4X+FzT9g2foUvsrimqSp2+KwiM
Lw6FBEPyRiP0mh3+Q7mKQinEb0FHKwYXLIe3be+ICKtprmAWOXS8iz6M8VGa8/Vl
Zj/c6OpKEzh7S+CXE+vY7hSLwsdGQZwDVpVbOGb2qsJjJnGustLkgMiQOusya/al
CucaouGz+NLddSRZBZbquNaVrzs6SXXzvGLQq/uYDdxDXAwaikS1CRnaGIfRVEH1
vLR7sWVRUbAHddSL6b52oTeZKqRoij9T3Tq+BhEMOe6FeSuKgRGspGCtwf7ZmCi3
SkeYSwwdspM32NergJHMzut0XqrLLFW3DHb8PKao3ZoW/fwRKqlG+05TuhG9Xddr
Dez6j6YUxjdsE8zfzWkwmURNvq1KgTdEuf2KQ47hQE2/0aGeqaNzI3iFeAsJtz8q
gFv1tGxpK9CPnmdnTIPiwsZnyXjzMcmw/up5Cilfy+KUhKp9doyT/XK9AQmt6x8c
TgDZk84n7zesmXBi54mbhtDBx6FuwVSmt5gqkL8fzYY4fNqUoR28XLz2rVEkXTCj
57kIhK0Tyu5rr4XpY0S3GraXMWYeW+rdRsBXwJJAiff3QyTimi3W6AI50oyXZU/0
nV7Vg5eLL+g/3+6VVrog3Rp2W4cTY+z7QZE54OcTYF4da9ROUx/ZLOCt9eJD7sNg
B+PhUKl0cYTnzNqnySv4ZwZ7Dgmb0VEfNwu2MIUv2WsJnAfgyFnDyHDkKh3J4pqq
ZxPeIRWEB6kVZDjdoNImrDpSA+A/p77j20JGfKMjr6A9HujYgMMBVe2Mx6SyEoyM
3OHzkD2KMF68Wz6Q9CkKve5kKwgHrdZkJSQ7kHshB2dfvcv2TzwkDABkSr0NgkFX
aZgOpH9DsAuTlG0r6g9BMnTm6t7QpH6w7SrhbFOoMQLlYZEkg/+cgrogIoVdZp7d
Jk3v3UDlv7GQvFxsGjELybAAaXLUlELGsENHHtGsV010U8xPMpDx7yejGXPTfVxh
v2zFN0e/1tbEpkurOkwrnofCQ5ZmbptdeXRvkLyTGsIxKt9RIahfZ8GXuTFRAa/i
43KU5E295UFsQwHUfb9/Mrwq9dQ13dNtwTiFocb66mP+MQJChnE9z3+BNFO43CER
OWXinspopJ/AVcpDhXTeLWM8Byl0K6vzKznxGoP4S6BhBUFOK4XKYkCgO1VUKg4U
IDJ/qVQcNY3qriYKSwhi+e8Bg/h+c+F4FBxL/dmIKWDrrz98/hyAEu4oZ9Ik0GKg
BT1ZClyjreZ3rNu/7hCaoI9hH0i1ZDoWiqosxKs+j/YMgBpV9FhlLk2P1T+vhOrz
5DnByb/rOzPxjwyyNYGQZ3oJu26SqjPepIN32FEP+rBsOkD16DthgWj/0G7Yf3HS
7fL/+Nd03KoF8Ji4Ep64wYPeHU+RhH4sYP6eAd8jLnOSmr0U1A5s4ECzQR0JJexc
Uz7/ed80nExF0/pg1YtwgV63RbwVgm4te3nAbnjIFfemoGNm6GhkSf3vMki9sz2Z
sxyWdjFn461jBrLI+gBJHfE59r0DsVWY/OIqzGCDqu2SP19iXAos56tdBvEZU9bi
t2Kzd5a2Nw7aWEfk7AT6B00DYPbb3DftTz4T8Re042q9bX1GvRXcpbuXxOhQlVcA
YpqD/5SoofGzRQi+9jtGRsZHeX7tbw5aC9y2Tb1LbGch9aIGcrGk3iXY/FNiwP3o
fJBhk0fPTVtEg0E5CmRGUZq4+XuyKkL3O0PM6nywH9Cx5fZ8gydd2Nl2/2WGoSup
l1Q2Tmt3pybhram/m/KRSWFmTwpPYqxzFenIDpwQFrYSMwok3YaD8W4KJtlplZEa
4sLjCWK+QZbfrPy4Q4z2TzX0IqJUtHyXF60UickaWPv4/hm9vDWk1AnOnUVFNoEf
1KEGQKwrCSXTEbfX2aqIPYhACjTdMLo4e7fOOC35J4Lgea/EnXSG9GZAYUWd3NFK
8zXhGAEnJovoVlHuM4CiAaUPut+h0XK/OHVZcTBfyw1pXk9zVBqPctsF15JVNyM3
AnQ7VitkW7TTW+uz+HW04eGo31mG9iuj6Hep5QZcu215jxGUNWXJzDqiphAl55Wp
mq1v3bA3TZiDA84NlF5Z0WFEldb/agK+89z3lXIJJudwc8FI8Mw6BQEBPEBc0k7L
Zr8sUsaWrhIleouaSkvTE4OK6g/3hgCKqV4SQXHHHw/mC0el/2BOsLRctHKzp9t5
WrhfVtvioaltNekflDhdhnMYlVdtCoVLC7JiiabkfYqcHWwgpAM0AuiTF+IXEZfv
Fa7IOWVY8XV5lBL//PIGquETDr1+yGQRjECBU98J27cfp7Xy8vaTGIKrNPUBk1mG
/NFBET+XbxFPTjxaNWNx3JCzypeuOR95ZIvQHznbRNib78Sjg6pRJDmWD9voxuz5
79Ihbz1Cj9PhFeeKKsUd5rlafR2t9IqV94EqBgu3vXVZW83y+oJGtjkowKW2OJ0E
DbZteyAVe1zY8Xf/s9kmsYgMlZ2+U39ZFwTJfD9GBDtVjOLmbrw4/pHbpt2hMaI6
mcS7RPxaRY2qyxqtnHsDLMa/76ljaNBQ7wRtaDhD0iQP/SVK9dTl6PzifGp+jPc+
4G/OS/J1GnN+leNrKLwXEcwO9PNtwJ+dbPSCYS1rJcyqqm/eykI33WpDxVs9fam0
0SX3JAGbUrwkGHxv/yOI9Sz9RyU4ts7cVk1acmqLHBUqvT4Ic4BvBhUrT4iJkzw3
yyP7uy3EgphsVXOVeABhnJrlx/b9JrDNHKI8+/FMbTQE8lXM/77duIQLm6FSeIjK
b8Xn20jhOj/KDUuF9s9DCb8IKT1ucij5MblUG81cpY8Th7LPey8WTzxXOI0hWta7
+1eNxSx4FWDxcEj3y6PZ9mg3pZRgL21v9gW5fOhNM1AsJR3EMUKe6A0GfRFhBOBH
nWpR1S3jcN2n6AWS+lknZsrVmIa9HF+VEFCpB+DqAL6DCQbgQX5n3mjL1Wme8+3C
BwlE+M1Fg1ijiRpgy+WwfRV+xS7ltf/VaMQEd7+NEuZLdZLAjHbN0dmjCpyvN/20
8qNpgCIfO+qYuQYWWdTxuF34v4cYPPQBoNhcT9pDHjRIjyQCEoTa4QwVvRZlZMrJ
N+rdaNUfcFex+1iS6GGhmCgGz0vLnCNntuGsZvKeboJrwlASAAB82GqXNCwaDtC3
rtIQZY/pUHmhgrmp28hlUtzmFoxmBF5Oj7kjR8W301TbPsDLGjJ3DmE/5y0eKXLT
oqPH3xUcWvqXDSgXqDPm2LhVFCDGo42TrBHO9zGU8+iXyMLB4fh3YORYpZPN+t92
h2UhFMFMbP+F6UHKk51BEPZgSeHyTY9Z/+BlBVWMJuxjcopfUDhqwfMJzsGpJ5dr
1/SQNoOsOx8kmmgmtwguDm9NHsYitC4SqlKzmz8wi4N0X7Utj/V1NOLZfWzs+FnW
ntZH5i+6WqnM7A5WNDd9FhIIHZFNDwmMviY9bdLaI8z9a4q/Mjm6wz5k3XzBaXso
oPL9Ya/FAQFxVzNgI8vAmfqNy8l8Nhb4tFRj0onQeg7rp0fMvF/Z6MIufgyKDNNO
GoH3ktCpcGFOuovpRjYo2clwKbt7ND9zpMINsxHglmOJnO6OzDM8D8mexRMMVSlf
b8Ed1IchVMiifLGIU8aSiH3E3UkHH49VhAGgvuA5boRMVgXVE/SN+owgL4eyHmX+
3S8eKLVf4xZNQeTt+9Fa/RM/Egddf3DDAZIVQ5Ubx3BPaPZTtxdoSVaFkqymoDfL
bXB7WF9rIZADXAWBkLon5DNp4k7/mrj6E+WpmpqDReqAx74ZUbrKwHDLe1XvX20i
i4TfL8Xq7AL1sKG4cULa2BSOwgNHltuqdnmxOfxz3VLIin+I8BaG7VnKd5Z8JjsO
GMsgSdKxj8dtRJtAg9NC/e9HsXNoohVxP1bf4syWbeLjItBLhI00GjfyqpaxmQ1h
fuuOm1uUCCBmQL/nfHvL4obiG5WJBJxV7QJKrNn145FOWLg3xe+HH/KNbJhFzP+4
i93fxL9FJoTRVEDdvgdeBgqv8TehNYAQ8XgW6V6CCKh56FNKytUDoHv7Vf+5H9kT
K8ufj+AzXoAOdjbFFbNATCF13o5XOHuAk1/4P7sx3rV+B2hWBPcTjb5a8nOI0o/8
Iz81/Tc37JRDT6ALFSb/4C8M1CII5Meb/h/dvNNXNoY0/OqmhdVk+r8s14+h8/Ho
k+OHlbTs/xJf2MPIwSwWaQahFE3AfsojSZiHYBH3Qlfqn6aoM2AsCfaD65GQbAyk
NduwJKfCnp8wDu8+NwzQjj2y/wmj9DPb/LjXr0g97uu9GrgRYi1tHQGkG4GcsZ6K
I0AqWTlQ5Az9Lj70eaaAeQd0IliYT0wG6/Qr3wMEB1CFtC5X8a/hn5s2yzTbBVbX
CsHGirw+xD+iJqwoaaLgBLQm8S7h3Oqz3y5Eg/CAVPTXXjLsYQY1Q9Uc8fJAWpf4
oklrocWJwZtzOEUOU7pf8M9UhyTVeTQ+uVhJwZJ0QZnUYDsIK6GhAFsKVaJrUmop
ilCmUZgw5+iXVsmKttmaGbkhHVidSFj7f2HyJhGvUvg1jR6dfbtAYN6Evu6xQwW6
R/cVmdO44Br+YskW/mlbroWyb85TuUNsVnk4h7I68LfTGC54sJPwvJP6ERRtCRK1
VEZeWeopGWxH7CC7IcXhLyDg687Me2qClVObNdFOR9oJ5lQIrRt9O/Bc3hElrpQS
tnqDygmtIYYt6WZhTVR8vSVsRSH6FbrPswSBGknnCW2kIej3dv21gTX0uoSj7K9O
ZzmPO/+Vp+wNlE2IRWgXMVs0Or5TxZS3TAdOJIP1gqJAlp0pjcL+MdsKBdSnLw38
4vcnKHzhliJLmtRDWGHnNeHNPIIjUFuKUXtYQSIwcov/q1egaZxFhorNeLRcz3hY
oz+PsyKIiffaQt6VTXY2fc08ODACCilCVj0jyz81RmfE9IS2RKX+CJGrhuyUA2zn
B8l+PjWSnGmx5PdH5KDnPIfxm7AX8w/t65xNGi8D1UjT26toX/ah8I3oPSmRmOLv
pdf0oLu2KqQmshii/B/ESWakmTe75rgGtcnVIJrxq8vlBPqiia0mgW+j4WpOkHML
DhtAmGnc2lxPmquNiP4LvNNZWZfNbCP4T00ycCsz5ITDTPZ8y1XGzeqSt3fOt+aY
Fw/LUmjmyuNIKA90vbLOaBiZg8saUsupg8O/xv4R1SbUhgbNK/xdisn/QAcOjgz/
UMkDQ8MbV/+FViY7tIbHF1KFRZ40YFh8bA67iXm06An73cP5F1de/gROU3jHkWTp
0Bmg3y8Vwd8luQuHAg8yQQ8qQ9z8XjplwB+xCpGEduVEtMxKcqgwM7pXNQkf1ZXl
fCNQXxb73Uh2UKUMlNFmdLxQ/MhVxa1RxtnzmBQvU/BI54rNm/YnugpF1YDs1gtt
I09DEnd5QSetleA9JEtC9yg51v48qzhIBXaV5D5SzSybkwMzJY37g7JhJv8cytfp
GHrYt8f9o8ViLWUdda1pr9pevUb3jfl32b2zjnBZcPQ9Qw7PB7FkWnlP3gDIDiXi
FVrzDelxxwWkHKc4cVWV5/GarwSja8ckZelj3WDQNfb8tf8lsCQ8GGpLCvJ6Rt4M
6ecXYOPH4WxO4d2HYETD123Qzeyi8MbIKXryDyV3X4Gl7lpokD93B/6EsIbpcWfj
Pp5ruT02GfOxhDIVxSkh7wAh+gbthAEIATrGffhDixeiXFuPj+HIx0A+UCAMs9aP
kBe+vO4xV0HQEa3Lp7GsrCLXg0EELrvzeAabAoA6eYa9Ec69QYuT6cXnfYYq4Kk6
RTbm7JI44GuHEW+m63BJTLnSETO+zl78zKnqDuKGU+Fvd176tDZrsYh09qBZtoXg
T2imGwuL7FHGEMbqUOZlhHip5lLj7/LkzOcnpks3V89orXazlVmEhj/1OqBQkivj
BEWRVM+6ZGTnB1rk/dx3mAUmbCoFAcQmM77XfNmVYcaLqk0fIGPn29BrI4pjkAiN
9JkFKU0nLXsuTe2MqChEEfjJ3MfhHiWh+A8csM9Qez4wbVy9tuOlkjOmZmZxPejr
lZ+tUqJJPul1mYrXCzs0xQ8YUSqQ6mL9XWQWI+9lfEV1yPgNAj/O/xDgvM+TyiDj
RxUlZ/bPCjVLb6JOirdRHL/NRQiLwlUgvBh1n8IbAdHOffG9dsKUoPxRxIyHez9z
wX+J8E9+P486HInxTIgOaTK6kPBH2qd+Z5Fb6BNmbeA+pn8ZzOO0YOj7wur7HJl9
XbXzeaGoeqsNVxYH9M7fLi80mpqqqdnam1wpLXy/U0ujDf8H1j4In8nqEkqzirni
CHD3/jLFR1CwTAyxcKjyWp7u/dWx/Hb+Kut/7K3XVq4wx6sEvrKR8S+71rGsZnCe
N6zMTOUHgKjfWfROPzBhhDABmt124bMhoKGw4mW9ly7VqIqrNTWTv+jeWxUdPV1h
AYFxgrAk5juda+r7wkkVTuG6aRhoCww1B5mL38gVMaA9SNgqDH9vC0JiA2M9vhsQ
c0MHZQ3AHds3Q0jwWUWvqu3T6oqOaPlmpwj/xL/WkwbTwO38IwhrvaPdT9L5SRwT
aMrZNOIjKdRim5Z9rJlpqTANK+wSCmn6ITZ9+TdymDu/nKRZ0Mee76Ua+rn63zi4
X7zlg28bCaQM8zIxducQ2IlRnHq+uc5O6En865Os357jwMXn+rxaYurVEqz007ga
P5Z7ibKVQ6a1buThxpyFoqM1NDD3FxjQTQ4bRgbayJm96+QTyeg4WJJXPVo82blI
VHGeLI4aAmOtl8iIVd3gBBaoFh2TCNBCwSRJWgcwncRe7wsnJkmIRwubAQEoLJji
uazcr0Dje9nPbC81Z4NToqcUueZduAhL87VbpDrt4Em4kip2RsSEzFUQrEX+4Wvm
WVs9eUZSevlvQUqp2d8Mx8QNQwSdSjAAftanNCNncjRot1UD3k98ManrmQ44Mg0W
Y7htS605VhJIg8j5T89q55LExRiTfBM8pNKMTZ7ZIvdQhY6NqLqenl8wCvp8TLsu
DTFDAryYL/jFqUFSQb11Y2FAxt6lT4AvnfavFoxpCLyXioJcLQKQ7+UQOEn04xV+
HfgJvNAN6bIkn2FiY4jaZUzd/qVzhtu0eJBRBDDZNOhEFWxNTPCKjCZ+HtwloZJW
Dm3FSEDi59z6BsDgsz6fScc+lghCq6+NYKA3Wx3FTWShr9tI29rqJ37lUouhVMBi
6/NsrI98OuJUjh/cQr5KNMmmAwMBSCYYDZjMoUI/sZTuLzcqNHNFy5fsNhOP4rmN
se6LaVcr+PdpRD37X1u/2QkOrvP06KIlMLMm1O7dU5dEHhsIBoSbSCtOp8w7LCRG
h44jSCySCytYdwKSGLms79rlfL7IYGdzic8/pmmnvBTjQCSUV0MoIAKRaObjWK2E
EaTwXPnURgwZ6YBwNNXab30nbXNT2JTLAh4BwDPSeWqtfGu7mr4hDGBc2LCQwBJ2
RZf57zXpRozE2wwLGRnZhVwzpB1SRzzsMuEVI/w5l7/YZY1HXwznNKaEfzV4cgHb
SeSOtDKrAOCHEknkvayEiX53tFz0L2GHYhWKf5rPLnmeFI4tmx6iIMjjBUQxL7La
/s2Uthyq+DEabbmh9TiuY3vekFTpn7xvemE+ef+da94J8u3EJJrIkJcC8KBcwd1M
SRb1DuAwcVweB+s1QHQj1uEOkusk146b3U26TOCLdA9TsM5P+BE+Vw/CXUIJJCdI
Q3IUT64H5tPMI8EfYV5Koc05UGsupej3hPlampuckd2It/LHN3ca8n7a0MztqvNu
EL7u/TILpSFUUyscWd05AAN/SUy6mGBX/2AUaTX/VA5H+IlWhB1B+iSDvSfwHoMU
T9sX82lGw1oeZehDHaHlno7xFKnsmsoCAV4lsmLwsIEpLvLp+tamtS+1PKRMBo8z
/bEyLqZYgAg2GU2junXDqhWTk7kmdAmyscU79UUMBDz5P5wjKL6nd3AQ5MvsWNQ/
lP8+sD3a7PcUjDxgjXcCthcPjjjboto2WcWcC+LdlE7sg4R8VIgoigbTB4J2nWyI
5GuLG1RDkeeiqnoiB7jX2ouBceydOT7QmIrt44Ha/OM2udW0OD/79WJqES426JQc
2Qa12DIC5aGaFL6G0zCCE6QLaIPSRhEQZ1lKabh4PGabv7Z8f2gsQGXSHxUdrNWw
MNYyOb7wiP/TWYiEYgP6qoApOXLiHRRB1ZdnBhNCuFLUDeNREUzRKJrci12Lv6my
350aecrUqZeOqa3rhzS6ulykiQIlLTQfjF87BKRJSS/A5tpHnP6RTombval2SHwi
cODbqGMbjETKcRL0PoKHPD/aEXBt2tWR7zm984XU2OquGRQePiopasPr7AGSzjvU
4Hl83N6MNHlII/SPRWFerZ9r5v2tk2aP9eLDth72QsjmeANdAs9GyoGko5SVzAoo
ZhZx4WXmnXpulccyqeEGrE71Q9p/TWRaR0rBIdmUuHAduEfoc3+/eBWn1lth2qGO
8u3wnNQC9Ov+xsiOkX0oR6yKfMj9Wet0Kymn5vR+bE13wrg/iCVAmUbAbYps/QXk
TcjuCgRZonJFPEtN+Smm9ICu4GHJuSNLsm2mQpy9cAHSxuSQAf5kponS0f1+Dx4j
nYSZHGyScQTTCtn9MrYB//BeNUiCiuyfd6IqUkQeFaJpnDmr/JicLR9ru33rmk+P
Nr64d+2g3PWsXOrNCKloofxVf0iAMtYwUP+sX97p0efHrqQw+aMmvK7OtDKw56J6
gyCnU7ZyTY7XwH2yX56ZfcQsghNS+BNuIkR/Spc7ChRswv3xtgvntQNiyZaDn5eb
jVLLBTUN41hLbqFcfjO2mJeBzRd7PNPlfTnKHO78LOG169vMcE8bLjWGAgN6G15S
uNY1bUhLbKN12f3XmiOyb26ZGstpl2Gy9yaCfb828myPLDNJliotpyCd2IEbSotJ
Oa7gh1GgoV4bfHKW1hqmD4IJg9oPycqe+hn4uSeK4Ahve+5cAIEm/fjDmHPiLVo0
XPZXhWOq8sTksPZhPuAsXnJpqwA93Y89GtjCF6sfpmnm4M9D9qCVbphjFR6HjlJw
z/1fV1wrQagcAt1WUjWZ2UpG4HrjqeOyfoUAsdbRbUYGFegDKCmBFcUJEP4pvfMr
aG1ZtPSZBv8WLpoBVB0xT25Fm68y/u5AL29lI5um8zIeFEBrnxAyOgrLxMDA30G9
NdGFUjanFY2JoDkAu2CoggI+FjP5T7GSGAJG5XQbOJM2gRcmrY771HLYwvmmYv4e
0lQ1NIWcxi41qwuOT3IC3AVjWOi20TEEsyyB2yz3ENghI1bHEd6FgzU2fOt9CJ3F
YIOM7fZsSm8vzoI7wm1FTxqWAxNW/a7r56myn2cLlp4Yp/+uBz57I1bBtrL9UhCO
BilzuAcdg4IRFz7SafQJ1ofWRnEMW4+dekqOzJPhquZCWBFIFO7g4hagFaak8Hbr
P+NsL0fzD8nEZZYdMYPaMhUKeXBI7vkS6AalZgYkd06kqIeA05vb993Lduic4qV3
Nr18GVKTSLAd2HXXNG3uw7bYL0g/GkPK/1sGUrYfEpCyxI2Z0Awq5gpcQQkWhDyj
tQu285VPgSoDjtkmWqU5qyVFqGUnrBxDMnKnsDSKazAxfNawf5oLUmB+zXbxRmzx
fYIXGQUEgor2eWBb4WWp8xXrPqFCXH1Vuaxe2ffQUsK9iZUUQ11AkiTZE9xok0xQ
4MzD5tKWs96+uc3oRy1DDWThyCpKwlCxAHe7GS2GpfMpaJNbS6lVIi+4GimzDUlV
9mFLkh2ZYiMbZCiYP8teKcTzdbqBq/aAotBpsWRRVxqMqe+v2ujqruH+Gm+7yigl
278PFQ01BkAUHka1yatpCJ2C9250SmI2HsCz8woN/8kkkCx5LRVexiBIKFK1HRWS
11kYMVF77aIL/wNS/Bkk/sf/Rquu4LDUaRDHvlS+QPNC5XENJPkextlaB8fJLMhk
qfzbb3FEDB58kzZ+1rjNTSCfyS3Ev2H6REWLM2GYoh7CQslqIpF9zw+2XYOAoSjw
mXC2LNxTXB7dQYBhrxqdOfcPgBd1WVD3E1XJkbP8w/rzFuxtffuLe+aSpPtsEq15
LqZf/a4z03vbkLEJJxClien6jr1G5mv8+ALdZkkiGnpCEnjb1fVlzaPCGsPHHMTS
B7m5dfyjbA65MZlqJllvfumijgMI3ddb+YhRRZUAtG58r9JZF2pLyTPYqoR/8k38
X+KEAToAQBB2S4VSaO7xm3AG9s1syjspNVMy0vxnJLKOvD5mH6L6wJxt2Vx2w/fL
ac6DNT/2hjrV4xF5jCY0NneIzNcTFExZlT4Ms88BMRxjflMD1Bz/ki2XUMYY1mIu
msAuKo5dnznEseDyoRXx51V5S5Fb34TVnr8MeUjdIVysiO0Y/7cE8hKWhlTMEJzb
lG3pYSdY7VQx6cY740itmiBtm3nihOxCjUvx9Gg0h+NTd2nHwKLQQtXMxqdFHqsr
U9E7HgQMKzJJy8UzlHnfc0o193IQkKzQaVlm5uvJUxf8HX54dh6WvDzuMQ/Zt78L
lpQ5ZOIwoy8wZl46Ywq/r2fpGVd/HpaJS/j5/KvCZ5OmvzLy6M+bkvSRthFeTnJf
s+0uEbJTAmBZHgRkwZZbj2RK9MecWAFN4Az0f4ki31OyT0a/bwh1xq9LKgs+L+Ql
kNGsD2xgUkmwYj2lm0KZPCqJHG/KPriW00+vwEZIzUDNi/ToRvsOcDVVCCTBQ1qa
gdHNWwqW6/7F5mYKI4jvbbGwXqZaO2VqWcJIPHJ4/mu0ax9c/sMwxAD6w1ZNTRO9
2yGzpll60/Y9S0GRemWklZ93PtsqxXJpYEYK/ZNm59wX01iQHeiDNoQ77G9quc4c
U/HMiPT/aLGzxzH0DQnqgY8r7Y0S6GI8G1SkHWydzCtR5lkMM2Pocolk2LuvDTgV
cj1TaoGzmAajhLvEHh+F/bOF+UybVQEZZ5ANdPtLELge23uhNijZN/Y2PEkoRMCO
h6xigwne+5+JDsI8/oMszdDHqO8UTJQIayBLztpr+npQD8gAaYDIZw2dMUxXGlJ+
KIMcUdsTEVSysQtAwsIOhetRQxzrlxHj6LVg/w4jVkktjdV5oeA2yVk3BCbmnUtH
xpTBGdTQAP/qZvlHmfnr9IhlxDPQ9EgQPxdeVqpcL4u9HSr7U1F06ziWFhXMkFri
3LJDMBYE68+rmCN0zsZkPccWHUJBNJYkSJb8pbPUM7esJDAkCLyHu+CqHQjSg8Hu
fgDTxnusEV7gZfQbElPSz1C9TaQAlAdA3ge2QizreDpxUapvRDez/+OQ3AIHGrsc
ZZT9NKoPKamoOJyDSfy0Y5KoQx0VV2jrN7SrJh/vxOxNPs4tDPhhGOXJbdo5p8gD
+aHV3/uu8q6KzZj+37v1SNzGPYBTzYcTdZ/DUsuSVbtg6qKm/WH5B+QHqe1ZtkpV
Dq+cSJj5Iw+yN5Ja7Mst4ut+AgsQe1n7i03lbAjq7snIIT5hZ/0KtRufx5dWCIpX
QWWZpLr5vHjZuxCnV/49u+FQJ4AeeydBKrY4qrnyN8tnIl8h5B4hIJyRdCk2gtmp
aIoR7FTPmv3GsOqD7iVoiKTRJKaI0S3FUgGSDTvJrq8IT8Rn/43RjM41kv6Mnlr+
MeJk6qTlvG4lr7wWRMXmvE4J5cWnhwlL4rw4M9iwRf6lfhhKrNHBekDqZ2W8mq1k
eJiHbem1xYtvG9drkgLP4TrapM9+gp0mCFKOgP3Vcz8MP9AkjgFk2Wo5e+pEcIHn
aXy+kpky5AI7G1Jkh1lVMmIA1kxJEbMHBglmLtHO22hKk2Uo6uUtMnVFaNZC8f3Q
9iW9YzBtzUJ0lxNQSIpBiA3JenirlLZO3TQSbVJrAgY2LZmtktoCR45L7EWlSY/1
6oDGKeJNBATqJL+SoJU37PfImsKEuTP/tFqLbiuEIG9TT7eI1PjnohWcOnTf/1lJ
3cCjAoTRQYlUI5DwnaxiaaIAEoP+tf/gmCw0oM13rhsSFsRso5+0gGW+1r3Xx/xp
xZkPld+TiwWwMQZP9bVxSgdC0zwjHVJocrABEqI94IeFpG3fDUWFaYi6UwjbQJNg
Kwlod5Up9vBsKk9G8nlqgEc0WuJqlgHQIrUhcJ5JhDRsA0loDOMTeGPFd8n/tHG9
m6wSbEdXGrUfSdsxycs3q664ajz+Lz+3OxIa5h0VWZFozBXf0BTeJMMtFSFjE/rL
EpB5ufzvdpN2M1tEoY3WF4abIfvnk3JI9exrQACMSuzzjblQAvaK7gewvcR3onws
4NLiRNhJSwXVAlRxrKGCNnSsBDprEqOa6E+lXXk3xPJQPTfc/FM0dvO9luOXPT6D
18VUpsK9xr+IFMGS1qlsPxXDgpdWhbd95QSFqQSg82gWssNVIbYEArh3iFCosrMU
assDwZzDnhpvFaqUHi1lKoyItVLIr0R+VLGSWLXFAHWZupxFopD8X7nDy9CYqrpK
0YFVnHbVuemkw8u7FrobzRQcXuUPQet5BumropUUrPiYAPHxQjnntFWARyxs2Y1+
MLzDku5FpCnrIRrGalm8leIx9eMm+MpnJv4MupZayHgi8ehK6SD9zmq5VwcDpJra
glTJPuKZNhSstSVCfYnjrb/HM6yGKBfahGD+yGCRLKOlMhoj59NNUIjDccaFqfm/
qf/n8wn8YBvvTzx3tQuW4Cc/TEd8Pbjo3Nqxq2qlrCsvmUosqqN5c2/IzQUaJpee
ykLgnx6weOKj2QwoxoG3bZFnmyu3AZJxqnaFATOIgZMUrVyGP26WYj3oWOqZcDo+
RFLTJ90b05JmNvr7Poo2gW4rYZmwELFy+EExag4jEv+JLVZttp1GFWY2a2MKeBnC
4TIolpL9SqfYqYAxsiXPJQ5iFa6JFrNWJjC0pWBgTgBsBKe7LYqODf0Yxzla291N
wD7gfMhZjDJ3ygyOQiM9TDTwQNqeHW7sJ2/Hpc7mn8K1ctWfnUnAyx7GbZ9xbXBs
e6L09voNTr+g6YNN1qwqGTMPdV+6xPT7CtTN0Z9DnLWm4IxhNbNjM/ThJI5RGxvN
ofx2NroRpJhnty/b30uKonR3BzMTJ8Dt4lv2Dh0AYpmRFMrkRbKPowU1q8+8drvV
RsUYHXkk8E1c95zYIN3ypMBoLznjqeRbw8F1ftoKTE+uiBEdAU3ZbJtrzweoFHDn
ep4naUOpsbpre/St4gFZQ0Hb0XbK8T/HycwPTb+l/42+SoG5AK6OuOPHl6QJq8T8
fe4lZfX4rnvn9afwHkiC353kkmTlVQZHe035gZ1ihA+stJTq3C6kzOPfzgzamrc2
O2RE5NaSsydeTw7d4jwTgP91Y4FSLGglId5n9e2mptNb3ufD/yt5XisV0uOblESI
Kl23TPf6l9TKj23nZyBa9PvdBIuibKIzpyReIRm6s8oSysdy8MXAOmc/odD21lYE
5XqXCF6IrV1ZTp/tI0h74OlURhTY7XR+omG9gZ4HIL5Ur4/pmbHaNBX1Rz3wP9Es
m2/MtZ3NS60FGc24+XORzo1ODp7CGcNFK+0KxfCzUQ2sts6NCS1rdcRjj/4v2/5B
o4QopV/3mkWCnn06NlQG3od/gSrRY1iuczSjP7AiJ6PlgoMW+aODX0jvhSUcvWuL
wmyP9BRCOZURrtADjqG6Usb8YK9ofYkicY0OC/iXRR6979Mo2hfR5PxmDe5JRQct
x8zrou+FRRFDecyzXZfARSNZbTr0WXp2A8FPvVTmVdCw8RgSkMG4IXL20o2R1NTS
bn+89DDvkClyhdI4CzrGjhTPET1xtVu/FWdmp/DOZxrtHjaO36Bl7UP22Sy4dTRd
1Cpr96p88b3wzTf6ZYslM/3qyErD80EKYhaqcqb9mhPk8gCy35vzkkZT9mCi0IJ5
f0eUzfD6dz09qrnuFSGpMNRXkPZG/zJVXz3tbD9fDi/l1+DSES+wMtTUeEvUAjnJ
/wJ2jMFazY9qmhx7bppNP+JlDZAEVYnWE88AVD4/j4amohOJtFcnKS4JbhrJhPAO
5R9CvLqqJgYJhXGsyNSUMemUbV0WdB3i2hL248Uud/cfIlDLyj7BcQyWlVCqydiJ
rMPIiokIYTU7tmClmoZnvbt4RAUQ9PkiwZPseNXf6EiyD5kQOQl9Lgjd5xRIBVdh
fKsEw1KzXfQ8tjW2O+DOL8CxxQPrSxdt9Zynm7izvjzOaSTJkZst5AveJY2R/lN6
qUUdYXURm+mf7u9dJWX0sh5cbcpbZAZSr8mCDkLIXkXCaz067rck/sFxZnbBYObL
BJWk9+m/rLzgI1e8Jto+HsUET8qUJJCoPSM+MZOu0eS93bZqDJgYUUEa/hBK3V7O
uYgGj8lko0YtR9isd7Vw8F8+T5FGxzsCUGcqoLXk4jW+c/0FA6lR4Pl1hUPSW0Dp
d54dmpXAVOMEgp5Cxw9yb/gJaX5IbrjITJeMUlh4jFPg44ZOlhM0/Me4XrnJdBoV
GG6M+C7V1+CvuZZRNDnQcWa81LNQ1p/WyyLCd3Kp8niL49pyR6uniAJvtqdTA83F
7odqQk+esXqk+Of/5KMKIDl7Wul/l/H+2ngaLW9Jy3hR9j4kBqaZPsH4X8rYdKAb
OXXGJKNb5acq56tapqz96pkiOFsX3eCe9xLnp+RJPOMJ7xjatIQ8NT9wyvwMD392
kcO0OSgpWmSHsRwxNyaOFU/MuV30HAMANVAvJ4z6OZT5N1PfCti17WH1A4eEDfpN
wjcoiQ5vHkLVFSzSdL1y3b9A3O8ie7EMTmYfPtXHXYyjRHpK7YXT1of5L41XWYey
dcQIuVSdOJGwpZm0tB5jbFAr0kbJH1WJ+DfOB4fDA8M/uu1B9VN0nE/xp1Fq53+9
T5gluX7l1NxE29ORlpsNU+WfSeayoLPO1myyZqnuBoNyQA++KGMQNpkjGXDYDxHp
BaLJoYG+oetdr1jKwCmUbNfK3rOyLJIIdGeX674jMtTAoKxE1RzU6OyWz2zsRNR+
y57Cqx1SOckfqPi/6yEzrww9RRTsvS7a0eMTSKmu6mcC+tUbQgUVh0KEKeo5R5ZO
wP5sk994c6E41BSV0XSoasegqQ5iCT0o3EYNwobsfXcxltlTu3XqP87Xuf1CKniW
P2LZcf7gjjKz8BOYbQVbOy+xMTOZ+/L1sm6k1TZaIRoywoCYuxEGb2dPUPBMCNA1
7OgB60fKF0Mch1/UumYtMTbq6anEIyCkfnPdDOaqJe2uqre3VGlbyJTscAAZLQxS
R14jZgkc1HQO/E2c+Qcf+bNOx2ZvPCd0+aHSQJjVJCq6gkfDKGO766A+Sb/jIJxa
3tyacgh3FNCIoBnbx5iis+ovwRCLvvj3lKREoYPBfppuX68r2OHdc7jajgCBo1yV
bMlXDmFLpJNj+lY61LcKjmHxeoIk5R7ZAgNJreak8jrJ69OaS+EPM7PCsYGUVKMg
zclirHkJT92wViQFkVH8mW0ZhbhQXy+b+dM7tx+WUQliEdWH/MC/cnBgt9jYeZQZ
O9KhRJ/pStWA8jZbEaQYBFFr4tSw/tkJd9I4Qjb3YKmSpPs4WmWrGP9tM30k8RgS
EdjNoLbuIWKkwg0r9gTeWkzM+fqaAJA8EhUi55yOAfybBg+hDCtO3BsTwTQvopo6
8jPdMUHrK/y45zAYqB0tQ7g6EM6FoPaXdgpCpzjaOk+if0MSp4/S+RAq2tuuIxts
o+bcJ+6YQ4nDrdo8StMCu3Avg1fCMDR6P/ODPb4Hzi21if3FI1Q7zMXzfv3KOIlN
Io16IFXOlVn9EfnsJa678YGx534hAoYHGMfg/CKtj1SZ8i0xQL5OPmdJWDybgEdz
+2O0ufMxg8dRP6L7QG46eJqQKmgN3LHwEGIS4ohKNHWAhnlsxFFH65fUAD76EBjY
mdcZFmv7OUcT4wOy0zC1uYGzueuqwhi4caip4h+tIS588OFLWfJIqeMw75c3yHuS
2QFF7J4pgY/MPgfJryZA7SwtXr9kqT4xYCfl8l7n/Eh8ZZE73IhV2g40cCnR40fm
KB/mI1XGnFlcd3jXjNmmijk6TGSs3Zhf0zoYA1gpDBvhP8OHq4GkqazylWwoDYlT
V0bT6UT7JSvTNhJSriemfTE99HOa76yjRK6p2rfiJc2wcPmjAyXLc6xegMh1X6xc
3lDFS3wNGMSg21PuBsHFyeth/4d5JIflcCLVkBSpbIRVoHTkTGy+kZuWl5zBmJ0+
n0STurpj1UCf1INh8avKOGVPyNARWw5TSVWAUQlhILK3rKldyeFHjNhQalwNgx+N
9+5sREWvoPfmwUnSS341QpAskOcuVNXwwrKZgeNXrEK8dQEjrxUDlEjNWY9zDU4y
t4tlqmxdxFUEQsPSETl42Cx8ygzjM7yLB8urLSs4Z+kne3+0afIdbmhBGNyDn+jf
ZSnx1tOAmbqtogtOoQXoYF78v7feD/DZ4KfOKCFnPoO+4acmiCCN00++gR57M0aH
hPRjNoQk9++SWRECp4v7tU5k+632mQlP83U8I//HMHO6kf+Aw6Dhkp2Lk2T010ex
Wi3AA65Lruq/ZsuB/7J/4k15KKGZQuxW3MXJ8Rh1g7k83zuPMe26hIOfW/ty7OPK
ZHFMSxnCHRCAyO71mp7+vaGLJHzsjYwc8chQuVZSOxLDk2UVhjtJkW51WHhtbtFF
neW+WKPKNX1abKt2318qD7x6Lg4fwvX1wxdSErDNykU3js93yG0lo26K6I7O1Enc
fImoN2/9NZulatB644FY/hc4XTjB00PI0w2/Aeh+Hb6WN5IcGOHoai/TCyUboN+K
NrBBEvUmPwoJB6ZvBu6nkJZs1FDPIRcPa3VzEihO01Brl0rM5JL4M8hGhT9xOfmh
qs4O9Iwi+Jl3HGg2NZqtelyRrT7S92wg3wA4BJkS7a0KCjBhQz7je1eth5c43w9M
IQA1i8K2CIKVGOyd8Mr0x4UKy+fe/lp4zDwylkcTlv7ETdoWtcDM/GigVXlxA9Ky
sWWJk2ycaWnUzJz/FEzpM10EE5JYe98aS2ZfmLT/quStvYr9sKN5jgUnWP4FNxhG
3RJ49A+SHIJN9TNsuYfg7oLyatzeR5DjWX3Nfm8OrI0+c2xfx4eXfxfvMMdbEwvY
4cK21qxgWd20flAgIxYcpF4Ab+X8BXiGGCgJ1wZB/WrhhC5ST96c3SQvTNEuwvya
l7gc72TrBkrRB6O/UGk3GIQ4o8q82uS2Yn7RwQIPMFq21gPopTxo8YfT99G0M1+Q
I3HBpYFaos07kErq02GEqM9sgOy5dAmxmNmuqfsWZE9Ic0k1Fb1e2uwQSNaaSraf
EQlU4fEhQ9QzFLCgnmcFCrs9VyQ/ZXqw2kVp+pL9ZSvIK4msu50H9GOQ+ZDaXuDO
gwUpjPrroWNgkrbiFShdezeOzFOxukpYiMUYxbNL6mN5xpX7vG6nXRcTuI6Mf2B4
rUVUM7AKEXo8nAfNjKXxv3hB8JjIiWpzWsuWwRqwBDY/9VqvXyCcthfVD7ePzggz
GKq4bbvf6LJfJUKS+RYILD4KXC5scHbdibPNfVoP1KkO2Ekno7+eBiEft5YhD2hF
POK8SUFk/+YFkbRiWXaPKy9lIfxkI75s3U4VXovRkmva2/oeo8p3HTc32Sr5nAfc
TX2FOEPFc8r0spydxmtg2glm3E+0+0ZCjmMZeavp8Y3yDXyGtXcL70n6pKGwGGON
f5+pDNJDAU0rJaYtxMRvaPSKTqTswvbypHG0Nuq18GO8kaZ9mygP2GQYdo+UFZW2
Z/0d8hJA5+uVm0mWfDk6ma2rd3le+jAW7BDwciVHiSDpS6/jRgijfriUCCjnLpen
fsgKFRN59pf7Y+EjPOgm4HQJM8l2s79S9mmMC4/DJ84/0bnONM27bdkbB6QS5f/N
Q/Yg/D+ri51bEk9GkJV8RHbpBo8TrSBhy7gzPabObyi4aoDoOAe2FAModhrtEeGF
7abDbxUShVVv4ai8h72Ubu5cgcjmOODRZ6pypYYd1ZuDUzDpycrMtA8EjMFGYFrA
Q9KLt0dO/YSwJyJ0lXx4k96QQ4lU5VFKxuzpaEWHeNS9FAJGmejEGD6VyW8qVD5V
v524br1AI0ljteuGgM49liO4evNdAmmMIQ0w/3aRjmkprjuhOyt0zkLNZOuSwrdW
/cUSdfmH+AfSR0f194I57stLxCeX/02dPm9FpegSJ2pSzaAM7hNpsWaWYd7VTqAO
ydKhNbQQOE52oPimcdq1G4ToC4sgF7RqO7fkglshxpNHuCTHk7j1nz85gbWRq/AL
qLw1lX6iubda0evx0Bdt8c5o/yEngVGiEjs+ziqv8ARuyaXGEPe923ivcVKNGdJB
YhSDJGcOJvr2fAxZhTxfLi8xzpVZ2KDv0qwBgB1QBjdnApDGCV/f1MzwaD7RjWU4
gIp6NJ8ZGSOD7JfYRfaGY20OMie+QKXeFXKyMC5aKreRr/wnid3Kjt3LLk6yiJg1
RryfAd1r1Bb6xmcuIoVQ5wTA7BNVOzl9L+U/oz0iRi1onF1Z9x+fiSwZ9h2s7PPy
RZr3G653lw9tUcWuPyUyYSINI2gPPGoiHTgDi2W6elkWV9CQIQXY5kmoOHFPZNfh
LANvK8TXpOSCP2HL9024CZKZ+fz6u2pKMnXgV8Zic4P8c/Slj33oV6qzQU9er9DY
c09Q8sPP85dFDEq9GzUF9BhnIMIBrOxOCp4kOUExG6we9OS4cjCHMgl2X/hORPvK
O8WGC6FhtyGnoBP+AENTaLLasQxBvoSqwFTd1Rb7eUaTgU/Dq1yJd/zewYCP3I7a
9OfsztlBFclZH4fmPx1mpDP4/lCKgmFkuncGd2JQMfjZDVvZ8CVoslWl/7f/692A
8aaneeIOh50VOTnCuRBa43Y/fvruE4OcBg373sG5s1IoLSTDC31ZUn8JHkyZniLK
iEVmcGOvOYWhkbH+OFACi7R7ZNeLdxHDU53ys67LEKxguB9XOgka9Ff5VOns86KT
nrnkPWBG/V31v2/84UXVChw78oJDAzTxRvve3guAQxVzC67gI/H7WF/HM6E1PJn8
pfL1vch0xm94k1+xaOiqOsShaHNvYnB99jobChQZbv7Yn0nW644Ovi9oe1Mqsc6U
ZXp7dKEek32GILjkz5dTFtmBRgc7aXWyOczKRpL3LgDX3R4O6rVfk9gIFovN1DZY
eKoAS/9KE0oj3XiD8X4Gk8Ss1LwYiBN2KCoNMrk5kaEXYDcWdnWtwHoMjADlF9un
kkbSaBXjrpE6o8e3XQICEEHgYLZnIdVKKKNIvfR3IRl4D89PHKWHlBJmZ448BXKR
RKXKpJwA1moaUwbWT5yoUU8fDzYUn+hPAw2yhpxyZJIEm5nA1WpimGhMOOl1RRrE
v8Neo2aO/zGOWMn0GYG8y1hY2hC39FB+rKU7OrHK5EW+OC8M5Tszrbxgd3eDSai/
6G96ua9TvkI4dwvypgjlNAZYwvw22MwyGvQaHOmNB+h1P9Z1AKXkeKpfmwukuKT5
AbuXtGdSZb2BzIQkvp3X87DKVtUgN1EZ24q7bDNU9foAv8hCgSiJkR+IgtPNqx68
VdVoQzHCeQpcfDVGisK3G4WTNNNTUVgb8HgheziSnHAFuH+YSrApzmtTxLdR/Zgp
LZpWBAFVTWqcVx9CTL0tZkkPNOa3ga/dpImTSyOAvFhUF0ZHFo57H7dhswsiEEJr
0KbjK5mOBF7wd0/VrkdI3lxmiGKt3O9xhHiwFJCq4kHAGXUucQXBBJqYvYQ7Noto
uC+GN1Pe4Hti55dbSaMW3z7CyFL/TLUQqb1RF6DOx41kJWJMTpu7wNOsmS8S+fRG
O0Dw6YCYiIcGhc4OCyQD1lHtgepRRPoNMA2IOORnS7wWUhyJk7hTb6grvZ8SgLUC
qJptUBEPjKJf/FX3wX038sX69vZpEiW+w5XkfOsZwoJTcrnASNvE//yZjlIePSiZ
aO23fereivBQ7OI0mpvh2j7tiDabxqmxjKQpQsMAUEsBrZte4NrV/psIBbIzY1+R
g0NIrA63DFGCnfHqN2dZi0jMQI4/gHTtZdeCmE1CHcV6Bfbfo8ZzP9VmoFrfNSTA
39rSiY2swYDOZ6dv1dsyFBF6f7iRAMGjRMqi6Sj5VgwzyGqYoZpL8Bha/3a6k2Ao
6BFYvu23YkE3X5WDxGUqbmsJNb+PSFCtzn3H4fVVBfFtCG4rnFU0/wbevZ6m9NJu
U2Eu+r6jVJII2b1bhWlXZdL7VgG/g0ryYpveWT9E2DBm9H9Qj8ecMMgQj2v2FHUn
p6IzMh+LAqKw7lHAPh0UJkGEiQ//LahTPuyxn00PXLSbnwdGunb0h1SsdvtWTuxx
Fm3mrEE5p6zfCnPmboTARqVxkEMEL5zOoPBZug/i8jIaz6r0CkdY+R65wXR1Ibf3
Dr4k8KxaWB58i+qP5xadjc885Y8zkSz2AWpwXHogKF6JHjg3VD5ASk6aIREytag5
B3XnywzPl4PyEiU2YFYPKnoirfpKZxQ7YaNzEMZF36bkl0ASeB0n2lztsBguP8NG
zl5IjBxHuw+fJUxOizG2Jw9gE3v+xZRAxMSKxQBkK4zywUa0TIpBMARfKltp3f1U
8pVSG//ld1J5YFC72donyA++zyy/t15rdrZkDpYl3vPfal+6C2NmEJL3lM0BHZLu
RTsWTkN5zmc4RihPo9HzbgXu9RSu2YAjlmvZhnN9YVouEsBGpRRNr9prCpG6FI/3
H4qmTQTP1kGdHsd7t0+0IJjmUB/TXIp+PnWZvFK6P16EnZS1C3r17W7HMnLFJAvU
5t9Yyyq1IK03oXtmVmFlJp/fUhYQOlx9A1WBP+57Ken+1oospP8RbmEJVZZbNm9t
FGJLtGzDEZHavdH+Xn3AT892+vTnNUyn8cRqX0Qi3BUs8hCFyAK9OaLeWUSZMQj8
ArlTpe1FqA1wQEnJRb+u3b8uFFOAFtAGCwOMJu05PNlgKa3VvHl74uH8e/dizL5c
cZun2yOHrvkvIDB0a35z3pAOgMUKbOhuqyvyamNGzuzJMwG26pHKXlcOveyLQhNO
qGgX8eHRW8INjwmXPyYrVArGeHySB2CfjvhelYihpYDlYq8tDUzrrSXjrlxNQr+N
+VTXz7WtqhMUdEuN/LIbgb0oug0g1vlsNME/qZJf8v1w+WLoKDlfRNANdLSf0dt7
FgyRU+96puiQgEgA8cAPBURYtttWnFu2BN8d+NUafVnbid7wqRC6I/RiZz3zJ1Uy
bwAdLI6hz2uwUL9X3AvhT3NzqpBsN6lhXrZdW1RA4vInM87XOHA5QT4TeRtdLVhL
ov7KVWgjtCZik0GusSnkRFM3atQnAvudlx+vMC+mrMkWx8ajOvFqhgKWiT0iOA3w
DsJ4UZk0V1BWJZN/GQwmwGZMTbLgJakfW7g4npPeoQRjzuCEypKeEUb192vvqlQk
TjIVuWHglTGkjlQgsIGz+N88s0LWnlxgGJcwgkjYzb57gy4E+yI5WjWr3LKK7VDq
pO6W7pb0XGBhJPB4pEabGY1dc055mPbwrQcagYNjrmPEj+tnwfXVDuEBEZnnXsnv
eYn98L01d8ucabXQxzvoC6gZ8BcXaGOlGJxIqWDfbQ2L+HcyMGkecK1zFD+sKWUz
SLqkuasBEKkh/iighbLMs+NKhZBwHe+VfHzbUVytn6kS93JuX8YQxsRvAlRC7FfN
zsNL9yW0mjJZLCexL1H0GE6CUXTkY6o09oqCIEYT5nhQnqegtxfoWnwMTB3Gf9ca
vvNxQm0k8QtuonBZvrrWNlkEBXnNGBNZL7ex0Ic0gTAnO6a9zy0W2xtkplJDQ3TY
PBOPww0LM0xyl8zlzJjESGxdM+AJiboVONDJ2heY8SzEZRukDqQX4zZH+1u3QSVw
6ILZvaTGbnm96bMjDRf+ZiBvYoySX1ouZxOOYmDq47zgBWrwh4yTjG6J8W+WfMkf
MCY3x9yvBAKOnyGIXLmcgl92yrCyFWzTsc9wAhjQoG/ANdQGpyuqvKGk/kAY2V5+
0IGEZ6yLyA+ADR4hKVrSHLEasZNSMIT8Wx6wzyV4HaGBwumOUGRV7PS9kkgAdqZX
CNIuvZcqhb1mqmxgdp6nhkci4uPo3AUf9FfGYAljf+Y37JVKFwhChHFFZxHZ/XaP
eReXj7hmFf3vawxv3EEVVKjQrifI0l4NWlIK+48Y+qGDPzirOhI7lTv3ZTPcI6ag
6tnzdaG8jV+dTe2w08giq4BFq4jxRg3ZdnnA3BILLmkMer1DoMVaDDfo5O9zyMk9
U4lnh+TcwDkJYxQ/YujlnAYr7Ld5i2SNLoubXxMaWM8kscro+e+21bJ9XLC+uxp+
AfkYTW/7h76rBD60DlcT6Zdbx+9T5I6yN+16Rd6YB7b9jhYHHUCDD5d+fpdts/ag
ToR6U1dTe9aLrsduhKWJXq0MoJe56e6Dtlx2VvUo3unPPqK+BLLS18R4FYQpyTtA
SoYa4qoxGvR7ITa/QLjpWvHFbZtohG/kolktTLFuHbb1FfHBYX05pdFUQIXaatMx
DtZGLyQzZahZEhQbCn7NY9VQwd2OFqtcbbnQcmOfvFlYs3JFl0vfMStysQhTQGY9
27HYG8xcdQSbSjvaG9fiuge8RevBzhR1X2KFmSBzw67MzP6wi2gxy3x99H+v3QQo
aso9Z+zRyucOHWy/E5oKRHJbiF0IGBErziTdVviL+WTewh1XpxesFpkcrFbekgZi
huovDMSUcZmQ9QZ8P5WjP9M7b5+DLWS6C6hCi25DjSKOFnUik8zJ8ih/BYudBobK
q+5dtKprpZw2Uru/xWPDjDByGgNVAfdRFEgMv+8UxhhqBYEsoBhMU3W3JDBVI//l
pVj+s/aq/FRHi302xB5QpuSZUHVd82kCVvVGyCkdGRITL9wnF8ozr/l+v8CsX1aT
AFimorxy1lB3eYyQtwe0g6mRXk/Ezl8Bn38Qyx9f+BkF0TGG3HYVm/CH3TpyTPwS
mnvpM6dfm/OqbIvxB2tWPUFqjcSSfK+wMagDRshaSbxZcRWTBX7e6PYVHL3M5X7U
Uhn+iwPlouFbNO+sJ8nATZ2WSJge4soAFymFxcsCIo4B/b1YNzT0kEuE0dcSw2+t
dFIwsN0w/wqVDeBZjxgs9efAmak6fWCV5VSTVGsBpm9BVhnAlci8HZlsC4xEOjdw
yqDfF+C9D/3sq++YUUpVsfZ/4B2GlgNf3fWwQebplTjz2YlqeHjhe07bLDMDGzpc
ekep+J9w+s6cxS2+2H0PZAU6bJ0c9x8OIQ2DJ51/46lbvC1jV+xQsMyi1/jJyNKO
HeeL9fsGYqxQXN4osDnluo4xddU1tSDubksjxBV4U70nGpLLPPpMM2ljkV768jfy
MH6pERm9vFjby0UWTyEQ9AvuIVKgGzrxZYaQwpJ1E2ulR9+wztLfQLMtdEVlzuKg
xC8HTEWABvGuhu4zPXCN3cs8QNNh9R0hV6t91yU6MBrVm51RWMTg/lZRlb8bpbCf
QgNIv5I6pIUXOCK6BODzZpzIRECwIyRWD6vElni0x0jigA+G8OYrcgHN32yARbUT
y3HF1QphRWiyK8Cx1CXM7blDswyh6y9pxi2PHc7Zk6F6NH8Aznf1/y92I/ze+jtR
dJC/3dD6cPGLQ6Qrnia+FU0Pkye2OHPc9B9I1jxTMI2+Lrae8qAZLhStZc2619JF
Dm7W3BLzJALZSXpzhfC+yZjGBq/2qILdMHFFkK0fBQV0kmSCLuxvc/DD5xD8Tj1Y
NBmvz34ukW2B7PpMY5NjZ9cAstHqWCcueSQ9yBfJleVkasmitJhlJ4WzXUOgoxF2
YM8Y1mw5ScajfS3CsGXEqadoYWDmeoCLtsKYOJy+iJZROsmSSP60QKIM5fWwSzOZ
eaP5s1HxLnwaJUt+4aHJsTz8gDsjTFDbKIrOROLr7PIIKvQN20yb7rGMOJaj4iju
ZJT75ig+1CH3Y4CHi+UrzAmTte5BKWfqJCjNNjVU9KUQTuATUIsKqnnUVdbl8EgA
ZGEkwwJ9YYUU9rziHykjbOXcVnS3DoT/a12R1hk60aWGw8abAKgq6qFYcQBjj8rh
ydhmVzVn7WfE8ypohCOeSjAhSJ3CzkZVB/5QoCb3ZMUgquiIBZEZqn3Noes/jNe/
EDET00QDQ/fWXW6IDznEoOJASgm/78qFwOedxg7S9sf5BUptMgYri/ygnh8Tqj09
PRfRoKW/uPQDLQWTc2QVkppTNB71TygKGPBymmlJQk2/8dqQkodYe4G2opJjzFkH
vNPQ2hYyrRWuu24JubDOLpRZgFW8o481tUYSehFiJxvKCNI+ev3Y2l7TdAmjbOPC
AgNFznuIzubFT8C9raE/2Y9ZatZ4yG/E5ymirOcltWgFBlNQp+4NI7cdjTLsB9SL
566+roOarNjXWQ5UGLuKNDdjUxQ7o+NnPjcOn1ErwFvR/YjK/lr7VH+YIZnHZUdc
UtZr6hMvcjmyxgnWtkG37MpjsyoDopxNWDfT3Nh5KBstrcVquIbb73rjmBDsFOM4
isy4gJkVEetW972W4Q2GYMq9Y6iESeotRoQubkUZ+q60O0+3TeQvc8EDXOar50e0
/2hGhxYxp2Bb0Pit2kinxD6EWmIEfXRTmiE1d9GP9NwabzrT3XYDFKQig7ZX6DoD
JysxImDTXWAsV8DLKUwtI8xSNl54tGzIFhMvDQc8OeAUIdjc9pGR4XfVnDg96QC+
FqfLIFahQVDbw2NZMHsVwrkELN6c2JZat/1I7w6KP1ngXeCNuo1aY2VDtVZpInxa
UNKKa0fcWqqan1ySz+wlF7ql3CxAAhB0LGoYsCg+HX6njnhwRmU/aJbphF348+FU
+GM0jhF1Qht9fV/a/xBhtHWLTKIZF69aOECNF+Cjhq7HgD6OJ33Lkq9WDVMBZze3
BruAHkspBHGV7RawZyAebHoZk+NKDyCk9fGhDUXb82mVQfqNwVnA3bNSJimny6hX
cXerTBs1DV0gdv7W4I/E+BOmnN2Fo2DF9s2TpjgUOyug9qKBMdZyTLG6jmaMy5l7
YME01hqnV7pD5tu9Yqt1bNSwKHv7ITZhraozWOve4AxAucqeDZ9KSXKh2H/Mfjum
pGYMFtk9yucH1StCQNP8lVe2ssoq9yt6AGRipoGQpT5onVixei//eUOtfyyHRolh
uLj5NfId6UXHJn1ujUdw2lCrDJdHHFlp0A+OeyR4HSM+UZ7wcAvY/LqW2GithHVw
rb6hhBAkuP8V56WsZiCVDO1t7dSLpBKfCYAic1R2imxqFeyDk6LXUmLtPKjtx2ux
r3wIGFZHhWrhWX4+cxOVXSIcPfzFZWbq81uQrM0xZN/y4IQloRnMibHproINP1jc
t2W07871Gz/D7TYf/FMgJJwQUb4UFZ2/ZHuLPxH+c4vWUHo4AU80nGb0IYw/UTiD
Pvr7F6kS7D2W77OXXMPeW74FKk6jUdtWHfappaD1Nw/IRZlIfDN7mKFZWjrf/vW1
ioWOT20PnnoGRzd0Y8LiiaTtKDWJxdB4vAyU/OC0xdGZqwzQDfq9yvvhr9edH1v/
dCgHGN3L+vqzZwbu7csp9iqB5/MmpOX3+i+/SjgLyb+sC1LO8eiVvjAIaohPa9z0
Hfpx7UstV02+kKjt6h1kJfcFatz2L6jl2o3WEOjDMk7hVDJCr6s6awzqZls8Is5F
yg704LnGZT0z9Dk3MrZp4vXmXezQirn8o+vSFEITzlbCxxZ5a1UcuOLPpp1cnt8E
8adR9S3Uq0CefZbd+OOsQsKbxvgNt9NLcki29ufYHoe7yIozParmOIb9RUZReV6Q
4HK0P5cv6lYQPYROiWSthQqrL+lTnCpX8BLrtBjdagwtlxVa8KUl+abHU+HjtRsa
10nYHg14LXKAUgD1DQqYij+mBMERkTnSIrqPMuEOlUV6FymDscG/paFCzAoefEaR
achctix9eIgCnLfYfV4cwhhJv+kaGcQ1tT5LMid4+rRrlx/aJ4gg2DSZUU8dhiut
uQ7M0Ljye4lyJIHgkpdZvOI3guS3S2GhPhGvL3b5/zaKuvYh/JOb/OO+4v+eQy8f
lzlBtZ0tw5CW1usbXsKeuNksDfC9XUPdfGXFCfQj5v1a1aqa4occa5GCFvkagX+E
BQcLHbHquRJc3yS8xmrBojYPuzyVpLLnIBg+3F7dj5vxP4VCsqT82yZQBaZxgzNM
WsftUzm0SIi5IowyLlsumdO++/JPmBH07WEhVPyH1/oT1heGZYvHYtLJ0nlpiQ/B
U92LBsI3Qr71bdn6MWns65Nb9g67eEoMOi8BsVq3AVjZJaZebJgHM9bcIdaReMzU
IScAF6pfpoGCji6YsiYPyWKzRmjwtWuqtj/QxTcTzWXUSgw5fVAjAeXkCNnOjR3h
SA4BuvaJgsQfdLY/aFo1J0Vbg8AwOzpkjvXE3kNbxTSFa+1MF1IbiwcpkgPhS94l
FwmA5Y3mHZR8TEG1+GEf3U62Ub85TI8myO2qhNp654Ls5VejwUSOrmk5EedLjyCy
AN1/2GJISLDXNh9MOMYSH4BqYRrKUmE23yxBa3pPcDbU4Ey7Qs0YG2R1VA8OVFJJ
IzIpD3YncsokvbHJ83QE9IRfjtJvwJkL/x/DBnaW+IpGf425nZqsJhEuHgC3IV7k
248gKz+ph1FRPjP4ZkPbsirIgPL0UwUnyKh6zGiGwVjn6O+8A+vpfuEfW7HB904b
emEId+6KHbmh82h9DxAoqano3bOyOLr8QQGDJcKCBItALUJ5tVXvYHalELSa1pdp
b6tmjLgtTvRSf/WxgYKUZL+bcPXc/dZOI/df1BAOg4G38xVRHMMk2rqhfFMDHQkW
MiHkUPZ48gAVdY4bVt/SdZyWG/LdH3VesYu5L2V7pNkuD0sBwHEDunSgZy8X/5AG
ITiOxyK45yl4xSlkS61EgzoGRZoG7qlB38I42z2z1E9sEClygvs/snopLruOBEfq
uay8EZKO+bLjSCg5/39Ep+QFq+9OkfTIsfOLwJkhmRLY0z/g0VQH4nfB6Lp2sX4A
sbUBgjKGhkZVJk/vmujTV2eq+Ba6uGRJtZq8KPHs0L97hymO/1TwcBkztQXV4tAt
VaJFwzj28ZJvkqxI76KBosEe7Wtietpid1W8TiG3e9qaKYw1ABtWrxHN018XrKWf
oX7eElC0TJHSCAkab4k9RQkOwE7oWXZWUSydcPSH5Y22rPdemX91mq0W1sverwiX
We0PWiCu8ufPhk1xXvUacaanf5PScIu8iPtqMooSBKOX/Nl9RYuKnIHJpqUZLyzr
2M1vLdUPkuwojNid+ND6iul870LYXV4RLjQ63P7PDbyO6z31wPhalXlHXzDLm5L0
aRYJS6WPUD/4oYt91WmsgtuQQChLVWt/+m4LpFcs/AJSiZE0ZxbBsmNcuPj7syuw
4epV2cFdNsuN7HlZEpBRqMZTk0AdvTfI+BQqqj+tOTA0E/FAfpt9B5jPOEjNe2q2
ArDPQqQCrKLa4ewMOMSvOgY7WcwMFMKRpO77Y9AqJhcWSWr/+qDuljbxWmlqw9kX
jgH3hAea2Rb/jWRbmrGYfj9BgP7CMz2mBnxJH2yMAlFaDhf6np5e+75l/IoTymVo
ognASYJ2RTntkVBJksIzxigwgeKKGE6Dhbk1X9fyuO9wTkh64trg5HeQF+MQZQ53
sS7f3Mn+ntlMNdQR12NHISib8Ns3AK53JWawRGJoBuaiEnoIECcMJFtQWR4GhvVR
2w1qLKjckQ2tamTmvO9vrSONfFAjI5HmToYLAd9rsXDOBlCslS0pY3Lr1rTFFNoq
Nv37OyQXP1L6dVzpLnoWyXKbtHw/1iXg9RRHJG8ybjjHo5ClNjnQzCS5NksWcsED
tVrMt8R2E0KssuYqud6ih19wCOyoMdm+3Ypsnc+/Pq46LCn+zlAAeePIRV6bri13
Mb0FSNEE3L2tpMKNFN93tS+wV7YEpXBR5RR9mXG13bDzFcAvIb5YqZtuMoIpyTQg
TaUdS1OrgXaPMzs8bJOn4SVQ9xP0APUHQsg1P1JuIbWjf4rkZXGAzwSFvAOG/z5o
kCYGa9jC/gTXcB604AIUnGOkNObBoSma5shEUnjGMEgiXq5zkcT3KyMUKTjRhd2n
oVj4Uu2OxKFzcxKjy0kMdlnXtHx5klxMWFJ70eS3I9QK8h5Saj+T+l2sv/a1mrzv
b9BgmxCy6Wqir51S6SzDZH0tjQvo5I48zBTifOzRicbURgSZiiaJo6bBausHvzhp
qCXNYT7XZdOmaQlqAWbdYb/+CZEyP97lQdJzZLzR0upmhaYrcQ8C8ZgGHbGA8u8x
7l2FZp+9wBqKa0Lznb5hppv892Dj9mghAuoviMZRH/CA/sBLEPQL34XJDh82Q7Bx
Nl8fDh+AWfW2TKGJHNTUctKFK85kuFugpNtNlWC0Jk2DSh9AyjtegSeb/TPn4WBY
hKYchS3dN4WS5EMESMQCXjyfoK7aTcGgAASTmIoKg7gIy+HcH2q29i1bVzPL4Pfn
RxZXTw996AYYh9d8a9VRpniD8uDuIxCosSbnEdJ9icjjPSzkD2zitnpQ5CYKd2mJ
ZYH9JrIqqIjL6/ctOz5vgFD4ZfPBp9XrZDeWRIUSrb8BDlkUR/J0ERjqZLgVOHYS
16HahjoWLIHqnTwS4h+yLVedSIakJrgjtV5oscLNvvt19DX7DuU2U8zex+fBlMB1
kvOWbPuyLRYZE1efM0YEAxU/64t8ZBYs5QH8d17C0oBeH0xx1FdAI1/IdKoKXZXV
4415U0vo31cEVvCBqzqMBHkAPbH2240qvfMHeG1eTveNKPFPz/OMjEzU0HvCgslg
fclQOA9cRCUiaHIuc35DOcf5Q+TQ3tzlZZsF7m1+fFqV/ZPSNquTTt2OZy1WMgFw
FT6DSz5HwOKu5vDTb1VL4MpuJ6V/y4EBeD8bElM8Y4adlgnn2Yu2jE7we03zZKpv
nCJ89TkTvFvg+ToxJ+17ZXFtuEHCfgt5SYyqaD2k19NZW/oJTP7P5X3a/OFcB7pY
UXe9I5m1D63shRvIhLoSJW66Aq3Ax5O7Bsj2VRK8/ct0YwsKcBsdRYRuLkHC/qEf
a4xc3B+8ptN+dhoxn/WplQwtWOTknJIxHVwecD4Dch75EkVHF0AAs1tvSHKw1GeW
/5zxpb0+/HMDfcV+eMmpmKrE1eisdPwE0snymjFOecUNfG2Sq3Qm4crgg02ZSIjC
UC3Cm1eXEaF/58ibughTO9m3rTUY8g4A4wYSRLzacTZ4CrOi4OWyDQZ3IKUsi71G
t+CYVPsHuiPAWIhgjnnxtgtzELel0ml5vFPEligCHNppzzqAEVqHE9zFdaNVuPdm
1J6UvZKVxVGEfiNUJjaLSsxnMKJTBbqTYzTFm/B37dSd4cDoV5OWO/61PCbxewmq
v4JlziVQl+xKxuWhjrs9CkqW4PaUgaZd7YsGKaav4bkuuYcY86DUCVyzd8yYnp1h
iduO8znvWxIxcOzjg9hQ9xaxx01LtnqdPWTdDfDYuNTMIFrVS62l6TxMBW7wnAYb
NHxbBA7kSPoqV95cZKEkyIFXfy0WKWtYbe0XVF5+lEmtlpQOPGSMDgiYDVR4zo4j
TmS6LERDZ6ZrU1JucewgQJXs9yjcPtQ7moG6dQYEUjdtB/pmB8AHCFItKNhnx6P+
hvc+QTIW7QjRetuhYXBfuwjJZ6LGCIzizoOd98312yroN+GKA1HWQDiaTm7oAcJf
DeS8soKeXOkAgrJGvafQyKe4DL4PYQihsgm/fgENLb43/641gQo23/NpziJwHD9a
sK3iPX4YDRaTcK2zbW82Is+rONMvZQxj+Wqz+FblzfWwC0dyzptj0DNhbgP7VTJv
8djYrvEST+Rp32RCt4Y5VPOP4r9f90fUDcEel58bMU27jWKiXa2zjmfDLPX15RFV
MQKDOMBv4n5F2IBBg1Kgrw+RIRozW0Mp8F02BCEBsUbSr6WSDW6R4hidG01onmYl
6RrYFTuCViCRUo6rc9+eZ1Q264gkfxn7iSuP46CStUpKHdrZtvvpJA8M67f7ZUq5
QNnggjEu6D8HQ6J4ORyxx0Gs7bOnk+pUnng90H7ZY1xtEhMEzxTb8/Nmj+az1u7V
nGMtLh0igJdKg/CvC+QisZtjI1a0df684jO3C+tsSnjyo5ozqiOu2MlCeAcopFSS
6cHg5PykcxWk5NoJoDIqfBsYK9qi4UzjdfIV+cGee7xHskpsHqShsPirc8BhQa4A
VMHUzXzMpHZJsejiq9AECZr+NsFOEDJjOOfuFALnhN6kOUVjqlBsy+Sc5fMaZWKe
8sHzCNAv4rHOKODGrbu5z2J7obeRLp4LfB+Z9zmwX//iDXSIx8hMsDRm9c3F7dRN
nJCzrpYZgE6hdLYCSc2jtpUEZVIWz2cXhjqm9h+OuQ8OJuU+2XWDkX3mFyag+fkP
rWk8ZdspY1LGcR23QuVCQ7dHRQwd7dHxIvBq0cZOOhKJCi9BodyA0FI5h+KeCM17
nHM6z8NYhHHf1YArghVQZEBS8i0/KS/p6WgI2GHvp8kEQpUuR2Q5/L2OSrTkM+Hj
U0i8vXc4lD+WWw+4z6TUnf/XwmK7espxIukyVSQsTzuBTj6ae0CitJKanAxiwNsx
c4rnOPN7WTy1uaUdPKILe7bjBldS8V9Y50KouNQ0PdZiSrx0r0QbILcF/RwqMFlE
cw1qOHa5jY8XvM8FSmVHRH/Y7U/PEh8pirOMLmxe2wICTkacXVlTc3EdXBeFdmA1
Cw46D4dms7Np2Q9AswiUXV2ptrsL3lTECcFvcCIEUsnXnm8PA4HcMxaYDhGPbZMC
bgSz71anql4WaBx4BNEprCrZnLNMdldJWRt6/EBkdLwlzSUTJso4mYvO04CMF1F0
GmUlZWyxxzRcUEOSJ6MAQz3DvbE0pq4iHwGhWZBOc3YVa3QksHWdwUnuGw5U1ZeZ
6Lo0gj+2bWolF/eSgzzvmfqH5Ifu62To7JzMBCGhv2fdDUGl2O0DpYSv6r+3zidU
XZ7iseqYT71SySLpDkBRZ9MM25dlL9W/D1JX6fc3zVhGQALVUACniILf26vtw5Th
TCYg0T+/wQKAL8ZWBpMbwwXFEAWzoL4vFw54lnvaa2oaKGP5NZM8GlvyVSlyVq5J
KKSWCZwwvAESmfz/mRSjikXY+bmNIWPklbxBAEx6CFRbM5lAFjGil+Is7wf+JzDH
yyS1Qhs1daPq6iEuogJ7vumQ5Sze1uRjLRBh1tomprYLbmmWULLisF+ocrSaivc5
71uoAUnkhhCHX70anfRft/jVI8mf66u1ZUrDhLmESyfxFgkn4vpMWWS2v1kThrLb
E9CnF4gbevFrW6TroPjEd4FeK/u6GaynJD3pMIe/hGv3tqLS0kpf4x7bv8Rwx+Ta
BNC+MVaLrf3SCceOZZFhVfhaRBHJ2dqjUuBXrXr9anQvGi3WoGAXGvCDGob5Cuih
AoYiIaptj60NhoQjUgxG/9oab/5OBEmxT1XOyGr4Y5UoOj/6rVwMRPoTxvSkhRTz
Gai3i2aHqSgod7S4MZaz4Wne/ilDjT6h0+qvUDUP9kvE5HMPdyqEZ8MCCdQOGzBu
Jxk4vt8p8hVgS546fZsy/Y8bhVtyACSAu0tEPv13MjNmq2mV/YA8JIQ7g6S5y0JE
ko+mi/lukLL5IVX2QbwN9pBpze4lPbbVlz441K/0OVHvCWVzYbgOQj2pNIuMQPfI
+rsKL4obrbz/8mimTUV1+nGK6pDjrvX4fBrDJK6Mqz8dH7ZlAjBnyo73v+aWusb5
t0ajyiNtz4mNSKga1NqKgRoxzOE4J1XJIR9h3Z6JVC7mcuDN2tFxPCo6DNHbeiWD
VPCBhibJKf7pobyd4QknGGhpOqbykETltiqyVynTlunO5dt+bvLBQ/kQsI3txhlX
0XoDn3T4sysDH286awLxluji/FTiopye7rAepFq1V9tW++fep0uM6pO4x2Q4Qp/B
y8WX4r0tZ8d/JnMKbUq0/enfs3Zg4d1ptkATujK3Qxve8iPaIyAkWM7pYt/w+b8O
KT+XInA1YbsqE0zCweRQJReQ0pQtRMkEDbmIaRhvBItuQoptdwerC5qcoW5Q5gPX
6n2NzBsDca65xgHD19jwirVI2xiMfEJYnV5WNdOXYa22Yv0QuXe+LNX1fCarAYI/
LcyWtLdpli5HZiPOz1wJ9aahi2+Aylh776L1WlATNRN8tdj6U7L89xQzl7pb+Lxw
YuK2z8Pyt3nKS2yXfKqFUFlJd1GMT1JSiGqaM+om14fPZ1g1klaLbbCzZE77wtP4
C6f3XruaX0gRZvDuZiAl6I3Q8kWz6QpoW3ikCjgo3Kh3cB55k34+pS8/GzcvMT+i
2vw7BBqsYeNxzpElAQmXZ2jWGsK/Q7IrmBJjk01rjOo1HKeypf3OxlWcSYHTvz+n
v80qnUC27SoJ8s7NdlHtzsFYNkn7xAlWwpui7KeAa7lt6ii1JigtP00jEcua86Xx
T2JVrsPw1wyQ77n/Mpe1rjGx+fmTkgN1qq5rc9HLXC1GLvvPftUkw5t22pXyqEH2
QLkjn/fH5tTxD0UpBYWQYMNy3dnVVQ9985xnL/aGwc1b2NdqfeadQkIrtDj9Voq2
IZV/5qPQYnOporLWZEWJEjMVmKM+/0HxbQFTfzSt2/D2H0urhMBYbVVG/wpByFqu
EOS9k9a0gMWpH97HjeSF1gZ8stirpzY7dkDRa3PCvkshU0gluTNNlrR6cnVbUN3+
Tbad/AWlBpKq9KVtBffMEFSfFCU6F/YxPuJvygftI0wzJpuXDUfuBFxU3qwHMmPU
x9x58/NWpFTzR9ZdOl4+xI/Ft0fdo2detDPZ4HKIRQaMuFMZvPeqQuRyw4UjPxtf
nv6xcCuaggFdQpUMl+q+QJmLe5mSAWLPcBUBYWf6LCliMe7orIjw6HrkHjhjMSoA
2n5meYjHS2aCeILt/GRl0jsexS8O8kMUbail/QD76EWqFGHYrXMHFD+wIUYiyxie
nSeNZILNCTGdQLU374otf2CH1+FM36xPK9AZ8IExhkUySAOlcItp5XXfUPqVC9EH
CilUOzGTY6mmMNX5XF0saafte2JNjUvcgBdDGW/6mBXphAjXMenKkmMFbbmwXR0H
GeS5LFXX3GZWzJIGn5VnXUNnWiinL7JmAiYDILg8elKIVWvk7TrGYsfUgFrXdfwO
5zsOE/YvD9/xkUFNTqJqQrUBNeYsmceBM4NIDffCFhNuai82pEGJf5Qu6v6NP8q2
Za+KKG4FRtj4ey8zGlwV2jpLkSXiyvVsEZrZAqdfdjFlunTlPaXjjUno88g/2Dfe
1OrQRCQxIHpfGRD6CDLvqE28+LbKR6B7p4a2a3LiUH9PlJr92+Nc4vpFGGuERo4Q
apczJdkpAF+f4kuSAT9Mkva9he4WyCZT2G+iJjFRY6bx5VDDafhbMXKIS/FK+Ikf
rSfg7LdaivTCft2FszwE3qQE7hcOrKKztmEnnEISeB3T91wIlLx+p7Di7oqZohLB
4Xwf4syxBKBeQnXxAGe6TOhD/+JvS9CPHMH33I9dTtV5CDcWbujjHal37rwrDduM
CIxrS+f3MdYo7KsyeZ0IRFZpEHVKu8y9Qv+iHnmNmVEKzqTel8oYfQokq8mWXU5p
V78ajLexctSo75dKJ7SJ0YWsA6412V+BdBbKY64AtlW6rXkj8t9xiiZNfKyWfRim
jU+sspEbKcmR8MDodjzXDswV26zbaIsBF26sCvga37jO8Hnp5ctxoqZnSAK/Sr9m
mq2NiL/+6HkXHFMoaEThQa4clS5vbUSfqz7eVqpV0JZklvWKE6Kfcxy86cyyGS5N
F6dJ6QHBxe/IvXL6AXCw/c8+PUjN4Vrgt3tRAQiYLEtJh6n3K+VzjHyoOuUubhih
FqmUzmkv2Dz0vY74CA7xj7UoG9TjTDU15Fs9byFYP37wH57s0oqx2CdiAsLYjeLW
+JFSNiDRAV5JwgpV2D6TnRrXXHZHBUpuEeQjScjAGqizKAmiiK+l0TFCFxSQ+RRs
143p/xOtJWMDuv/YuZZBuRjdQWMng5wiyqPp349xxnardOrLnu5GCGOACmkyNykm
qzZp9Z2eljJ/mImuz0BfWzKlD2lPT0IR1Da0tjsbqT+AHCoN3JzvzJaMaxCbOAsM
+wy/GVMcNzoKLFoUfu7//MP/rBmLqnJaAThjM/YAir22hFPrNc3tEWoGfs8+PujA
vWPKp35c8znJOj3Qe8DTXAudIghxyX9F6OjS/J7b1vWsshxStlhNLGbEN5tJJEfU
CcX2iEpFGUDKhjM/zvFFIGQ5bloUJgNBeY0tHPkGCXXq1LatT6GoInaKVSVDUBA1
Bh87xH0R0g0cQIcnjnPmVR6FjEuwGiOpM4SK21jUV/Z3it4Oamm57ejis45YhfIn
GpdObSwZGuDLgqlKFqAry3TlAxONWTSK8FKtl+BUCg7NNfVStUaalxnDeHK3yrK5
zj5sLrykxz7eYXDKgPzCdISnf3odipNlXj/P6hjCjWcYKgymlMmy2rCrOFEe/CFm
LeKS7QTAmtCiB5fTJYiaxbROhBTZfOePtv06nq4mBpoATxt9XH+MTjnhcMKmB7sO
GX2hZMEkpoBKR6+KO8dhG3vwGPKc0IPIqVmKpFcDjR6lJObqLWTOPXpZKAPMKJTr
wBKwmJwSmEcwAO7SH5foA1UiVaj3eXotG2ShFD6S59nLuF9J0rSFXiQyRkFDnLTu
rPKnnaHfGPugmu+wll4vKHzz7bm4Am2zqLLpQz3h6cCVXXmRKK1psWznVJRtvF22
VK+sluHsGsDivO7v7QApMDZfYNMnTnYLvUJ0KdGvzH+NmR7OY8uqBM242id1185o
IwgGuwDdpzV8QEovHNuSz8DtYEXLIisX+BVZiCrRSdusUjNmJA3OHGuauaZeyAht
+6fvY5lbzITGqvBFekIoSEtEvQAtwJY7wRsYOhTf/HOcoEXfnI0w4R927VG1zbFA
oHBRLLTeeBuL5lZgNwFeQ7m0QdEmhcrX3gyAx5CVbzSy3kLCku5Ma/FDTHup22wj
+8uieHQP/NA2YSpMYmK3Cwr44k72mn4K076JLEFbJUifpNFCBl59mGaGtjXlCmwW
bd7TgPccVb+nMofnfHG55cpcQ/9YdCndwp+1kSTsQc8zunb+g/ixM41JErZ/Gvt/
RoBWp0BO/jA2phR/htQ4PFTHOSV8SSxLKW9MTK/C+DytZnkg68Iqd2WxerookTEX
l0di1ANTzSvnRvhL1i21f2cfH5F2YPVev0jLFVbtXXzVmKCMsIMmIX3wZRC7QRIY
o0j5902+ScmMX5gmNn4/Tw11yyRRRkySss/3qX3pXaGQRc3/stGz1gGjgbQy1UxW
fsgyIQkFRiX9rM5qjTS6EGTEq6C37tE1c6lcHpL4pJ/THY2tNR7Pbz5PfX9L8p5w
x62i+8IDF/0J1LCTW7Lg/CSHfR3uk/1mbIV3LGRwShLNBXupIZmVX1fSaIGOdqUT
dnF16/e7DN9poVgMYOy1iQGQCG7o1pXwPwpnxnPMQMOgdngwkc9Whm5FWsx7/1tK
M6SESMI6t7JkCrUcBrzyl82JcY53RT2LyBYyscpYP9BE8w5njCifuX1usxr3U0PF
9JbEe0HZDvKA0aJvTO51Kpg9hKgUdD9oHMx8H1cn4Fdj6uQamNI5wfoKbpkjSJns
7AMvKAk+7h28P8TPcmB1VCTAxXo1mcnt/zRyo/DiMou32l3KVAb8kASWHlkYGIrk
EShuUWaCxtCSvXn2PbnP2WrHOyjtmGYdJM3ualOA+NLpIvSz35WVQuEsqw9gvLXM
qz8BsNeobxDp+vF5S9tT2i92tic2fnv3GB+qsJvDNCDgT7kVvVVQmDyiMsdkZIHL
uKH0TZFJqnTolhUYSeIbTXdKCI6wt8nncBs8OQV89/JAr/HFwNYZWTld3rp8XgdD
hK26OXUme37q1sgRbFzeKJFrnQcDaI9/ZKnhAyYhVfxqmYi+DNwx2frbatrqMiIm
P9amvLKi8LpwVxBzKzPEhYr/gZmuLOP6tjWzO//s3+pBRIudhwWUCYMGwOoGaLNa
SRW/bvJ+liOjsO/g6t7mcQyBkR9TYRC4RgsZ9Mqs//69mZmIgrSrY2mswICk10hA
BlB7gWpyNB43o9dRCt4YnsW/ARvnOrtTq+YIpZvJojDiIcrlwZRU1P+7g0ydmg/J
wLU+wVKwH+dHN2VtAlA34P+LPCH8hwQQqOsG2WntZC2hGfYKOGhr0MEMm9RQVtVv
AJrRpif8dHrGyL63G3O+rAjxt40LVtF+OlCtRwiEL7RJAC9f0U08r0v3y2UoWxDa
Ql1fIASEPMBci921zsWUDWQ7SKuhQIlpk+7dIBDj1IOlZNQTKuFet9A2zoJrYYB9
B6zdHjDGYUi44qoyilKO/6UX9uNiaY3zGy5ovQ774I7jRbKsmbEN9J38CT2QpnCp
fp+t6e5sgnbd9FPcRsUtQErb5ZFzIjzez4Bvtr6zrfTUGP8G1gGSlMT/dN2WLqTO
8ElqOCGY2MpkWZLna9urClXxVfV+cV9STi3FuUObzpOenE7ybA6VukaJiWeNCjyr
kAd1inT7eBomBFpjfbQ1Kv2/0H5Ml8l56EK5xUh21eISLgn2Dy6hmw9Znw68Rxxr
v252Uvw2UIw/VyxBc5ysLOgY2deIIbGUfXn6CGsDMlTAEmyWTzw3ND93CpggBNyc
Vl0aI437qxHxibv0kzl9eTSvk7An1O8cYXw+oMVp/XK+0QM7SEVoOX7wwr7gY5uA
R9lR7v48d8AO4w0oKGkFIKNi4/+iWQozpI8t+5NliDxzuHzgznp692dVoqM+2TcQ
MqWADbvbrU9fxX0XBePJwXUzGYYjRl7sk55jmKYYBcfzNJKCsgukr7ldaxhr7ccR
zz4oM2zTWCvKsCJOjrdJ8egWRVcrX3Vsez0WRODL/MzwloFrcRMZ64euRUaChh+e
rFQP2hjqqquMpFpFx1LcMzysXv3jHKPx2r/RSWmZCWoXwKpJtXjE2BXFXHJEwqfs
qXpcKwRpDIpQndo6BRu2wntoBeyncZNL0EM5bgtLEd5Eill3fGF7tNLLQ4kj+6cT
5mSuzwr50eyeBSER9gQdHFhT+mX/EvvkmCVKKsyQehAUwEOaPimIRvAXUbhXBzcl
kpPHx6k6uffJwV3/8G6paEDZ8f6MZO86UgZFqioDyNE7+bPHJni0p3K9CzU3J/dc
2T/wHlV/HvEYbj51sqz4FNhC0AgANmXK/TQut7iuWtC7jLrB7KuM+rQ6JEL3vCUH
y6wWC0iiVkTGqNb1wPB3IXc+nR81AMkTpR+tbRb93LnbEN3v4TEu1gX8ULSoO7Nw
e37y7wucxWi6f0F2qCMTFsq6jd0uUadhu3SnXRjwrAUxZXFR6yIZNtYwz/8skNLL
2inBtqdFCgheNStXRVi3S06EYVPk9nCCnInxK3lAxuqpIZk2gFT3NmEx8LBmMKPl
8WKBw4YghHpJn1KnT7eGWGavN+7y6azgPtkS4C4og/31MnT0VyBXoUKm8T4F3DzU
fzvsY8Emje8cn16Orf7DPyV3iX90NQEVbAMRMOAo9vxyqSuHx4ha8z9PNVNnwTCv
wYFt8/Eb2FVURkELDAnx5ISsMbjJCQAJHrIacvoXIA6wIo15cufDIUlThFUGkMyu
AHfKAp3l/Lht4JVdWkXc4VLcjGcjJUc363jUrlWJ0ma29/DunAo9MRA2lUdXw2IG
RJCVvSNzfD3MezaYWa5fQBCklkfJBHOjuPTITCxkkL1tyswMLP0YNR25KhsDXMkr
ycJkqffLwz1bsChm8gTEmngjblUl0eW8dUlEx38OBnQWB/C750afG8WG6bkTMH2E
eCyy70z2326Xi/NUZ2AIgplSjqFS64acocTJQ+7BjzNheNaC/OuVbAnsOhZHX4iU
ds3ornTkVSneuQB4j7Ga/edf9MlDyvhxqQlZh3nb5pv69G2Nr+izvro4Vai2Vtiz
l7IpVRjMkJrkrUgkLJtMXv+prxnxTJpdxNqf08vwhdmfeobgJQ9Htu/731igXRyc
1B2t+BHcIiMxyB+WCnvMNb79OdoJyAtBRvsgsEt9vSu+2ObFjAxKndBRY45gIJUs
gnr80y7hpMuQ2CohBsP7wR3hUKYqDyauixMwJYiGf9uq+PUvmvy8TpMBfJZ3G3ZD
v+6ML57hPkR+zaGuAqi9AbXqhulkWLAyzTnzb3CiPSGkKV/HfcR0aSbXlR4tNNFU
XA+wvY5SXex/lvL9utsrtzS64p4sIG2QtecSkBNeKxeLmtKfeQWOrj8gaPPanhcR
dmRKEmEH21N+v5ntiXgFp0a3n9tTUs0RsMFKE9NcE/FJmKDNTfY2clPDPzorLzG2
OjOgGr2Lsi1ytiBhSgfAepJYbtkMhEZHGzzDXJiMdXXfbOgw697stKbyPt95o+VO
bVXo2H4Xcwy+CBrGLvud5JpjZF0kAxZ3Mi/RDonInguEwGNb4db9PLw4Ow71W4A1
qllifFuKVEiBclRn5/jkKF0x4kTKIvjSJWTA0nrdBGd7QUbRwR3b4HOu3Kgad8Uy
TPGbqkQ0tMPBVH+Kyx7yJJk8aVPqplH3nKtUW7FuUQoNSsPKagqoeNTPgTHNVp1e
u2RodOO2Th5zbm9FPwJz+NcvUMsCox/70CWGD5YMf29hRf23eLfp+2U/24pkNGq1
phb73Tg2Yw0qbePhM+iJmgO9q4X1HfsO/653f++KmG9Z+M9WSSxKzi2uwYj/PpnO
sy80+6ZVQ0HT2tJWO06+lD4K2VAlIqcEPiArf+di+c418j05izhqEFdkQp/GjLQr
YKTrUoTV2taxMGmAprkHZIUEGAbUp2jmvBFRfD24Tk90JIxIG17ew7+4PZvKDtYE
EFIqEwyNSk7WMw7Uhc9EQOi5R7B4oikM0cYVEozz4GreqUR5ncxWq63G90ObTJzm
i5TOqIxjN8ZcW67XbRARAiLcZC/T3ZKKoBolTjUaBv6gjJ9wEvUuIt78ckg73FZG
5u+IbS4cHuyTyGnGrrmLiy00PilyG4PrArLxFTK3PvACy0Wd3DErTCKvUm7592xe
v7YPrjdI+3tjXEOVtKf7A80wFtXOFJWjFGOqgEAmDlUbER3xfyNXRTl4Q1sBLIwX
K8mjS0539rYE4Xnbbnsn0hcG+GUUbu3CmMHVJ+YiukSf2pQyqRPlL9jPKNYIKGbF
wGC2pdliPDVC/t6x5kTUeVEBeHjHReO4Py0PSWdbWJfsZTahhTwyA320LZdKc5Px
7gqnT4suUqYgeIuuDogHgG+X+Gs2utlZ/3kimFYUKEPPIOOkoow63xGTMX4hd7Qz
nJ57eBWdWpRVCEDbWctE8t9+xrA3WO6Kw0Yn1k8msb3ncz/z07nRYMppWkMHXbaV
cMPP4pJHJWa009GSMvxVvNl/GFM30NGCgVvljiHdm3Ol31yxdpMxxxbRqX8lgYFE
6IIlQdo7oxbhgSqcNJDoWy3zEVXqJ8mSIMP4sXjCbWgT7tQzQmICRTMKg5vTRMar
R8sV3rB/3VjBRG/iE4qq+w386l/J0/vvtWUNOGLQzAq7RKs8otDPnX9Vj2ujJ7xs
d/PKj/ajnWwyJBUVABGH/NEh+gmRzfTDylK4JtsWXEpDChnFWnNpuh355qLiz8kq
ED0dCWSXgO7jGwT7pXq73SHF6mZWRH0L7FGAgoexAEEbiIntCUrJzQY2otPsFs2B
IF9AzIgIPFgQXho1GfgynHvBQgNP88l/QWjivXf9kc2dlDBJxRz1Yk6wQVwniFa1
RF92HhDF5B4oock3LjJaEzNHIoAdOyIjQGxvaYlIzAC8eVV7Oe+7LiIuDq8quye0
WOIisE/HOqW0q6553sTLORb2qfDLBe1LVxAfMntwzC6IsxHHVxe89sBNYS3o0BRq
tDNaX8zj+MbLu5B8Yk+UVanSCghsTBdwq8YXFkWeUY7tlvAQCezt2/R8grPjNXtG
HmWSMxCjvuOP/GKpS6fycgLtlS3AfYx5f0EHfxcGlz+IrplPDoP1sr2MebcdD9d5
nd485NJc2aKkANksMS0f5HGB3XjYHV1QJBmuHCirKyndYK4FWSqXzADW4vxvYRuh
PoUAmF4cEOzNz7Z3VYesmV4ox9CRndsWUl7sZoap9zY9sxUV8pEWjmIaBoMKJ/3c
WHKN+t6rz4EiWiozCQdVAIf6foDhxtf0N7JLRSLA7GWDwiQBmCIlgxJcmhLSPkuU
pKi7l6FTGnYTTed0I2V2dkR+C6pv6s0qeuuEg+mqDcrKcSQZUjvpAyo2NHu+hMQl
7s0IdWdZyNx/gpTXw0olGaoUzRf+ZWur25qhu0E72ootPQZZPLAZzi1OFV8e0fWk
awzht/MpuTgjvxDiAVO+XK3CV9NO5xDZOGrtEG8CSSYFGJfXre+oC7sc1ou5fZX0
3vYq2ih0ltnhpe/CmhjbRAS/+CzjhBhKR+KrUZkPHQaicg+VKhPs5KxZqwmVFCVv
zNEaF2Jj2rErGHc35pjGAQhmu98H5XmyLluDEjKP5tQc1GgO//qINjqKCs7KG/uy
PehFX0oX6ikVOU02bIJ1HbYeaVvILTsdL5qoFJi/V2QT+vV/C1JHkw6lh0C4vJ5I
P+1a/kTh81GUbdRRHPZq2MI0h/MVyjInx/kOc9Hy5uP5jF6brhpFhf/cY1hbliMZ
wrgaQftxSwR3PmedOW7EQi0Wa/PFAPRIrq294cRX8PYjraB3wry7O7XXSIiKOYyD
u/bx7BT/815YLWv1Idguxs5gXwkqQ6lffDG9HeTH7+TfgABKQKXiM7FayWdZRLDh
7maTLk2q4Sukm1rqIJBfHEl1NlDVnLDORqv4VWQdx703pXOGqICBGYKcpQa0Dw0a
zL5QGWvAogI0p3Ldmd6vKgf6rVnLr09XHXTtGkyddJw8WETtqCyGy9YoG5M8SglL
hDU1CDkjJXzQS5HsIDuVif8u97JnoyCvPPVDZtZxIzBrIEn5GH/h/gJkpBFyiS12
U6Z1WAHUplXdGM+rI4j/8lquhbhQcGR16cVPI+A1dpnhCjmfSHUmeWUwrqVIvo1k
ehC/43e4Sl8pGaIm/1e+zje+691HJ+ltVV9LFHfVzJce6XDVktJciIugOLwiGSYW
DkYmEK2nC+iPvZILhFNRi35DOa38T1IP3T9ONA0EBJBbWR9dum1F7DggLjZ33vLf
O7ewIREnqDkCkfdR2kxa8Rc9/j84Zc5xaoZYny8jjrEdOqRVx/OwrT76h7HHB4E0
vR8r5EFH7JMFNfFFcO4BnrWFEM2AAPHk8LHG7R6maV8FvGfclXqiDL672to/qDuB
zSJdEhhJKEHhyAhSu71n13dibjqF5wndTo1Z3i2oiWXDw0zua8/ptQPFq9/R+okJ
qbn7KeeNOLZ+hn841Pf1KWuzf/LHl9RRl7XssO93WL2HWknXCh6VNH9jPhWipfxi
6N5s8vhdVmREhYsPzVBQA6I5spAjd3/v7ud0PzDG5TZB8/7ImSzhzQ4V/sFWtboG
7l8aefeZeNMDyaDXcLg0ET5We88aScgkBBnR3X47InAROzimTtGIi/txjE9yfsxM
lxE4AJ3LUrjtvq/UxrUAULnfKMJTIVs88L6a3JFcIApU3/lYJeHcQAoDZjOm4DW1
ZNtHyWfAC5eX/ELHm8TT0Vvof70kVzAaTit/UVtG+XUWM3w5u8JSvuAKrw+z63vL
xHfhTNLoFm6+1bvta1yS8kOEdj95M4I+vZWS9A3RXXE6S0CM6+dlpCs3yXFEcPK7
zDW6wvQzM9jFHel5C6W1ElVzmqb5EkIEL2iDBo5fm/wBTCsFHKfF0aiIRy3wlrAY
jJ32ZgFu6fidehleOfp21pG9EApedHeHO7KWI7dskwLJNNiBu912evmulJ1vy6U6
gDIVk1kfSW0pDmGbx8BOuId0TA3c/VPqZbgjx6K5JJXy5Wdlsz+vSNgATnQ5B0sT
r1hIZRcW7oWANc6GXzDdwbhbb/DF74UN8C7FnndVazqSJLPkb+cfgMEO4g+nI6zP
QQ3USnTC9NNrUo3XOkiMqDxBFXcRMXNdOT8XvKg/3/E0k3NS0HROqjnpd5d+8cRz
+uLJ/ktlsTH1JDv3wvJ3sWZF+HVYeIi18gPtxw1O9yQI29UXSAi6RM6kWtZJX2sC
5ihT2zHYdWgkf2F5Z1hkOHPmaf6HX8oz/Ice9D2KCycOzADEicrW5miVqn9MKRq+
KpHELeyzJgxLbhsRUHM98DQFH2KNXXMi64490v2Kz9bvZsTksYUpBzM5puJ11qZh
ueXV80VQNg45cOXMkfMEbqqeMSizsp+YHvDxGjnMCX3yYrEDb5ZGcNeY4i10hrmz
Gu52R9zuFIfgwKjz68ZwGSk2G0vO5mU9oSBNeDvRXlL9OP2SmWC79FCCBph+YOQL
4S/OOTe5+N12YW6zX2G0XAa2m8IDtCK5IZZe9VzNJL+wmkD7j4r3qcbPnk/SLYSr
J2YZ1pAyGbg2m3LC/g+v2OmgrPU+r39AmOoEeJCKVeNYcDAmZNPies7SY+F1XpWJ
Vb4B59GMkA8F2a6Ul2LtTqp7h2GTfe9EoD5AKjqgsFJ70fULaIUDnV6zvD862Ewd
iL6Csp1uuQAKdswyE8R3wOliEMfFEb3i90XwnQlNmlYY3788VCdh+ceXcrPrEOxx
kw9Kqsj6HSg2KW2NHdOa77kXsZpMmlPVaMf41esQcPs5J/zRlvF9SguC3uQEy7dg
08QENhXVRhTsM9OZQwzXve12UWfpfonK/2gI1WlCONi1umDo0wzLB5NOkZYZcepb
K/tlYNsrEjnOTAmAMPqKGAh79gHP5Fx9tNEzFjkSl5EYwrEm5J4Uvt0XY0QgDfoc
lUsRwvZxRQlV3H+a2aKHOIdOb/X/gy1l3GNoxeDyLdcp2RS/c9aYhtra5YCVlHir
/5xWWHGTNRiz01OGYAnOLZtHiEDjkLiUJPEPi8DrX/d5tYuVgMpvR1tlFShGk1UA
iKoPG3/I+HKb7bUfwvj1QgphsX18wO1mvM+nF0rhzgTseBWkjX2jkpKEmtL5OZlz
obXG0BA1ILcR7D8bM9KMeCk6mylOOo49R/we8Tnp0zrBp83UFnKMDThBFNmf5BYT
7OtnMCHP80+QF84199nd56xJI3GHvUYwuHpMt/4wl/2K5ECKI3KsheMyetnfkcTf
uhH27HhEgKXq+cw8QAKKrBns+lFbRmOzQSjncPO6ajXSlKD+llq4wmMOYT79t8Yv
R008nJYjNXms2nIctyMFK56qCzbWzDl9mbGfWi5nJT6XSBZBFxg2IxIntz2mkuMH
4jdW0L94k1x0+r4ujYS3DA9b2Ro1hYNcl7evRuSMLspgZZrOgA+/10AdADNsThFu
SFzziyRMI1QtDOdKMAzaHTCZ4R7UgkA9JjSuhznvVVZJBS1g0H/qmRcBkZqZsGJY
YBKmKllRXH9xEXhG6eddIvm838EnyVjNpkEP/+fBGEsdY8ePvw0pDd48/m0IiXjy
eHp/ew8xKAuW55q0OQV6icT51V297EM79uZttSA7GR3yWL9OJjyZ0c0ICHzrnucb
Z2Zyo8zLVeOhGrnYhMslgarBAsBbgZlZB6uM01H5mrHvhTiploZ0GLEuEiTyJQNW
yH6e7X24+63pv9GIJId74geq42242UdBoiZe7+fnZ+Nok8nkG7GtmIXiwz+3/xyg
lurzFAEOHOrsMCAFqV6gu1ERhX/5eHw2L/60mMbksDok5ah8FIi4y8/epfUlJv2j
Fh/4q/Vo9a59w9HN9ANGHHmSXlfxhzdov+VRyvlUlV7bEoGWtcdN+vkkVvFJsWww
rNAOcw8yD/n2WGwHWdG6KeIXpE6JScuR+tAfeFMdeeQ5vQ5sq/k/+HU73J/iQWVW
wy3iswTRC7EBr4fQuZ5DAACfDiSILBuyZds0rLIMxWWJIlqoLlXgQsm+4k+biBYZ
BMJBg8Wouyv2h5UQmTmyFk+eGBznm9jCR9YbNeJPb2egWnt2cgJFufRweZ6HF/A6
piQVoZFpfKo9CzeQyeMm4mjxSne8VyP4LwS6kR4XAVbIwQH4j0VyDvRgOeBNTYWH
F6qrzsdUJ/amoQmvDfkAGG3xZ3o3b0CKjC/BUYNnERJ6EpobQbfdPVNGluDYjP4Y
xHHTJqLBD/QH1Z5aljtNEtRH7pTnVKxN/sJlecGPpkraTXB7381eXJEgNrzo0+XC
ZUrpmq+JYND6iuhJRt1ZOh5rmPKKknbRv5z5QDKYDmTAsMMkp1pooIguxp0l3Xyj
LhsgP6PjxRYm2Wfdjkcvl9mRRnfgaSfhWc2vmCxDSdG4cSSAe0KTNZrjjW662hr4
7sSf9viS/0Z9IVGJb0ioSTYzT3hYJWI3KJxolF8kWrs3InvKmTxV/aqJHcoYsC91
ey/yNrNpp2hAhyIpplpT5tAOo/CGA7Rs36pw7qWFN+hbiwTpPzGOCIEOLGoRbWSo
+o0VOQPb92+y5EMhtnaQ38pO7puGELajwKhzPc8QslFjbC+3/9QZOo6VEOu35suZ
Jj8Y6Rx8lKOXwhWkRNWimTzrE5QVrWT9yrQAWMpsa5W2YRLhTA0hITW8ApeTIa1p
TVvXg6h1FeBmx68Rqhzj4SE5/whwqOpRnGHyMkV3Ry5KsY0qnqcauJjczGSb0dq+
EDLNtYSnVB8m0jccXbQrpIeB9JB9LrdQp7tLc0jHh48Twd6gMSUiqHP5LbH/mPgK
CqC0xURdpcZlpWruB6YC67E+rHIS+PjD0MixCizIf4zfMNTXl6Sjhn+bW6nJrWi+
R61d58JBNrLEkmuWaBnM3ia9U2lh8T+FdNU09fWeibFCFAzi64xnRsTJ9PtfxS7m
+qSMt9XsVClmPbKK0wET0Bd5fQBfJ5e4u5LhkUei4dxDiAyAU1v6hcb8KsWaU1at
9Hdu6XpONFMR2brIlYSIuV1A74g+Jj/pEfJmhR+rNG5dz/WGO9fM3h7Z9wqnR/WC
hnwkKKaUm5e2lsd++7Z9dMT10aAzrPi6vVb/7x277wSmZYSc+7jbd/T4xyubcqwy
vMcDzEok0Pkp2TpQYS0w2wQ3260BwvnWP2l6qQFH+KTqBrnLLFDvlx/+4RDOJcR+
UGoNIteXxb0z9WSEjqlFx071j20vid6Oq9/EIXy12X4RfE0XJwd8Yq82kN1s3l/R
vd07ggrxzKdpxFJqbD4zk1L0Ed8DEzytB4EctBqZxJKDr6ykWjRhj0gp5IUsjnTf
qNcv41AXg8NK6KWXgcavg1a1q4mgbSphApWHHz6EEIAqkq87AIFzmmIwBw44Zbel
8dKdS9i9WkG5+tzRyo97S2fG9oqO5bAHcaKW7WLpXfmxj/IO5WPXmHlwqGF4GTQY
rxuC3gU1LDOuWcginNtviALLjqyjjqMHAgG11RxxzoH39dcNA/KFHJXVE6hVXyYq
iiJuanPsWbY6kAUqQrw6L4uIry01ggFfDXXY8beI+n50Dgs/cRlRa6Al/D2HC3A8
5+lsY7AOJYD1r9B1/XBFWPpMl6w3W3+U9/rmb5g6660x8CzUSvJyhG3OFD2lN2eg
7JEc/t7wNOz6AyJM86lpCqVBVCQbk5wikP0C2PmiwYSiMEp+L2Bvozd8HOq/4Xfa
VKYa1HschYetAZNixHxBmZpnKCajinXI6ZyFGJvP8efZmycyjA1QvUOIGmoF/Z28
JUAJ0laDYvfcdClk5qbtPLkueBpfQzK8pxoz45sDeVINPgnIaefO4fi8FSCkd94J
5oMN4MykWQn+R7ou1mj95SToAPM7YSqkjCTDHJx9nfQSzOscFpaJLSFHkJmturEa
21EW2zL4/HmDEFvL7KbdHmawBr/3MSIAVIPOsyvDEgFYYKJmMoSSQVB+oqNmgLbW
uedtMJQRDTSThbhGjmcFs8wtzr6x+pwVmIs9wT62acITBZm71FHyke/gmRTd4def
HDgey6N9zkfD6jNSsjtATEjw7lQxV4ozCg+t+qKCR5u+llrhKeB8sohAXOOw5rQd
5/r6wOVjnOvFvxJOFdil6bXbv1szOrJ6H93ZBSkqp1ZsDq2Sw+W8UhxyBJsNC9ob
ZWv+RzEOyl7/ZGgB5jJZkNLzYlZLGSrFWMcSS0UQrkoDyeNNPe1fj90Y5FxaLJAQ
FhXEPhgsXPT+sdYAAGQB9SYDqCG4E5MzbbY/osF6ysWwExFg5KyoXjY0uKkkktHE
TpIu7i6r//ZzzWsMyi1LUwPoASX+ale8fHHuuAf1IoBn4/BIH0VhqCNuZSSYddut
GaVRJvA6iZ2wT42wStNLy4CWJFzWablLcMjRE5K3e4o1piCOREu8EbGB5bQ3h7Cc
8yEkXR8xtvBIRHSYecBWuL7RCu5DJYYlh3UdkTCnEmzOXwDTz+bH9SS0c3OpuDmI
jf/5aKZ/3nQaewIYx+6eO1fQ7LZNqaUObTA1nDF65NB1W2P/juz7cbBVg9wnRPv2
AE/BBuYFoJ+mkhwOjV8Tk/OZQcTj3UB/XfDeqiRnT0BOfl3VOEzcFRSkLET0akmF
Ra4qLudtWCRGWM2nR/YbmaoLhdYEtqAwKYWCNHNOckI3bCgmwDA48aU+8RyQG6NY
FuiNim9WJUQdqJrYzcf50cJqgiuG4M3SmaBu4PFbRUgq7C7UqH7hABU6wfa+dR2d
Yr4aQ3MCAc/ubkC1O7L5oNskj8pSmQR6cdAZtRm/rMacvMui5yul+FwkrZqNnhGH
hEOTft2P8wn0DA6Du8HszhOSYx638i1cMC65OoynzSDW0FF+YC5QSW1MZoHIKRjf
WMF1lDJYF3fgr5c9Zth5X3TOvpkcHcaGxvcK4li3lfk2DZ1Pj4wWzHvvlYf/ALu0
+qZ8BNCObcZNEDwBfibFiUBaxyehdJYoVRoAMxRhzoO24K9yW+KIezOmuS1diCNw
lmCe9ahe26FgCNfiQy8LCcP+zRMUfyAMm497+8t8ZG1B65hcNxTyMkSGts5b3d4U
YPhxiPn0qbYAv1u9YIbJqcodbqC3I1BXlZky4zkCh5BY7Px6NAUm4HTBQhDT/V7B
4PT/ouBWJ2cbDfBUD9q2y+IaD2fne1RXg/4d/l9Ttu9CZJxvehnYdeZE0Y5y8XaR
BvMqEUm9MzNW102eU9QfRXI+QjIUAPdSKxq5ntrkPZp63gQyQxCzwP5JbaJfT6dF
eCeWa5vWQ8KZ7J4eOlqml8dty406jSSa4egW94cH2WDI6YpzicAHeZ+ZKnq4F7zb
7SS03Njwk0yeCazv3mF1eaT3UtY1hc6AMDs7YBjYcwAicg+RtuHPqWtpA9nC1YNU
bPwetfH0bJsOUH3rU4K19mNIRx7abTXhjhu4Vq9drcJlwL16Xpm5r3kVI1fzowaf
ugj4Om14NhXmTrch8bz14X3BOGMNVor/2zduYs8FL6YqnctJNk5ELs1HIqz5+LG/
0iZhC0pJrKFV9qgyauxzTqznEWhW9G/TFg1FL1XfElE5xN2miGVyta8wgPxR4wMc
dIp+eEGJpevgQNU6rCg45Pzp+PzuEOYfOhhUtUHo++VhYgbHBI7pCqJWkfZFLk46
kY04NI6jBvhdzpgklm81wPCOfgxptb+OJUF9WmWF/ohGMuqqVy+MtPEqTaBGCtOv
62zhfSNs8vU7PvguqJNbd9sl+//A2YX6wJoS1kAyDZQRCTZjwuEY6e+nSQ4gf+mi
ThZcylr4ZojRLPRZJ5+8SD7l1mm2HHKvsgMHxTUAzhambH4SI+F6XHMic2vcoBHd
YNzWTlCyKvuZgwtF/i/SJtJDSMDZV0ybo9rdRlx2RdV6OjcvcOISoT8Do3h9PS35
x22KCh1Pr3jjhsi70CA47JZQINiCwuexrwYaw9TXk05UwqNf/MUkSwqP54T174jD
hER9eLSle8ee0hNATHLg0cFDIpTaSyxRkUtk9uHArpIst0eu7ulfKyt0msicSWPr
o3ExhX3r+8+AoXJzCD8ICkJdtutwGn1/YTs11Ugc3IXnpYKna5ZnEKwuXDC8wMp1
6MzWJsDBO8Y1kLayswu0GMXzEa0Avql/BCkEJX8idW24CoqGWPBZmAWnVyMjlQvF
Pxut5oxJsYwftboZ51oBqakhH5u57TxF9FJDPdW19g1S4s8UiHqL81JVcKhrnR3U
lOP0dl+O2LMAvXSgGyaZk9njzm9ufOAsPdBAJA7GTTG+8lYUSFqF/yyti14QP0aa
n8H2cfoiJjREwHvB3mtWOHAh6Ub9adT/63E9/BHG6BWf4EqGLgYUUCammrYR5pPj
wWtgnmMNyHjkSxREXfRWJVO/+Ky+aC3ZodzRBcJBGbPaP+yNx6eL8kJGkWlwi27P
iR5uz9wHh2A8lGopTRsr6a4He1V167N7bTZJbKfch/Ki6EU/eqrPd4E+ACV3OY8I
Ppty1HBpgjE/yFOVWc6IbNrfIN15Sk2GQ4xvLVxG6EfqviinS+KqCbImSaC6rSD4
yvIgmF34n6cMXGZypnKpnIBLb1BxtnO6iGH+0xygEdfI9nLmkD5TXj6iu+sc3dx/
LKaBn7glaHsEi/v4WTopywpgTPxc44gFht18MQnhMVsocEb2gJv+TodRq4JPNWlv
QzGPphN/lIMrFSwNxIujdoad0jx/JzGDWlT3uTHZyqJCbEC+EPx+ct/b6ePgVHcB
ULtfRd75XeFqaq0pYLQxRZN2WTTtYDwERDa6IWWC+l1weeHWz810TRCTonZAr+ca
eWUCP8KSrehIrYcsr3rxM5X+D50ZBeRHM29gm30Vslucpyg489hkocV6c+xG5D7b
rDp6Tg1gCTe+FHjpjy8a0Gg113GKuV1iyCY31/HdQ6gm838Ama/OM8ny7XZ5Fq97
feGn+FAdktnE7MzIg9shvV4vP2LQGD3iW0PLG20WKp+xvDyYpHFCMc/oRwCB43yz
lHXvduK0Pn3ZQcICdAj3orHy+O3OC2Gx6MNiYYhaqUpejMLTYtwolnpdu3YT78JU
EimIDE4aolEa68+t1JXcfboA9AzQRwmT5NdAbSavE25EI+yVNM6sTtxvNLMYEToo
VBN5aIE2v45MOzhheDrfm4Ft3NO07uMOmicPmBNzGwOVRW4ErsPabtu1gmSJ8w6v
+AiG/INatJCw04KQlOdE5QpyxMF7Ha1YeqmSy6jRKe3edCzLQas0TD8TAwk/0L7k
2SrIah/W2XWbALkJLeoU7qNgLo9Xe0sZct2l+888RwapDo2vSfE/DNTbojh0exHs
Vfd9kmZYdm1UA+qDhiOTY/FFBMlJumZGqNr68nQ1fPxJpjKGVCYHoQV2bb0YXNXx
TuCsSRU+DwKSHrFtMD2jVSIwnWt+wyUjjf1/MgCBzBGYold18/31sP6POAnCiGaZ
MVnIwuLjNiwYB/ltrDNhy0KjeqF0iiy7ZmuZnp/TwJxP8vSHnUSceCFQzLarccuN
IObn9JKaH6msJO2B4VKOEnSwuwDw3jeZT+y2XCbMVXdFs3fLRIrC6uhjqp/ZkSop
Dw5CP8zDzIfcIcTIjj41jkKJk8SleTsSizUUFhf8/yCk2N4vYC0xfWvmGLBbNcOd
f8gEj8z6HdbULdFmyfNVtR3QJ2xvlYajFEFuYmrZjwiJuoA6QCQGRKCNec1GSO3t
uPusfYrNdbYEscUi4VTVAoFBjIr5r21eEG4EL9j1B4oADYS34J2ifyqtpXTTlaQd
xqTbpr+6Uz2BLpatAx7CIe8WOGMQWVxKN/PU5ef+QhF0+1iBkdkXUmi7Qx0rjt1F
5s3lIga2+tb06VkUaMrGMBPmGAuJMcSMY4ZTDqwU4nclCKQ0EV3GOKDpyvPqIloK
UD8mI2Qfo0zIh7eu4K+O0lLFryqUt4M9IKea0zrwTTeQ80FEzeNHzJa8xPRAUgBi
6c8Eors7hMHXLx+QU8kGYesyeltFrGp17Gl0+nfYFB4wLvMSfpktlMZ6FHSMjjVy
kfsTjHyDjzQnKfb14mC3Kd1QNw/G80C/Y4BC1Vy+pZ0APn12rnyYJ8z4KHDXZNOV
4PGUBeWKKGpAWBIh5LRVX01UCaPFEBcicKNAidLXWiKg4mQh1T+3estk6nYcHn5+
bRxWGvqpnrn3a1W1by7ORoG+jB2E4GkOolSNTY18fuUTZyHuAHLurc4NeIcEYZ0t
YCmFS/qZaQJL2T35jObU9qbOq8TmyEErisdoHqttbvDkGObEu2P1RMa2U6ISmG2r
Pp9UPWbdU7TsNX7O9ELDLpInpoZNKPvZzvFPS7i+6YLsI2XFY7ooAorLTnX2eWGp
lai3vklqfVj96hxyK1by/6w9dDOCM72xV6vuKT6E3nf0bJqS4tKLKkeLtSrokZOD
TldLY8uLbaw6S+4jvEewt/02AY7YbGpY6gGOebbJX701nL6xgNRzbRsiYiZl1Pzh
jXT1jNcghAiqAsKkuhAtptOluGteWUf/wZxV+EUyhj0J89TPv8O4fdXX8JNwF2RY
XAquNPlf51rwaSFgpxAIgy6vFs5EDkwW0QjPQIaX92ik4TccR2T5yOMQRCOGVQtZ
b2+gihknoiLfKDplIGemRZChe/r3X8lHcSx6xkGWImuwX8KOq8jUMxj7+rA9RyR2
m703QZ4LOpdNBtPC3dG3s73dOkp/iEM4pWF0F3XVAIGc32WH2QgYoNwoQoY5efyG
BwHl9FeeNHKTTTwVnheCxshxyMa4tocRsIxZquiNJQX8/30dqLJ7heP5dpn2DxGg
/4RD6pqiy6luVG3BoY2n+m4pJaR5xAAXDg2/kyINxRoc/Oq5j9B3nf4/jyRBW9kA
Yoj40nqrEz09nSIHWkAT+88kapKJL/StJuxSZtPqTaSQkw51GcMr2hVbYhV0Ibgp
2bZWXmytsZmqzZf+0NfGPtOTPE5VOfmPZH5racTVvyRbpWHXR4tPvNj+AXUnmEtR
f+hBanH5kqC3gQPwD/C2JvD4ZCiwIkSZq9l9eYCop208XWdK5hUjF9rug7ZvUBVZ
dbI3yi0mMuGtWFYTgLh94SyBwwEHFrYxNwz9JE/15L40QR6Y2WdRmNLepwiWxzdD
l9poqQ1CWqSJ1uCuobGKEnwpsZes9zhF6IMK3xDMPFn/jCN37YQOTQpC+7FyH7SZ
A4nOoOQy7CylOT+GUQaf9dQLpmuFYoiwVtG+cLeYx5LMpbtNb+9x4oEHDB5cDr8q
tqw0QKATFx+E8/fpiZyMWeODjiUxl4kAYzZQRGhmwTfz77d+yRwOKJa1NaubQ/HO
0DjAHPUY38GShrpufG038iZxztDWbhTxG0Erz5QfgWcOy2+sQkfgkn1omzqkrQO/
7bEZqEBGAtIOrYCEOiVK5LD63IPiJdDtjN4nmTRuf0OR2VOZvZQCODF2mX43yiSP
0wrwPZeCh1GQOgAMDDX7cg90O4HOamWtQPPVzzXGkFljryVmTZGoM13CS1nvUNCc
uGp6RjAcx1jmFyaP4H/QkhEvBG/oqFIKjQSY/lo9msvpR+nhrqpZtDK1XVs9xY8Y
dOtVBXKp/xj5Vak4dDBlyMYI9YcoG5p47eD8HvSswAtphlw44iqghqDMPRwUuLFN
/Q7GjUvusRq0mZY44bkQIiexAgZDO3XLqJnGHHd7z0aQbkCsww6+VOHT+aLbD96x
eFbfa2vML62PI++XA8QXM+dbuCXgs0jxhrr3ZGYO6mitJRsQWqmAhJJOqrj0usho
U6V9VpSouvSqd9oloPC2iK/miHgMXU8WwvQuIiR8eW8v6ewS+0cp5AO1IZa31WoL
Hw3t3rRB4hPyRDOaQAsedZ3bEQqOFKHixnSCjmilCJM3xeJrBABPRDWSrctQ/Js+
3qWscVbAn+2tpoWqK1HXjT0WRb/9Wen3txFXsbDv1eCVBFDt2+c4/lJu6rOzELtK
kDmupak8+a4qsPUMg/C/oe8t702Bv1XH8eK3vNLhPc6m+FrQbhAV199GmXl7Zq7A
OPDUuvDODLYZqfEH5r4Su0qUzrxhKRNwT3e7HreHtb/HiZUwyzG0o6Uhw6UuX+3E
thQBUzi4bpIkbL9O5m90Y0nXGOYsTzG+kAEplzS3IMKtG1eB/1oXiK0JSMLntuKX
Udc16Jopaa/BksEZwIW9hNB/Y3/5ECVWxyNGhqN43UP25ql842Ti58u0ylFeqHQP
jWhaipZPvdYzuiVOvgS7X9px8lk+qEfKJxxz0XN1ya6Np/pla3XB92/XU+10igSn
4ULdwGUHhkeEVXvmHmQL2HiTjAFFr3M3Afc6RAjayW5hf7KZwo1eqKxjKrCFUNIF
tAM7CsUxg6q5MSCeT0nyQFR5Vq76jpABrcs64StB1is+3fqzqrskUjbiM1hGEMZS
0jF0ibSfvq2C3IcWIX+jmxK+jMMk8l3dt6r1BN08uIMJZ5xC08d3va4MjK7vRrLS
XB4coljp9HbPnH8SYKHbqohMOi+Ji8Er7MAH0kfXXrKkqsgjNf0RNtKy2E2n2KIy
PmsWmB8V/pFweszmk4QIb5vawb/f95Ep3uEbM5ZghsYnfz0gzu1fMz/3bGaHTml+
kjZ2bE7GmaXYwUQEftTmO3cQG5Po0IB/JuY8Ik/AzABHWxVBEV/pyLRuySlR0Ks8
SN/U24Yzp0NDyIRpSsXWJm8JczalaRyTtdBZFYbDhV4qkgl6rRGjL/QvwkLgv4Uv
Eakbn3tmyKYh2w9KrVwEEZZhvJgcFo9LajxD+PvKTf4m7AK3ZJ5BUC6o8QoD66h7
A2Lyy7y09DXEBe5xSAB0Zph3xgRWsbjaUkQK+YhrxHZDXXVDZ0ml9uF+Z48TL0gd
sUuddXU3Rw7uRw86vE5ZDWoCKFxblQ2bSc0G/PF6JlusYrTabQX3RY6a20oYYexu
oodRVITy5HSUEHaCPgQ6kIVxMT9y5DAftFYfzuWktfMALNjPkwxBSxatxC/I48xI
pp+Yddl0rENNaxCicsJMQYYxafdOf+FkbCw4x81kSNWB05XpFWPkf6JPzgvXbqpT
1eCrNRRKMP9qMQyGIIvr3exCNgAWKKRQ1ShrUx8rTOOyPltBFSq5NRet3QLjQtK+
HwORCzpOLZ3VXr/SLkUuIv1uvwx+TL3DA6Hxojy1AOfsj6Ui1Io+ymB6FPnS/lCn
WGmFTbJk7zfpnytcxQuEqOsDgUrl07u38cFJKOQbAWvozjqryVIWNB2B325UzDRu
95/F+Qk/ggVZhcYULWiccMkXlm/eRcuT0BGWAVMdpn+RooUXvRD+Ix5twssaKfnC
A/kUIo/r/UcroAVPnwGCr4LmNbfHFijIrBtqFIsyZYwWzTa+o+t3zgrHuyjxE3If
eMh8qBpQDWPjs2/ColiWR/s+ffM3pSQBqBE0BwWPLtAAliauCVYxr9xkgc9TFIsG
S7UbbEr0mQRyw0621mmoX7ppQIYj86G/7nDBOlTCFuL5Hn2+RcTcaxayvQOZWwhg
5KcX8BU9uCrmJmZapjETrrJFOuSYGcT4n+ymNDWEvzuvT3TTxzTgr/soTKDcmZun
XtM1kx2qERcCU1ilvMmO4TBnmXv8xDxg/8OXZQaR/zZRHlzIeEOaTjeo1VSKIj+I
NHTU+F5estesU117dKpbPBNBxXZTgXi7K6irjuwn5a8243tskWRmU758A56bK0BO
bvgbBooMaOKC8eXai/t3RmPediha1ilCBrlXpncce+qK5eYROWsZb4xn+qtp4jxe
D6Lc8Wrjh8S154CVu2rNRcC10a4hcNyLXk5SAcpU5JB93yooFZq+rkBuN9m2RVzX
Ty0WvYl3JWF53sVLDNlwW5FZO4/ykGYx08VgjRgPa0fFzcQf3A4Fo77qsRl2iZK8
2V3eJD3nRvQBsEhlzH631/4IPPw9PsBuAve9oFs75qTg/5NyZg5icPFCgv5QWUHg
hS8Zudhqf+jdhG7vMUZtv0fitNw+KHbe88onlVqmVIn6ZNeLeJC3IrhddCmXjtLF
B5QJQT9fM/+c5VR76HW1MEx7iQtf79LCZYIjYVAFLTcnnxCbBX3gqZ1D8er4Vo0h
41ekdfA2CUSN79A4dLpMqMbtghYhTMK/iTK6X8/hsvxD9Ybfz38bfXncUuigPwv9
R51pUu7hoDlC/iK9E3QTDCO5/u048W2Pfp+tnqs+hkzNkJZyXf1oEJwfsqXx8QfO
sl1mQ2538SNb/34hUA6s2EcyATtfZV2J20vKK2XgoodJZD62b9Iw+QJ6BtRxL5wV
e3+/oeuKOfY/WfHm2qh+EYFDxr4Cz1T/dx9q67VWfLQkMun9dPn+DiynBVQNHitx
u6SlBvNchwHLFt823ZcqSXILgf7eJWRv+OfhQ9HZFbfm0S5lPKSfzdwUuTE3xTAQ
H76/LT7PqBAVud9bujAltI/7eTA+/GHDagqcFb59pQMRm4BGAGl0+L8EaKS1KRDn
eJSO8RUfwRzpclRCcHRie7mRHwQRnXxxDhNKv61iRSr7oqmTGiHEtf1O2LbbFPit
pNO7krSeQ3iocY0rY59sL/7cm9UpY/SXKDQJBfkdRvmoqiDatwzgLIb6WtcJ0rOL
Z1JzVyFuDlgRcMsjkMih4hOukqbrPtGgZ3nRJD+8sgipSt+th901gtOHIQhvvtPA
0DBKcnVrfmX1ji8z2Mpq2GleTcuf9T9HQq6Qnx8iuMIV1PiS4v143SUrZfV6AacF
k6LzWmqif1eKGDF2wb6jsXJe4+KBDqdR17aHaWqoGxLotqFwqHQZvwGaoipg1d3o
tDM+aW1oML34dc31UZUMh3K/umtplkeYB5Y2SMuojyTvsgiF/0BIDid0tS8t6b2b
kupwqf1a7zf33QjfyHFXKU584B6U+hBsowhdo3W6DdV+b8Zm/0bF+XXV0Ql5VqgT
WqxLklvUarAPR6YW/lOUpkotFChD/vvPY8wI5CLGtzD5vOyAcPzm4YRFal2DEt+M
tE2dglLjYXxsR08ZIdL5EHb02m6MpO0eKcLcNldrAbBE0erYBEmU7Ye1iTF4qhZC
Hd9c3MM7snvjnJj0L0v0e+ETol1WHMhXM3H9CdgXBRxMkqSIN6a7wOWI6Rd0clZJ
BORjr8JW8AhtJou0ewcW+YMSr7xLti8QUkhUMxsypuDZgU5wZQMvULUaC9ANR9Rt
3CfOQjn17K0GynA05KjfCGezKtP4X06u6AyqqIrWNM350zLLg+h3CFMbwONGUxGU
13t/p8xydZ2xV3819CDQ7NZnleiqMVW5RJusrLcm42eDe4Zo1qcas6/XZZFruWXn
/hrQERXGjf536MeR1iVqMcSYvIAov08Bf7sZMB2u0ukjqVSQaoklvoUS0k/6RsLm
mOowQjvh1TpOkm/SBwkjlT6KpNHxxyOuXFaYdWumF1rkjtku8ExBzveWFoKsAjAA
hUieMOE+XsVVburaflTiVoNZyZbiNnGEtkkqKGzw8z3Wzx//Bjzpo4+0ZY0zH4az
ai3E9IvC1w6LMipmKc6Rn8kPzp6I2I7zaWu1OiOm9sIpEthCU2PvA7qvsD61ZkNW
Q2QGCXIvkDCu7UJzn2hSuxJvJ+oJeK6gYr82L/sNQhSNAPJo7RxlLFlN0IRk0YFl
SLRUZFMbbW/17mf66aIWDqxqIW7cGAHhJaJ5e08bhUc0K+7Sb9rPEZEX2WlHPcz+
Wzlhc3xdmXWSKn+1JBhevxbXyGRzvvFJux8+qbvHXU+tI2HFlCM2uT58lFYXk6Vw
vKRA+/lpDZ21i/V4O/HBtBx/tnaX/nrzVsXZTOHlxVnJKmqOjHwVyA2dMsoKGMQ9
8iHH6GLw1OeEARQknUpic/amwITcCANFpfH6KfD6UdAKpdWJ1mLIj20x8bdvHx08
4cRsKOgSXGPWdBwAB5lPGabYKsXE4Be8WjbnX4ZHAvP88hpdLmgIZ/tnlzmb8N5D
9nsboLdOjPCxjWIBVmCDKx6czwYw9xU9WLF47fkUckIr2/SqIMJ5FkN5rdRNs8nd
UKv3HzzDyELXyrvWh6oKkupbzOsoVIqhYLId6j7VrX3voaJ1TbBb5IT005mHaoP1
Aal/ZVRE+RoGsLDyaEUm6XkuZjj2p5YEtWo+0+uaDm1xOZAKcRPPeXaspEfRzkbx
VTxkBLqbkdA5YFr8Da5cESZSNQry1uPXCb/k2LqCJ1alR7ldyt8PnSkX7nwr1Tm2
xWBi1sMdGTh5Q89yiu/gCgg90q5Kn03Uoq4jxRKcMVLvcZAvxf6eaYNcc/LMK8Iy
LFDjcVwqA0Iba48iBbbDMBiqwOfUP6RK47IHuiIfVFwy7oEQ3fGBiuwcnEcQS7nw
q+q0EYcb33czpRPVj+aFDRjV1s5lhYcA9/Tni84w13u4YOILCWNMLWE7qXRdBiYZ
y91/3qpH+uiKWTZpqI0+55W+LCW0aP1F+oYlClenX6SJV3J7fd1X9bmvKQFKrToE
6UFW2XxjbS9ihz/u+uR5O3P/ffUfXXnBDxodsvFoAU6OoRbaDlvvhpXpPHy2Wxa3
Y5Hw9XxQ15cpHF1DW9+d6m+ACOsgxzjYWpiHY9xgW5Nupq+L0diyUz96WvpxKedK
86G445C+1QxQ+muowzMgodk11fZn02I7d6e9ZYDA2Wn4Gf1clJfvZas3B+B7/m7s
l+CB7VWbZ2xK+t8eW6icWKMHdnqDSqb4dqyZizFQRt8v/JvzZZ5VH6MKSa7kTqab
+7GzvsowoNEnEb57PjXxtxyVDKQh38ta6Nj80D42zGw5qBWn5XOY6Lyt/dHZKtbE
H7taprBywGWbILLgwsMXQeEgePHND+kVL87OAK5d3mJer4qtVyjO1GXuC9LClGL5
Ea2qV7az1LKoA+8mriHTk9O40ocFLoi25o8EJmBoPsHxL47UXb0ZsspetRBxmFaL
82gTQdqwvHRF7YttYuOOrDAWYo29Z8YR2+v7JBFa9RxMC7OcvNtk7u9F8L7rFad8
EcJDFm6enJW3pbgf4+tdfa0HSvoNMWXGNcUEDW9vH11EWTnoTYgvQfW0DxxCaiWG
34uNH4/q7/IDUsGFK1/wHiug4vkg0fJCRKYaJDzdOc9vIJmXs+WUpisjboZBPMRg
ibJTLFVJft534ol4PVmBSnVRBiB6K/wHamJBcySJa9RN9i6T9gHDGDSPrOdNEDln
C4+lJa2s3WvskH1+8p+XWtQaU7xDpKlkhCjsoewz/cz4cQfmy0A438Ntem21MRla
1sQ6eCmKVOJbPytMFoLx03Dzrs2AIVt/aPKNZkeiNexrS8RMPKYRYYEoVQgWwpAJ
mr8LZtPqSMSQLUS5o6nmfYJoWCPiyxI8uQHpWoZ+d67a79uQkt9+e4XdM+QSOlJp
NatRv8iPQsm3h5I7Vpw6QNDfpPUVISzWrh84r9SueEsHXKTGIBbYnq4Cm+mpOk0l
BhFpYWk6d/kW2/Y6cJPs0x9rlUIyHhFPWpcAmvBUSR+UmgdyrZPvoOuzf58tygXd
NDG58Ngr2Z1ccKYo3gur+I9riZTcFb4fv4AqZ4oZAl7o+qsmOtuHAR8IvgGectCJ
3fsME2s9/+vtU/q/Tbwn0ejh0uoxbk+RSEx8pJOC6SKzVxqSkkknk5xRnNeCAvwF
XuLOq5UeJ+oeFr/ulPMJ2LQRNNO8GUPjyntJ1G6KSjAj3DWrJYheCbsxwSWW9w6U
wyddANkXS1a4364PtBe3owt93n2YR0D3PbaB5KeR+DR8jex+eomertVh4+SrSX1q
Bvenvags5euD+DKuJP19FF6Glw/DGrEpIzhglV4oBLoQKDopt+w4csEffigzVzVe
wwejY84DvHoPVYukceEoeHDEr7LMbIIKAKYExbZo+g6qmJf0niJetQcA3fcZ6gyW
Pw9YW3ecWojRwZkO7H0fKHTfBw9gh4gGIapKJp11gAuLEzjeSSX0buGybZ9H+0Fc
sBprTwY4oM98GWeTf1r9NN3y6We1MfdVzMrs7c9s+DCD4QWNPzR6Gqc9sqApF3lY
JeaXhkhMbRGUavI4ILms2wrjRBCobALzlj18T1KmVtOJ41AFLaYSOQ3M2QgSpIMp
BbPow3ZJI+RnKkCPYGB3QEgpKcAAvF7kLHZZoNmZNXde3vQ/dg/Hkbrj52VaO2nm
SlnwnSNtzxdgZ5rUdsOnTS1VQ9+9ge0xZ1UpuSxhZ3uDCBRuJWmjOONmhL9h4VoV
nxT8ZMGzuvilkvhp4ruqs7ASoAKthH+dEhLBabaN6ex9LHzIm2/8mCOgdwmHZnAO
6vJdqcXFRYPTJPe7mGGY8ee+yyX92iYovt8Xi/qYoBpZ4EpiK634/Oin+7ml20I/
5d9hNFiotMl9EuTUHgb20/MCsUjNL3QtQEjEFlyM/LUvrxRCz5EEacbYAdIG7qZN
9AdmwgGeqR1yQHYkrW0Hw4eAYzFOYuTzzRxMDClN1C2MNP83cvYxoDRWaWomgQ89
DwGgLtxzG3Ca+n09aok33hypi/0D4sbp4bs5qnvT2oFcVeXSV4riJ/676JyiSixs
SSaWUvV0hZTzMLvyScH54duA3X7KsVsQdjuJNPEGuLxvuVe6dZM10usQVJYyqtiH
R7PDbuauzwjV757VuyD2hVmFC8pLoOzmH2sg2BE11e4bl3Li2s0uAfAM8u1SFkCr
GeQ9Ngz11+Bv0DWMLPADPz6oP6Tj1utG3dpJIltka1l0WcBg63n6s7x0u6p69s9S
atJTxOFaFItdTQjHYtj1gkaSvFJuuIqMCUT3TptkYe6S6+sTrq90YvOQIMX3jl1A
haJJcelEvZwIohYT47V82ELd3c0dG5Mw2rWM5E/bUNkGBXjoiwZ1Xh7Zlm8EdOEl
LLcSmcrDDqB98Te8jgUciveK3L1YWEG1x5tMKl0Ouzw9JDSYkLQ7+SmwPObOgyml
NdEBneEnaSaLd3QgLjdDQhBo1jZiUOqxg1RJeUlMT7KdO9DTEeiDFFVyQXK6ByvG
GmXUKcbIzNvgaXYqCKGckKUpovH5W9m0cgstcVcIMrVsAvxpDqj2W8UvMnyQ4MaK
arD8lX4R1RmGx7GePE9lxV4P3xss00JHfQLQqwNZlTLDvEDfDELU+ME0SlB+d5UO
coAMrz+DVJr/egqiUTYgDpJhH19fDWvYjqUZzAE/23hP2sp6vMLkKJnF1UyvijIh
VA1s0GG6A3/YV6Ke2XfQdZvEQdhJzj2Sq8WKyqWadyqj6zSaJrvykidILoDEj1LJ
VYHbuIKEIGKGRClwlLfIqBneXVB9ki1Cjria4L32zlCIHw6F/uWk612lxOwpQZ97
8vfG4kkOOGrP0syqnc7789Pzz1AnjK7k3jlu/lDy1CHUfJSCyMJQin6MaumdOqw+
Y2k2Sd9tcs5NXHPwp1NCH1W14s/cD6UyiXObvejSa8TGp6YiugvHbt6Wow3qwyr+
cgR3m4QtnMi+wQy5H1ZhizGKLLc1Ed94pOIJzxy9xoeSMjpYEe1Dl99NDUJLpEb+
TYBI4deIf5vekUkpIobtsHD4ipnFTWgSZdA+s48e/LLdxUbjH2xPp+CdmJIyuygg
jgfOcpvVp2CmC5aMMENwYLbAZJxLXmr9+wQMrFZNKVuEYW8RHcrkZ4qMeSne48w5
/fAmcEnaaLvc+aM8UqCKoM9N6APflDG2h1rCyD426rxId66Lok+6jxkR6ViZ2C3y
AYrZYPMskBMp1SNmSzmP93V+5a9UQCsm4U+kTvAfXdqQ5lX1KL+1vSZEBwAYrW/+
PFO9udITdmjtqb++s5ePp4olTWuE53vU+PnSYvePMypPPRTSEj904rj+IOcTRbLC
pMGQ+PTNz+rH/0BTLyAFNFvgsuAQEor59wNYlVJer4uiXLH/lgaUrAAZvvvyavEV
XxxcqTRMJNdjU2G+jL6ZffWTadMhYiUHRPaYlqKDmQaZgAgSDdWiYzgheD5ZwOX5
P9ZoSYySG/YM/dzqWZUYSVWxdfe7oHDINdpl5To9R8+meAmqCuTb4OR+sqwRHwvr
pHVZA/I0nLR2PpWahrjIHoRSSiYfK9SVpE0jzRISXwSp5PHA8Am+ZdmMP8vlT3Iq
6Szz8LZCki760GqG+s9ULFN1c8Y6CEUQqXL2O03rOkIYBpvtRyrqHGTB6+dS5U3v
fsw0D3M1UDayiakMuxq3kn/XiVjRXSNfNQIGXBXArjxvC28uJbjKBTbYrWIwxcAy
xhYUaKgCDyQPdOJC7OKwSf8OEVXpNkIc+yjTNwXRqBfED3YLedsSbNvdnYIqVBbE
rx0SjtT5me9u23OZANnWq8N2DdOYxG+q4BgSaX0YaSQhPP+H8V49H4b69G79U2MZ
JcjqyhEVUheLXfRY6ySYTScsLYmQVhvZrCMw7C5o9Bl6QoBbPH5rLuJWSkkA2Zab
b0ofhAy6Hn/kGgr5Ol/y/27+Xqv9KoSxGE6Brh2WbavOpGGt8DsdhK8ooF1CWqzO
4b7v4rTmfvlSUDUHcKCsqM0ZyrEVVQi9/3AndbB30b3uwloYmO6Frh7Kg6t/VFzq
6Wi3Ns5uvGcsoqtYiCFpvHeGikI3X40EvOTcnkUJHzBdo472whoXYgEX4LM2DpxU
kNKmYTBa31dinM5a7bUlbPjPGUU495gsSO1x0DZDnAZ+Yj81JCJNAt7EbhCgDAzP
OQN1Wk56fYPtc1Dj+x6h88jqZ9ECeK+CsWo77UCv+eSS3na0A6b8b7+VOYlkNwBu
ANmbYc2A58b5f170sscX/8t7Px9/smUwRZcxZu3WOlGsdS/LvO6kgjy8eCyGpCMU
W1HKc6p9gM4TtbP+ffP0Crw0rXTsmPmKOsBvY+ldS1dAmD6yrOMU4j670DzGZwOf
EKh9MO0BQrbirK4RRerFzrkl9bq6gmmF4gBzbfPr/QVJGUc1gRkWQ5vfZ4ZfTemP
2wxlbeChvnRmKzFyy8uAHs9lz64tBL2eaTJwKJE9fzMva0UYIDcvjiizKkBlkPIM
uFULMGSRcX6d7gBnlRlqUe6FGacWIzZsR6GmNqQoo0UL1Xafv3Hw7cHEFsX24sjK
VAlX/X/LK1EwSgj1PAi/Xb0sX5UsasCqbJBVrbGXZwZ1La1OL8luMGRecbxyJeOE
WUmsELuUam157iHe3HB2G6lB1SwwKEL9tmQP44++CvppoCt+FBn0SGOydsfmI4qc
QTbFttm1oOrc5gnNUeqBV4suxPC6JDWCutg/j/zWLd9cNA/KETM5CmWicbzixN+Z
vX/n0JV3aqhZv7xFHfyBEl4XmDdj9KdhNs+Yc7O9bROYBr8P0KKN+IVZE824S1f+
RQRvwFKtZIELNGUiIFSEp5fl9/uVskyaZ3T1x6fXsTmvz3S9PwBXO2jz4GGQp2cr
PFIU83qKsImbQgbvJUQtUxVp4G0/s/+sQx7FpZ9zJy6mTYyPpehg9H4t/TwQL1BD
eoBBGO5RRSEOkxOmuM1R1XqJMlzGZEXC64jUVLDeO+StS8olKGR7cqTiYk+PVC1c
zTPQHXElBTNB5ZQziCTKsdrN5m7O/R96trbK66Qyn42SkAvqOOPJ/NQwysWWO/Nt
LYGbBRzxqsP+ga0EGnU5UqY5NTFOoNeOtydpxg5m0zQ/L6WtGorMMIF3s1ZgXO7J
b9CdcWDXgZ1eeZxMfFtLpQvASIX/zeIq0EpkDrdrs+PC0ydx5zSmuTC/t/u61pex
nzKhtUB2ifDVnpUdCwP3C5t7WQ6LxsKsnSEF42/FuhePiQQiYCLUp8OFQwdA+Xmn
9nNkjkm8NgFCOsfWmxaBDH45i9keOLv14DT94Ayw+97GyZsdNhXqISAUFRucicfv
q8tWxrDYk6cwZKhjNSjy5k7bgno6u1SQ5RkXoV6L7zyhu5JvfKb4E9obUQG58gIv
Gz00XWjuhv8kBCMna54D6JuGfjcBYua3SU8ut9QHtxNuz5jm5qOksbrXSqEq0uva
zHQZmy1wzVJfgI20ku77xNd0FxSSNc3y/N3XSDkFtvLp1CU1OQE1o1ki3H8kRld+
ViuDWNkUUKZ+4bhqkoHtyt4yuk9dOOuGkmv6dEvdjQA7AgPS7vgzDpgVuG0N3BpT
9o8yUCYJQy7zccbPyfU3nAfx3MAEWRxCiH6pfVwI6DAdvu9Ry7uGbyi6ztqLdbve
7Hb34biflBjKlASHy6+pdnsganZEdYfhm40pSzZ5ZR1XC/rN3UmAUepmHzz0T+OL
CzYwIq7Q9PXNPfJkOcHzpyTdHizg72R7D/MzrFgssxCPCO6dtIGAMJWypA9YvDTe
D5qLEMQEp+0HCqJtrRdhTDR/AMvMWnjf0Tbv9/Agc0P1glj+uoCbh+aRxcvJfKVK
5yq6emSFFBv2JewqiMzXUU3pU5lh1qZwWKU0TbezzEpSlu2viPZJnzNAAZcg10dr
gNdtL8fLCDqp7Qn5eFskdhaWJSJqqubwsaXQrw7xZwvfOKlceJlDRDqj/xFHTeBl
0BPdaAuUwdMpNUQwYlwu7MA66ZkzzQku3uKHq5qIAKmwWWS65Z7ADWm1SLlQ/XtE
Lu+EHS3EqX8J0zvEQnrDoB47KO9F+B8A+LhGegM2pXzhHaSPaidA0GzOFXE4ACcl
cQn4RGonK7q8DuSjQAakAKcfucOZkSdkFN99sWLqR+5ZyKiP+SRwRpgIw4R1QVuR
hApwggjhZbPWYQtR8/9ZVjCQn5LifwlMBdmnbCo3bgI9lkhzwblTYBPUDlyw1wyZ
lfpwGvGCYJBZ/UcbqRjK2jxy5pGBr4MkdX7StXB6W8DgN3bb7LLTEgEkJwCG6OMU
4bUjqCZHYWNV+QuFwQuZE6T0pDhnSHZWJ4A66RgzvKUZUv2pkKjUabEE8zpkUtpR
GjE1ktWu5yAa+0aAB5y1RjmA5drQ85pWdhZIpYC3mwNjPgwXojWFaxAwD9mL2BP8
NONywiwxZFX5JwqeY76hNJlbffeAMC2TqLbfrqnC+iLyByTGPUivupoPZv4v3/07
vltvxq+S0wgFFAaya+UzFA+ht35NCg5tAzu/ii6qEvS+GxNrmPGmjq9wlAo0cg8p
2d7Tj57XXetlIBkohev/00vlfFj4+wbnCWypScVHzjNL3HyHJdswFhdE76FPyPZY
4nY/oZ7E41jrPDJjJd+JjMfVs1hrNuQA8WvQAXeWgppjQUcMRjWmrbxGpwMObDui
6k6KdaEOyFVXFuR4kS47s+HgghXGhsqW9jSe8qP2V2sW1xfhwP4A6F+EyjVhfoxE
itRnbqAM9UsQsCsuMNx/pyxNY9QJx8+fmxKB2OoPpO2v8LWHSK/QqPD7bgGWk26E
ZNkK7Sv1QAG5XxQBDm9IA9T0Qk6TxKBKSOUrIjP2y41yPvjd9Ap/Cs2wHRVtGTED
c4kw142WnngABVkBFKuUzMqOhSFlbxEOgPrlqAIX072QXRTQgD/ADFmHRNulzxSZ
QYz4lZx18qeb5bqUwoUYVE2rtBoruBTFvylHUfjKE0vdkv7T7nFSvKvPI/7nCA8A
SnFI0XZEvaTdacnS+F63fSlHQ1paYDqEK0hNoZwUmuIo5w94mEHr4s4Ca6OEECIl
ApBN11zD64aRmCF5Q51q2+v+CZJcB9iVwydr5uWE3GyfzmnuM2kVmp5LtY0BexA1
EvAOflyDLfBwaM6ZMj9FztKIT+xN20ewXs3y3RMAkEB0fNl3F1jNlDqPEwtvHDVX
NuLH5+JPtuweLTeZWgAEN2aHteZdf+p6aJPkNfMy0yvc48gZT20uUdJBF0ri7Ahz
ndj6OglpB4M6ONU8jCKNqwzhUISzVeE8izaate5OgAnqIWURZQEzl1NSkE552Bjj
oivQSEe2qNFGakP4W26sYWf39iWYeLwR1gwo8y5puC3NxFG+kIBV3E7HWVdxIU1Q
uGj5AQkqPl0InhbymI3a4/Vc2PSTuzYIYmRSZssP6cpB37TWNq8WNWyBDGbPCM9Y
qhDUSYJE6zix3vparcOCmKbw/QZMtpbkk445iy+ufVki8ZxmRDbH1cryzE4wR662
nCQq0DnyCD5KS+mQ/GzCNr52OWp9gpyh34kYft+ni8evX22M5RZuYtiGaleOnxEC
xNyAvwUZrEucKIlseQvrxK1HoYNVSDls7Me405NkG8j4UTan1iHtmECDbvhrW3HN
jtqjyEiLyQyJdm+zVkrrvADHRwd5dKjF/GN43ALJp7Fk6o6CKr9M7/2ZC+P4nuA/
dgAo5fkI5+IzAKVzm+aZHpa6S2rQzKa5Ea766w+YNziNm2CEqnLQgMc9BtBygQiD
HsHo63fMJx0XrhNoExjEh7odlXRB3HOdmiK0M2XAFz8lCP8jtWQpWH+AN97JBW2x
FaasAYUBqPK89ryVCoZmTK5RPyvxzJ/PMHzCKbay0GlBd5zjYKMctiKftjJm/kBm
lxNuw/kldNy0BrkWXk4PIQEv7wrPgnKxfjJ9QnoaxR8bkR3t4/Rq9L2/A+Gdfjcn
Tlffl6TrVvUHd3sdtIrGDgliSj2VcxmG8Ox6L7ei+Ck30qD0M8Wex9kNqmebkFLI
/gBGRqr3rUiCclLFWDuY0uLBwxPGZEeYyCgpV/MlzY+JbQwsoJ2M3aD02QRMDy1S
vbUtJswluBK62qHynAiLVtXKEsHOpM8pW26CjAJq6FPX50c9ke5R/ApPaR6HexNS
RHi70AeAXf7AdTyQx9FsYRKqlSDAZwsellip09IePwP8zQbMy55qd37hb0iTMy5/
cIfmwzccWlXWM23ooGJZuCsW4LZXwizsoC4qkXIAqqWz+KeKlZdp4+4mRYBLfNEt
RjYazvKms4ZjtlBdUmEofIJFTVSGyziCAuGwNPiOdy8eXusEpt0u6Bkms9ECptES
QujVFm3id4DdGoIC7+h3G22fDzVFiJ85vjkrJ+ZP1STKreCDDLI4tkKRkAO7tkmf
9drbZlLS3MVwqrgeLGLR9/gQPyFZCDPaQdTHki2r3lhNRMM9+Naz14k6YJyPN7Wb
AebtqfvCr21sDbUw0OdvCOmiN+yfR1IcLtJ7jgeD0lY+iTqbhQwvYEyo7hVoKFPd
b2kHVDyYrUb+cZ1zMbySDcwiqa8gaNJLjDOZoGR4Ho6dGHizvQrBk6PAzLt/5QyT
hLgoPFOkS0N4ICHccVvq68BFDWlroWhua/pjgVhRmoFq+UXSHwIEoG3JE1/ulNMV
rZZbqNPMdIO7JVkFvnWDK6H1qMBwmQaES5g9vUVve0PR4vr02xo0EBkIBKrIiE4V
8ioArOX4ZA3swf4QRw444PY+mzJzkH2maKUCHlCrJduane2TE0nY2cVLLmbg7wlD
9w8T2N3Wt0neWt5rwIbvTgx3v+Lol+aaEXGPzJQ83Nfk8DrPXGZd3hPQaSpvBG0y
dz+e8+F1Jx8Po9QlX8Mde+xmp9MBCTK2HYJ3bku8Zt3v241nm7YkhY3VeDS3qTBo
AunYxisyzgA8A9ihJ5nu1kvBC/Q4JeacsGzdnSdYzpeXqZwESCQLIwR7nSTRYbSy
9lF6SNkZcEg0LDhHwPZGdPXTyI1Q6k8I3r22Ur9/0BkWUOkS9ZkGv9QwBIgPT2cY
WMZW3bnNMbtyt/dKxcotGZUPnGJFuuxfe/7ziwp4y4JVlbUGTTIF8eBNI5MsUPEV
/EkdAWT475ynN6fXfgERbHEmpw4erg3l1uQNVUL1IZdzFK8WrjZa92+mLyQC3qCr
1Po6OxmtwOTgP4lCrYagwniUM9RCatVYPJiJW0XdLEiTVb1lEMKxPcjXWcaAmKVs
2XoEUiV0lonEFXVpRK3E4pGsE/0ZZPX+LRMEZ4gKm8Vg3Yi4VYXM3ttzXYsJ6Bvd
3uK4YwyrX4GGlIrYMe0l7rGyK2DTDEcKej8NLhBiI0bBiB2XL7jd2WUocd+rvoWj
/2kHxsDuI+167KOxK5o3LHKebH59zG+wPeaYTZGO1SHz/uesNo3qPr1VIdkvx8io
UUlQcXJIRW6Ydoz7ChNQ/yQMB2xJDhh2k6jiU97zjwUh4gYEpop0MI49rmOK1b6a
k4q6iiVrfpdjPC4q8BTzWEkx/dnSctvZzX19pIZE4rwwtzSrnqi8pHgRTw71hpwX
E7Puv9i/jAZWcWrpjwNJ7m1ZOqzwrYmKvDSw1xRC/1BfgW5IA2KSHSaFJnBkZJEV
pkqS+yTvWXsHyZIzSNNvq6zr232DemZ5CdvWX7lmkkxEyVmUo4jTtSYGufJ1Z4Nl
WFEHnxGQWRpqRazz2kyVDmhSbaJ6S7PKM8vFYOcT2bFz8T/dsqnQS5rSFmYx2bRz
TU38ERXcM0NClwWBejhedVGalb85hFgpSM+9gw1kqsLCVDRls8uwDjGtvO9enfaQ
q+2TdETG9rBbNwDuCkOmcM8C6YBJm3/BgF3kqbCvNzyWQ+Je/pWypBxzcWlY9xKg
soY7hxjklDA17loLKO/v8uqQLj5NjoEk2XqQFTBZxC5HDvD9RgLN+a6+41xhQFrm
uMOCfJtbeKZNW2FeqgYvyDXiPM04ECvFr4ubMlj10AXZykdJWZee2WpK4bLylrUt
95GIqzmMN0bgUeokb/vGXZTF8dhLbj8GhNphNE0KpXlTtY00vhCqL1HAC+QFrL/I
uqToRA0sI2E9XyIwH30VfsPdATrdWpt/XndxJidf9tTFt7dZcnZI4xRsVZigZVhj
r1hvclt8TV5LRNZ4Nq7QbwMn1qeKdVKSsnnlZkxbj+jfOn4dPFEnmJg7u6RFtD6E
jtUfTg4TamJmHC7vdyqA1DL0lE8MfgxlXV1aqrp9lTDmDzy8mKrWLkQMgstuEVCA
ZskQ1CTdyXv8AgXjxUwmpQtg6bMUWvJ8AIZQ7TG7qSG8xGxg4efs18hH0OPLOpwg
DRraA03sv61AeDvf3cKWvRP0Ba/0ecDjWpgJ1jRWmn9YJRSk6F0KKXwKuTMWdNHS
3Bmrg6rrzPvyGnUgrPxf4CescfxOV0sCvaz8ujaZNa1h9Me3k3z7pnO9ETe1gVgK
zZLZJoZlLtngj39PhQUsum/jUo5fLzNKfW2ewCIAOXGOxGxSv6ySyWgWWab3L6y5
Ki+1wW6Q7oori2sz3aJm1YHuQAJDRUVuYYSuUjlTEZzPXW/7dhVX8/DOGl48pK+f
H9uJDIWKAtvLl59IEZ8DNmH8Ph+g3LCSIUXjCMq2240Fd50Ura54TWZaRfE4RPrH
wQdegkxNmNaoyyH9ZHTLD1kX6wYH4nrkQQEHojPLv0u170yllNoClHyaGelxA18/
drvA/2rB04dh4dM4G0tb/0yO3yg6DZGiOAieCXMcIAIL1B16HaDp/kZ4O/X5h6TD
RjbuVe8w5VPgrUj3IslniQ5rjADLdREHvzwqdlWf2pc0aoy8sVeWQnkai6GXQZUd
tAD682Y7RrDPv+qW7yTtwKRojzcu4qW+an/QBXeqcBl5Kxkm+7tAZLQs1lreYl36
oMQbaN7Mqi1sr5VFhJotlyuSLfs1JD1M86wNHGL25phOi+Z3U0eQYhHcb7fYqnA1
omKCPJjlaYC4NH51XHJaJeQnVVbNM98gf5oa3VjhN+KEYNYNXM+EqSBjpFJsAfu7
cl739aBjdQqEMs9YIxk72mp/GHvO2qKOIVMK4OihiJeU6Jb6zltrKJ+sdkoxdfPO
uA3Sg/PXwO3CQlYgMwMWt8IWcOyGjhGVJhnvPn0wnGoWRKrAprLP2YlhIAQGI30i
Zshin0+K2kge5qSZYKUpELoTj8NpPbVGOmjJ6YUajkgSgZvDRCW61eJHcVbxda14
f0R91VLcVW/ArUUd+2109VwDvNkMaYSRQbSOcKAC5Y6aHBQAWsexPHVVk7Y0eeMj
0Z9BogXD3qAvHKoZ9nqizZdiiYvgGQczf78B2SsoOeQ36Py19TWDjQoJrKWxrj76
Yioz5NjpBDWB5S4fyik4FFtLZGrmXkL1oN41ffQwDnX8Wu/4PWq6DirMqkTtTlu/
7LiXNLd5sBb875bRPmh1p70Jcm4Z+ASwikmhIu+g0U6v2q1aCeEWGKsw+6+6UUCL
mZVP/3M49lggUQFlvD8+EfFTycm1swOjn8CslMsZWxWIeScT6esXHVTaIrDnYg2U
Xvh4UxXM98X48k3If7RkyY8W5bUruoht6R3QmOu2HECPluWpgS8zDXcVzTl9OGO/
GQgfFsZlieEiAFzExCqcYgJe+m7yWuBhTYgkKttaLBgDRlL5ClSB5GZN3zmdMCvn
JDFlmnaSPjwukc3K6/wLzpAcqRHPPV+qKOnkT56R3cLyjQPvNfX7x3dgZ3HhZbzH
cecBG2MnQu/UpdgDnqdcPIaBfSM2g2ZNcy75J26zveLoMeoIVNqmAZ/JMM1Xfo36
IkzuZSN0L3C8QDnlTdM8aHyqFjuYWw/lOqrSCOtE9AYLDjOvuSkBYzY9FPFfzcPz
asRIIfPtF1U07ccCpBw+tSXDHM4Bx6cFZcId8l+FXOHh2qF94FQuMPQTRaPiGi4m
kqialzzUCYNMGWGq0hkQRPgHihpJbToHv1KpUPdbGYk+dIFbk2Mk8ehwk4PbuXeR
yf+EpAekMJwyz/mB80k9lUk6Rv589F2rwo9x050tbxRY+cL3b1NbaLPiBE5QiUmt
Wa6C9sK/gWgx1IWkC6ZB+NWl3hRzQSOoEUrFe2gXZcTCf+JW28oXOMARN1Cle8Pe
hT+dNbpYwsEX0tn5axO4Iro9dc717oIim0IUxhCnTUkfkEHoiVcp1VZWtOmACK7k
Z0Rb3NBHHhxgAzIOdEbd3cmSU+1OjRL/OoNouL/omLp1pV5xBQHlOxaTvxXXD/8H
5BCMSp7XbrMDQkvW8rEMxIODYooCcfH5RJyX4m83sVx9XE4Nf0lig1QTq3okb08o
lFII/942lpEIbJhbmMQRRVFH7DojTfKltoe0wPmDJQGQm0C3V/L2YdOp3rZsk/2q
S+jvn5Xlh8dj6FBQ7CeGEB3acoq+fBQ2q66bINwRhw1zfyyRjXvoE1DNloxe7rLE
daKl22sKh3Kn+zM3dPsPPDGgF0dvqkKtd7BF36O18h/timGcR1WzHhGEKRlY48Fn
wxLduj3Qy2G5uvuNE6Yo8TFGeDyeywwCbRtIYpdkN/G8rdmgXSYbq+FDQfeDrdpl
5H4QHEpNINpmNm5hzdH+dgp/YrnYS4VENDN1VeCLtFiUfPVbI9oHWfkdg4iIlaoQ
A1m9wlnP5zUBPhjBQmJt16QKxpjxq54eqB/I6NT1Td+O22+iwwhCIkdZXnEs97fW
qOvVjBGr08Y2BbH/8UDiKsuwrTq2lYTufEnB5I/pnaVf9MFagNGMXj+sIZUcZUAA
7RTTlM+7U5KVCAEV4CY/4sIoxP4Neoqtetx+Thiv8tl5luupXh+1WGMuVxQ+HLq4
SHyfYFro0fTvKzhBakFtuLrR67xDYQQO1Dxkm+yBCO9rgWz7G51AsRcZ0g1RqMr5
T/TD+aNVo9YmSVvnDqpgcJM+BnvdRC3CCCVHwPcFBThDjmJlHHNUoMaj65NiiY6v
0cMx+4G1QlOxO+RAGbFpPXIzZQ21mrRv8+mGdRFGotl/R6Vx7rPE6fZy4fWyJ3A3
/tJBbN2HCPB7VmJMxg+FAmMbA57skFPOJXwI70c46j5TPNPUw8gvrPjnqragUqS3
1r/AkI19h/WuxPWHwq5P6ac78qgA3kd5QDL8ZV+qbUOwImKM9g/b6DJaKLq/y/uh
cwV05aQArDddCDI8glGouyUY0HxeJx8RsyIF/yjc6aizLE76LksOa05P5aIQ3ET/
g+lZsWQGRKnumQI/bUspVeVCb92bSSHCJIcpQcCZ1I8+HWeBuvsz4Wb4QjARdbI3
W9qqzBeDIIHzwGhCO9R55ho+7ZhwE7pOm3aMFFxvL/uFBnL7m6H7joFWXBTUzJ9R
LUQN7Q3MPYy0d1HhM3WE8a6AQBJBT1OsBXf88iS/Fh78RAGU4/smXE5zR1CYdRey
Yl9ylLeP2Vpp3dpr3IUxTEm5dc6MdWSDQsDlAmUwyWrecBoBXKME41QnOaSL23QI
uvc8hYjP6JKpC/qZP1HG+VkNZIdWhxvv9mrG6nqs+IWiE+vxl3RiqEdaxgyxuz8g
I7Ci1sQZNB678Afbj4IrgtuC47pub1OcUbKcm+KN9qXnHUrQ5sVyfXXuoCtpCJ7r
qN7CFfbfRI23OdpAvTjkui0o6MsH0fA+42q8RLDp703+367nWbxnm9VnERS8pYUd
CmNaqTeOQZUgKl3/PmG5FrcbQ49e1uut9Ra7P2FPNjhDq7wj7DuL6QDpKYeMt6MX
RnOcGtKcoYRi88Y3eSmhKacYj8INWa/PMmo+RtZ8dL4VDjGzeJzlrPnCXSzH9Fpx
c55+tcdC8ptYKVrQ/xJvHn/XdCsUwC7WzUHWxDWNicYvQR976kRLYTWeWOoxT4ZT
LohylUueKVuYG5lF2q8SLQiCl6VqS2D/NqkkGL5scyCF8MvRrfyAuD7qI9KltjrV
+rSyqI+eQWVMgtG6IlHSzBZyB7Wx+f8SvxJMLQ7SvtIKsiImYI1ZaTw0qViTav6N
EFxHVoEZ2wKYRXMDDOydSGaFap+FI2zHYg5x+1w1AhXN6D5d4sm+H6enK+VeshdE
d5XkYg6DOMDTMn1/Sq2qO+u2CnvCw57fdQo2a2TTWP49kLz+3u06+zfY0Wb4sXR0
HnbC5wIMjeCyiXyEWTCnldiSp/pftrr9xrWwIFFhOvgX5L2arThes38yIEQRzlfL
uI4ZyJ1DtIQWeLO0hltSUfJGMg648VHzdx/FcqVDVuNL9kmBfM4xJvmbQ+RP3QTO
M7+AZtXnt7UsWXFZtCKC5PxeGP8pJVXxZ/43Rs56b45MvUMN/mpGyRTW8He+mKA0
9/mh7K+XQmZTHJJgoWPPHRs3t5kIDUobt1BQC0MH/Ea2SOlMsVKrmmvf47MpVZgg
XZHKw8gK4g4cXqLz6VSvwQrZrobmf2EXZ3zUCNUZzJI08xj7Xf7to9q1SDw2hk06
mAnL9LxsN2vqBDaUinUptEzJ0uXV0U3KpbRXtiGde1VvI3pbuilYWHbG1DIzLoQl
X326QwNM7GLXB1vrhM6ubWKGOPPmdsHrzsys0fWKfeHclsC7qokXjZyFXlm8v47t
W5BVIk/FVjwk2x9KsSJanwf4+D05xuPZgsXheN3LKIOQAWLzUKo4iBeDG0T0JLn+
ZIE4RG2QvjMfcg992YrRvDJECXJLhO0It2aqlgmiGPWkjeaUa5HH9wND/eHvEZSh
9dY/GAI7hv6d7jSqmBkwaEShfodxd1J4Ds8oXtfoDYY0XdHColbKPEQaIrUOB0+W
JYoecN2iOxlif35HLi6pbTD7ptZXYA1ItxkjJ/UYa9qHQLGmoHooV8L1YVeO1qrB
RGI3Q+FmdwlZtYrglFT+lE/Ex6fHqVxJHJEBtVj67q86zEtSTD7FvOtMPT4LaCJs
zZd2uw4uk0xeowP283h+V0uqlWn2sGunfp7iVoeyQ+2hINHxJsDnhwp7Z8a8pYsM
cmBenQmAfQK53CBDZ8rtKhO7syu/jnTTA1FeuyIdQ5YRF04ZzPdrsD3p343CXucu
kGt34hRC3YLx85Dqs9vxAh8a07mQ2gJYyRZvLCH/6azrBHAr78SjhJ4Oz1p4ZLJW
yHzeU9nAZoMs49H1fNkRjy/Omxic+nawi+f2HcondoZXtu3DTt354doSfRCwtAlU
0uhrVsy2nO4FHHoVdQfrqMI7ES5ALA/LFHfU6R8f0nMuc9/zbcugXhm1lksTNxui
6U0Q1kG0HNtvPbEF6ZgxYG7kExrXZyiLaQrAEi5RX9J2L3QP57iOeDzDbdYSaW2z
4Rx1xpAgZ9jJxQ4nDDGq2qki6xkFAZnJxGclb7EOmyXOrt8ftXLwTj0Z5BRseDbc
YAVtF2AczXy2rJdsHrlwpySiXlGxeWO85hC93IzNwmE543arJ9furAcR/CSn0zH3
6ejg53bn+uDMJNxs39ADaagJo/H7KZCeTq1LUFt56dF9iGm4tBPYcFU6r5RKzVL4
Q73YhyQT7z1KoJdF+lW4+FWc4uHnD4CnpS1zIvmXWbV3co10vSZbKHJmO2CxFcP6
fwZQWEUjWrZifha8321tYUjfEKP9UUWMzOQ7ivz1kdmyUyqTZMre3k9glPVnSxuv
meIOzwobgslIMoJgMf9HLy8As9Tgq7LNibf//ozNdlfbllAjT97Gu/cENyBwqdKP
nAoCblBWQHYkgJbCrlHDqP2r5/oeGp9vb7T3EyhNawIFF0RakGSDGWq2d8UxLEGu
PV1smhch4V2tTzPccg+4ZIFgRo9VnpzOKRmYRLsllQhh7BO7NsErB2AOrUlq2zbt
w8bR3I0QFFS+/F87/xQuyDTxOCJOwsv+cSb33k4i3bp4C2jSZ27mpb5Vh9fJl6f3
hIvZwujBak+fSduCE1EASN5Fw/KiSwYWGWyoL8r7ItYJftp1s+DIA7bbw1DV/zn3
/TKiu9AmCch6xK7vuk3RVVsAPk6cAD2tkz3lhBwpyayotDGiGDo79hi9YWTbSMEQ
w0/e8/Fk8iDrxKXwjjAtv3k0vK533rlJ0d+edz7S3W3HATYR/xAVidGNfw/m9v9S
jpD6VSCeCZsngbRbeZ8I4M5+3egNcoFcStpDI52P1jcRs2gE4za3PtRmVmCQwYG4
kQ1IWMupwYVj60Uo9nxj5jgvLrGG8o+MlJ1Dnm7cBEYOwY7VcGclZy9uF37SR8fJ
weZeh4zYl8IbSHIpWSpIGR1R5ucGcGyUnz5GmDPSJAp1Gml08lesqOFFDbxmmnyM
aJ4xkfIfP3ALbUkUDmPT4FHZqiA/ZqISaoL0xy00G1UnIu/x361NaurjejB8QXTy
vTVC088aiswMEzcl2nKvLenXUNcg86JLNFNq/9q0vnuVuj4CL0WO5qPYJxVl1uzz
z1JPw8GiNxuFmEWnG1MF7Cc8BXO/B7PlM6drUM4MX6Ix+OT6E6xO4OH5BFxM8zVE
p+qFVsYv4h+Yyc9mhNRorKwYIacqChT8YvGZmp2WZSNAqOU7IDbS17A1PZpiQSOB
ycIlhVqtWfnH9KGDZ0T0q5RTA6oUCIWZjJ8GiIA4Az1RRcoqH2tIDwSm/OtzqJTR
Wda1LS7CzYDHTh5kT4SkPPzcou6rVN/4Ll1vXjJZSc2gKeuDbHKImsYkK3u9h18c
l5My3WjCwTEv2UsIlix8btYdffHpWBdGU3osVfnAh1emOOcSO6olbjphf+j6EZS8
F0lXqJcPWBg3LVFl67CSSbrd4xaQeBdS1zzAae//RYRMMUM7G2YpRm7FQLNdK/Xv
EDTgYjGpSmpCD+7fZNBhZ99KZlznfgeJKUSMyBLP3wHiYbXkVxPe6sBQdCkNLYaK
cZXM4Enzy8WY5rtkesbWMxXdGhz4N+yV/rYbUJVEAQbSQrTk10oTebjcupZS7Puc
HzXTc429t67WCV7/aIA2GQu4Hz4tGRtcgPKwuIhhMYtPV908jWgsGZ+1tsvU8+KI
9+z3wnKphUMyH2iB3E3osQTTGDaCQwEXLtMouI69fILMpqpADZkE80zMxNP6blqo
I36Sg9/JgVSYdmXgpCDwK5Vlzou88/E5oRO2JSOGmRwqnYfTELOvFEiGlXyYSxV3
W1YuDD0mbpp9MqdkGeox3epY5pei8NXw/zDzOrF8S88b8xN/XdY8BuM/6ngpM8FZ
SNyb6cLQWNPtRryTNaOlsWwdV3QUymlQQ0Ba6kIY+XzxMLaRx/WFyEXJ1K4jSq9S
55y+qFv6QJcDz6USh5kahKdcYaDFUHWNk2dulRnhAZ/9fLfSBRGyTSR9FrGqKilw
hWiv8hT1C3xiWBXzODo7QlkahODUUOFo5eAiMshEtIkc9ZucuywAFKR1FaZVTEZp
BSGXFL8Jpnd7m5G5mi1xmB50GX9rUSmcZYHGn61De/wF+wLsoQaQytQ5DzcW9oFq
JeVnI8JW97wAKCbIlGIUmWWlctqjmHr7Phlq8mx3jWqKgoYQXYkSuDHyfDlWW/pT
pNzOCRpR4rvUZEa2JxSMTAI0pyN2ee7IbPs9sopCMwnF1JXm+9roKnVgaGrky5pz
CvKsqFKYox+pUxpBxFz8W3GrdGzu42maI44hddezymXW5pWhKD+4UreYWUK4C82C
LrX9KhpP1pHAMuKE0h8R//P1D7LAhYXNLXJn1oYE8bLHTibDaKOF6CS3wLyYFS1c
Qq7eQDMZp8V/Ag7sMLwMbKE4CeB77ccIqvw2nTYUM0n054egGf6iJQkix/ehQ69T
GcVvMu6rxTDHfxWHYFoy8+DFsPv47b0qU1cFp6GJ0v+z7oFxDkFTNVO9xuSwrjUq
TN+JsusS4gGQehZ8MQeWd/WwDgdHFudnlhVmbDjZ7GAu89twhDnEkKYy+yHrRVp7
rnvQGQaSiyWGNwv+bAQjCOZX6cUKpYVrtIAeCvTAWPYTwRnu6AdipH7t5718lLIW
1i2a8mXUITE9/ehTM0mwbQ2qcx9AxSLOFEmYmn83GK/yGBuwuP2IyqNsHsTWzYCK
bwPUS3Z0MxLkYcHEAds5F1VNiQAibahjThBA3AEvMjeaw9uIgVYcd8lJ17sEiZf/
dOBOnoaFhK+UybOH4+zG9MWL/nCi212sRbF2gl0wYBdXyrIYp9WL2XdWcBxGAUYQ
JmnrRYFtWRWL/8L/CfOaiNWI+9UwWogF3e/7GLAJAFa1ItumQzX8sN2/m5+JkJkz
MIarfvMTl+1HVxKfwrbXQFVt48ZK7SwGAb+X+3VSAkcDKH1kqSqXyPB7A7a1Ya64
/GYJOdt7/h94qfbTj5TGWtGdoTIUk5eG1NF8ZcsJbNyk2C53YrMhPK0Knm+b+1RQ
GWWILLUA2N7qPdvF6tJX3o33PdApM8aUD2u7OQviQ4vW5L2vikpT5j9umdYlEUnp
rMJWIHjT4/qyhW08x0u20EUPfUH934nzriQ/YgM9z0j8KGFWAmLwOeaRnkJXA+f/
etXLuxZWU02lF4FFTDPSBcfdLfj536qFYBO2OVpZQy2Dl+fI5ULShIMsvNz7iekz
czRIG9GTykBBskfmCZKoDwuW/qgYCslKsdHGHTKMXt+jm6uYqejUUnvJf1GYGaMT
jzTWRGR7X9EKYkRwabMQieWEOAXICNG9oHbDJg+9reLDT7gDCRX0dTz/+oK2KIQX
N/qaw8JfQoimeNZOM+hMhJR/DY4XR8fDc4Ya6S/E/mMjGntuqMCd66ie9s72e+Z6
GOdNvFajqZb4R912e7w9lmt0UOeIlCv9pVzsnwdd43iXTGewNY0zAvV02mKV3OLI
cs36Ts+WFP+9JrUDtiUT13uwtPtoBMal4YniQyOGR+kQO3X4ex5sh5s9yh75BotH
Cy68WhkxKs1YErhOzOepgNZV+SkML5ieG2RyLuLBtNb4xiE5wqgUgdXLyaX6gEQh
GH5tEaXaDzZlJ5eFL7G/1fpcNOlJpS42NQH5YS675rSP64DM0lg+ALvHM4xk/oAJ
K6qMI1toG0IFKvsKrvCR7+fBXZ3k7/jj/O+fWyKqnM3WxTiPDBcPZLAxg1+pcB7Q
Bliq8iAIAIL7cL+tYxSSkNE/TBuV4EMwxceE5RB1gZS7baALvvHAVFfhZkQawI4r
M+davr9N5kafoawn//T9rqjsi77nzQ1CeXRhJ5uBm7kLd6AcRkpDz9ExV6EyMJFB
YZUe54VNcM9zCAfzCqJ6abdHPGTuNA9MqMwEZUhHAMDEvZpHGKQTfzbIc5ncqFax
i2q12HwTFKahRKRHymJQIUES0ksGP+0dPQYIqxTdmnDisK1LfqFA7dzZUgm2YTkb
TMcPst04F8bCJycmE1AKmPLX9AYiZSnatu0FPVuGzsdeYEpPQYkyNtk12wN2DYY4
EPvGQqfqQdOWcmYWCEDV7XV/oQTHhSGdoWejBZgaPDzcND8BiOOrlX4ltnIcHm5l
W9muD7Ta/VVzwvYxdOcjeKRY4FgptG2SW4A5CE2F9Pgxw7NYsYBPKgIm2riSTHLr
kUDAkYIk6ETbCjaHzvzSZktxk3qUcOGuHlydOxuiqIfsgDcS4OA/tStYuygbIQr0
JMkw37P3U5vUNFeyIKs/E66ljjjeL+HoGcje2stgpbPtMxHL8061BnXwqmKyx2qv
rubZW3NWik6jQGLfKdKwSbvMQV2T8XuJ/Bc+MIcVambY+7BqxX6EKRzY0esvVatq
NoaHJJWfslhDFzNy0hUGWJpYAI3yVi25PEVWaWeU8nXfY4pt+ff5upSvsMDa620k
sXuV7ZzjnSGyoQeIs00+wXhubzQMehWD+8cRmjIwO1Nn5QlAeC1jO0s9Rk3lGRxf
/PqldlWMNsUOoWPQsDRaJC/DW5G+0jiNgpJtyWey+tYTB6H3ly/GD6PZt2mol1uB
+so3Fi6G3tMUuHIIirvfyC9BS10Mi87d//0JTbXv41GytdTTYOPkRep619IwlvNY
Q3M1M9nby0amO9Q9hAAFEfCyZ7suiWaz3lfGnc+hPDbr8jfLGkr+RxoFsG3G7H+D
YKobxUiiFcjOYUAKRj6OJNaBmihcoThpEQEeTTYPy5h/O6uMJiSqGbH3t0SqA/Ft
fm0F2al/iM3hPguVSoue3o4TX9Q8EYeslktJFhVHAcRp5BmzKBgPW+dPKh9otIHB
LvT5EuB+/0Knx4ovEsHgH3DZ5sdbcgiFLStuG0ZZIQ3lAioRoQCxR+8NelWSS4fI
MZs3RHgFNAZsM7Y+YYueX5t6OAhW0pNChrL2bmA95hLn7PxjRYTOlDCD+2weKTH1
qUJ4Ih/zoQenX3rebd+PKBzz7LXxtMWsy6S8y06L7PKUfMdtivPDPhuqFDcyGdFq
4XOyRR+5rZ+vxegL9IlnxJJAzu81G9W/YiBUGTYrKDZ/+G642OIXa91TGJRX/jib
kdMZJVyNTO1x603rlloQOQzhu+mcifWT2fBmqxfVZ9MpXIUe4MQzMt36me/fGnQv
g3T7etcGjmG/Cy6dflRWBmfF+NoTlAk7+LwsQfgaeOJOz7fnaywLo/mDu5nY7/0u
fx2nHHGJpna74H+E3KuHNQy2wmqL9plll0Cmolg33Jgrrmqy9i+s4XRR6s7xkmoG
wuwVyKCVH0JoshBbueT1GfHyezVw/Xvw08BOZA6EV/jsDV26bsmSPmHVh/ca+GCG
DJmuwdOzl1Rbm183nYrs+WZkJweYVDFtXj20Sx7sAwcYWmCRk4hBfsKkmOm4jq3R
UxbAb8CEzrwiz/Bth+16K2HrwxE8LHKrHwtC9PkTGoGyYa3g0O/nI4+0uwLHfzCp
ODWe8AA7WHGU+6QuT/NRMPAPoFDGIdD+iCmnon5q/qAe2hl166Iv8U9Zl/O+7HEl
9NDRWmCvN+2uug+NhjLdqwDbXLAezXLjXj1OFM7RzsvnA0v1+xjtFES+1XsKTdsa
i8TCEtUWj3fB69phoSdnFys7tOZjAHqG6DRqUW/XtzREYHfNj3WZBWIjWLhq9t5N
stSCGNq8UT3f+FA+4M09KPTwRRqat3rmbUfODtpX/mZWPP20AcPpa2ADvFUXq+da
+NDmc2ERcKzCnzlhHdh28qjPeEWvpHSFhU8PBjfKhVMx5iFffCbZ0toUZZZ6LLzD
4HwnD6mBsrV9uhDX/cFzXJTFFcDJvrW/JIoLtoyJex9OeKUMHiSvoYwCFGD0Egqm
spdmy3xNUCt3qwDWI0BJa/5AV7MRh8+FLoHPlOTnsBwz2S5i23ankHEQAHwjcP2E
U51A3lh4e0+ZML8tUBPnjo96Wy2lYYduPNH3Z1sJzOrCidUCC/ZoJXev9cC4cVK/
zwpdhjHmN8qogXW5R8fN0h1wVOw4BjtetjyBVbIhgeGFinmtCnNoSYxmmAwZiNrV
bpAYJh4zjkVTwS9OhAhtn4iblQNkMT/nMu1Rx7uJoQIuQtIukyuSrBy+RZorNEYx
NpLWsxCoiZN4QSnJ6HKn4/hmVVS8Lxmvy+nNsOqDN63mT/x8hQyky7ZdDuddiAta
rV05eNBWWBxXTmb9XHFqkEgT30NwNd3vVLpSYr39Z9zPJrSKn3tkPRuSSZI6ExEz
QiTqBORuUFRkmQO/VMUbZorQ+LsamaaYwfn60hRAKcytqLZzAJdzXWF8Iv5lAMnO
0dZrLQCpwd9K8BBpCFLY+7z6CzhcJ7ZYyLxZYawhTVzRiSd3/48UOTRS0eZQmcfv
eZTU3Wn3cX0fHnw4331BZ3qigx8EM9KYtg42OH3EGHJA/ZbDD9t01ssMZ9ASU6Rq
4A1Pq7kIgTh0T4ZPw7+eF5wlH/DTdqZ7NWGXAF54LR8vSZ0JAvsz68fOaC1WLaVl
dhAe0Xirxa2wvaD1nAS5Ou/zl96YJI7pkMrexDQhFTxSjdAgIOVk97I+q++xB0Vc
aZLK5SE5wGIOdrloc0MHZGHZmMeC2UdFHOwGWSNCvoclRe3BOpztNMVNXSJWfzHi
PBIAmMQtUXgn3hRf9JEiw+Rxb0N0dOp7OgUP2N1qpFa0P+z9vnvYSidGCjfgiozr
+OgVN6KY1n8m/l0ycZ/+tIGdVgv0fplUBpttVm5Jt7rbpKnx6uaxJ6c2tjsyv0Aq
VIQsqE2SEgFi8yRsesA4NR0FmjrVABqR9/XLX9LBTEmKBemL4rTkHv2z3HQnvDIR
+InuoLiRODao2dpLshF3myv3aDyKeo9Y2jB9lZdYXIweWvuPZTvcwyldzjeKxhmN
KPXZ0fBuLYHA5Tti/h0f35IVl8qMaURFZsJZlmrZlkSOKuVKTUZ6Sm4MAm5vyPar
oyp8zCegNeUodLIcxYPF57XCnmVflr6OuCQF4UlVVdTxMFGjQA2TT8gwL+M2aUgu
PhW0rL7VU6eCzG9/yZTbE//UfmAAc+J4sKZjhQuefl5RF/Sx8wSzM2K7ngF78MEx
MjCige+zlBqfwYluPSpVhArig/qiVdCcxs0mDlM7f3vT4nxS0sO5BCWoDmHAVs3t
Hs2+SweNZC9AT/zm+InL9Nu2ji2rZMiF9RQyIN18iLOfOS52zy+df5c1JaNJOPdF
b40oAzh+d6yQrZAP2y6seUwfHQ2IIo8qIO31UALjrsc+Cst/NqMIp47Rf1pqjiKK
jG+/Ap6vF7SFlOJ/hSmWtZVNGi8GWrUmkDT7oqbDHkebxqCZ5ExuFz4Zi44sk32b
UBrVTL0biY5L1SxjSwCPclcQzu/QEtE3GhthN9OdCtDPhnLrEenmyy2G/+LzH8zB
8O/UgYACNIFVQ9BRcWAwNxmp2fu1erXhCwDidLAJAf83ZMltKAS4qOFcCWsqkMmQ
ZEX9UI8ZiWpXz4anTanIje2ZOy74BXTgvaMXnQwlAyqdU08YUk028D+s5YxUFRaH
CvByrR5EuBOAWHiujSKtNx4ZKezKrznhZf4lC/e0UyJvPYkOAI/5Txp0I35Q5zT6
Ii7weYGh8WV7bi7vgToOvXfYqeKhtDJ6dcuaGLj+wZJ2ZzDAaeogWMKRcDur+1Kk
FudP7m1bRFdUJrF3ISBpKte5UGLUvPVIWJaMJp30QgBrV9jW4+C1PcmunG4pvbxb
QQBXOVpJW+xNguvlALUfCgjcmH3KzbclVjJDWqO52IkP5ehlRbEiRvqlmxfqM7ki
m2mWEAx5yM8RzcgCO9K9zPixZl3g57OfxIVctRS0GzL7XzXbKd9Jo5J+EdGlbgQy
TISRdQyKxxM2gklo+7eefVx0lJEvu6ILw5yfSv7WRYotbO+A0dMA7+if9JxFWXIH
GWyywcTjl6cGC3+DLqcQRQwJ+2I7/Clm8pSGxRh6kJTlHzJxrGVgbsSXq3afuW3D
ISF56p7cw32gBAb7YqXzNiakq1bSxsQyu3UEqNBvuIMOt7NzHFrzPLk55zZwm9sy
960jKbBHCN3Rr71DJ557F0vrrES0ctkSws8V/gf5rJdIkNLytFytFoxqYjXtOl6v
HMAD7dTI77yn2BvffopGDyjHliX0X7sp0bkw0habbdllmS5EBAI9zkQbFB007XsQ
0Z1keTBONiKtvmsKlgZOr/348TpoH6moz1dfCXopOJDRfFu8DM4sbiNWKUdeHhzK
UxSHu57SoqGaCOG1bZXK5An4gBZEYSU4j02bD5naj9VU+vBp4p133URhyrWnK/ea
WHfe11yttOLLZgndj+pDzHArftc1VD343M8FU5gHpv8V6NN18lgzd55V6XOFYP05
NV3XtsEUdVjOtOxLcM1nja2cczLSco6qT6ziFcUS2sy/pgFpcJAL/9iRR/mMl+vi
CrPAgYaZ6zwYkSibtyKW7RWcIYtg/s33+l5Iu283LjFKAM1iMjKvYykFQmMf7rfW
t9dgfAEMPED97zsa9P3X9HVqZ3rIl7GvD4bYDaUz735kxnfgdlhczV5/oHFTB7bQ
5ksGAy1BBjfHXXpOagkuBQ3bXo+43Q60kzaOQfabvMGpSfmyHcXqd61+QWyV5ybY
NjUjP44bQFS5skKbKshAyqxcVapToGXQ89igLKbKNzaUqcMltVnMrE5wAiJ3KGpC
NHfAcvQ+C2cUlF4dBx7jJ3GRL3zENitCCngpgBLqPOI7U8rKvUcFd0+izMpilFFp
D17drht5AbKcQrUJ7wBi7ncl/StfYx/8JhrO/my+bFdlfiPY6bImPj/LUvBDMYm/
baUZdHmeM3eCgIevI5VLOyN171xkWCTqIlIO0haVm/ieo9hVK0fHIxxd2BPi2rjc
z2NmENDX2cvvl6B9RblgVM2ebG5Q6wuXKvFPy/iTlILudt0BtqeN7hmluSxl1hP6
N9qQoCrKxMdPzljzB+5+DaYbRqvlL2R5Xro7e9+a0jul/hZT/fzxyqf6PxKO2zj4
uAaHrRqq5xl/j9Bm38wJFMfdxJz1E9ni2O9ME51pdDKCLavaZagSHc7d1s14AZQP
izYHfmC29UMBiQraTKvRfnw4hoxwGceTBwbtin37SAuuzwxd3EIJYYOJK5R6A24S
PRW9R2F8ZtdY2rFliDWspFczH9S4+MN3hGTGuqcZ7/JSpQaEPCXfeWEKRgOHjiPv
/qsNyziS5+3S4Q4fwXnar2hq6dDYrgklP64c8TSNQeWENtMw4Kpt4qn9DBr67dCv
KqxttL/L1TH0ZWeKlqOxmfTbHeMCNX6W3iMGJtSG5bgkD7Ga3O757mGbq3jfPBSM
7d55/IpH8lku4pqjxU7HERX6KfE8JvGCRnjroX7cb+dhj/UhQppbw9IKkAsrF+fh
HsY7ZvJVH2VHCXzML39E1vr9QPocD8kaay7M6cAFqE7dG8m62p8xD5GDMRgGo10Y
AjZ4JJfeK2bGXTGnPPgTX1Ysi2D2qw3DLwXOxZrercJZh16uRvmp48tUETCR+g/Y
5pHY0RD+uOefuIcbpgvrK8f4l/o6yt4HLiBszE1uhQFSW9zFPCWp8yt8VmoKCYne
NyiIrGhr7UZDnP4CK1IoyozOxvyr8fzSlWSb219TzVbD9SkXBRLh+OYWn0zD8uh1
8oop7O92xvxVgZQ8u+YDRFyfnYahzVnONEHZtb01o2B0TVhDyU+kMKPx+lsiS+AI
5Fp02LFMQhSEck2T81LKyzxQfNwOJmHrkK3pHvx7MEaTYxoQnVMz2c8zKk3OHi42
fN6fbrucJhCPek1HUksZCHRzxnlIE53VlAd1IPTgfpjX2nfQmPBU+ojSPqBxONso
lga17h7zT54XKKFBT3CiITMZr1T5NP/Mex0/m0jp8HYtalkYIQiJNvCbOPErRDqd
hkQ2DxzihW3r8tkliTyAuXfoX/oUjoeE2ASmM+hKN9GBIWq1r4njx2TTyW8We91g
9ZTEpME4JcNlImXUoqyN2c+x41GsbJPlgczR/d/C58xJwxGhEYK+CtJ4DC3F3Me+
wxIawE/IbS3FA69VJuQ0I51rCPsYVEOUmojKpi0atlJ0RgFRwQJ41LTV2CSCmWDD
ptpSBBzs66liDQIe07HZP3vApb6BIXWarUMUmyEnxT3a0ovPhdwXOv8Qow4NV9Xw
p3JpPQXibT9IbYm06FBh8VQFYjfdBeBeuesXj5vBB/trnI1TLtmroFkpqPMasPrB
+ufkHcVmFCSqniyyvF7cSYkyVmleuVX55SVy5cWd2CX3l5wbin4/jK2ujxiSiXvT
WBDU8oAkd7Wtpms3K1tKzJWjvF9Z/ZaxnuPAI2A/XG6eNMZqQ1rwOF6CpT5zPtwM
UwD8fCmvsMtP6W/JgQ/gRZJjBt9rJl1z1cB+ksasV4rcqnob/FLZsEqp9e2MFWw1
cqzOBqJRyez7YlHUH1xkl38RkoNI6rrdMmgPR+Zin2o2IB97sOLFN4Zew7s7gnt0
uvKvbuGkWgBW/+9HTVEHXgslbWYv8O4RCoPfq8qUeTOGCrNQSgrWISKeYOl4Xne0
6rYpfAkUlg3JKAcH382G1sx7Q2ilF4vWz0oz3dR5XWrlM8EaVz3s6B3IaK2qOOhW
f70DbzZ2A40kbzJQ1lFjlNaWCkySBt/YYkL6jmPibBagQ7OCHDCwX8+q2aoyVila
6J1Za93SwUoBnHO8dOk6w2+ElZKD+0zqB1ZXYHjeQkbjVqrW4lV8pnFbr3ov0vFg
FYx47+GQ9gj1EqAzMIkRjaY3CjzEw0iR8CmHstLEcK30WwMjDdKoEelCy94+hKrZ
hBOrXCl9K1sjLNegJ1SrB9gPju8S+/b29PS6XuZsWAWXJ6oAInvAuvstD+mrYYaJ
m95JtbpcL3PkB7yHFqnrXzrLqUZlu+6FFRaxucK8Ifpbmo5rb18PHjLLrdLLIAu9
Gc4yDgfm6nit52ye97kPjPKi+MNzHhisZ6Hsp1bNOf3+u3rYgXdzJSD8a0sbjc3C
hD7OiAzGqLhJDggyPoNJRhw6ft8GFd66YkOaAnTUd8elQY7ny7jiczYP/7YhIN7B
pWIHc3RLFbxum4uKw27Tuiyi7XrfohY01SQVQkYlN4pj78j6FfDBVVnZr4jd3nlQ
/0uOjnJZXnVuCa61Eeo9rTYLZ6lbdhpVvGamFNskkfuKHaiNox95GxO773svrmvV
+eOEbaJYAbHTf17cYsDyTAgTA8PUcf/ug531lQ1Yo5n+JV486lUXnqXnIxS3kF0X
/0IpYTYMiVMvmxkmujDO3HuOeBew5ZYEBd1AS95/uDdJY/Rl5STc5nCWsYVHM3PC
TtfGbRM3CS+cCW9IatukzUCwdPceD/RST67TTpUaLuvKfPJEkAbGGQyfEvecVZyl
/2X0eKzf9+RbrMX6eWO0nJILVNZtAtTMs7o1uaM6XMaWKUWT1fF5oq2jlMpqQCLU
Zr8R6ePWa/c0UtEAq+UUpM/G1wp3n4daIlVyCPsafDMg7I7QO6nqxmc9B2f8uztA
1+V13p8ulDC5ZRzY8VvVxGVjOIcgKxbzMpu3LrfztO/NUbczWmLzw/yWgKvAYzDc
iaHPPE/RE8S8MTDRgsDxo6T4MCFhZ56EdhtkVczCk7wwvgxDtrxc02ttdS7f11P9
M/AJ2nMPSCguEypAuwwZwwDhUH2uq7Dl117plpmPdkSJabSXuhCYncgPCAj0D5KT
MRyBxS3PBLd1sQzEjXjEQ81YQqc8emsk478zojhrrwPyc/aqV8jdhWD+MM1peBSE
t2f4Xs5ZOHKscfHWrYXOVZDErW8BFgJ7qUQ5JmdLNYrYMRCST6CLKEjMiTMyLOj3
y2T45iYAO3MJfHvNjNrQDKb37OZAXig+LUUb6Kqi0iGNlDdYMcXRhHiZo0HI/R4h
hcrh4lLAd/GdIxRVdGec3Hh9X6NQN/txsEgxvNmDVjJyetipgHsPisvspJakmLMI
bxwponwgzZs3dtAf6fbpI2wKv3yPc0pgsj/sBFs5pzVoSFHBsf2+17gB3gGKH8nq
CEtf1idRyIqfC47cjAcdTlGnM62sNLMe4RTGONHfPj7Aa+aLWrbitibSCNSv8m5i
Icl3m+3/En0NFUEcYh9/D3z8gEU1Ljqt2C9lMRdDpJvrQ4gUF3MCxZSDk0rvqk3H
NgAbpev3rrv35bzyJhoDgYWvX3YCNrAOnxZneWkN8EHqZAaL1FAyH/khSC3E6Xoi
iojG5itiSs8r1483SCP6fqAuqbe8DWARr1oAwxD7AxCpUbBVM+zh85SHv8lDVqC0
MF8vDvMtEvbrWAoLGHTt9BV+gO09D3fvW0X6AvSXZKbYulOhZBcukWNcGm3Yt4Vq
FKqACK9tOl5vkoLdkqbyi1zdcwupxM/QK2rBI140gf9E1IjOFgbAtJNnn1ZjKhhl
w7VFlc7ALj26H6fbKVLi/aoQ6MwYArMNb0zqOJyX/Q/UZYsoEcQaZLkKQmZ/vjTj
DJX0qYukNS0zvfss0fU1D96hR8h+KZNgAjhF5qL324srQibQJ903AKAWGlX4mtbR
bkG1ZbVyMOfCLhoIOq3oIZGyJfFc400Ym33oX31RxXHMpBOin+Fot2CsUK6c1P+r
y9ZIUONzuEf1VicoFeTyr1u+0m5UW/ZxhM1+zLT4ZLxcBrDYS7Vq1tgKuciI0y/h
zXbUq8qdFz1FFlPbAHMvErmPGvcVJcPVjLbEtCsl2cwAZe7z26A6/32/HcpLYqHt
hSqIbuMtOZ6fyTwiGoeZsTo+m0HjE9gfkSUyfHdsAh1D0Cj9RlgEVjTcWcyLRMff
tkkh/Yzxu4iYMOu2r7laD981dv3loWBCFA9knsBILo16wMXQudlXlSK7vEZbxW4X
l2c6Wfp4tSmUpYDotQyw3j1WUSwLP/JEc8Hi/r34zj8hvrYnVqFhqegRDAL2jXjS
sMk3JlPyNiYvto2npKTvND6OohfnHgipdxAn9Y7WoGiP3aeRy8ntPaSn4ADlT/z8
r7/yfpf1wO0I85i8fCAz1FCuVkVwRGg0UMw3goLoQq6tkx/X1kl7A9ya0njaeHPC
0eJZkgpL5avavnazzmMk6dvauOTSxlke28nTqPGgTt+h8RypXaIN3FuBeOOPJIHy
6dxfRsoKcx0TTXlDQ3Bzux4ZzE5/QYUDAOcqtJEgaatI4nQgMh7/7ZNODhe9izP3
Lh3WdH1OaSBtc2/RiZBGNdhTF/guCy4t8X3BaHZLNtHWznMN2wuWh3XQZ40Kpi5P
rzxLGUahv1HiE2TlKQZU7VP0G0INXh99nS0cVwB/Iba4COHmJtLFFkOBNuJ9k+TY
ENVpfDI8s1vGCVFMIFT0jX2MBMLzUYWI2maOupwg4KZEdTwhnKpGSe2BAa3/qZX3
+veaOTRlNKLvsS0sFr2iNgon64/NiTA3T/SWcJN/Jd+Kzd5EwAMSrt9dF0XmlLAA
29M0S2nzjThgl8/qXfr43TAWfHlcDSa/4W2DtPK85bxEvntAWJX0CcqzcOxxSrpH
V1c5+9Rd5ujoA3P4Cbw8WvH/F+2udiLLUMXWbnw2rRQR2Y//zEXahkLsYNQmKMzG
7UL2IF4gRfSIHoPpFpDwcJbvKiUv53b+H9GBNngZltk0ENUse2GVAO+6BuTou4Ro
NrcA/21MOcvBJyAdQ07b6bq87CL5rZAKq1ir9KAqR5QPevk7/BODm8PHQ1esk1w/
1YUf6cAg9qSIGzjwjMc9JnTZx21nPl/uiv4Xvpi4GOI0QmOh0Y/ZjAh6OQNUlcBo
D9O3il1osCrnT+4I7a1AiLZAGloXEWYxNXXYUtzpBmBeLRa3bR10v0ADnm1XGhE9
cRc8EkuxWJKZVqrkObFH2W3zIYKuKNpp8AcEFR4A7X77+qiKPTKX/JFFvFJ3xXLv
O/z7vwh7FpGk1u7bNJnaDgxVbWnysykZcRk11OCuFeL6tuWkma1M4AKD90rFHMSD
7IFt5qycRi/xBg+b9KIX4HETcG8sy6m/Sg/HoRPiafteVWC8OgMcsCyT9l22SsUJ
RmjxRQQLoCuNLnvOw6VfXfRka3cwqSthrYbOuP6NTKYLnDGNHSyf+ZJYLqkVURf9
BEWd3wLnYF/61yVMbRcgpjXeiw+smn/ItAYbAOHh83T0CJyYLGLHHCavZlOdSVIp
ZNfWx1MAwDp9X6JLozbAJwPcZ2FU+RqzM8otstUHb5SN0qIIgn22ggbCT7hPPGN0
oSSHDbTM201O7xoLLaIma5Vsk0I69IEF1ZelBtxfPKBSFt6GFkTjfC6zJcNcxmEg
WEgbWDChIDWvIoOLoBa6BPkDks3k1nggJJ8gmKAuzdCqO6vW7QUQAtxmjE6YPoo6
0zHhHv20vr4l/iz96iy/vQcnsGC3f2WXZVNciHxQ5sZt+0WrjrWY0tFczcxEYnQH
2cB5htsjzpAqg4q+ju2teRC55nOO8svH+gHZrrtLBmxsyRWBNJqiQLVIBSDuBIwu
pjzQoOJlyJsJ/PoDrzLhniTxZgo+eXKLIjTRBKd4sMrUhS2NmK80S8nFrVhNaM7H
RoWKuT0Ru6Pw7BpmiuMG2ENuuJTcPt57XYEMDgwcnvERl9XGnIYYPUgNLm6KE79T
mwlCmDxw2tJVUiKwpgLDsFeJO5wAMcvAjMSHPUkwa9epD2/TskR6xaSAk8PAr7F0
W0fnPn46M92qkVFulVi3M4UhbWcO5JDUIRwIjE/S7ztsssiJmuTx8BPY7/Rrshg8
Q1lGQI56BKnTnzZppyXx1NaQNblOdVnyQG5I5ga9Uh1Gn9mOZcATuE5pkOGVyezH
+ZFc4nZL0/n25KKowA2Y7nphWrobAWM4ldKHudI5531oI9+5G9HegZ4fgDORnVKX
SXfiu9TLwJggHVyJ/VdUfYqP3FATjJ09En8nrQkq/K22IXj0aHeOE1omMvdNKYzj
7WFfyxVTr66+Zn8+2rGm06+ht0NTDLPARY6ExEuUvbbHMn6I+wU/rBOpH4LQK07H
KPR5upTtSaj0xotSdz5hflvTtK64FsKtpftw7zVZN+6CsB/w1u/fmGcbS8IzsjVk
HEvW5mfVEkWE5ti3/T8nBwVsARK+cOV4b7S6zI6SXky5cTGYzw5KSYBs4MvXI9K0
S6QYLK+TG2n3iUfs19YEAMadN6Jct7GqOm1kdWeVyvFJWRlPOyN7FNHSIB6a0Bqc
/QczdWgKIlSzckos3ZpdRUx7ZCxVLoewQreJ12QDL5/nJH1tXvRn+V6elcvrF5PA
J0oZdkpNGoJNPQnj7vAoFmGj5t9FmeyWxCfn4rvfljINjw9VutVZvD1xLDeJo3LU
4QjZcql7IP38HOT0uIQ6uHp7Ejdilg+d0yn9/Msc6FZ9QGn2iyms9cxoFEobsk60
+R4fGPA3vs1YpMXKVuJkx32NGk/2R0LAfHXyfu037nUjRDZh105uQeCvh7dSQUWp
+zSliYB8cub/eM0FgqA6Q130AdEp6UcLkqSq8si0f4Yg+Aqvd/uVE9aVYocdVtqz
X3g8JjlGfw+fBKHBQ5VRlHsPEWXC9uaA9vGNOziviNQAeEXCV1y+MuQ36k5UdAA5
gnhLPP/f4KojUkFeC7Sm3jjUUGVpWyvxk7Iq7Dpt+bRRsObUjhO6qLynKFO1hZJD
zl1MZhRWoCaMjqIxCr+Ly8WeSJE6LX75HYxxS8JrEtdjUo/+xqfG9SM/wz2LgYtO
BE7czR/xOmOVLh+KSZ+ao/9xp5p5amIwEka8rP3Yx/qk9oO5bsdnxkIOXN5iZQrB
hb3HrzdH7IbDEMdXWYB3y8fZxQnp/jbGBfUwBOt0YhDGrThO3+XxvqpCRFyxvA1q
slQOE6MnZybexDRJz6Ta5ogwIiDJvimJlyw9ukq9SNBrW83vX5BNybqtBwXtsrg9
C5FHhD1RcG+V4dosPzlNP5movq5LejZFS83Q1u04Z6HMB4vgVUZgalnJA1gJM0fj
Fa99Xo7FU75fL26MyeuzOY9JT/Q4lIPfREHD8O1EHA9Kk7whRnnjFeQ3PQyW/i55
aiT9t8qgdsORAnRaIzS5gmL5U2+v7cYngtzteKnOmhAPzyga8B2NbK236kQmAawm
43aoszwqGf1GiWHRUrdt/zBYSNHrpQbf8LPdK+kMW32aihQ73t8Np0tY6ylAZydC
mHf7FM2+2k3g79oxFbSx2Hzr1TVAnIhaRY/C9WLVeqDqtfKr1C4Sq4UUfkLJ3IRb
s/JXQCbGEz1e2W1Nm0TzKZyOPU4mifzVpmpk2fUoPJTYjhvvgAmY+dR5FkyGJQmV
KDnNy0X/DfTAVXYVO8E9D+y8iPtDRdLgtCwH1BzZLnzc1GcTKzFIoBENbfV8wgJ5
Pht6DVTvtj4sH/ELgQK2JSCMxYXzPTMBOfnU61eQrqAmKL7tFsI/QnhSPUdY4y63
3+8QBrmhpVqDkeqaFD1iMxfDwq3cWJtrx62R2vt8mFSzoUR6khADDUeETCA7a5fS
ylab20Hyifw42CW573rD5w5Dbe8xbEjuKXSOYbk1t7Radj2VXxOvQg8EV51cloGY
/mcyqG5AqjmvFJ4aP9RJmMZi1m5BYEu5FNI8uDFdJY+T0Zt/YOWnwux2AzN20z6P
51HIz3kA33aRSgkHwiZB5dpOhUf+CK+47oOGSZXlehqQUtmqXOakfLd3GiCD+8F5
w87J4A8kjgxZK5xag11riZ3u1FQNU0Px1wvyRDtniH9dHD/KpkVGebtufMEkn849
DUxY+AoIeZE/LZE1pi6VcanxU07aA0++939+PEzsbDjpeBN0kAEhX7+mYftzxbLa
rsyi/PVGBU170JExlHyOpZ4a5ZOtL/acbbPHkP4xHrCi4OJ06vDpXSSn/7G/+3Da
VPd8PQWlrIJOE0A7TxcB2Bk63AZEb1pguWl89nG/FflbJY+PtC715WMsnI/adxOZ
1MAXEeW9bhk57dkfQHljl+8T8mPoYh84oYW5ajKbLfV+DpNUrRfzqStTOKz+IqtD
oGCtTLPMCwJemb0L7Q/mCsM0F067oe4KBJd9k795F2N7Y6p+GGOVFqVV0XjoLQPm
Fvl4LNiEc46aegYqsbaEzDaSLi44MW8PN1KhszH8ZgAYFlQ4NABAOpKODbRgnfHj
a6/MPmv1nb9NjApXtrqf8crdoBjE5pd16Aee8RH5E6Qavn7indQkzT+m4zFEcM/r
yBWVdb3VzuX9VXB3upUBj8OeU6x+pb2aMuO9bfNCqz8j9YsnICCiW13EH7kTlIDh
ViuhUthk4jdFYKFjCTUODcZCGz4AaYKe/iPOHnoNaW/qSqLj5rlz6RfxeYwsbka0
z/j4NehJ39sYx18HOBJPgHGiTUlqPsV2gsdWsGzXhvgsC9DVWCTf0rBh9pUCixhq
y8gavgmdjUVmfcRIK00I6OhSqqz/C3UsOudX+xuC6lQgWBCeGqinpt1VpyD1wSFK
h5noLE3wcKyaC0148qkLvsBoUB35QSs4DqSMu2kF0LGdLuA+tE9OjkcP8zC0Bpeq
Uj7C5wDL6W1pSwNcs//0gaiuiL/6bQTezmPqPAhMg1T9YQyh3xBKgDtVlfldGFyX
NcpM41JF8jGd4xcXjx1qeVaI0JRGB0xPiq65ax6yZbQ1roH/MK5CZqww3DB3jJ+b
FSfR/vZx/P3FvMzsAocsdWjQBSRBG399xngERVClNv5GvyOT6qs5S9OmK411YK0W
WbIX+IDqihVDkbt4mI0GGRqNk8eUpuvZdOK9iQvfj2TcwwzrUYd2gO4PvshQKrsR
4D2iYRvkTtEb2/e+NXMvLkxNaIkkIa0yNHmRjHinWwhic2MMn/X5yOQoOF7njLtx
BWA12vlRHdeiWK+qSD+OXGbSsWoZC+gV+1/uCpSuJ+eLrd9PYv24B5g8lu95PeXR
Y0Fy3UXb5sEdDp8x9H1xaxE/+I7zCfl+8bFionHiXwQF/Gaxdg/m0/zPgzo+zbdT
+Gm17gWRPVgQfgXwUESY+gQqHj5tVf/D32wh57vC+En47bhaH1szfPRev8IaiVbV
OUb6NPtnJGj57abceoaXMzXjWPLIZBabJPLDiYnFBrShuQ6FIv+j6kzWFVfxda85
4cuzlpQBhUU3qpElkBfLgrbUS/sOxYaCncuYS4yKL2JolNKAJewNcJjEz2XwsKwO
4DQNqVimVGzcGfUIwWtxX4x0ydEuvKd1Eh+tnrtZxY/SltMlDzIlJ3p+NiQki91u
aIDIP27qd5/MsUboBwdkJnc3WxRQeL5J1LQFgN/2TqTffb0avWNVoxGEWRxGqAFE
7yewdTc9KwtdjEkXm4jy1BZS54u/sUqWeqykSlhr0sXvVqSjyas/Gdjq0Mv0qDi2
Ei2OYk104v2uvlkUciRj3YkegiHk4aVKL5YIBKccWhLaFjBB5HFXZJVxAk32x2FT
/bNd9tu8dtqAqFtEUjtc9ZaGAVLdIn7p1JL1TbBte7g70eDvxXAEfTAYFI0LnN/9
M6W6LMC6Ngx9PrY2UPCD9dqfgnPHu6PhfKWr/Nr+sjx+h69z2AleczLitbFk7EEP
Yy68QYph/sLOO7WgPNs3q/gRymvwH8siAz1QY2L7fpFzkL5Z2I2JCZrTXYvNtIZ8
7vzRZRymrbe9QXagIeuLG5q3Eo9VPO44Jce9R7PP4zZjF4uKTbCLBtW4MxGR5daz
XxHtXOTWNRDeiIvQWcUUFLidw7YiMsTB9q/FjRxuSLTEZm2FY8kgx4edA7QAjXN1
0bCtjS9wmPf9nPhLIXr+riN1gHdCk1NDEkNGrrekCr8HRb/U0cor9vGGV/LELq64
v4lt4SkW2R7RpaXaRDeKNnkCGoXUVwfxDib/Z/2MZ0aejTIvIYYGoxoiIVfh5rjo
r8wv8apPOsbgEozgjA09mi1ygq2Ivd7G7AtmzL3AffC8pa7f9EnRPfZ0LFcatGmv
BAc/5jOx50gs6Krcib4BfOHIFau9qKyX/6I/H3bJZaBoNZExlcqFkfhSRsZN5sSC
6nEg0defrVdybJE1biHdlbiUSiKXqIMyJxR53hjc4BTK+u9pzOhpI/BKumcLOI+O
EhqFk4qGNCvGED5zheNYhv3B2wLBFo6e8uFA9kXqg2bNOFHZpqOywAFt+2A8IqZ2
3WGhmusOVsKrejC5MWPxFOaCNcD7lsS9p4Ac7NWNxO8OVeEcZTVX9kzIgDXZkXWj
PCqPhqhgTYMOdrsazDM5VSlKeIGPtC+pcxkMglQErccEFoz230w/iYINNergVMOe
BiflyUP06/EPmEL0dVkdr8eTiGS0Y9Jc65K3Poz0TLlEIX/JGyaCdUMNCJSyKOtU
H+CfLHJh4KjbBpNVMtYfH51tpe18SgpklgDZB4e8CV35hJmXjyXTtiD0GRqQ0XGV
yhAEzgjRgV1lUBRaN7uOmK6AC6qoQE8LG/MYSzAUnL3UU3SqWdndByly8SXflDTP
QK14AInnXSfbJf2ppzCifBPv2ErJPJV1tO4IFvy+bC4nZ+DK+LX1QCnq4dLNuvIF
wWbAMS4hUIEkVHyKF9e3RjPKhdYBHilXFsidFOWxKaxULl3J36ynVii6ziwAbfkx
OvFneu/HA5zqHhkOXSSf3qY3tHn4/qL3J/xgwVuJ2+kN+aRgZxouRsgWgs7Ipmo3
S4Krt2/g3WNOf1BwOEDjmsei7tgBaa1Mkfp0nGqRfzn2L5SObasOtab2HzgW3bTS
DTISrhKfsVMgcrl+wQ3xnLbnMMnj0d05gLkrZJ5EF0h5oNBuhuSug+2NX/5n8RIx
5jHfG/0mJvRbczOxbvUUvwoa9JFjJACRSSEIsqGCzFgDh+v1GaobBvjBal1vAzR6
nTkKBi4TTj8KAprb54edadM4RHachYIEsFU79gWh3eMIT22NLbF0AKB2uY+uDp7Y
Jf7CXyCfIc8SFV7OiiNDMrKplbzcLbaNi85WIl7ERaE+sy3GH/Swk/udRdoJXFVw
lueBg0qaz1HGMcxhYYFuKrg+Pf1YL9nO2ieBVsOSDBIK7GQ0v1YcU3Gx8OeU3TLv
FQCu4ZJldeADXy4PKzibwnDMbgQ0FCOOLPqf7BmlfjV/wn1qnigO8psIZAvijbbZ
9seuRi14TjKVPh//lgcAaVXGm48cDCOM4OAciezq5xwPB3XkzojEiBy1qc59OEXw
l8XkPEcD63d3LIym+DNYG5USt+r+ZyiFubXdxAp1AXKyfHUnMDSWZF+nNaWFwIxU
Ekyy8rhPXRlG/v37O6la4jS7Y/S8LIUE2oRINxsLx5QJLSBnrEIu3+ZpwN38wddF
YHY7k5P9xA6zrsH+l2T5caZu6bLNwP4xNqcycRf1uZeysZSxkboERYLrndKGtJ1O
wCqi5mz3qPsZj7oG6r2t1z8gIqUQSt3nZf8t+EXCgKDIWOfDot0/rr1ZvImJl34n
CL7UldEumduK2OdMIu1cYuxm7NYy1PlPSSKV5Z08Aue3jkncnT/l9HvzN83/xJKm
M8qXVgQ7299isJC9OaEaIComHuZ5rlxK/9nKImAN5IuEgoSfyw0PEouZ7t7QPGJr
/aTrfb4MqUaeo+eD9kUMCaqcvRTlE/ebU2vWwYH3PKxB+QaUD/4dVjp4NRQawjmV
dDdrBDAD3qqyTDYlKeAGVSxF/sqCKkvK6hX4D/Auea26T5cKd9i4PUO82JCla2IN
4OR50rlaLrcgdE8ArvrVxRjkbcRAnjygCeXjJMMz2vv3XOaTb9Kt00VJmmRY7XN9
u7Qr2+llUbmOUnJNMOtTB7Vnhe6MaS8qLhM5qYs3nxumr3XZCi2dqcovPHhJAaop
G8DJgBHpoxLstI4KxjLeukzoJ7Y8khnvqG4lqoEV/yj9j7tG7iKxqGNDVKFG/QY5
gV50qChcqFdofonWXsyldKmJMCULB+8lUrWZIQ7JETsoubPedtru17lHWeB701n2
dPQjRfSuBUczGnZiccSKqBYkD3pyJY5TIApmp2B5Zop/ooPmOfX/Php9YsORDRTi
HGOnObCpXLY4vPKC6CC3nZgqhYSLILByISxHeeCrKLgpuJxHFX5Ogg57N5mo7efd
lFpF42z1+jXwFpOHkOOGnZxZ5QCdQHSCZbZ8vJlHfBF3lTiBVlq6PaeaGaN1wHpE
XwE/9eO9eIe1fw5MsbvrcVAaIOWGOQyY582AcJvQUJCPMHF4eJy3a6Y5K98ByjEi
fv7k0CCqgn2cTomuUDhb+rVoAorkjOdXLb5qTVwBrUUbAw537ECNW9/floAjoYC4
hVicJeVSvOTwwcb9yql7IWuxwIW+vLHmTFARh+zlGCi1ZT3Vm5DbebmvfajKKsAl
HQIDM9qejef5QbOP6M7U5McNTXEnUnys+FD0I0VXHk2PHWYJkHJpBg5FbBxkQfIU
n4mDCNzTSAHXPFL6aX08wAv95k7farxvFIwDDlSWLyKGEelLgZ0+ODxGs6jXUzCJ
R+AdLrSW/IpL1kmxyTJ3Rj8Ft8+0F+fCzohUccwb+zv5V9kG2rIIfYg/9h4QCP8D
P01/WdLy4gJl8oZsOoKgiJdp3o5GrmLBm8qXaSH2TWsjhKBFzO/eccyeeiTizOp5
dWKt2NSN25jrf0s5Msmqe6906ZrwLpvjExVX4xcdSqLi8HtfaHLz8rVkouloHXI/
q1eB/U5OLXnv6sgGvDvRXX26oB5aTTObDT2grrnJl4DLeyF+0COu/aEYdbsCcjXQ
rvKcRVv1W5vXgR8Vk/JiOCijmkxKLwxDndrXK1zmk3zxACGWPl59oh3XM5oOeep5
fLE+tvPQwZfqd+M+YeP8rkHw6lW6n8mdK7wzIvQfUo2KhmhEerfbMYQxdCKnJL5I
/iWyASlrZYjLmy1v+rT9WnlJWaGLBo7LX+8YWr5Vg0dnOu0jxpd4NlmoH76qh2wS
65sCwWlvPLzq/jz/vQu5j6bluBGBTChZX0XXPv3UyuHLDM+IUIchRtoshqhKhNPH
4xVF1pCFIhvXwibGrHjFm9ud6j3Ggl7Ebcn9KzssHhedoyCyeBna2n1Wlco7T1nh
seswBoTgujH+Iqh6yq9wsi73spt3o8cjMtg9l/c2HedFsMngUT1jdPhCfA0JqCxq
Fd8TxQFTnGfGUyy2ofz2YbunlUAQYee3rB6AwfP0DnGneJn1K/V2733WDCmGgQUm
+7UorbeJIGDEhx0ZtOY2DQ24LdhnonFX/hlKH2sig/IhbaXJb7w/KDULCnTHlE/Q
Lbhp3Xr2MjDKYXJVE0qybl1+qKGrRgQGbu3Ng/yFlmdajdm9h5jImosFDPQgRPpS
nhPsH/MbUPY7PLGHC1Ww6CXRRePgSslQjS5z4Lyqs7B2ivru7cDzKWhW9ByxTeOL
Fy8IROWARtpbxl4etuZeBupoILRJud9R7O22KcT3r3H3RGIWkdhv3DXmd9IZWuZF
dSdUNIrz1/rJdSpSAI5xS5ty8/3jjWtZS7qxtzEn7m8/B6oewaQy8riJpOmRBMiL
JlntsNJVoXQMIUCVUVxM/kM4XKT6OYvPI07JBFEpqoK2yYgFYOE4/xJ71mnkOLd0
0Yhx2cYnX9to+0DceE/F2cexWYrgrTgFtjSks/+6Q1jKSIbdnHYYEkKPKTIqNVNI
d7cvA5wG5CYLQSnHZ0BNMhNp0jUuQxtIcZG2fxT6TAtOmUnglICfMhARR40/j0NF
a9c0NhIGOAq49YhlGc03XqrrK7GnfDFAecT6R7m60olW0YN1lLXFbkzSMrQVsTh2
OaURggTh/jnI0FKioZOaPGx3uMyk95PGz/lKOUAUCnnqovXtUo0GPpVU2FDp9u2e
+1AcnwMd8YHUS9zl2HlGVyTR/iDvPucP4/MZxQeJDvEJzIfg54Gc5VSckUbVP12Y
RTCLYjtWng/v6sNAS7cOhAtqP4uVL/Zcf9UM+YQHVX7OKVpdW4SAQszXk8kEotES
6M4SjqnqNwIT0wQ3f9S5v91kCl9Oj2R/Bg1VzHEc2GIX8C+3RQO7rGRj+tTwqIFM
oFXDtfnv8TKkkCWZoIMRJAAA8hiwvZYLPXTN8jEKp/tHSkszwkp06pupsaOXQRTi
DLjcit8s8ueGrHHSio8+5oi1TnlDSrKxRUQr6wsEO7ipTLbskddZxQ6DUK7/JGKj
NWr51qteijkuqoRjy2BYFyIkO9YxknIqulMC3wEN5GHNoWX39OkHbmBmEFs4qQw0
E82NeSJEyF+BztiHwRnbp1cBkwvp15kTenk1DdVzCAQ1+XR2u695/TgM5VMt7mQS
VvScURQ/EQpELoVmCNZzamDojcGnOHzCDdUNoPi96vQHsHeVlxIM3XmSvLtM/4l0
2pGEUs7KmhMVbsyqwzpEXqdK1cuhPt4Hpetlcapke5nbBD5viinK/yjGRueuJSjN
r34pcWKEWErwtDjhQLngn0F8PfIThlaYanEaZabvOkmC8OST4Tai1UlBLOxgvsB8
rmTNAW7qgQTADAmo4wY+3crHRfzqgTs7hWFFdOHjBMXX61r/Qd3riLhwH2/YmPe1
FEIGdPBpJwlSqGFt/x8LQLQYDmVqb4OPtYnMWW5mnMKhrVvnsRpAVwWRSTfgrsa2
cKhfo8p9fF2ohLWa1TBZSJArlqkmj210Htr8eMFD11wAx+/R3XNdMjc9G76zEEWs
CMmZsb+5vpxaGHK+BfoSC+LUnPdLy94da+614hYe72PlXFv2cWsGMCQwjPdnQIKU
j2VidsYOyHPaMoZ2CrW8eNQopWgTj4b1MRZSP4ZgsyZELDpfWka42y+aOTbgjvwE
O6ig+lBrqi7o8zODhO2745Et+pFMYtlKSxBkWg+QASckPR0evySgGndd4+7gRSLY
bL88KEB9bs2kWbxJWA6jnd2fUdU9V4Vmqemj/sOrwOzzr4Sq44FrwHNAbxv1iMcr
bgPDmhKMhBqpd5z6kzXRYKTHjDG7kv/Atgv1FPyw/ZMojALtt18Pg5LduLgjE4oy
Hi8gXChIYxiGnUJ/sY/VCaMMrB/4bmXwOlEOwrCvPaF6BZ9Ca9I1QnpQNCyoJe+W
JFT6z85pMqYcI5RyqwFXhHeQVF3CmsHqaTluabkaxE2YBRFvlB6XnEamu7zy8NT4
ebm8yWvENjUWeOJh1qqM0DJyHmuOckSGJcUhxmxExSoSkYfi5qvQzcpl6ercVoSa
cTgArZrWSIl8ruLQ7CXlIHYLEv1N12HfzzY3yDE8hjSb/obiokPZqYKVfF+6W84i
ILRcw1ig5S1ntBJYxjO2TZrvvKqaXsZozoshog3gee+r7DzeYPlkA2TalkYHeJN/
hwzBeJEKIquhHrI/79cfUfe2K7iAVIKzRIPerqGyNpWDDjIWP/t83IoEnlhSqQX8
wkM6XVKbnvCu1dkxxvDT/plS4ZaMCoJsQCjoMp43dDGP21R8RrkM0wRCbwyeN60D
koEaj4u+6tmIjRNlTCw1WLvDD/hhrMN3Q/q09zejPPYCE9IfTYiehaoezgQiuZ4l
+SwN0b6fXObP65HnpX36KoqX4aVgOH82kKr+I5FULEU1nQayP7ULsj5EHiborr4Y
6wj7iuomzxAdW1MtLLY5K0nvzfJa7Q1oEcrMhhY44cPBTlg9FEEgbwVk3me4Roye
cHKRBqHaaCkR377ZILdi+qPf+yp/s/99mbnF8EzgRv1/ydShxO9hTegMzAek+Ryw
jBoXzN6sDcBIOEbO4laYV5ZoA9Xd1onlRgsUir6+fLSfhhaFMX7uHt5LgZEwMexk
bkSQfbPKtx+w9mksOGztVoBqLm8jCCKVPhLJRgyNcnfyOW8nTz5CADHa1tzIgO5n
lqFCj9AS28faJ9UqRD4eF+UoKHGo1rEZ20AZc6rNqATOAtvcA6N5GEIJ3aAhh0I0
OVk3vjtqe5axR1UoFXO0Nb0QSNoGcmh7v/10GRXEELBLEnmMLTXWkaU+fNfvDECP
v4ZmC3kLJ4vpUIxF2NNi8S07rVPW4+gbDsHME5TV5adL7FxslT0/u32ISQMe1qiB
2DDajw14HkzWC8v/e3Pya/q9qCMTuHNBFIvcnOBM62qKcMa0lJDuafa6W2kynOmM
mNCQmIpeZDX6mtDq2V5lVZOueajDs+JKjS7lu6fMxs9x/41ChzXaAfVtTc1uuxSg
dS/uMyyDFrk++KG8ey2yf5cumpA87rChsPsuYZxUM2kF9i8Nj3ApSIYe76yCI+nL
ME6UDUzsNLGy6a5UkwgCYmzeybDmFMqxPoFjTB+wes7MlKrMlWLrnp8A2EHm6C0R
NkUvyVB9qUh2aZZNjUcWtDOsZCX3Irv5v+sfxv0Dp6WrzMdibphN+TFC0qXavjxp
dlk3BjnSOzg45Jcrih60oB2JZaALBtJEiFHelqAoregQb9npEdnrR2C+a0orB7LB
BrdclaSb4q51mxVmML52vt39JGrbXPFW9FyKPTElGnMQnJ9wuAXM5m1pYN0mEfLc
5mQQooooFkL9x/q2FJ2HXZs2zFX2p8QB+wjWK3a2Vdiv0hWjKCl5zfEykQBfbXpw
DmZQw3vmVZ62UUMed24DLJnZorJwuWmjZu/AmYTy8VApkTcFfjs1gT4fBLJrLIby
G7NQn5s6Zx9WOZ4jD8q2s2SDt0awaQbFgylFQipCJ5EkHdDJf7A53kgKYebU3ANu
nz5wf6LQd4Uq/qinhQtv8qcq2bb4Swl1yuXRtg0bIM4sFEGVEgqqT/bSqc/JRYtU
MYiCDrqvnjATgAIJ6WjXtwjBU0bSkdbLyS/k8eIKUIhmXlCw9HkiBNCqMIkOVsPI
NoWqlIOe98nN7hSSwd4wMNEX9PSKGQaHiUewPgNCy16l9fkEINIZL2fA7lVPOAFr
qIr32w+66XaiGmL8373Y2X6GOKtEzd/j/AKNvj3ZWOCkJXCwW2UZDxbdN8g00FMN
mB2gvjghG3ps5prmNlpPT7TBPGteY1NOggvQg5uu7QsHEfaYm7EeSikVWNbq77OS
iR9G2hwK6hFkaZBARoKr03/Eb4PxucFVAuuFV4vf3g1SyeP8OLIRDc45JwSDr792
fRqOVglXqJ4edXmgIdKn7YdkIwx1qCi0xvCVGBKW0sm5KQSCK8GFbjNWt58v98rl
/vxIy2M14ptH6nuneuAFbZk4nXjJ0Jru3ozRXEd+iuOrNVK9OTnELIQCnMtZLuPv
AlBDcGw5hDrR797ailK8StpF0yZlqq7UQpgoHCYWlrVH8c//fM06BrLGEj5xeMQk
dE0iC1Yp4OrmeuP6iNgaYHf3RzGNn8bLRXtgIvpctH/FfLJZ9oz1AbiWJl6Pyo0X
ZtKJIwdt2HEzNDpV+XpZ5FoWMHtv2o4vRoZP7Mu6sBk1mlMQOM58FNdKgEBh0rm4
AHzAnzRjv6Xc2oE2cE2z0qChDAx4oa1ge50plMA0DMEBLvxIsMztxlKsx8WdVPIW
PtWlPlLy+Gjtoxa3eH4sBTWR6wuhT51+LmUw/LBzrCjRdmss6gGG0H3m1BMRMi42
qmMhMS4dtQb8R6FjOWjbJvFDiROhWvVSTpXpVbjXS4zeY47k3sfrFSpQhfTR8ef0
+/xVnaa04z0bjRfLjSIwMdZC0IEef8wrkxA1f2/59i3WWX+wL5ASsamefn3delKb
NnsYUrSZGk6jrmL0L3l9MH0Tqc0Kz+7+qYI0UUnKFB6AgKj4AA4JGwqcnPMQiBA7
HjBOIVd++dYIYIYwbGcEY2rWP6rX6G0Dk8p/a01+YJa124OOv5Q4DiUX7TbeHCYI
J3R4S0W59W30XjdinWLKzaB376vC2LlvnpkPe/PRHKtb2udrrEFGuSwEXPQ3Knuo
29srTz1qv9by9xiLy56jHIXIbXz4g2tZMCkZBcRz6opHNrVYZOPPGAn9cvJ3FGCe
n978BuzIuZUu+j4wLYUG39pzYWHLpPFMfPWJENLh6eflDHIWLNP+lzrAYtr/kvuw
Lz1GZh+H0GUJk8BPTFKT77++DoNFtm61uevRKVpcXAcen/Ra9ThBb1Acfe7pCIRy
fkLXR5lYGPeNPxUyWiooRg2jiOw2r4q+FlUQizVd6vG2oSrXntql114nAYeCkDI4
5bKUcaRZ30B9JS0mHSpWmWVeWK6WHtyajxP3xXNNMp9CUJTk/9WCcfw38pDChVhg
j7UKqPRhCr4VCWVcSA54F4uOB3YJPi8DvgttyxS5bmJ1dbRokYpmHhKIMGJhuTyO
qcSXAfUc5Rr3k6eHcW2XQwIVMndFwaERd0jgtJiXCsDjyfEiqwSxreIGAS0nZcll
vi9RU+NS35FHjJJl/wHMcaI60Dn4G5Qz0HKj4GKHPq6EksELgNokRGff1IZAULQk
Axu9ijguO5CQTSoLiEzoWOP7NnDiBwXaVZE6BNpWYK+dwhTokcaYpKvmQF0iSPpZ
VsWkWuCarLQfASAJNARStKZc5BeRwErQiefZZ+/QAVP7itddwdA+KYeTLUBkA2HG
kxJ7EjIg8FhezaiOZ+Q+JK2dOa0UQ3WSic8OtXawzRq7+Vb8dKJ8IIG/RtWhWzuI
NI7CUVWNW0lFZctB6OMM1UjCvQ/OW69nbM74XXr1AaA0iteC5PjNAlPSd3bQYjUJ
fFro4e7/wqTvSJUowfYy3Ptakz/OvZBSiMDN7LZlZc4X+9RDbK19VZXAX4rqnKCH
p4jG7wnlYNhNw55G8lS9GfEgXiXcsp76l/l/lwoMaD74gBkFIYRtcWV6TdHDJg49
2bcPrAbYix5L54Dk90dTCjaooaySWpOBiiKwjElnC7g1CO9Np0QPrAc+fb0tOKyf
csL8Ald6eWeDVZxRjyR1SHBqnojw78jrmDmzhg5En6IxhXk5bbxEsAi1xHTk8itP
345B1k+RXWgiY4zW098MndFtnxSutC/DBog9x2uzAbwVGsIl2ipNsvohHFqvUnAf
0dXpNPzbpYV8E2pkAiWpn/inn84PRrNWzPx6+8Z6Zj/IS49ZfLj972abGfUv8L0a
BOxe5neTS08GbcmCpJWdWD/ieD7VtKu9OiFuuBZaUujdeyeI39Ue4Td7svCzigAG
fiEvg3t5TH+b9L5OB/yV3VpB/WoJwLqeKc6/JkeD50BxUwPrlRhJks57FNP0im2+
o1Z3e5ghzp3DcU1TCVGze4oEAAqZ2G9c/RzU5rvMMCZtSQMSuPZQptUS5LxUS9em
a4BtzfFM0v7Tidy7BNKTQ6e34IjFyuoNmLcfF+vjpY1dKChesa2WeJkLmf+Y4l3+
f1hupm2MlTBZRW7PpoiiEl+74cfbyLXLPR/rWY9AtILMbujl9A+T4Y/yDwD0UkhR
oqRNQDMmPauVnrltk1lXoDhFh1P64mesB9wdmbAs7pyyWeO5WsKO/YVyhXzznLyE
cW/PHfLTRcjpD/L2509y0Rb3aYO3Bye7q8+pQUllXaUBjOT4HBcfmJAzczg3aIer
DcYQ9XupDum1ZXvhnI5B5ufDAXwKMkAb472PMP8Vbf81Jd7E6tEQ+dNe99NbVSXJ
t/A8hUPoBdsVjY7CUaF994L+jiznWKB1xMEcVfs34gKOGSahvPVeBBdr6bZyO5Xg
QUqokedKRQgUtCcKHJmYjJBodP0hB0/SJ5xIPhJp+1Pne+ZFuR4gLOUTdqjQnizs
URm/guvzufWHmJjRAJ5TTNMMruENA+L9qI9eCt6zIg3rQ3Xm+5THkPOSN8Sh1d6j
qcWMJPm4enNrysobj+0N8pTV+4NeZ/YVz4blngxWPSEVelQ4WvJtPa/vAFQPMhqZ
eXw2RNZa7sABBQ8b7mVVDA7K6VEmnci4EqKtugg44Enh0gsdqLg5uinQy2w+XP4Z
iKYIJJEoX/CmcBcK/hDvx9o1uVPH2G7RDWxydwgq4/gImBK6dCYA/31IHzKKTrZQ
LgYHie66nPVJ3gPpUeLvFjBhAjdhBuypbiEYI6L1UXrTe0/XutUSsa1MAnZvkEWP
/KT8SIxAhEgWZ+OCyV+N7wvYtU0DFRwAmbyl5he6iyrcoWr6xhICabB/5yP9qKCI
X6roxECXe60rmeJMnR8S3cmCeLml5zLJj/AcCgn15Cd/w+XFJaFvDk99ah9yNQZS
S6UExOczU5xhVv45hqn9fyuW7hTe1TIjpnXslyh6SSxpRjdCGKKmTZgPmbEWXbGt
HOy2hZAVnSbl4HLqVirOTOsW/YmWJydu+XA00V+f7AWiJRQEunJxcbxkAA8aCt7m
fXLBRvxXZaTffG5/e1oXUGvCTgDWatGWfBareKsA2NUBUlxDnr/RnRdTq6Nv68iF
L/cdw0U2fUk5ZUdnx5maGnEGgA3D+yfFhbBgR7aUBa5CFgdO3QmwZmiatVQMEO7F
rSpFbgp0rgxGV7sVjGRl3fMZPvUTBlRa3/3x4n6N1MKClqHTvZ+oGMDVP8/njgcL
JdoPAOmiSPhu9JKeyNTs20ci/WT3BM0dG514Y3pZtMtIGvOOTcjKrTfx7R2xC5MN
WIVooJoXeCH9rPsM0wYGJYWhodOlf6dttJDaW1SULAU0oPMOpDSqKF+6owBbfP23
PY9fpMhjniv+WXbfO6BqSM1VBYQNqYVEX6eya+E1zAqxtfrHBduwDs0ehwZHVzfF
GX5ILryfc/RzEDPqlHodVQtu6cujcDC8c6xFWTU3Ezv2fqLtKH4Gz/nn/FqV3KtU
DfeVP99MalNB0uyaKptWnOx0YPdipffSITNT7bdvfS+XY2XaXF+b+Qp6ydo10U8W
s9heaqKoPvpHVNGIDcWwGZvRy+n3np6wfMHWjKla0A948y0fVgGGqDyt8b2kqC4+
ZYrucEk38/csIE9YlDAbHBtwvvXnLrgTX0/ItrJRNTjebuF2pG3lzJ4TujZ2eZjD
K8kEVAh8ujVDxsFmwrRGRL+CdrA6TytX0RHscCnrUWAU3Cct/pzy6d/QAWGGoY6H
nvFRIKJEzMWcUMGQUtMCen8ZvvnR0vdhiRCjLgYECKaFpigFuvtNT9SYvdQhsZjf
Q4lORukiowg9UCq6Lw6Ol1zrz6dwVXL/uTAnntKk5hAdg+CuqUpUbcUqM2R9o5vF
Ev/EMo/uORQo8YepNjrg0TC2DHLbqcj4fAFS+dXQTISf0iYE4HsfwBeRlLVMYjaC
9WQYvHciGIXxsvS2UVAbpUOWZ9KRFaM39s4nmmDN0tgH49gLi5NKd1OMc2j6QmKO
ugKvVzn9xGENCiDHJ5rProdTaPQcEACLQXcmJtH8GURL/moqPn/t5AjbW6ZP2oJJ
zdCfcVA0VtZgjYuHe9RxOX661qZe68fl2eUe8TlaKgLXkLgaU4jLGHBWRESrcz3P
8U8Ft3fk5lWN5QX1zd4HN4JP+195jaOWn5GWJNM9k0FgNS8m6EqJbKMgWXqCA0nf
T4Dbdc8zSfL3g1biiM9LtlGsFBJvX6HdUcfvhBBkcgn7HBXwAFs5DyIwE57X5FGd
49WLNAkh7T+bBHNIl14RxnFbR6y6M5DjWMBcjnbPbxP8CELYBpBdJOAwJmHQB9Fh
fe2dwE6hkC36Jl6p0XWfVeWeWGRjeXfxAt5RABde84d3Vbzhgl/p+DJY6zKs3XRu
wAcvR45+KMEtf2KmZcbej7s+iYg/oLNkYC636x/Ya8wNmzG7BXKs1vp3gm983Ig5
oJcCP3n94B8o4x4gppRwTVcDTAWyZ2cnyGRf3mN75nsq/fTVTzoNGPOw/0Etpp6F
b58vsvWp6kM9SVmR/2/CzqpaEIshDfuRuadoWC+XyIjtSwqB3mXrl8iQHpxcfKWS
t4QyqKuxsaBquIIbVF6pg0dWFCgKX7nbTfLqAJtoH1JbNoxkOWEFwKUA3yoro2GM
YUr4XP7YP/khTgZMWj9YPj4yaB+IukwUJvr5kBmMKTC39vnXQGRGvv9kuyMwFJXx
UlxExL6FC9qN8xVRZGvDtEB6GYZm8DaBfhmzYFZWI6pOdTNNBn6jfkYQl3uRT4D2
RwiLN2XRtyWIj8IjhMt3mPZUXimT7Ah1GZEJNH6c4uszfIv/6WYqczrA9elrZUO2
32eU2yrrXLQYRf39nqwuKFchd/zgN98x5o78nmfqPC648bu32gkHavSkZxOGk4xP
nVIKINVU8B7NH2Xmhqvcdt4yUIFC5mrfBQvWaXMozefG5K+Foa2cHnPFCWBrTsFL
mQ6iOcqGLMYpzdqRJV/nVdw5B9Lcj5Mf1RVc05G68UdlQKpuNiLemIjmsEcbZfvJ
uRdYm4AghjgUh4O/9JNudk2kx6hTuU5OTmi2vOQrqQwrj52ZgS1d6z5AuyZSP9Yr
KZW4q44AvRIcbCPIttZbxOv6UrsdcK5jHrI1r3B+lPq81p7zadGK1Q6ZKGRx0w/V
r+Pa2ddCiIMfitL7Z3TntUe3yazsxwP5sWK7fyL1jfNI2xQV9xhialaRUt2ncqkn
OBu2+85VyXQMFmIYv2p27/egWZMGxRy/PZwWPOfAgFtnjnanjm+PKYxObdE9KAgZ
rCJ8EjV3Yre0Dlz+UHAIKdF5fe23BzRwzKrgiPnsJ03tET1v9aXNif+BuRwqTliT
IU9Xw7/jblY1kZ/mwsP6Cdaq6kcfMXbrv1zGnNIH00MSV3d/hhyIbeMps41nElb6
m30G+EE8B9OwdZLQPqNmxqy+xVo7alb/andFhNME2zuk3BD8Mmg4GHV6u/WVZlNS
g6g/QEnDH1MG1i/X/zsCtXFkjvjqbut0MHeHoEGNPgrpvwBAGi4NLhF831RrXZhb
FljWJCMcEGsZ9abZg2KX8rqyrt7q6QFhWbm4WqmWZC3+WXBtqs9p9uTy/On74qfG
/bpxEnUnBrXbFsmnt+IJrLd2S1f/7by8TLpMeasb6HeHGUJSOgROfhGCbpjGjq9a
EBZOpOtgQgOMqPk8hYfDqn9gcWKF9RgNeFYF7zuxNpa03b36ywIvlaAZoBM32Sjh
MMV1rFwUOfuzcHc4aQJFPsoGC2QaO97xf+WI/3oCNQBkMCFR/etr/IZjy6601EKD
dPt42Vk63OwAWmQ08dRcwChMLhY5P7fJUb+YTQYzrqKzObmz7BV3pxqlSh2wc4x6
4iaBEye88cIWIQ2qep++B+7sz9Jf9giY668oVPdtw4Fpv7CV2Lg+w5TL8c0IFsPk
lH9ds40mXyYtGYEk6pDBPGf4eV1A2bWaJLBnOahKW2Av0arfGhfy/A/sqj9Ksu5X
nUqDCOx0datrd0LKH0+QYrmYO1BE2RPHQmeKquDWr4F6+Bpuj6iT7wDtB8NGCgCA
YHLfY6fY7upz20bP/WWW0M7MUqgg9qtutwQI/EBz4DgHwyKHzS9Y8YY4G8RR/bTk
Lj45ebNwqXzgZczXAvjAvAk7t1qytuXNkB1W9fx9w9K1fQcBnwxFDbUsR15qxIw0
nirD54YHTfjj2e1LDvvWFrNkJNqQ15m2HfpbktqZw1SrbX+1o4NUi+sB1E85jhxb
K3Wq5KsmsN/3480RKf23rCN0kmur92R7yPrz6eZtGIUIUivtysAnC1uzdu0kmRsN
tCbIVXrk4U8sgWso5eGoptJxrcrYOCqGp5QMta0XqxkWe9tooMD+cQ8nFluX1i7n
4doZiIeLRuXZunDTGz3hABZCBWdxB5KGtseexgW15I+BM2187M7U096iCQ3POZWi
JS8dVzUUmiGrwnhOSCzByuMX+oQo4+fCeLPH3kkWP18QjYF5uF8675RXQ0zobU8N
xXPSAKbLZGtem9j7Tia539BpQgAbNadnxTW8CVIK4yk3AeZ9xtEf4QiHKz00avVD
UCRN8n8R+ERbrQccoUnPqcFPp2YLdr9kkqpw2Z357DsqPOJz38TGrPQnmZz6aRws
Lo5ZcBlnxnxbPNoQ4uThzj9EscI0mm7toZZdBomBxnPfJ89tPkagQYgY7NULXl1W
uMs04+/LcDagLtVfCCoKT3S1Ij7W4xuQG+jUeoF9zkyQgpXlzx5O4YDBT2Ppp3mn
wkTKk7oREYMzIkNDh9gPhOlxKgBvFzxLjwSicgCtaGP5j+bqr3Q3D+jhVI3qIZ+d
5JwWrLAcv39jah+KEefy4g74kfg7eyMQsIH8vQN4pk+5tui4mhkQ83d2qSH5ab4c
AHz9Onre3BstDO0BcvsnL6exTWe3Ut0zl1QnBI5+gclgxxAilHYrGWN3kEdkdLJ8
k4lRSNDyKirzrrnqNts9Vc+2raLtY1Rmztk+PKbympvVDX+Z7KTI+yGjmqATPlNd
YDauusDRLESXUt7kQgenu0E34y57wuQ3yYACBsj4x5nUciPlilMz9oBST6bWe4xD
Q6OPckOINq/qAulrebVaDow0JO3xXLCXuy9nmo8zhh13KDvztOgBKpL6E6vsPlpi
ZuO4ub2BzuIEzrCGJhp6uPSNhfNag8QKgQyA5CIwIGe7PrgVHhGeqt/ATwxvQ/NN
TAldMXKFjS+1kFF06jptxZEF+SLx3Ic1VRQdQc16fjbhHipA1xHDHYDNAxC1TWsV
K8XQLOjHGxRKj/ZLZrqHKJCANmDXG/4Hn9fRCZFaSERWEeVgIHOlhtLgjR9ClTtA
NlBvQ2EEJZuWioLaG6kJ3Emtz8isy3LfL76q54AEVlC/IGQDNn2R9gP+VLZiiY1F
M5ZKuezdgCQk3EQd8S/hJkvWVrLMUxd7dIxJlL5NdkMsddIgiQKcyToFw77ZAdVV
a0X4D8nLRojHaYHPrmC3WeQI7yc1coz/fpdgq5D7gSRrasKxS5R7bBwNOqbHE8O0
tD0z39IQGWiFUZk0588acC+ieu4urRl9HAvC5YXN6n8pof5dSVe0R5Ipdjpt3gHd
7lT87bcbgpRk2f6gqMMg8xuyUEym3Ugv08KIANw7mcYhMBer+ejoRYDwDgEYX0ap
+wLUWxJ7BtaRYu70r5IYu0GJ6w4itQV6vmaHHtb1Y+O5oZtK9ZayXSHVn6Arnlss
RkW6K/s9vu5rs5xWOUH5dSMU664wdeN6Zo75vvYF7ZMAjoJ0x0YQUFmjtsHmGvVu
iDHL6nEItsl/Q4ddGkDkJowDUqdAwVmCKQGGwbGxAX6HtY3hRI4tZKpTY0ZlMvWn
GSF4dIXkUPepAw9Y8dtPBVX59S9f1oKNFlVLklpSWXlZ0xCcOmxw4Q0HWk/XBrZb
prEPoX7Yq3tke7t/S5BJWWo3aFlT4qN9ySCUjEncMtMELb5mtukYQtYnF96Rg13T
iKwXzTuKn1xM1WmcXyLP3X4rV33sfU0kH5Q1vPfh0Iq/69VB0vGYM2ruFm4efwsi
9NEjtmQrFx+DcJU9QMkRcnng1nMSnJUzDNl5w3hR4ms2eejysr+B1DVqy/qUN2ki
i26FfBwViZhN34DTvJgJskJbx0ZoCFmJSxTk5Z8z2Li316dovtaMpKiDdjDy64Av
bUsaq5GWgcaMHso4UghMAeM/zULQ0LhHr7qxWrgnrBDBhAPVcv50Nf50dP/KqS3N
UKaCfprTRTgdhJ8xuQe8Yh1O8OJButzmEbnLGcDD5kpcB7jpIJzNtke/iYUoOSP2
qc+FubzQGbPaWDiqFf8fJwS/+eQxNkEoPJSg6V0JcQnGknmb3iBGymEnUYb/KwmP
GP6muILj4k6EsHUVJw46D52E+IB18dV1xr28m7hjYW0j5H2cuGpAfKrxu6KylZyW
px0/ISqHNWCCImdsv89Y20Mjrdvpha71wb5eZ6QyKgRjM7m+HGX1WlVaNxoWVA5H
mAbP8R4ycBpbPoaouTLoZAN/aBsOifpDzv9x2/tvgmRv9kEnmzMbaGA6tF4gqBK5
PVC640IQIsIBMM5Xy1Z5W/Xi38YM6jcnwFkT/99wtiAjwvNzw8CxTpd0ZPgUEQ5Y
BztYcuxsnqEbEJZ6aES2fW2Px5ptQkVgjuOV3wgFPS+PJgDxwx0GMIogQGHVOIvq
ql7MRn5A30492KtOsoVdIvrMZ2x1f5RiMQ1qVjNW6uB0JJEUe84ojUZGZR6nEmZi
KKnFm34OOshoVCLyZF51uBcxnBs9sClA3Zpky4MZlfLt9783VK3kup/spS2paLSn
4AcgRldIjcLecF7Aa3p66F4A+gjRuRuFRMRIE067OzoxVBdjFcRMvgLZjnGoBUZ3
Pcj7bDc1TQc8iaLOwn88vH+UTqFcPoGaOE5oLldzEtzZL3BNAoaxAjF2/Qlbftzp
lMoMPh1O+zKT4iVT4ATOCgAMrwkXuege1HRtRlj4NSPURufzgh/AGiwDqL16ESn0
3hZqteSdTd2Od1Ox/jaOFDsWD2HB620AXfxKrgbUlLxcihWBaMUn8PoC4MBSM3K+
1fby48FfanM733YIfGK7t2TgMn09URsfxtJiuZJAmD+fiHj06BAqeRsF8iEi5KZm
NqVHSZ71lAd5aqGV5E97GxuLiA4RGTOP9oaQKzuDUALzGe65BBekE0sS2qrA6RJB
ACm64FDkXdLnO009k5OikZbNCasvwzzX8OAiTVfrl4K2hmEJMcCv+krSm61i1u5t
TWdeQb5uwhP8vaORlaBl47Nne77idPU5KCN7MpdpPGgBk9dlN8cSeqJpF6eb7gGt
f3clrR7F32MS7ODBVAXZNHw4LxdP4PbHKyl/YmIiM8dX2VKuOaVM0dXHXSEfD46d
v9x9j0ozXVLXGjPHkD6Rh4V8/v1RyPaQaNy72UbD9asGRMMuQBooW7rLKdAg0JGO
syyQ66Ot3Vv6+GeKsrBPoyQu7tBenlb1hkwXqYDX93rkygUu1yxcw3moXA4mWY7v
efK/ldKn7VHK3U6jf0SOsuOvWPWpzlavJux/CYcvTAuSnZdIfKKkf99HYR3qMwqO
CKP/ExQSuHRTipnWRE3k3EccXq8GbXUvEbCxWkNvBRWefPRAD277qrlaz7eQpyGQ
67m1e1tr1VU6hoCkm5l5Wj5H2H97Ll6SLSc2d8Bw+Y6a5cx7DE615XBXavOSPdjh
5YGyLoFdPxn9dgwbHNE/qy5th6toNmsshfuUrVwv2ZVAR4He50KMZ2gjMFdISdQd
AXh57JNwNAL6enSkRvl8asczF+MdOZzUkq/v+qvcZ7rf8AZ+VwW6es72yHGWSKDS
cbBTzY3vG7XZXdkGoYdV5kozwECfz85vF+ZXJZDoRHnGXgYGRg6hx3j9MgUT23bA
MZ5jQOOpQ5VhJgMxf9i1tyJI1YLEOBaE/Al6GrC2q0SAFwSakQgdnD7L45QNwS6g
SU1Q6ZOw9yZEpi3LVs7FvtcDlpqg2hod8mductpURKCY/0AHVFl4vexLE5PEPtas
j1w+E4m6SzNUMNuqpU/Y+j84VrU8QotwA9iaZKFDmGyzCY9AZzTwTekGT3iCYqwS
QJK5jpkRkcafA1UlhsSrUNt+CjJTW0UnJXpR3dUbxA8eW8MvS95ULYtoj8Y8MUwZ
Mh5MdSNEFs+gvwIn/H4eAWUite8JB/9gqj6aFpd/eKvlS47Gdc0uDCmv6idP4OJ8
fyTwxdTo/Z95YsSdu83D0/2JWnd4lD3+2ttM/yvB6Hb2rF9o760VAW2Jl9qLF5j0
7qvVbAICtWaUE9O29O71OfaBj2aq7Tg/eLG2sbi3Hoj3+cvzyEuWOFb3wFWrc9y2
s7HIHG9Y5DdQ85pS1X6v7/5oMdJQmclpksaETUYVqav4/WECdfP+OQPh5UN4g0wk
Tg4SsLb2+MRi2uW3YoQWAqcTlnHqSmBlAiujLu2STASCFMQ9khvAkifqnwOI0zz0
Qn+kWDxODjUUxCZ6ImQ8ERtrVzH+neym9tu8M5/qfmafSx892UwQyIQ+H6V+dFMr
hMbTWITjmJUPnLrJtU2sSKCQ9/OMGgCiULvwi79WlmpL4Hb4xBb91nwyvRE2JdQT
jPj1IhQzq820vIsYip8m4IjYw3fmspRKyMd1AO5W1rtnid7meI+j0d+NYwCikiLi
NW5vo7uMLWcFOLDtEYq29OxNyWlglIsyIghng2jfD2zO8tprN22YtiaTPd+Ae/Mu
4hXrpHbv38p48iMsJT5Eti1rHUqniMv783CO1QiT2KMcDVnXKtczknEyInHWrMLc
h+0i4yRAoOMmzhafmnbiybFYKbY3+gNwx9OuYBQqVJL+S1r//JkkKrou6PkR+T0d
U2ECtaoCDqZ/X7/RREmoWww0QoiWcWFqpuS/1lKYhl/9KFHhqX4Sj3x7v+QBqt2W
tOIfp3dwMZy+Ang4urTHbLv76rzPfwEKAUGB5ByVjeQS5JtJVP40bVIJ1GUqt4i0
tq2OJSyEeT6Q/2TrqoaGnqkDWxUA1uFLJ78YkphOZTgBx3h+5ik4NMeGeSqAvwcd
38HQGaWGO7afx966m2g6kuQHwtDWZeRZiKg0JtJQvIRftTmS0H4dn854yAPvAsDb
rW3g49a/qJj08Y7o4098NXpDqQ/7nZotHUpZUp2WbDr6tBEwPQCVg+XUtA6Mk7TU
kCd3FkSX3LCOO740PH1tgR1PVQGXi7UlJRwqpqUQQFVT67maptoIcHrZ1t2kCDhE
wZCMD+wRRRlYFbzZAgwRZBH51FgSURAkalGLfJOHrHABTC+5dSIzwmTtIc57DNbw
b1W02ERLQPlhOJNIEfv5y9aTg/aPMlhzCdYfQgRPphkyjKvEP77nNyJOkFY5NpVX
r5QOWJjs1WXtjTXerFqStrQqfFkYU9wjKQhIwyIr/ClrnEyzn5svd2EvjB/CuYPH
akAFbhcQ3avPKcJ7Rn1/MxMhNscPOgpYLni0uJF5PwADDrXUUyUO9lFTcqOkOSdz
FCDjKydNMbsTmBOcTrYjiTXsKF5e4yWbIn4C9wlfirE32Ns1hecqgYjVk2WLyVfP
r91X3s4baYulZdMSiOanVBHRrTYyQXeL6YX+ESIdCSpXPDOfbkOrnBXa4jeA1AE1
uWmhkJEY0h0FbBvD82o+MDrcjq1rc5u3DgfSTfFiAWjpSnTCC/93BX0Ggp3a+MVM
YMKh0PkcNvch5yY7XdBAnho7jU9DLlgSuFqp3bSp3ju+dUMibyXPed8uIgeaeXb4
eOAmpNcNz76mGrLD273KDCgi3tfWJ7xi++ibHgBoKQfs/o0CbM99XXMzaC4FYFcm
+MZorb+zCRjD0NOLhyeUMJQ9z+0y2GcRZuDG3k/CWArUbFRqIYj9aJRkPcZ+fneK
zemDfqIE5mK4EO5J/wh/Vtv/cwdvjF734AcgJtT5liRczXHBgpjHVADlnSI/zLzh
3KjQP3cGjbWwAbnmbKl99+pY9oMIpEbOjirqaog0+Xg84qoI7b1JywqVWKCx+JJk
JQT8bZfSj5s4/iQXuFsZ9HnpgJ4HnQfst/kQDEerGHjpIlEqua5aexx9ZlbQaA72
eIynER7O8VWIdkiedcMIaLzlLR6ju20UMmKzSxf+IhabR+nPeihV7ANdod+kdWNj
C7I/xYVqcqBNe/oQtdFC4WXFD7afMaLKJ8iN5GZ5ccb8dxbMJEFSIu2yreZ+WFux
QeJZmdA8MIjLE+k3WcNSsFteO6+OW4r7fgP5P9wkTvnLhI0mhWDvyMEbj5U6/hIO
+GGDBohN8kDRZkrokYWkXJ0tPlJdq/xw2DqeAhOM3MnZLRhQh0ZbYE8W30IjtHvo
IEYFaRVKwUzC16BKr1MYXHnPbpXKkZgQG60RtnDVhxlPzKySlsIK5YvykuMBQyXy
yTLukuyhrp2QdUe/QaID8FuWbtaL67olSmhUs4TooHA9W020vbosYU9u21L41Ril
Nw39/kCSRUdy/pE6GiziLcXWtQlkQaZGfsp+DVyk/4QK6amH3t6Pq1g5WmOWZt1V
JrPoRc1Z/mE3NtiCPugDwx2yXlf0d6jk0dnBYICH/Ua0INOzu96xM6izeFd5G4VG
xm0jazhTqNOq1LdfSLNXMrLLrEUXESQQVM16/hf3RCEWzTsfuH1top3+0M/UntRF
npFwjT0MbdSasiRVWjL5lpsM4am9gRd4bqFDUk7t8Z+/gBRXCk2E4XUlw4YNw7lC
CPOjfVJKkQ0JKdm5Vg1FdsUPv6MPp8plUwurZdGmLuk0AuHTvG14Ys08YDkOY/ey
rJzXcFlLU3r16/1FTQfVAfUFnLDPMeSWJUr2W5d8XMYCB31Po1Nk7GI0nWkGwe5D
0bbyGKuTAQyaUal6WewOyg2xkAa+Y5seIZX7RtR4M15dIZ/XAkwGqfmtGlWHg/bE
kUYmf96BpV43si3j+0mvOCGzdvZvlvu3Ojcf20MlPtUyWIsN3yGmnyM1MAQwGoTN
HqGS7rjvBBt2TVNE6yTlRbSKLuErjQtklHnNb7aV3fYLqIV6snj0S5ZxkL3QQLWi
JFNd02joUi+PXC6jtbfr1vI/wVPHIXMk+B0q9lB6P3FfV42q4PGGw4/oPIMi06gf
YyPBdmw1t6JaW5IMWjT0hYZ4k5UB+mKoVvVcHdtG9Cjxi34xucMtu4MQM820s5Cj
oiTWLkxFFL7v8ES/PqG/wZ9J7SmlT2f8VywzqHtyWAH4GsJduRuijgsqyGRlBAnu
MFdQtb1JPTDurdksb8VW2SiPjdFtLaSyP6K4tmiW3rrwxuXIFGw0Ij6rm7C6T12W
91MSo0CnNTl8v9gdH3syM9uBT3GMZ6uvCsMERIPL9gnEImC0WVFb4G5f8hX+oWuJ
+f/q+vRQ+yfRDKadaHUi5ivo5HFp41hoLiR7K2feoAFnbcp+yDChSgvZwDtvpVsR
hAhpBITmON+4dy8kJ6zpLWDuqFhA9ofk2Uo0LuMmIU8u+ccxZVdPI2PkU9vNDxOk
ChSRLKdxVmOc7iBNt/5HBPbWkN8bsWaYmCREobZEX6pdeC0vJ5at8cwaXTrINYd8
4yD2x6n+Q6est7LNAEsMXXvqE9K0k8x4UYX8IvD1Ni9qWzYJ7cGhNWN+8Pw/oMvs
ebBAf8Be/7SQQCV8aO+GGHpY3O3Xu++tZGiR+6O0fkWLk2ffwV2uosQc2E8pgwDT
y/nRyZhAYCQfGevbGLOqhDdIc16erAb0PrPXWuXzzIRiSQUGKh3kFcAef+tM3hlZ
duAYGoAXdjq5dx8RQDPFYD3LIHiI7Zo+ABXQ8JFYParG/Cs1/RiFZ+EZ0a59cWkk
sudfz2jBOvTNI7gh3BtbTEcgJpz5nqkARiXrI2wDGxEeitsV3twlWmK3PUc8b8TZ
SRcUZ+tLmnPDgeY+IovKr7Ycjxwd/tToeQ+HoclCkL7EvgvK5HRBQaKGEM110bfK
8cw49A9U/T7w+C47xv3kJP+VkFNx13Q/t9mUOT6NvizcTSch099Yx9piNb0tzGcy
oKGYhFIj3C24qZHNQtyY+hsMHIQ9Cg6/zkUkv8uiTLE+R5R/MuIIk1cvcaJ+asjf
fvBsnTQuawGJx0iszhC9seY3fzU/3+58gg1oEupFt8I9t3M/PhsqiUeQiNYwhP1X
fXXKzaYrN/WZ/OGoSY2ay8Kv0iHmvSe/GZnQQuJAKJ6HlnYX6FONQy1qb+YdMQTJ
hXR2BYeCPUovA3uRM7fUz6bfPZ1ezX3rjeU2oYnQOLfIgAKkrgigjQeP+Gx1Lfrm
lPvErogZBQ4dp1l7A8CIuxPhfFBqNdDJ5hagfUMywwK3zUgXovrhjQ7cdjn22eEx
mlrRstzhDjSpOuCLSgrnT9rHLVtkLfjMY2TWiL1LqhaMt48PeNVJO9a6oFxAYdfx
OYjkRb9DDnhHxOCDul7pffnJ75LrDBzQehEii9eRECedx1vIaelCn7J/uGd49mkb
Wv8WKA8grf/ypAPI+gzw3D3YSlSo2oSRK+1s/FdrfFhDUWYBjvf/aDNU869RtM58
V9oqDwAIfruZx+As63pTDTA5iy0OpnxdvHF++s4CpxSIZ9K0w/tsBhk+V4/7CZ9b
ShzJK3ddoIUb8bVdyrMxzhp3Zw6iSdP+liiKZkkvNQCMaLwV6hP2zHRdRKTnchwc
71T2nm8vhlUAKZ4Pj+YeF/2/s/3piJMcPJoAmtY7sOONNDlQt4z4xDF1AZvCnWjO
ogEqlB42A9MQ2HwH5RwY3GbXLNnqeYrEcM82Q3FPKa512x+keZXXCi8aY438b7Uc
i0v1XCXqV1sTbbtgQbb9F+QHNBpTrz14ML/72EJBk+QatDA3kJaTdYt5v9PHHkl0
EMlMedOz5t4s2IbDBWugO3ChB1diq3df4MuM656DjwYelpssYol3HfyUOsrkoemi
EEKWILehYSPe+wyzCRB1nJPlGPOyqRpUtBfaffZ8IiQJp2npPsP0a/ZLQ5YtwLXK
6v8Dgwmnnx+RqmlZHhQhn5UtUwdrQQnd226kfqDxtbtItSLQax86JXQGN14Mimjp
UzWo9VYuQPhYmjVHHNR5c0AbJ5lk6EGY0zmzMoW+WL5BXzjoTSoBF+EEAphHi6I3
S0/EcKTGED3swGwTKOOP8Cyj99Ejypwv2V14Ml9Qa7u9igQS0zb0fE5RoCzZlGat
fB264Jn7jseWmjMG5F0AtUVxgO6i61NWuz5fkj5bf68IImt3RMCxwyzWwTEv09Sk
xYGoWUZQc7fGDKifMkfb6TJzLLM3PSjxwKIsamnxuNdOgpVshzor+YzP0+1yfSye
lstvgFJ5SVP1MM/mY6BM+ZVJK5TYd0+oB2w95QE20V+uopxC+vzINICAB3H6xJoU
jz2ZFiLRZvYvQGkVJBO8OZ2GZXYX+SHbFhYxvSkG9VgpLkH9NzDO/n8jxTotmk5a
vFtk9Q9ng8h5hOs0VLE1J0elm6KnWwT7mL5ejDZTivKVNKwoXpO63Rg8S4uZo++a
tzNi63/YdoyQYTE2gPSJtjEWCFiZhgCLXJAmTNZOiXfYgF+5DP4VRahyfRAx2NP8
krOCLip2CilfR0LymxPGLy52M8UCO2KHZh7F4bhj0ld+JDOb/NXWO5ISGryoG5Yd
SSLS7BMVla8qFI6+z5aVZdC6XqRx6z4vIanwkoxVLJuyDHMGLkOVV+uN70e3p2KV
AFzUzMoHqxa8a93HOVHUSfH/AYhNjrHPNaUe/7JWG5gPQSK+wc1Qzly0V9hnpzGr
g5sAw4OLIlQOD0KfBr2ZdVaGKfBn3+oC+0j0Q42gJ0EycOG/njVLUYH0Oh+7VWhb
RoU4F3Z0Ynm0S85VLLT4FCv34R+RYhSJmKbcGplhe1Q0bC8+HIgL+FxSF8HFGQTT
u5uXOcCKswFCsdYvxda4QROjhRjOzwc5ZLx6p8oboiI4nrbHd44w4nxKwJ/tmeTz
IPnpeTWJi9BzMqjpa5mxiqud/ex0lQK7pTPXUQ4mJHYJWR7Qc//7aWZh4AiOBitC
/mnhlx8kiOrihEu/iTlqN5VygKmYzVdN3nlT3Ajk54hruCYKKP0CXNM2MbL7HNGd
/pWeBdxM9boBIVElXuwX9Su19i5XQHBrUPcE+juRH2iOoafHj9CFi+8nqeRE8vH4
tWQw4znBJUiBMWd23RncbkEFBlrtI86PFz3dteWXkmVizXI+uDVtNBxnTSlIm9qE
fcaSkj6M25KSaZH3f0ESi4bEH5sZ8cd3erxh0CU2hRoYu6AlZvHlCrc1+EovLRd1
DiGi6bKBkcYC33LwrJySSnpQlXI7HE0k+ENcAc7QJfhPAYudeCl7MrkyLczz0Z6Z
xtUDnsTB2TXtmzeU5TQvHBNFl/zHiV9884wg932DWrYLWAaLX3xxNp4UNzt+AVxI
9rPdMHZWh0Ax5bF7bL44L8nrf/VzK3t3fhpTqqcdkLbXqZJlmzth/apfPYtWDSSd
GK7pvPbscDQ5+C+a5ZLs9cFga3HHWI6fB4v8W25T4/lnxsBcmHdvbMGFvcA9oWqA
cnexVUH8vkbEp0co1mObetf5D6MF7lLIx7Kn7B5SbnbTN+w0/lTJLyoUpGMDIOgW
kSBOgGBvVS9Ei+Frd+XK5nf45HszLYqg9kqfAoyJvL72W6ZuHCpcsPfDIeFj0zPz
qV1UE7WjVRzVpFSguD/z2xsfxUZcp6r6mV0i4E2WluqHJepZlVauiZd1/3GqaRri
GA0JpS/oZtRAQyvnA6EamBTlI3Tpi0FXw3/sgTc7NqXcNy9UnjzAqlKH5bDFSrkn
LVNbTnYbFzqTCpY8NOmX1ZfGQ3ACYw3LDlFDR4AVVhpHvx/SHvoJCOnZNfy/naJl
bRRE//Uc4Sd08xFGkzJ44YyMV5TmBJPGm0kDgKcKCOTQKA3hXEQ9QIyMm6lkWdZ/
7yN6K2uMPlhLVaz7aB8utmkWTs0L8hyikKAi+DdcTo33YPpLPeAPmC26yhMmbwFM
bFeN6lPGbeLYXS26JFCndmW6RGSEbrQA60mkCWVMhQr4HwMzJqID3hZv3kAwOttg
p9SIpJO4rcuXcyy19Ox6DBY6uDisrvEd/akp8T3r6GmlsHY1sFPDNGcSTLYOULZQ
svgUsNqB3fWx4+Dihu+yp+U2MDn0utPGaX3JcfvCWuBTA1pF0yGeGlCs5s4ZEQLk
cSZMIrTWNlpMrf3dqphv7cc+ck10v6MgxaDcPf3N5Q/rxJViuzpHeTl0qILMXdmp
0QXVoYhEjfKRWG2Z/pZL4NIoF6m5DRotRNPEHt4JIKJ+yl19dQmCcECWr5gwtzrP
1wskdlicemn08JOXcEypDuhKLHUN30WIeJ2kojwf8f50h1fHuZyvveQS9RRJys6b
deTctnUpET5UFqHnh53nHdUmLlxYyDWkAE8svYhoVTipFOms/c8o8592qXbPdv+7
YQk2w4fxdxBy3Ndk3bkctPPxfGLP45mglU6tX+6k7zm4XPL4NeQzYVmPneTjtMnM
Z6Nk1pTnAPAxmxGaxjQSkwC5cdWKO2qQySoen6mJY/2qTu1qT46yWxfo1AWnP4Gn
guDx0JlqQxJaio/1ftzr3VlgniDh5bMCZFHT1RCc/YKwKkhmQnlbnZewAq86ORB9
dP6IQXZbMqHkPY0HcPN1T1JsvjlaxTJcCdNwAdiio3N8pOzOEJ5A4SUh6ejPtWqK
NkJRZnTJzABNu4tYtLR6Ex5LFpCvqNNnYOgbKLptDSc6B4VbG/2sVRwxmUL9B+I7
T6e962YjxpxyceC8XWR6UE2bPopfmSG74C0N8KjW2D+mBTD3QOT9dcBculJtkWmw
7M0enUMjsp+cN/dgu/dROIqKw+0hkK7lliI69e9MAXVfn73QMziGGscKZpA0S64G
mi7Krqv32bUJ/0/a+XBQsrE5Wwr4HRcY2KxENU2wzknZytsAtEUfDXNLqBvTZleQ
C/GZ3U1wBpgdfGuVQWRBn1rXzVg4L2iUAQ3DAXLetheLpvnaHXNL3+p3y1L7GD/H
H8Ym/LbdH2iXLJewI2J3VQQRwlddMebPqMaa6hQ+ZHtBIvcj2m5zjIQAuMWoB3Wz
4XmqVCXhnXAjlUIphr0NTstPMS59WTmkt1jgjyXChz4E684n1oH54It+Wts4sOK8
NTpGIMt3t06BJBSFlvRG6g6V2mmbHFS9xfUgZGl007ta6j67PUcNPOD/c3/0yY8I
JOQqib03OkaDisDSmds5n1F3GynMeLCrJwtg/Mzo3i4xBuqDq2/h2hc2TpNLYtdX
6CkSSa8hFI183hjQRmYvH8huCjyY3HrI5s7IHsHAseiFAsOcs/s8pr869k4lOMil
vsJlBF6pmzACQdfmoAEGJ7WwrCMFit9BGo9JEI1kQY4gBmbOSpXhNDijsIm4942u
bUu+SEXS09qs9VTio5cyr1WUlm1adfQGT3J8xvpZL43oI26m372Ev59/3p95bUCC
bl1M3jFwMliu7WGI4m54PsHVD7KADft4jmAODbS2vbrRckjoeqz6utgn4mUVDK00
WoZ31nyZHoXaed5VVb4M5gFunTdX+6qaUvEK40jMsYi3sI7M3iBPPqtg6L/y/UoC
4ZfCfHaEYABkqNumLci5oYSbaREHRbHo452aF3Ga5SPpDmo1XQEvIfOSM9DyNzj7
nZaDU1WlPjb9cWlJVf99v0ju661GMvSU9Y5pCJwruVDFpzO45aINoaHvWVnQR5zt
rNKHZEjpVKZEcOpLI261j9l1Cb22qZlhZls1K4ufZtJZlIF890Hlz+whQ2naIBlJ
VYG6OC3lcq/QEmviLz+JlVBlEOxwGQhV5kmifdxH3mNELAS5f1fdnazcehaIngLd
MG7faOqx5azRRB8S4n6ieSNllJyslXlI0u90EG8q+GNYl3k0JooO+WB5QmvW8JU8
3TZk2eNyduoR+Qy67uw6RXM0zDjVU2TAVcCUjM2iuE4aMG6hsb6r4XLBupUG28xi
ZbOLZNkU0usbViWe8z9Nvlt/uGNh3aYAqp+tUuKkpEeHKEuuf3pNAqJSvdSR15AE
omk6r2hA+P2U8ytTO2vOdyQhhxeh11RelLxq54eauSEVR2rDe34A16APo/+xaKw3
oVmZ0iPG5SqiOazbEBq81yabkwKlWoQHfwe2QNVkFKH7JP2rS6j9wA/dfrlnhS+x
VKLgVu4f1SQ6Jt/X+F0IOdKomnpqQcWWvv55r6Kfiwh3Tzf821FoLV/OEXeVucQw
od0a6lEAY3BlzB2Qw2tNN1VvdqRJQPcftItkWreHy9EOK3rUxEdzzwK1pHvStFLA
KCNC2F/g3VV5V+UecU3zt34nJHF+VL1A+/2U0lUKiILAuazqtisdRSRv7bL5fugH
zxrzaHA+Pk8rRBZsYUaOhO0aMuZJka5h0n6IrRHinia0L+9Stsg77aIlwrSkz29c
v8Uklj8Ss7SdhMqgttPVafFuruY0oU83lbHA6sxFPcvYrCJzNjOr/VVk7+lKybJE
2mD6sAEHT4EF9IaWmy9RImhFUh5ySKEVaYLI40YW/F3KD5Zpw0Im/sb13jRzxZBz
/gh0IKZYorok5a/yYvzYcWLdvUg29hKEqTpR50xaE7776ur/ByopGGlOqEn9qeWG
V6CbLDqo43Tl/0e8mpCIvejLkWshmSIbbv1hJTXxVLDi5htVCWix0rozociehE/f
U1XU5+PqBo7so5zD2xXg5snpLYeyPLxK3u+qjovG6wD+6DKCarGUxLXwzr2oPPE2
eu0SIvIJrLshrkiYNqLiuhPhVGvzQkM4ZvhK2zsCuMIlKPmBZ2vKe1gQIBJEcG7r
3q9LihWW2lnzNFgrSyxGjaCZQOlK2E2XRqZco2DaHUzmPgQDKtlf8A9y7GmviqL3
uUst9+H7cp/xi//1VTB/oYyYhD3vZQYILo91oBvgOZWcgR/N32oAu1b9ePvaEQyp
yNCunceQApeHRSUuJsYD8IY/rWKaDsUwQHBPpqZYuCn/CzoSKLoL8r/ZZB05HfEx
313IoK0oVT8DJ5qjry1dQrShG1PN2iPk0xiYDT0UkMtDCF0IR54KxSBNtPJttBG9
KtRG1Xkri92qMmepzYu+6/XF3oJzvf+XinitlXPU1VLdsCadUzDADhh5ZCXoYaib
LIThjvzOr+RLUTI2PJ99M4DGNOUy9JOUJCVYsIZ+VChTFh2q03USEnEHQufeK/Lj
UpXWS6l4XXgdWuw2+x6moU7crRxXQzBcnjuZry6Tj0e/pvdqAnH1sDY6CHBgs7lo
8/U3PF33+kl3sNbbyc1WoGcaYVM7Olb6aJ5HONhqIlpL+ILCCVGDQujZKBl5yNPC
g5cBpEyrk8pS2Ltrks7amGC7KdtLdg41Tdp3tYz2ny0skeHbAegxJ57zgxHWsoQZ
Vimbm7Dx/HAkvkxLePpNhNts18P1C31FZTQW6+3BcDJN/4+6HpsacHp4fcu28IvY
qoFuLqkmBZ/dnRp5nglZ4IXf4qzrFYwwxS06EbzkUTjlTcxIZ7+v3rDx2V7eP/i8
EEhzpZeY3biaMqA+ar6ECehGN5aSz1rFk45EiKYDdvTL56VkWfr8fNPFYafgUKaX
pqSjjVOCdMPE3hHmDG5PTJu2KPXfHgtfedq0AIPwFL8XDNeNV19pqsslFiFCE115
1U/kooqILuZx4qPxZDmhIuagZvbOeWV37igfJih222X83MLBPbRHsohfkZYvYkGB
vdtWsdb0kpF3wLfuZpmR+n6Gbhi1w9sVXd0D+jRJ0Msuefl07KlSVIw6vIujK5zw
s0juDGQb/822Qir/3VZhJtnHdEkk90NqiI8RkyradcpakpfyvTuxiqWLTm5prLPk
lS1WQcXU5cjZLyZpfEG+bYtlmORmgt6LNEdmZZb0neWGSgoiFc7Pa22W4Hh1r0So
k9ji/goZ+abYIn4KB0bqQqLgUFVUM6LOtEcoB/cbtv2VPefDmH/yy9/sSonomXLM
BfxhNgF4ka8mIxBiPr56ufNbavoP9N8eEbadw2YO6llH4Isl7gPI6bFNnQbm6EPO
bL/oC/Lb75NYpIFHPeU6EVLb9vAw4WPgwobnuO5EME0NFP1YCSyp7dpm58K3J2FW
nZVRrpCNssyqetNKZpEAHA+nMVx4D/muaJPAXpoSnGSSgJuDxVfM2ElNe08Ysqbz
zI+LzuduMXqSYYihyilD6tieCuornT2oFDGCZA59NMH7S4mhi4qGL62l/B0TV/vF
3XbO9AfBqYUj/F8LJegeWHxhaXCjFqmzYMRNCi/CdAGY7GDuV+5udrRLVQeHpvDk
RoTYxvMwhAOOPWEk07jyliKzcwzhtlLvkvvyW58wTFvB/DnSrSD5w60VvseelbuL
t/Wv5G6okhrr8G9C+6P5fW0gNzdaRacrvZuC4NcACQ7Wx5hCnm0r30WTbnBbeCig
ZuVJXQoOangGltukiFwBmt4ptM+fioBZrHIZAg39wxrjld5ocKNm5wLhoEymJYZ3
cHJMWXsCFgmZxevQKg3bmRsWM1+cz8+zJKfNBTEhxrS0/b9r+sSlEoWDGyZiKPFl
5NAWHv4S5EuMbh/CducrgszJZQhUxnTgIUmJIciTtqErfWA7vNomJndwCG9Ws8eN
Js4R6EVzIXQkIxV1F/4Im2rQ2cNbblPyC0OnHmY36qJo2reFthfwe6czW61FiZ5C
ro+VUfKKvISvd+eDiSgFeOcT5kh0eXZMNn1AjcvFT5linyyxmcX4Ax+eC2SS1i1b
xDYCym45/cg7ipuyt+EROMbAcZ/gsgi0G4OSg+qnvs9MdzcNChTT+8s2bwwo0AJ2
aHGPhJe9SWCx47UuenWkfH4BTtM2D53+uKEYUgZs9VFiFAXrRZkw6jswetEd25dw
HCEGkmqO7lF49JYuNFyeWFm/QYc10G/N5+lei2Gd3XXxwVcCN8QmNXWTaO01gEpo
XpKqVz6k65HwOCFvmB9ZnqhSQBKA+XKkutY7LkEm6qShbZFdk5+hwouwzg3xrKDr
ybJ8+oRqm/4jXtS083YqgoEdME5TfO38PxSZlm99WLOdRQW28t+cEUMaAEeCN/WH
bdgymnYk/Sv8KR756Vxkj+1a0dZoUiDSQVcAPxScEWZpCdj7/MwjjUGLnkxC37R2
LPLa2JfhpXBiEqRCZB3jTMTcoK+OIlzNr8eP7snQSPwX5CLM60C0Qba8JTicHW6k
/tMKX/rHR63eLSSgBcmP7kRnL5SxNZshGo2gIDYECDnkVc9ikjfhVHEAm2l0BCgK
hU6E81uYwVfNon5nTgk5UuRwwsgQvyTCgB9CgxI3q9W+PbZCfzGkjf0t1rTTHRsh
hEAUuG7ymsjdpg/vlIie9Nj23M2R1gfpO7rfj0qpTT8nbqkYHhAOCl63zzLXjb5h
qntp01vwu4rZjI/PHIKbebjhoUtvrTuRZkPqhdTeyuevgHu9TX+MIL1bf/lRvqcW
5xjEctyPNWsifSG8xbLt0ZDcjg+FdN1GdSyRbAeKddQD383pmErWa94QaIDZYrQU
zBGgNj81mgZ1AgqN/SDLVDE/U9xoYej8HI15V4q+zIs1c4oCxiYyu/YZBh2NUmWo
z9gJmsLVxSRChv3sFnHFqG59IV04Kq0MPWIVKSis/5dQQgQG0T3xfMfnxeb+bHmC
YG/Kwtr7Gu6Z+LbXb09CpHrCFGCCZ0p7/ZuX/ZYmIDa1MQOfaJlOv/3PN511X3Pn
2nN/qU0qTv9xqOA10ETVUez698ddfc3ZCDuNbcB3sfYUdw4RQ7r2fZ9KDLbMcjmU
oyQkyTgZJRhmpI6XPXk44FM2ZVToa34vy69dEl1+JG8nSHHb97aElU2eajbsuJTR
mMVox5i+Bw/T+jjhiGT/DSkh9d6xqvL48YoSBUwj71tm81ubelXt4YZrv19km2Du
KiqMQ4iDm/JiApJWgFcxvu8thPilhbt2yFYh54Peb6KU5fw1E3YGr0w/9r2DVRUH
eRK6zyjZ2DM7Knomn24yiQ7yUeCf9v8RdFEDXeo9ZaiSfREyoGsddcFYlWRJbal9
BFxndEVHxG0WY8WX33NKgRmSHeevhrhKTgPQqjr/NN3ov8xfbRkf7Quw5hVybZK5
yKQlDktmuBHyWWCO3Y71dQTZiJIosynCWWSmGujlU0Kny9JXgzdITEpMQr7S6D9O
BrPra89wt2+7VOkQel2cMgUmL4hWHSi5+xVZE0K2+ylGr+b0nS4h6GNRN+asA+DF
4tErr2ubb7KF7nmrrg4Kw+Sir55emuMEUBU61hIwHtkHRgOXDmb+bbey7HNmCSJD
upp2pCtm3+EhPAo/Lk2783ki7oDj1LH6BojC60cgWbw2EuJH5j23kUvuRT2nQFUO
IP/UQf3cpDQZ/laqOMUGO+F+Nwyi9q7vAosssqeVACRJ7OoAwO+uzTneUMgweQJ5
YZ5h2WLSGW6YuPIgz8mLn0X7GFw2YDGUFjItXIzME19xqo4BosFTLq3JLbQyb7wG
AYfUAjovRY24VKL9ooMm3nzRD8DEvzG8qqvgXGPeGpYm087q54pzyt0EfkVqNBUc
LO9V4zMDNWZXgrdP/fI+f9hlE5okrbNcQzCjdlO91ff8qzVXxXPZIQauhnoscwVZ
bG2YVXkpCtdVsrHw7978cTzTEb+QAtDR55SkcuNw9KpBE3KAeoSbFQUAcEi+JEs0
5O2xNGX9IsvLZobdYMprLuRFkpTwoikiJ3pLVXlAwTaqe1FkbFUCD72MGXuN0k2H
ENPEx86u+EmaEoIq68hN8AJYGQf1rOFvl+l1F/qHNtPq2OmdswwLvYZ0At6laoIM
qqM2osJzTy+A7//7VaQFWQV9O7UkMHANi2hk+q3KwfyF4BV3KLgui/iJdb9rSxvm
sqSiQ/U52CjsQd9o9iewdN1raDS+wmm2V8tifhsrrJKgeBm3jVeaeirl7oRycezN
6YetFLuvIXfZCq7DbDbPWYJSARPgcLYQwvhpfOY+qK5yR1G/zPHssw86uVpWsLE2
eyYk8XKd1FxrlgbJ7OFQnBBKzwXxYXRylnXFp4WuSR/r1YG82e+eysIwx23q4kSz
waqXM6vGtKV05974LdqRmy6Von+oo1wce93jG/Dcp8BgiSPR8SdoqBgEjd6sVdGB
exZKn0n3RdNo5NJ3L10yDjf7NBQRAl3g8GoAPwzJHj7O95C6wjfyArAE/VCXnnjj
P6AQ5vYicV/qDKrWhmVzqVa/wYGVmf9U/ZdGEpZskwwwGNt6elUJ/ukP27J5oq1V
FGYU/4VID/UOI971DIP2YfKOUwvyN9ktFIxiSlZSvsIR5h+UctC2+iGl3vzDmX3Z
3C41t7/+BbrGNYCu+1RXS0g+j5SBt1zq8w5DeETN4wi7rLUYJNGn1E4u96PYkSJd
Fzmow9VQ2UjblxDUz2EvCw6n0Kq1lT4nefFA+8931mMvrZimIwIHjAmWg1x03TQn
N+SMnEHS6AomOPIoZbiumZJKn840adBGXlj/OZTMsVdjF57sN6tVVKkg5R9r8bfm
7UHz/a50rDsHGJFpWZnnOzxvNfKHdFgkzH6KwPfmsPt4J3T6p3rZP8CZpLJSbfs8
UofyJmS64CAVRPEOEPwui5no+y/HOJ20fh8KZ9HUboQhYUfp0T5GpUSSTu3N4gd1
9yLMuSq9zWGRKhfLmqGInVYUUOHAbIbYocingbeI2NuiahiCTAeTGkDC7BtBkayB
1DhsTlNwrOWUG+RookY9POI2NeDdc63qJxi6xe/gV9ScRHek46Fb4lp4YEV3Q+1x
hvvqs2dyT1ntWymKkMMR4wCiO1uZ4syiWBYznK17Pa3aezpfaDTZagKzTunCeX6p
rIbALwdjh+rrxWH/K9eZp5Wen13CNh9MZfJSzxP4tkn1JtRe29XM0yPzzVRvILDv
4UeyMwAQjlb5dOZ3rvrOwi08CPJ9qWSDC1zJLTDi3fh7CXqaTPqEnBJ4BtKNHTzN
hlAcY9Lu0FXWJYxWYuE6m5GOkHQOEXGfhWLaPFGl7Q/1RGf/W/rgJ8V/djbODqgL
pyIFABaHlK8Vk4pfFv1+0l9rr2Rn8oHpHeDpOxUQsuRIbboY0cKLgfowLrELU9ek
MEbPu4TJST8AIDXezsAZq7YgKySOaJJkAxHtlH5PkYfd9QvwY2fGv6sbPDBxUupZ
Au5sAOrB3jc2C5h4U07zgD2iAl7iS0+4klS8QmcTVvvGETky332t0IQFqsjTTHbo
ShpJoPiKQEy318mzHflVvblrO5AIW7tPuw9EpwGT7D9VzHGgckoXT/uUoKtYv4IT
qF0NgHXsULQmXdtkQkeGZ/2aCzdgjPVZGApR+ncNEqsTxxtQ0h2Vju6WrCDfoXio
KpL1m6fRzQeFeqjILn+ewXa1UumRwolLQ70L7kPrs6cZ+dWdTRsrgSJ/yxnC34zg
xMdgQCQ5uwQdgJhxNqngppqpWi5qKzcmJIi5oSTCMbUlQMf60sqDKZm0FrIC+hrX
iG+HX3uEbcNajhqz3o4GCyA9gEZc5D89vsb0ksJWimUlFn7CO1tNAQWzN2CoBdwZ
aVtCQfPMQJby5+ss+12989gb1s+FHiwDWmRrRJyKASKKZOXv4ig3q90cWrmLKfnB
jTaV9U5mlJ5rHZ544utUvBHXcVz2uF9tj/0MVd0JpWLeD5Jl/i9nIqqez7hlrXCZ
iV/Ueo8M+RqtU9h8xpOMVyz82IZUXTgrxGGzKqC+N//0bdcD5PYxdJmuxvXLVjHf
m97svHR+OTTs7lCls+GR/IYIg0VJeKJvDTpDzTYg+iQYXw98joiFo/pGe30RoGQ0
SNQrDbA0y4IPRaABZO2cvfD49P5aZFZVhcVmFXTSBYum0ekmqDwSaOXfa6rf9LLi
A2ODQ2rOYpwgzq8yYDBj0/2Anj1G/yvqUQogX3OiGVZNUzi/USxTPZW6EYMleyDh
/Fu3KOGKyb3nOLx4Uf6yFUmAsHTeBMuxH+wFIv3EdhIjP96meIzcUWgX+OotgnT5
ZfMiSxzv/ogtQCne6aMgr4ZzD1FAInjf6UV4YaBai++CCC5/VGkjWZ/lR4bSE64L
RivgnbRpCZTDQfH5o/5utJ+RlkjwZSM4mBCzjfjW8D6e4DX1v74Ms0kBXAb6ByWl
DhxgYsdP0Pyr9zUJetLjOST6bhIt1o7RTClr+78+Ym9QQ05diODbhcCPfAMWU4fz
XRMjgAzqrki75nsUud3o1oARE94ExlWB61ZtcSYTzmeK39nMTAuq/eWEmZv2YvEP
oMRDpH83SDlx/o40rF9C+VLjV5Q7v573xGheejARS5h7F83fsuRQtrWj9GBZBpU8
svlIkEIvyT6Zdxehq639Mkbo65Zv/bCMnZH1BDV/k8RPxYpRv2Y7YXXCiHUhqoRI
uns3GS+vTcwhBq2r2MHRp3p9Sf3YdmP/StWSyB5g4Kifa1m2dsljP+hB7aVr0Mcg
FXiVxBegku9f8jMty6Sy2cMqwJ0RzxvXlRvnsHyXb8SHaAkeNOac/Nsjm+cyHf2b
GDH99AruLbKFU+QZI+NhIaixs/0xw1Or0olisRDy9LKexzeXyxhaYaRaMFx71tui
/AQq8a1YIKB7//EOypht80hEevoZ8wMs5RTGLdhWdtDpUArvgOGZFEEWdWr2S5xa
Qe7S5mbTjDv7p12LU/z8FKVjviBF8rBAqQqpEqK3jc6E72dNW8LoF2D2xASaLLfk
AJtXWEb0TgFvTCcNJ6EEYaf+fVbW9mYTXyoNxjtg0FJQMew2lp7ca56uo88yzy0T
c1PI3OPl8lffboJwJPmV6Z0zLlVCAPVEKVtRMRqPy8YvX1BX6VFVIqWzIyNZrwzl
6cD8uZLlLz/EaDpHDzctQ9yZiwoI1YYWXUQYeSVp6VVRo5nQeAfuy4Jrpdtqdjof
b2F3zUoJZ5Ox0lwc5vtDe8F7On2ZOMdUFtQhImHH9pWPC229J0v55WOyiullwZic
1IEFBc0DCRbZsohbkfBk3BDR+U2nE6RLl1TN2IYXTtisFbGdd74var1n0a09sbBh
lLs4FaxsCrqIRPmaydWGrmCMXsWGAbVkOrK0tJ2lqjVnwxohez25MhhSMjQ1MLq8
cbFT8DNbljs/p9ed67p505UR9U0nd5NJgnvdi2YtWOBpoRaPINsXuoaGWD1ZgRJg
KNgKPZ/nX+PVHFxS7ojb5/7W1Z8LZH8uF0n4Cd6mY0tbhzRaRrsHgqeQukOoCLvR
uL2eBCt+FmTuXFMR1IJIh2cRO60fO71cenQuGaHK0A0Di59c5HCQDGdWahNwFrME
PeUH5gTKkGF8uUMmotiUAOAdtiHHPmhvR2f6FWedfQhQ8UdV0U2RZD8mfU1TLM2X
lWRiVNsjQKJEgVv4TQGtHVDfEE7vi4NFi3uTUaB3InxF9gEyaBwzNH36GzPze2lM
z1Csxiq2KMLodp2zbvhzM8cp5Pw88mSJaxzsmSsItI/o+QpGxVpx7XSQQQDa3LiV
hMJt9GdZ5OYcB98UWALRG4tUvcKMSo3tgNihddUfPb0YKDLuyj2uafe61TNK642s
fHneeJu1Dr/iUcSNm9+h/wbDPJoz/0WyePZ7NuFLPygB3l1tAfP8EdPKNEIzD89m
9GB9lKd9x/gseII9vSSXDohZV7QeP42u6ZWzZ4eHf7snVbkzg8wj3h322KocPkOa
j1fh7Gb1UKbPZ0tNm1HT6K2nBalBrhF/9VLZzhF/fDwZFScnUrrknpeAAMgVwQM7
oZSpng+T+czMYzF1spWlsR8NSAcFk+vwVchpGZhQ7OrofXz+EsRL2sQEqZ1MQrFu
4jLNjW7dHAtgphvuRe0xNDArPoGJWraatA8kMEd4bsr1DwMfvwa+ifxZM3ZWYfKR
Gvq2S4+jyqdcd5HdRj2ewz6htaERYmYzoTAwhL7EVy9EDS6BCMZvxB7heJpBnu9t
zvM9Mch3vx00NpNbCajnOxcjJz9SNTcjDHKQNtl5cadeqVUi8FlpZkVwuN86sYXD
NkxH0qPVclXjx6ha2RyzvM11HvJWFLmRP0wZk4ieZ1dGolhmxTthY6O7P/A17psY
XeKeyhEE4sutGHPsdFZ7bWW7q+4c8uvx9YOPdzbEiSB3QwuxPSGEgGck0ip9VPFW
zrMLT5lhkKSWviO6BCPhRE0o4QptR+zrhQlI3T+8Jq1Ey1vijp8NsD4JK5fQDMLG
lr7QpTf/tJYUKjMS5DBZ08EBRRegzJIUCWj5yM8dylZ+Jx1UxH612ZU43/dxObCZ
ReINE+Km1cjhOUiYp5xubDyUJ7TxY9OwzRCMhaV+rjLHBy5zmBXBBCpUygb8DKo6
BAKbk41AQ5ZrWKu8jVn/cf9w2Iu1I0c0jBvu93ljEqc0NVvCWfckJeeFnayP3MLI
OMM5YRqx64SBfNBfgqAAUga45s70OiYa+JUViLsrBqNrVBR8uwqXPcry5xclSFFW
jxYIO4ZU5Sx0lds/nTIL5DVM6bZsrIipwKjdhWP/efBoEKcr6lZC9dwIfpDbKtZC
HP0bTnlXlhim4k4ICrmweihRX2XKGrm6hmp9gts1ol9USlX58rR40RVQRVodKqUd
XkwVI54f2YwpHxIVlRVRMK/eUI+TOuqPK4nX7xqSpeNWfWXl8kQEkNEZy79v6b3o
he30aM/8qFLtO5KHL2de+I3bwVYyFJW6YEO8tf3OlMccdJY+wCwnzWTAxD3atnPK
Y49COjd5nQWQ/Dc05KqvcWQhDHBmX5ViqF/tcB7BLPqlI6Vd2WHJPCj6+txcxejO
fEEN7jXxyNhy47ZE4GS6YUKnLOPN83dledsQmxm4y6DYXmLRw7bP9F2otGFXB05S
wWGZy9UVAYXdc1h3hYHzJxYZpwNRgzjC117fVpnGP2jxYfswobV7qZQdL1OlUY7/
azR1Der5FoRfnA1NMOkX/nFZKRWqM5U5GNBwvv5d3VFM5cf3360B1dItgkNSb7EN
JCspvUI7toHhRe9l0Gui1xmE1X9ISxYX4lRTXZ2+NKE5aLxrOTQsJR9uSxnxMXDP
XUFVcw2pr5AePYEWD2IIa5f+Vwg6oqyl0ybZCQmhhZOR4I4f6zbJiUwjsln/TuQf
VkVkarFtIHyWBc1FeTOl5xGf0Al/FWADrbU70oc+HDWPOt45kxiOxdAy5ZFN5AWh
9+Ns0wr1/GUP2pulzNjT8LrEHyTyetNjoXadwwgnVu+TVCbHnmOonOHOOSWIcfEQ
8FAyifG7xKLg4CNIsbGSI5eiXqmUwnW2q7CwjbmTHodxbm1EvQrAVL8a0at6DHZc
bcV6SjVAUT2cV9/0eb/NRVavHXIkD4WEyxHePrB6NKXbsUEyxHOqmWhKLRQKQWT/
pMR5F5g77AnNsXtTzbBz8CpZ0BK7HRlHcGtb1aGnumR4JVYo1bFlwtN7BuCpzN8W
qUV7eCXjoYoLpyO1yyaYyD6ank1rP1W92afMA/5UTww00UT4YQ+wWsh5qPjStk2G
CmTI9Sw7rQF13/2chfXtg7Z48eNkyScwvk3ElEX7bCdhzSE6Q1fmLoQIh3xFgDNn
Qim7c3DF/IPGS2v+fCjKnlihUiW4fBd7Tas0N9eG/DwmfsL7iGRjMxRX/bdSkxOm
psWw3gXrw2ODAZt4705AtyhsbwoJQJQyxPDdoGUoCYCuIAq6BF8lX2CAC0IBYOTK
gl6/DI/Bfe0FnruN2IfHQbD5Qp/9cP5qHZ4xyoX40TtVv+pVtCBK65ZCKQtKQZ+F
Hl7M6gin47o14xYV8HAhraxGIe0XFiDt3QTd/nJuIZOPnu5x2vBA2JlGfDLaCdBA
m3fJxyiqcI7b5VClvXwR2EBbzxBRCSUk+7+iXsNpqMIUpJH0z8zLmN9FiBC235WI
4/EZteWIU0LfrlhVKQt+ZbCPxupZKwuP/o7u8MCnfazCyqc5ckqGBq4HBW8gYIBR
2z7QrGHyilhO8Aooumm4+pZQ7YdHzJtwlZnS4GcakggBmRo6cnEOLM1zCckOmt2L
o+sO1NTMi3AxMtSRku40+MpBH82AtuN2AEoQ2k5TextUWr6R/Y2NUzqhfwcWMja/
ChVpH//kx0/r/0KXIM/eBaUxsKihGHlg29Y1O6O2ANpY6FkccFSNuK6Bk5mvLWQR
kdPVk6U1wqcpzf4C2pTeTrVSry3ja0XBe05RUD7c8pJrcMKsaRMwEv/eFDfdm63N
Ag+ilHL/u6q5+xAf/oK3R3XkjgJ3u8i48ck8kw9TwDVhwY/ehsk+F9jzE4nJGs2K
YcWtzVjW4erSKPxZL3QuRWmRLzfvMftwVjhI6pJfgeHGhoUI6jOhD8V4lpTddWbf
S6/5nRO8m31RnDWSzMqouA2ofV7Dds2rmBkVVDF2WKeEAXEsv4eCpA+mSaLo5+6R
9i6oWLONA1Ejsqm+aWMxIxNt5zQdUfsXcfWR9Pjm8F3m08bt5kLdu84kaYH9K38s
lzOexCaFyw0BXEHOaJcEsIQ/fvPAE8EW1gon743JuGKmkxsN+UK+BzJdvGTek74J
DZqm5mLzDMl0R9t6CX7huDs5IROIhugH8MfnrMq+MbY5IFvSlUW8/Zci4UkxSb0f
6sx47/f0y33mpAeDR9kpJMkFUMggT4oIo7XhBRHNPgUs1J/fK2qYlh03EH2YGQLu
Pe8T3/bG1r3A5/Suc/6CkeJsg+ibv9U1jpYQw4fXRF3Q6u09UHPFkxi1vnmz2U2B
lYtNceWbfu4+zLCDiG6yK1bCedZcuYN3P2136ZnUbgNodSYv7cp1lvAYSNpAxZyf
d7VntMZ4y2L55fQDhdAa3rmqMAO51NPe1YASPBN5Z3eM6mtEyDy2n45BHYukEdIm
WwSFiCzpM9bJ3eFDxbkC7jHNG82Cmk5NfdLfe0pvR+37dvWIfrtTQ1u6ckA7sHHX
LMbLTKKMRZHI68o/MeWqErt9A3rhkH4hfb+9VgMhgtQVEw2VdHop6RMkLSN7swoj
omAaU5bOL8zPB365VS1XKIKmRK1sYAK3J2kczVwUVQp4DQtFj0PctG30J+EimRxO
AVTyZCyjlF0P6Qn5rugLV4QCnokL2gd5/RIdpx/b6aERyn4xudqVjmMnK0A+xyYz
URHlvIsBDN3I6DOsdePyO19QYQMWOnDRN0FgKiuSEQb0gk0BabnjP/ggBm/g+jIu
leeMawNqxZV8cE8X+bDG/nf0SUUqMv0zlCVL55XMQianCQqf7XyGSf+28ACLlT1J
inehsQelYQ+5xoXeJSiA/G+bZRGk8Dpog+i+0FW1AXl9rg3FnLBp440oINBH+xc6
SXbSZoWDxP0sPiVcvvMoJZOjmizUYXP/CtnM8Knt7yr4HUB0icVHdQM8l8mFhT8v
TkYZzs5GLXcEp7DFqsXYn02e+fLRtbmAwbSDdnV6mD5xTxhYw0yvFljSs1qGSC3d
OYxio2ZC5v6clWX0HutCEFdqm2aJxy8IC/8lY+qyVEP1/Cbq0TNTxBGGJdGEhfUq
epOMZna7MH8w7Tvr3DPdyQQ33FKEHfVedd4gD4HgLbj910Jw9wXb8A7m8BMNIRMe
Ap9ZUMsyKdSRxI1YUub/pAAgjIgyX7T8C6gv8raUFKRib7olUvdKxBwo4FAfJENo
AUBN1ZEd7HCD8Ni3TtYN3Zy34/uG1qlFYl142AnKuFDsZP3SDNinuVkscWY4xsbx
H/m/y9fOa7Z21A5tJ+zNZEZwhnUmlcg/PCl+IUN4K29CMyoEQYVD2kqvZ9Sz64+v
8grTvCVltsShtZo0OMK0v8V8aSZ3RanPx4njtlhmAhxrnxAPOnMdFue19glpdcji
1cUfUvyZhrtp5tqMtiRXbYQNJeDZNWk5lnC4SUl2VoN4M/Qz6Y6NRlctxqtRioNN
oYTxRdo7XxqIrgiHs/v09mSlzJ4A68K9FCf8IlBkWFij703yw+FZg+IfHeX/2x56
L5gawZPTKArRlGwJaw5RVpskMh3w0DJuWXOdLYzv3iobVbLhho96XMuBEYtkAFA8
5d7tst8k8VWGJqbvNtwd856IPDWUx2GPj9uc+FmgqDHCmekwEr+b9O8DH4vgxRQL
BUthA0AZ3dIq+tF+xyGba2l/Nyojk/T0ujVc6tqHvsEtAmTzyZJyaxZq+Wsj7ZTg
YKmHAFkM/xJYnXTRrtc6Om0iV/cZK9PzuNlf4DGajcR+rnYdVKhK4E53LY0Y9iPf
X8InfmXg1bz+OioBuspNnufoqbt7Jc4hj+2aiMdttiavBs+a6iRm2EgJl/cds9sc
GrGnWcWVPG9skLBUi612cf+EpI5IftO1qkI2ClIHq7xDKNWv9Q3VhcRMqXLWjikS
2mGzgJRpnVDCU3UnDIQC5XaE99m7HxHfzl+hQO0opIOHi7QcutrmPDYa7LJZzzkz
SM8sej4HSuuVxyoIB9/x1jiorNK8LeeR/KPjG+mBZ57mrpDPsVK0bxYl96TL4v2i
6NcD5RUzsyvi6NQu505zEc770t8f8/AU3qkCdbl6SjL7v3PZNNqwk6HumbPW/nop
vHlFVeIJPAyn0mMrrUqGmWY8J9J0YgNZ/XiXcQ3O7N5RkqPSH71T8DBvlSNKdO3k
Rua7/AsIrYIIuxUYnb2UfLX7fsaKPhJw6wd0kyHO/MO7jyMyfZmL1AA390hAfPJY
3jVZhu9TbvUJZeHNfcz3Vfze3B72M5cPEEiKrKWgVqIhENSF9nwZE6yBjYb3UOEj
IXrQCeYaEto2nnSM57aJ5MApzBuTPVUQd6czCD0X2GArUezATL0LGdR3v1sE8HXn
YngJLGrJQreTznE1VSSKyy+dL3vBlrjAgD6D4pYneMFC6CBhXlsaUTLkvpPJVPgt
MYl5nt4sQmw2g2v4z/r8baP+Bm9liESIQxK7pFdzwG1mZUoZjaBKKa1kd2fbvOnW
VV6rC71wL1JuoYeJ7wxDYT0VUap3GQQNl4t/d6r//OYpFdiZG14hddUB7frxlS4T
skkdmzQN5fy34DQNHu/V1KiIV62fYn0By71Djteca8U7QR1g4TAibNbw+dHj9A0j
9FeNQBZWK56A4FWsZbSkMTqyICWGrWoglyGLggSABr1CwCSGGt33pckC9nvXmJio
cCAbIqryw3iZkOtNY611o55gtT8f47BSFZvi+xTjsu7E99MLsmFo+jEjyUavvLSS
ZRnLhpC8vusEUjBGQVkdQgt06BI5WoadtAly3HB+omDBh5PSn3zHQhaGA708bl1r
XQVkUZE1r/1wSqcLM0IKottrhI3VZ+h5hGr8YrzS6Wo7wiZyuvU7NEr5ZVUkwSeM
RXVuTPPX0rhcYTbUip0iLYk+8clzWgb62MTbqKK1y7d9Zk9LQF2TxGFuDZPwrGqB
yzJL/a/5EThQ3KspiftSM0zAqhFBXvClSL3eGkrOLxaTXbVCqQAPvii97Q82tsLk
IZUH2CnqvHki8vDbmaSfO1QLYUberLh1CxZYX6qp4klFhBO83wUwFmARZ3ZNfzc/
UWn89W2H8ifEvsQnFVU4izklsSPEoisPJPbxWVjoYj7dLu0wW+pc4nvlru4eRxG7
EOzRk3rOyKBeapMEDRq/ocBiElVa/bhbrXZ8benCAynrf1lIm10chE/gRMEFmOuM
c9dROlOv6uRJDJAzBdPFTEod4j3kdG0owgtmOURwbmbuqPkyCmnx9JTJRtvtnAjJ
Fk+She3je5KwlUazlj9vUB+5zQ2f5r+qIk2X0XAzcMpIP2N9c0bv1qx8r8jkxfRs
/l92WYNzKDHG8HjrTtn33mUlIMFbTMxt8cfVYr+Z0CGvnSGdgNjUZlHXKxgBkR8c
cj7oE3/xdh+Ls2SWLkunnN8QlRA7nmH0Tx5gEJan8Gpw0ZZREfKOI2j2f5iGwnSs
APeq+kgSangivZjEpAjmXDbL/QVVyayook15VOmkxau2IVhe8hq1xr+zpf7AC3l8
4SR2GyXNhquhAN381D5AfkUm3WmxAilgtB7KMDqIIhvm2ViB1oPvIb0fJ/Fi7rxw
oXpQC67x1uWageOBJ/UU86MxwjDmWaigf0K32pdMTp6ygAHw+giU7R9+z7b1xU2W
s9RnI4NukdYbA0SGrkrc2E8So7hs6Oq/UOV3jISutLGv9TgdYktffeDXXD5SCLlW
u718ViPkNLz5cAQqFMIXu2rFkx8T7xMKEU8mHXOOZkKCDWY9gnsEzGKcRga+vzp6
60Lakm43S8UXG/QGspgxW9aeDDVb5WuZnRxNA7mcWNCMReK5VIoc+siIdjr83alA
/NSiDM1dTcv5tpi7A50uNV2saHnZMjMTyVU44O6Jwt8uJAeRPaRWSlsU7QrEyAXr
SKLKLS2/SXaz1lftP560sRzUjam0KzpZlwtDvP0ELk3dTHQbm7+/qDTEvuQYGjSa
YWRH3+ex7goVm/4YDGsSJ240atv5wjl64vg5wia9kPXBWWzShBGdDlIMMFNtvawv
E/6m5ko3cZCJfE8luA9BnEQSFGIw8bAe+Ia8HwoqXul5BvELYFV95BEb96QNODbQ
kldC1drxpep06o4Z99nWlN7yHvMWvfjnaY9tn7FSV41JigKt9puDxVFvYnsf8dwQ
831UsskUzCTh6fEALutbOyioyaiO6KTwRpMDyteE1ZlYXlIGXz1t7lBgYjD/Wi49
k6ZN0brj+vjHjQFe27pAdIuWIUfOxgs7jlK6uhVuy+35Qog/L/ywX26KVm9VlYVP
jUnhvJOJcqNyn8IGk+S7oZr2g/2BqPWLlDy5OPuESb1zFB9LS+44NdIP+INv8sJr
dwcNu7PE0lRhGFMaNh3Y9WHyYOMARtf6fJDiylN6Lkq6j68YcAhjDhJErKIVZD4u
LVgFCRKkhaisajQ1RXHM0ZqxDJ8kAov6ky04jGwNLO5qaQdFDWuXBNrSB549kNMp
KgmQz7wplO/tk84Ued432PtXrMoGlRVjsQLV1MQHH740jVrGkMHdsOlGqcI4UfbO
ShIstaOy4HgsoBPXkKSweDR4j6qXKzvsCROC5PcvIKi9iOtnaOP1YlxslVDzp3EZ
zgWUar/3Tx55+pLJ4D4eSxIwXU9RD3YKf0H+vP7A+4VxxdmWvdVLTzJUW4/huKDQ
VpkUl8dEJ2pOXGp1PvlSaCP8Jf1VCwi2+fZcoF1zP4+G0W6aa4p9HDqWDDCl69ix
NjRPNxCwSHa8Lm88ByO5FmeTt7hp8dMk3cpZaXDxKSZI6oG4hjnwVxljzvZbbsuM
mAsgjWd8ikZ7uBJbavM8a6uVqUbZ1FHdQpmvr02+bsZVN61ZfmTCIl2CxRoPGhh5
1tuu/KQddC+jGHSdee6p5DEsRGax5ftVi/c12RATgCft3is8d67FOWMGQYhPnoR6
vvOWr3cQyNqNTBcrQ/S0qOKVkDUf8luV2QAnpAsFRHRJwpot4vZkkEaw96wCY3gd
kd4FbXYT3Gq9nMHOZbyJgFoMqClEknKmbiRwo62Agg9sjhgqZyLeQjN0RKEHtiRg
XfiuqkPjirDQDs7weWFSyx8dD25FluIoZSdhJIE2y2/MlGnoGaeDT+E0DXUxDJ82
7Bkhqv7hRu6/vETvFQ/hUPrDbtjmEBdY8rUGcwXC0mA9CfwUqEJDqOos42CTjZDO
cFdCTZtLbALZK/tsFfSk7CuZDFnPdZMx0zY3sZcLmgS/R8ahaucDW+4PLZUVJDMG
noJCN4gwxDwfBG0NQ+/h6ote+790t8NdT42FA4nH/eHjM/zbx/Iu0RDV3abxY1KJ
w1FVUZFo79WWzTrEv8lUjKdvbchFN+ZyIJnFak1iBz6wYNGVtlJnGxdxveRXgZDz
PVn+vcIvpgwrln04bJMmfkkTmafuvgSlJnVfR6wNcai4law0/tSIDtmz7jO9skna
jiIqPhfegpf3AMbs7WsGs6rYT1NmR9dLjLarr6s1LbfKV9KPH0xB7/CwDDwN4hHn
ur5+4yFwsq+yVC9jlVUn5SoA2iOxNHYfsnzC6Mi/F414lf/NLXH+PXMxECWzheys
B/1P8AWpM6HGlXh4JWTi4wxHM7Ou2gGA4lIMf4MwltpUPD9mnuL0jBtFPrbC6l3t
/aL3twSQTqw9/dgDz0IV5trT1pbgX6+XCtcTq7yNTOPSimCPTIVTYZ4tDu1dJt/G
QvrFkj/f3v1gwaJL/657JuNRRKeJaaYsxT0/TcZ1elXUSLQGpGfebYNMqRVfqwPw
pi0xZWbBVrY/XWKMrAx1BwWQaXiDlkrrP6+l1zT4WOJFAYGWh87V9Xs3XKWkgSIE
JMjKbL2tmc5GUZBarW6RMZls0egQjKI6OogsEwZgpF60zTjJGixi3Xeic3VMLP4I
k1szRcjCbLsDZvb5STmaOs7e5IsViOt2V4prOGHV9qY83oHpXR1kHMNId7N5fbOs
42RxTIlUb/INdyG3p4IMI9RdMBDeawA/IkSJk7YJEqTBP1DUZJSd/7WBVcvZgaDt
aS7pxHh6oPgAD6UDUOj1DQg1lS71FCJEV5fPk7nvT7wpsEyVnD9Gk/+5P1+GT8eZ
P/5VVD6JXQrC0X8QOT2AfE6bA1xyJX1XDolOBKTwcS8z2AoXVuUpt418fneIewEC
MOAp2PKOkie1joNBwxaJoBde75ul8ZKFvq55n1EtHCQHwp64jS9NVVNVN0PyOG4k
g1wpj4mQ7E01YxAw53n7546OkUJFS7+LRMwRAe7VXXFfw6uqOpgJ/BTXyxUjzAhV
GefzLwhF+D5CVYajRWHj6iSsSa9+OICcirJaMn9LgBE00I6S9ybpQrVDOmJ6fVf0
dBAb6yUOywqS2wVB/LiRXegiCxbnSUlQ7Ihv5ApB/k5PutaV02IkJPAdPs0Ai86b
pgnh73KC+u9u21rLZJOkr0ND0BRHVUeZVHYThybTy2MgX0K8v/9JyNpXb3hsNpMa
HhmrHx2KHW+M/rfi8B3QpdfsNe8mmGEfjlYDgCN9qW0V+h0GosqQrmWkZzOkzs+J
LpFeVOJp50sUdPTPZ4XsJFLN1gxghRIgTLnPHYeJ2r5elrZP2abWAty5WGGITVx8
qss1VAF3XOQ0RxzhUTlOi0vZMBRwA1fY8TVN8BLDFP8YghQMyNXJ9B3HYtfEfkRq
cGXfQVe5PigH36UtFnJiJTMpGatslmBzc3hbz59lnryucGnxn077XcqUsrmOgpGf
qoUTeFT8erEALrkoQwFD6YqEkvWcAWNbYg2DwJgR+eEgrg6JqPWhyUTYMSVQBSPO
hyxLTL9+oRJRPprqQHV7Web24VfXzLwj8yq84Mr/yFoQ80WefRogJvVDnuAF+oX7
B/bVED+IRwp6nK2yxZOkwl9EiXctlmOYPg/w2SLT8cXcC3+poDGakkbzG1sHlIhB
Zfbgsr5Qog569O9BKJHiXftTrGxsDrkaFTOy509vqelKgJATOxREUKWfHgG0qQGz
iHq0EjHlflfApKIMh1YvYL+JjYiWwdWjk5vOfNly/zjNOgUvhJoQ8n9MVLXvgL9n
WWWajfdfYRm7jb8UXtU93Yi3aznsFXBr5rf4c5wU94g9YTE6bJDIX4FytGe9W/cV
phBd4L5CTQSSljzWm1IFGZDqVyf+XLjMaX+5RFUGMnUo8YTBJExgU4J3Mr6C0ipX
Yet3mc5lCVUdPwfsY9GAvzslGiZh4iLLAUIyyTyF8vO1ETFP2418/HIal/U4vG/X
UNZYLMG5w7ZswRfgp4HGjGL4dMQXAUs7dVr7ncdF0YCHsUS+8ci4inMu4+tDpmEf
yfc/P+XiTBXVOJcZkj6V9JOVbzTA33W3lWSy05UGYBsw27y1tut0UBjvIKjU3lRZ
Fk/uahioesQB/DFEGlL1QjSqw4P9xEhHlAtyc7REbezmnUeKpy0tnVk4/BlWJx+b
Rxl0scWesLenef1l/tV7/zvM+hFF2VSQrFT5KytE6zqxPdzje8waNbOPUdXe/+RA
5yVFlI7AoK3+2mo9N9LISDid85PXZEhOOW2Z1S7sTU7H+9SfFV14Do1q58EuZehd
XdG5qd+DFZJE6kNdIOwEd/5NRb5oafhbAxwrrh5ZDAR5sUfs3jSZU285Knbg6xDw
H72pTeAUXGgLfZ1oevge+myMEY9ndtSSBc8f2saj3pN/jMya0zm/yBXEYhg+ehkd
5lFHOwpBtsKfp+NcOY+hDXAnInI933Lxp3ZvCk+LG4QsXHDY7vyljaiucx2svm6n
XhIuAIdepAKbFM0BgsENRkUnG7P5WXr8SCz9tFJKZFw+MY9etqXkvghI3/4gC0mR
eSBUFMrs0ycdUripLg7bqnUv5WSTcIQ4SFO5buHM2BEEZzZBOEJXg7gRDkyvwsgk
DRoanS5mNRT2zoogZkn+fnid/Cv5efEuZfN3WbFKP6oDUxnbi0cJSHWweJly3G+f
RTfIR4mzR9cSY0gWbDJvospTHIJ8Mr5BabKvxk3IwgPhtSD7YihTsZqgcFNX+aH7
rHdfXz56ddh+ahop1CSaJUWCYmiteXTZ+nNYdos/uib9BjypNRFxN+GTL85CLjhs
X8NI3MnMucw2WnNvUQMLo5KlW9UJJgJeRA0/HtpdNuWRDxyOh8wLAYnjIztX244T
FW7a5T15H6shB39Eq9Wa5dTGHf/I/KU2wEwbHISYlecPRwbuS7p52L2wmC16+xRs
R6Fr9d5AyMMOe9oFEn0Avug8EY/thX9mFfndV6fgaBIL77HTRGyaG7A4uiYJ0tjz
9y20KCWcX5itNTzergoWAP9e+pF24PSyaDo1sjFXHvZlnQdZCG7lTjD4HLpBrC3W
H4q0IVRMgbhvlFcfn1YteOunPheo3B8eotdwW11JEGPG3DGVJPXw3FA9Dju+2fM4
YVIYBzritLhLCqUTKSp4UzpbI3RogYYpYottI4cbs6uM0p+HHxWxYjHrmT47W3EW
ZUbl4ghZz0r5ERWNq6IuuRwOgAgFi6LTnz1y9uoaJ2ITain3ly637LlFXncnU0Fu
zgz3DjlfGNqB0aSRLSfIWpm3lc74E2h2r/019+EDR6sz6kdibV+0RjcJXg4arbK/
EHtGdPVS4eiSBW4R5W/M03yduE7UmNOtC5eT1JX8XKFrFgjSrCW6/pGMHfL/Ib/g
PsLoYcg6LMPdGOR0EHMBfW7XBoXWNR08nZ232aqM7wneQzRIMaHNL1Mugjr9Bc7N
eTswOg1jWCHmglylkNp+OaHWy48x5aqw1jwocySatZrPW7vl1mF4NSA88zItWsNI
mmGuq0bxpDJ7vkF+2NWqxOwiMkUEBIIqkq/bxJwfhsNBuNi/aAei/PCS4atTcl1V
9zblJgxrQo5sirPrPY7TCu02KVJ0C2nPc/xTUjIhoDqQeOYcggaUqNFmRu8lcNSA
DNkQBXs5nLKaJZBVOBuqSTjcmbDrwCCksO6iibbbobKbRorMlfMdIjG4ljFsJvcg
jcfwOo+cldVGsHPa2fBKmT/jnWRrhzzgPl8EnML0AOp2iDr0FEvk8SLAe0Z1En78
ql7SDLEC35Pp1CDxHwLfQqFnKwBk20QWvhr05xjs4Y1hQ5GQepR9vzTjMP8fjYvJ
DbwNhb867pYoe6XlTe11HErh422/+clEs95n7XUqTU66g0qp8ApJEdgjDj2m1wLF
9l54BxKYNC8EPM9m0ZLS4x3LW4FSS7I0+d7KldEZpzv+lqZ0JFeqgl0ZSu7Bmiid
41Njbvg9bHxwRDIgM1ZbrNEz6iM33hKhs0qO7Oqwf1QHHh10W3uJEb217cFv8gQ0
kUFkeJQbVaDuySWwWUsWHDUv3rM8Uodb+gxW1oONkhW5V5BlhcOfQZ54YEq70aAZ
jgt6pbU8Js+r2C8fXiJHOa9zLhK4GRmzf5X7z4Ej1wGGClK7rArJvbSRJaJ/86vx
22fsLbWEZcR6xF7w7IC+IMRINBigY0LyZAzGJcEeUTmmKP52q+3Ff47BA8+uDtl6
2nxmbgj4IdZtTduncTp/B2abWvb8VhrYTJwZhThhcG6/tmm5U/ICHTACS1DZ6Q+f
2OgpH7kW3HJuU9Cgvaxg7ZR7eSc9a+0gdQRl2TnDr/spQynR58BXVXJIICBhbf4E
OjeILp3x4M67hCAfag7yWzK8OrL956uq8eZtF8eFRj14+VtHZQGzpdL9NQJ+TBQ8
Tb2REpK5C3We1EC1uKCeZok0GT9nBm66DKVDLjkUenKiPUQU2rbcwSAhyNZHk7Q4
dIJBi2d8jspCoAkh0sPdrWcWCPcPqaCVrCY5OtHcfxmiLXyh8K5bYeL8lnYyjcej
DLkzfK+nk6DUkMmry5HDRfXIe6cbSJaOUdQjI0XZ0bQGtm+hcS8MXiqDrDxB+GkS
yFE1yvF3USNSfxmb/EEuEDfInU9qtaZaa3eLfa0e8I9YS7r1mJLtTV28XNPz+35C
H/LtaI+MwkBE+ghOcbNnWPCvOBrZFyOLkJvUEoNf7ufUFhzdjHB/ttb3Mcf4yJd2
hPhpkxbE5gJ71z3VxeeF4GYL0X+fRe7w+iO7VaQ0U3C5426bQjzwIujymrdp16dn
+U4dLA79L93H//zrw3WyXOVU+yGHFqZ7YBIPmWoSWO2Qq4n5LC479O8V7/xOm6kz
SmZNBU5NRp4lIRaYVCftng/HV4RRwTa5/pzmao6EJoNacfITyS5KlmUFAV2ib+8U
tKrkjI00bCq1pWjQPk7luIxMUeLX+Z2iUgDpyKNLVpjcGX91GYusedkbiZlVE+vZ
i3kAKVUr9ikK1VrLOUIomemwdy1GN3rX6aJ4DlO0FKMJSOk8VDa5YkwEKWb/nnI4
sPMb1R73oJwyiPH8sHX94WnUbifnce/uQhqMmcBTgaqH5mbK57Bk+Z/f47SRaoFD
mELVxJ3vVPOHFyaORP81f+LA584N+/lM74qPQfWpGw5CM/gsLXir3l927BSzjwRA
4BZDXiS2A4CKJor6rYaRVGr9oUcinIcKsJ0nSJgTVbz5yKsbUvYe6Q7Jj5HI/lfD
RiD0wHOYsl6SWzuUds2yvgNomtpApIo/hWe5uTbOs7q8S46MWVk25yOrHOVdCHM3
4Xw73DCa/lcU1JExE31+FXC9Rl0OY6XdG3iQZROwLpWtz72AC2h7yZsHDm2leJEX
ABTD293Pvvd2KdUjHZF5Gr13SNT4mlk/oeYKCmjZlqq85Og45nWjud3NStiTL9e7
QGBBtmFiZ63EizP37MZUxKb9JC/Suwm6dwemg3dfqA4birZoYWtFHxZertqBpXQY
9V6NdpwUTYZYljR9z6YmSjY+/D6MWulq0FR5eNTaySs340K0SMVjA6OCjmflQfNS
moc7E+jCL7PlCYJWrllrO7Qk4l+ysCOw5o463wPnEDu1oaqBNS3TVxW+XFhjP2/k
ElWIwzdKu/nv6iKUYb7qfGtQaSTRKfKJmvmZLZyH77/k+c60mofwXPelTAV2GEkl
5KoOBgjYEVwP5Zxh7W4n9uuxeEZfjxXY+pFnC0N5aZEJZKx7tm2hNW+HRptz9sPT
ffx4LsHZaLdHyC8TACGJzyIBq5k81qYvphpJ4GPOGO2yqSC9d0Bi4GhnzgA7G0O8
KFElhEUezJKyRF/gT+h0e1yRKpxZcFA0DL8u0lOA0Y6KFvr5xHewcEUS/e6xLQ/S
7EoNqr4f4NfPQtrqt3jURU1cub1QMkvM/cn6cOmNiBPqefayfQkFdINFeprBjSLN
ADVeBUeeia5pAjip4EXjKlkWyeGCBol+8lEmMRlOdR8nq5EUCbwG+ZM355ZMZZpX
D3bUh5JD/O+ZjfD6Y6/W5Cd/6cIJOL1deFYZk/s1j5YetRB0j+seHv1qnFvn8ttl
XB30F2oR0zl5MTfbcBdwXHGgEVyVkTym2FTHog/p7dyzkjUn8kRMKbL51kdVWMuh
w4Qg5x2WNHX+IdHy0h2QnLJNnO1PBTnLTeHiTpYsQCda6SOWiztDqs+liytL4kpT
Owbw4yMpnt2QMNJ6L7AUE4p3jr+bAHkH7alTnma268GHUp91+7t33cIJuwrqkhlD
724U3h5PhHvtAkxYO62qHX0VqMCRC6ZkTcBUN9g8Km95vtiAXvwnwlrBUoZSAF2W
PsfUHHAZlVruGMdt/1qAF6r9aeGErnnpgiW5OLoMrr0=
`protect end_protected
