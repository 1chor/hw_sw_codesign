-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
hRWwqxEpID7Qg5vo7WSd4/drlePBC6lXt3hHHUASeFjCW6MalMS5lUUkS8iohW3C
nAdz9pFa8lJ7YURpjw4vzI/t54iznvwkf8NlDl2WMgfk53U47O972bwGGRidsQxq
zL27zCPeKjU1U2AT44FPOYYl4scJYZYZAGzBdyLNuZmobye3ILeszA==
--pragma protect end_key_block
--pragma protect digest_block
FjgwVr6dFeoDqzZD2w7qWWavgoo=
--pragma protect end_digest_block
--pragma protect data_block
cj73gHanZa7zWZpMGwMGF3Ze4QBQBUJL8GBeKUJ/k1Stj4+YXhRO24lCqfvKamRj
PZThjyfn1k9NzIfeuq/V6hVynGPDVkNqrxouozM/n44mWNHG2vYj16r7BwAGrByU
yWi0+lMOrrvC8Av6tp807DLRvlURq9jaftu0cqZJACoKBbx7M7CYZtZbBw5shwMw
tAiZtWjQ3EfJV6fsTZaEiqFYRJ6TByZF7OJGGzTBASAv4OgDqIiSosXDAko/PAmr
zGg0zhTHN8H5QAp3KFrOmAtpIIzCnRSo9xxfQWPEjjCDVU9Dwkt4KA0lhYgoX3hG
hirl0cy3rRd2PI+0Vp71dg7BvMEbDvo3o7kpEB4TWEbibJlWpUrSuByJXWV5rQwL
k8gCzLjS8HFqJ7H+7GtpSzDoAkBmT4SZc8+jlGWi2LgPeAmYWE8T/cxrGkx5l/PJ
EZPsBF085i0wMQhhatAke2cLnxN347bEvQSvhBLlRzCvc2d8EvzeEifkfP1lsSbp
iIbCxvHPIJbQKTuYIbxugYq63hn/kC4dIsOYVIzyEysA2N8UQ3bJu9Rtr+PqfCMu
aYKD1RYMk26y9nqfUHRb1lVj08JcGNKR3LIp6IwiR8rnXTG2bbxeJMn/lSxjwLgH
gnXNTHzdCLVEha+xHa9s4BAXv//L2XRi20bFQV4kcHeX3OS6iW0LQ4yd3ZWjgP66
ZMcswwphDf5rCxowvNgFDTPP3dAdTYXeocxZR8F9hhyUNw+0PD4Kaz0qopZxVHK+
jIaxBeHQ0J6EGGQMh24RGCyzKGq3UMSKd8tlH0zEwchMvYZ6dv183kOPW84EwyJt
dpGeX+YNtFLMI2iLT5GmoPTkwllpLWZ1lb8C0hCmbY8z/D8nI0MRAZdbKm2KHfnu
IJTggKthKa7RB8j6bt2WrZmQB5RPuR+noFUoCIeYdu2vkIKQkWHP4Keg64bZIaBJ
17FalYWMeqph2XMAxCs7+zR6Yj9px72u2PArYrr3vIeV3QReRMAdh5ym0frZ+jdj
2OHu/KWJtdCcwbfa71ax8J1ejJ+iyPZLsUf4EuFklrO6z4+CG45JBRkNFTLH/Gkg
aUfaYuRKdSfgGHr6HpLv+YTkGqWfojh8T5K4MIfqlDuxefN/SqibP43EnZ/n5m7k
ea43SC5XxfLKNsaZX8uLN9coSSsa8d/0h5hyXr4qkAd3bNPnDzlN+UFdgdlsJe8T
NZCT1ABlBUXuji7hM2L4KvclbdqOwCCiXjWXDbLgTy16UwVcKCo2rqofyv7sq0Ow
LB/nhhRsXHHgF8qN3iXO7hHjR81lhYDF/A0wHkKHZ5jtT95+Z/UybSO0IoWI963G
3Q0/S414canGFw/mm3Mg/D23hPYZ5skHamTlDYqypKfV45WOuvzrXBhVdSC9ZmF5
WR0SE2w1DJ27j5L3Fq3v6KeOej7fcMWrvLWAe2oe7lKPB5sf7Y24B4NPqh2HCSBz
h5dqnBid3h4GkE+5FqZ3W/JyY1myUadvx6fZSe3yE644Q6UcJCdIWyJ9C4qY1rMp
Q2w/KSeSTKiaZUKBletQv9P11VnwmM51OJKbcUNq8f7QsX6m+yOOo2SS8K2kKGYf
XXAf9Ov1QWIrkJaR9K/sPO29Xh3H1zqTTswhvN4RO2SfeAlS9xuEa7TDwWJyXAzQ
n4gQWDkMRRzbEqxZbsqP33+gxskhUNYP5L17Wfu8doA+yhQZnnm3VvTjUHiR0fX2
ROCZSzvTjsVVXYRaQLeeZPSOjkDeMgoXNEAvlynQ34p5JWbVNxuW479zcnqcTnsm
c7ZYOefEz9WXjWIwisMUfH5FV1Ayo62cniug7RN5iIvQIN5ELejVHcRIorC0jo3t
oTWjrp9bTWF+kA7HF2Kf4awkalXjheVe6QREiLxmV0hWNhtBx+cH27hdZ7NPn9kA
ItmFfdOCyGm733lWvIw6ezs+lQOArcV0c+lX34ORuoQDHxG/HQNc07WCB766ty0p
3NLyYzdiQLlAc/6QVHxqx/ZF9TI7mly96/7EXIY3gp5qXCUdbcBnzi1JGC0qNy+s
cZjLi7IQXyf4vM3wEtDA04icyTUUQdV08GG+EPE5TUbo8gMppbLZ6FbR0sQwaFSG
B/0+YWJS0om37YME1M86g7kAMLnxk/ccD1B39/JW1L52ldWGulhDjZhVV4XgSMTk
DXIy86LJlrKKRrIWyFXXmL7OeK4AWBwGkXmh+zJUPmfLBLzhM2MHrbnnc5uJXoEs
Ag0m/hL4x5+TRE2xsdqY32BRXlxlTaJEn2FztWEjRHaZXjikr/CizqFPw3bqsg/2
UTkfFF1XvQkYhwACVXbIXSZO7SXBUqmwH1JP+ivHr67ED7BezRdzLt+z5MOqtZ4H
Jggj3iL08uF+h2Nv65juyL21r/gGJ+gZSdh/5P7xWCWUvtHc/UW81e3U6do+C/ZX
Jfo6lzhKpQ96XsgmpTQh3o9zzpcCWm+pRCZcp9YY0EBtfuBWr4j16cKCYX6tX2u3
GwsNvOU01Ow8QogMYwVlzkyDocvg2F/nSlvIlAfIt8evRZ1B+96w13nYefGcxMyw
lihYM3IFf/lYL7fqDL1tejNVloLX4ZQ92MOSxr3TljI9Iu+JYHGTPx18sGUxwzYv
GasxCuZSE/mzioJ9FI4DSqVVdiabJnj6n08EWWcJIgcvWu/jN5aFr/tN3BfRnIFG
RVSRWTEBG/KHrUNb22ve6QkleCCj5KcIZM8xRJiVtxAVXSYx2LEnl0u/RVvl5ZOV
pEBymJaeKm+dKYN8LslpNcJAXBId6jNYfiBCFqhrYP5Rjuco/Zi32J1aB3eAeacD
kt+lybxlGyF67WbAMLz7SAq/WcWbay9eBs78/d0H/AWtHYum7KWh+fJ4/onU99je
XtKj5JxXp9osnzOPJMK5/2UecxLozCaZ20nU9hDkyJrrJlkiixNUuabzwYu9OYR+
4T/kRNDwoPnLx2QTS9cDJJLx+s+M2vOSO3ywwVElP4e4N57AUssO+4QMc/UOZe2k
puyUGmOHqAQyGCV9RZHozSzFxPUC3usZDSXmnOaHYOr2/L6p+GyLgBhYIpY/XaHZ
fjxHeC0y90cTHK7edwtJ6gjAUvalebwDjHBb9eNrsVHddJh/98bP8RAvIOg+PBgz
PHsL8EHsvwdjooKUzdHsVXKfWJK8su3P4gvFPaNKRTYSy6Zk4ATV+kUcvXNKAClu
GhcWPcLvlPna95zt2Xlcq2pWqcb5S1n8+JKe+JfoiR87IuNNU3t2pbdHnC9PfK6w
ivyLy2K3UlhlvJuLmuVNJc6x4BhFTUE2fqde5v8SiU6pvDoTJJmzXMrOlRw0x7uw
Sav695ktFIDSZgQh//hkiG72UAKaGqUqp/x6VyM/4Getfp8nFsN8t0lLU1bpkdIh
n12JTiJyUIbV+PdPVplpGe5/Zh0WPYXgzgILMmuehpEBPZsAd7PezRGwDWWqCMC4
YhKang14EdWX4itoKodq4hQTRei9hgY2k8z2lnLp69BmrHSH5LAYJD4BUE1YCNID
t0KXiImsAolMAXC8BM8ofYOftwbGP2Jbv43mJEw2TwH0BjM3tYxhMtyVyM5vZ0g1
eLL/5yTVfIp9XJo28DHomIHaVakyUswad0SJo+2caNp/kMn/Dcl24zliI3wvro7Q
YQLSJWt+mV5Vu5b6EJY9w1LjtS7KUCWN1CAJq08OLDl7uvoKRS8xtfRbkf9rOQF/
pUSNYKklNztsBY17+zk5yzFrBbPvGctEHgzh9ANldMcBqMwxYyXaP4GpiqYVYSk1
zRYa6BPNROMeQa8ZdETuXGg1x0O/WpXoTQJ7Vb6BPSOElUFig16Gl7fVQIQy0Y/a
Fcf8PjICWPx3auJK5NiBggxZH/pOojn4n97o6uEgzuI2VsuZbX+4c1GmiYI/Na2e
A83jKVOHl5NIPm0krb9SylNCIPjchAYc+rOdn8G9jFIxbdYTewaVxdOaoXjCBT6y
xDjd7WnxQOC63zCbJbwyUd1c+lnLpncRbbJdAevrjY9a/RkWNc7uZOI81/BgQKA4
+xh1o69Qv7UtaukbvaNrnp4/k2uTUdbHVMXqwwPj0jynkYm+oZXPTkF+rWWcKydi
9mYfzQLEMQ8uVHfQFS7poRmPFDa7lrKNITgrnSTs9zr2AlZGCf0tmD7auFZLM0vr
giO72/V4Ga+08mKvQLK/slMpPqnLAvv1zpyABGXk2pfo+N8kdE8qflWwNC5YSd7b
7G1KJ/YWScikuRzsm9X686qkSJGwflIO1e2QAfK5awrfSg7K0LtR6KN8FiApgsSf
nUoTmJaBocjTYXtNMA/A2wRksuWJYu2NdGgxXFTGiJpeLN0o1S0i3llu9oCp78Xa
m7i68TG8g7b9Q+Eo7PUcN6qGhpJin+UyTW2RJQspgMXyO+gJoRk/vNRoEPNYOKci
ZPZQOIkkewVnUaGn67OWUee3wylPxbV3HIW7xHzB0JHXpVKo0e767VLgbdAsZabl
OkOHqKqO9kYpITBEAoTdHL5t65eGl7Jbd8l65QIN2rkiQ+xk4oYUEK7SktCtq3is
nvX6/D1xo+SdzUGdbMRrPlJ6w0E2/de4nqc/m5dS0UBiM5P5Z8WdJmRlPcke0ncW
dO++uJ+w2YYGx2APlZq7p8GBlLrslNzi0LXG8xbsPBYeVkQl+xD6bgU7/ydEgKYc
7HjB3V0fPzKbQgxk3w1I+v1jYVY8CL7ME/qZlnUA/nqof/nuulHNK5nU/3b4VOIU
aXfOl0udf9YRe+rc0Fc4A1OjM+KaVLnvYq9wuO9l1G0mf19OwN0+T4SfvUjdAq0A
YY748Jp+o/1GVmN/gctZEkQGJqMtd/WnCPgDTH3faYEPEIgCD0DQq9gQaOGVmbQz
0MlpRdFRuwZsS4iyVseZUvVpvOniJarsueA8Xdx2KCGlvbgaiUr59sdPI55p4vSx
tieo/mOfPjp0LF1i1e4MaXfUJkJrf5KnZQ81dppXjOkHxv4uDqQWmp5G3ywVBukc
Z+Ri7blkGpMDfBSOAAwygQzRw37Z8+zY4B3ClBkdQQ5TWt9LjrAaAiaglGaOPkT2
3XGnhPmKnXzzKb5jQsgCQB0mW7ocpxyXlkqZ7Eoaf7wuhK6TH67UhLIjP3Kxkr45
shA8lShvekfMzRwZpoP13B5RzmRFHrYu9iMbhw1AHqvVnq8t3nOG5DTTmh05ggMD
UZHLy0w/Eo/vFTfbj0N9JnZjz97Nq7kuForvfQk5wur3/b5D5a00UzFa5vKpjgO0
e8su7Ddn00nOkx1A1VzuYtics0Wc4W3KkfDR8B3S6+hZogtly3OML0x208pX5h9u
s04vlT3GIXPojKDR/0bhqCHsNORDZEDiRqD/6pYuiJJZEqCLftsgz381BE1JRcNO
fobNOxcKRJ2REHl2QFas7R0axqbeKGibdNggdxlXaIHTTHJ6KThJx413gM0bV4iG
BOWISFnt2KI/M8UzdwvZNZhsRugJ2tSf7J5OfCjtHfEK2ShfjUNITBjPxkhSDYM5
fk2fZxRgraqMtddysgvLU6FJpzS6mtIzBjt8fqThHIVEdpxjWaFeOOs9wQ5P93iH
qxbmQGF/W1IJvT9Gkvi8k8goc+BgP+OGVsah3E3Jkuk7w3Iwyc7FVNnH9NaSH0eZ
gULqua3qNVDlOvdRuompILJsnerP/iZg/NYijsQ1eJchClxnFZRmv7VO8rsHuC8u
POHr5oKX/wJD5bCv4zoLh6G0qbI/aw5ZznHnSPzy7SnurJwhPFua9IgdYXdHhsjP
D1nvOmdvqgoiRSlohLUb5Q97Vhh37xBlQ5umlnINC+gSq3z2uruqEsMrqPeP24To
Ox7sFAPqMaz3X5SWMY0/K/Aosn4xBsvJrJcseX6OfA7268r5q6qWidC7lP25bc58
xvTTU0rEF30U10lllYSii7Y8xhq5ZCeOKJp2fPGHxGo3biNO8KWhGw85zdlWkr6V
5OywphClWPQnDTntDbalmByECjBxOUEaiWEXT/ByQf2AKfnvsg1DydIiY+ENYVTl
mZWa6uIOgQYhMP8oZVxjy+57DJg9Q39LVbq+i12ibU8NtGRiK40cqD48qVR4OR1Z
5UMpEKrTUydf+Mi0972nCPoaLiRm4+3YM+3c9kePpLYv7UaKKYPM9IRAEs5POLeJ
z41oWGVX+QXkFZABJuqeb/XeJMrvcq0FZl8IFFyFp9TeFSZGovAxJx9VQrud3rlT
LC4YnB040i+wzgDLNWyXmsSPJiBcEjJFF1CcnfR7BHw0ipOqdCjXV5GiAB4mZ/Zn
/fFYpL+jkY3snxUQsUXvC4ShcOx9leWH7Hn69NJFsemM/J8LDiX0qM4GA7EzVhMD
lv8bAHwWly+BRwCFz272OcBGyrzB7WxiKt4vTIUCa9x5RI6NCQuLp0rjdVOOhJIl
IfxxBW1bZh7FQSc8dfuRPYuQD5GtYkx++BVRqv4kasN90QN6CkdxTTIXfLSNw4ro
0TcVGZ97VKojTYxCQh8ubIlF+tyFXR5QU62E8Q/gFMEtHdOaszQt6XWbL289Bs2Q
koXyv/78fekgsn6tUkAS+XmHrG90jYJQo8WyPTZXtWFg+H/69AJzOiQzw2O9d2z6
K/GuLbgcJoKF1UcQmQN8nnmEeLTY9WxMOeI5fIJmBlwFcBI1FqYdrf9MhlsbgjQi
E/8yGk+JKyEF2mBGU+Ua/k8KkI0yQckqQrueFYDjXRFB0eyWbQAL/5jDqFJfjMmn
VPdci67ffUfiaOhrbDczo59TiLZjl4cCczmV5M5g6ALXXvG+spUJkrSOGKB6P0Ey
peIbTzOWSUjB6W5tJMDwZQYPTFvnAsAfBTQJdz0qoY/PniNnb0/gBiXhdex6hNhJ
n+S4HlGtebldEqQFsdIQMigpZB5ERbDR6yXPzmFOMSS6HJOfLm9JW81YiwJjyXAA
pYRof3vYiCt4AL5GJgdfY2MjBsLNayrBp30iP57PpCLxyWl8Pipuw19MKd0IGgSM
jSmsvIGaFo6l8SNwS2hHqbyglcdEZiX/AqGzagj8Th4VGfZusjwU+satJKv326nB
ycClSe20ZEdFxJjI2MDbYA2kaIZRult4fYw6K9y74RgpRJ2GPicf9lUMR1owSl4C
3BO1Qpac2Ngia90ofXeltSTmpQFuzTvy6PaCSVEm1/zTVrsCgKADGrn3otlTWt4X
W4LjQk4Qv1nBjIRtSNlAMVWgtDN7z4PttFcpZhRwyUR61Rz5QvxxDiLdPZ4LRpvh
A6gcl+eHCX5WImlv73UNGIJ6VGu71MCY/ksKjHzLebK4a2VUtIl4k/bY6pMt3KXP
+WJoKHc9RPQWz2Be0Zb1TCp9vjraL31cokOGYyPv1q8NskWs25nTNQiUJcCHB2tN
w4mkoECffuykY5VoEOm10wYpU+PJz2k0RWXuD75jOpByCI0px3nYd/4RPvjQVbXU
IXk6YbA6rRcvcCqrrOxpePx0sXFmiG0iUhFi+GFJO6XTegZMn37/fASkFSLy4kaU
ko0jprO3qhBWtl3EU7rE6Fy3R92cq8gqH4XcbXPZihp9HZWI3VW5E+DnupkEgt1n
qGNYx5KRVQTQfZAojw2ZU7l28YrhPl2EqpQSezzwKyotN6dOUGYt0Xor3TWuISiv
5xg2HXprGM62Jjv8+9iE8WgJqG+xuWOofQBkwRGtXcDikH2ow5UXEUrEC2GM6ptX
kkCzQKeym7fselPCOzz3Aec2w3HsNAOAIH3IP5lfe7ZzFNXYtmFNU4rF9eEhtjJ8
kCWjsY18vgSbMKrdTjwm1mpZG2U0SMSpNCdL4ho/viwkswCtRjcdJcahauvFa7CH
/weIFuMGwXYBlCKUum+uj9CUpcUqiKPnN6ic3CyvZHPilf7xhGg1Y19JZaM9yvLm
G6f+oTr4vLgl+yZ2RKKNK43p+TZQ1jgIrQZ4gqsi7V862nLa9bsryhwpNcjATvcC
I50zKKtLREjQ0b6R6qeGKGb+WNTMpfRmU8uEfDXIrM5/lXHywJsjRZaba/4MaBk0
YSthi9hpySNM8u5kPokgHyplStTLzpT+apa50NR7moSTV7rdP+CtETIMuC6YfU8b
ztqOroy987gIZY4vUFPB1B19hapHPhEvzbTXDjLmjvThbUXCdoonqBbHy0QdcHFj
iDtv8i8v1d0OC2WY4pIt8S/ZhsXdE9DFaJHex1CrCMSbJqx7uw/GYB/lF/c9esX+
o/Itkwh4ZKUDk8iF7DYrYW2CHIjtk4uM4IbxS2qmp7QDen5pvZ5WlkE02e2Mumg2
QDrhuNkvMz87sS0NTYWVa7jj9NMf3ij6s+4nBlXLzfN44WLcoPXtw/cqPTc9tZGf
UQxIvIH0bqvkHXS5KzhjgXfULm7RU7UdGi3+JYKeRcBubPyf3VC4+N+o1gb2IENv
Q65uW49TlrGtMZa4/2uR5aqGrfqlhm87P/UgerT+pjFGhPRMsBnHmCoc74pDgbrV
e+9SV1A8kTY7Bl08jHAWn4Uxooj8JlZfYZKIEyQI+87ipn3b8carJKdyaAnJM/y5
ii/ZcT8kUg+IbLIkLskhyh5NycA3Cm/J1gx6/HyX0VF9/Fx0Fb/dlAFUatC+nL9X
RczFc6YD6HFF7aaqDGW0AwS6vbr9aj8PQ88m4CY8h0lDR9RwLxGZKud9xKL5RQZt
6tiwGx1SkeXYOF+cbnLBkXTLqMSZ13Q6Y5zjwGZyhf0UiAtDmhjAfN5h8r9ppoIF
mc7cLpXZXkOfpUTS4q2/H8+/jyhUrjXItgKGlN0GSyAy/LOEHdEV0cwuawUF1G6C
PCZX+WGQZdVVSxS2eIoHSce6/nghu6fVJdpw938/sP/LIdAjyzGARvNc6fA5fDvY
+yZPLyp94kPlNBJXJ9DAkhEU3A9ONccWXqWgX/I9Er0Mm///g7fTBlf6TmzAmUv1
EHPwveKgrwxIXUHewO8XOk6NHi9rga4j5H0ZZk/LYwH0884W0xw6kGg7dRV1l1V3
JWK8jOsSlrtZzS8oA06oRwjy0umD8G7Isx+LQOM0m8+0ctiBp/3Z421uA/b3HoPS
EhadgJtyZfHTuEl/WA+Lvsi/RA7Yrq5mq0yj1vp+wki0o/aKbBd5BVZ9OnP2Fm2I
3U8ILTe4s7NVqtJpIq2v/T1ueCRcplcydaHz8qkEhHeZnLbpxo75fU5qV7pyGGGr
2iTf9xZdxnHSPXlVm2MBMtj3Cc2mNQKs2S+GUKG/1TztKnRU0+ja6IJgjVLWtAwI
9hxAe6vRez8a1vh3702x7KWKViLwLUkhgNDz4Uq37dKBDJHMMB4eOmQWp9ehIn5f
V1hkBwk0WNSlk8B5Inyi91mhWwYGZ4Z0wzu3LPevEkACyRyD0uI6jNrPEqwyKS20
V+GXHllZgAEN8YnQTDRlhFbdJ1f/irZPaOOws8RRF1LO7oMwjZ5D3qCFxQ3pV88S
EmJHQ9mcwqeTOUVQsfORGz/VY882etNTZNEQp5H4QuDf7fKBDnn5ZABiQvPetwFb
y9MTgaAnTDbl/KPMo7ZRb+ItF1ZWGLFp5bplt7jDAP8loWcXOOQZ4/gadCcDnqet
kdOOUGp0LeF89Dnk0oyKoMz7k/K0elRd1ES5PrZxDsxJs7qngFbjHu7XlUli6MKk
PLqKxsZH4kiqzKx9XbE+yyS/LJNS3t9+Ils6gVoEMxQQTRIawV0S19v3SMmDsYEv
aiseTSgJTxWIXtjWXIVsCLWQOMk7irV4T/1h5C3R4x7cgJzuoCjLEvlxOn59cRjB
yIqdY/IQ/VMbTkW4QPsHHTU/gS94rl2QE/EMElHJUdfoRWoV8WpvZCDQ84Qc7uve
5DyS81ZzoezQ4odNx10dDrKa9gqyB/3FdEymV7KChNNe0PcIgDiDwFPsRdmTohdN
HRf/q1aFKrHRikKCLtsyfQRdiiMHKYmvqh7gUGgMKKlGqFb/4lhEIs89FrdZVYHv
paK4XCYkv/rVgJt/n7AbcTMoSoH3aC+5VjZT8wfDzWOPRYmOijDB1oPn+DgBr6Iy
ieRzG8JHsUBYWIjKR0PyaJ7fYcB45PVliMClvM9N+WJNgETTJT80/AjoSLk8Lrfz
fd3tILJGOj5l81/5r4cj+15TJ8Un9e6/4zA1ooKMqLlo2HxjFyomE/wjfyOAbEwO
+LK86vNkTZM3nfWCF6b7crKlIWGP/xOHpDlks4a9U4p2QRjc8rUKL/37IkxWigT/
22l8IggPGAWVvn2cj2nv7KP7YmBSlwwi7EqaLkp1Ui7Ef6CIvIehJb5lp7H555ho
zCgpJOTRWjdGtGGMJ5tXdiwHc1BooBFc+mrh269SdTLHN4tbISQPSlgJl/8hnHZZ
Dfm+m7EQSz6Vlmc240yebqDTnvB9LZEEd5/4StkXUosYTV+NMl/I0qXhsWunrJxb
hVi3TwXKe3AdPxG5Ur23SDgJSCyFnynMDVdRd9OIgLsWxGxaHfPtQDRNaWHcJUE8
8n0den/Vn7v5oHHxRqmOAVzrKuO3U7qa34jcC730KGa0hEcwOpE0BWlAId9JeWZ9
sbdtXcASRcg9PtrxcxD7g1fAZ09ZWMxv2Vl3YdG6xRwmoRNFwvkalmupVEupGFmg
L3sZrS/zZkKi1whGvfAauyYIt9+v2/pArwcHP9EEaP//LI88QE4wyP2j4FYJxnTx
QIgSffEb4PLBL1O5HDkfKToCcSV9sjp0FDOCYfQKmaPfbvTvRcBGrREv9K9OFMI/
S6IguCBHhuZFSEhy8EqS6RFrdnjdvCnf4h11saeaguBtAf7h/baJ0hlwDTd7QdxQ
IP5W9ai7iUDTpIjlIK6J46G3QjbpSlRAAxcnwi2H3OPDfFdc83nsoWCOun566pQa
Sy9jc1GBdW7LnT0+SWnvuf+31mvfUnz+f5BoSowCOCWPNz1bDeZJ/HCx3EAXad7p
i6mQ1+imlrOgkum9Y4QoiU1AakmNG+atWSBYPFgCLfNhCuagfRUgG0hLnq9CnP+i
5I4rLzj81Utzp2LPUEd7zuD8XWxvZERuQY4UVTMT71/PQE+N3t+k5zmUVh/yExmS
iXD9ayzpvLzGZnRajoTv8WZGV/oFNPfQC5IsGcOL2xfNOa07ms9DFpWbF7ZSxXXj
bhW/yHyE9hf5pTUcdquJzZCwglHmI+2ZGGI8s4EbgTP2rot7LL8mqCc/LXvafAKO
2PWr9WTaKNgzk0c6PhicmefqEA/HhVqaMhJ6+IKoTPJu8/tQmWsuuwBUIveV4fQg
eJzz1Ab+4LNM5SO1o8GQ+GpvQ9tvf27ynKgra6qpBQzBeCtGKkoqxYVcYnvTzx2R
K2T5ZjbKPNrxvWHjoRrJzNvFGns3UkUt3lop7HHizt78c1I5yFbMix1d8ahbmeq7
8aZH12gpSS9Fg+TdaEAuhj+VIOddK2z9imvNUanYl1GJIMTfPuITasMALzGapz8f
DGwElxt57T6Lois7ClpNcFgxmhgrX6sVKzlxGesFiWJ1SIGRHha+qseumqszNP9/
LSZxqg/8R1YcOjS5h7/FD0sveCeoQL597bZUT27FYE445TMVna+wMIghiei77QMx
BQTwCPzktaFjRPMksW68l37F5F/60UMmD4iFJy8Lb/lm+zJE1HQ3SKl6DkaHybnW
HxKtZ3VM/l2BVOAddSWOTQiwUTTJGDcOuzg3CWeKSKTPDbxJA8BZHZPSBzAiJCUX
Za8gKIB19JSSmvzDQv35sNEfgCqQJcoUOhbJ/IJCx0pkloAl9L37Pc/myqxGOT6C
6lJ/ij2PZI7YqisbT/OJZWpIEQHCfiKDnOqFHzGiJRxdrCxalZOFEWtVD4m/5UEc
dFK9ZFI4cB+pogeRz0E3n1oTBKyPjLVDvP0AZSHbHHILCeG4iHSpFpmahal7BNVf
2mGYLH7ttjtjepILS/hIcLIbaELOiijoovTf5o6dumlbTXXyGK8ZiccCalzLTXxj
45J6tIVzWq62NVpXA2xlz20Jy1Hxip4ASiRCOsLu231SPqKMlf3IOTbff+qXM/Yn
exA4imgUeQ6O78VEUBo1FCZzW0U/oKK6xJCz9yXlj36yUzc8BReymRuVZdfjtleK
bcro26grmN4Y3feVZ/s3s2ySy6yOR5nPjlLzzqnJiInilsboR0TllpjPaRPl3tMQ
jx+Xg/zD6szkPruqTpXoH7ktT/V9SwbtmWRd+0AGTCPw5lz3LlLGK7m6VrkMk+VP
v/KvwofL0nY3S5DtWlr/8LCm5kzuCrb0MHOEsKlNdXJ72M3CAd1an+4XKfrTN0Qo
z0xeZqcQ8NxfiPZeJEhHn8tuQT1pItAWBQzini0L0NpT1Dc2Y+yZAuq6GwNNK8dV
G5fmuWqHIGOURnEq8dUv4pkwzetiHAz7oaXXL7PrxrkIXMfMkLBYifWD7IOYJ+8T
epGPgIx+RiK1xtd+jKjMUt69GRn6lfXzljbvC/vWXdfFOPWb14JMCplxk2HMyCrX
J6qpaIw+SSUAlUM4VgbRz9rItf6MKk8B9eRVr9POuqoOcTswHukxnED5pdCuOSlm
RHW9sji6RaYYl8tVnPQ0JRbykfAS7C9MwRwN72iEjmOcfAC3IJSyTGm2Xw+3tRgr
z11JSIvzwC5DI64WxFA5jqsBKcUu3H0HRqzeEodL+iA90Ub95y29ESZIUJzwnbBX
xguOcfAa1bRmPoGilsgnVt1yyLIvr9wqZ0vVP1TQTunAHjt2ZUu8GRjFoBZcKP09
NvdQZtTMeW2KF5PPEZfYRA4C5MZOvSRzxESWZlNeebiG4RmjwCHxPGhJoINRFvrf
mbeHsVQI8qnaobeUbi1UJWSxyAF1kdoN6U9yElt0lvFVbNtSx6/anu5Duvn/tRRB
ddAY6mNoF4y2aLL8eJSuTsm1xbiWts4xZT0F7L1yERgP+s5kH+DIy69AoluwSg8H
8gtEST0m5l+EnVMSQBuKBqyTFjqZDpcAqK8aI/Rl/4emalrOZKMS8s+Rbt7A9rvY
baIFqBFi4eNvUmjqnAwcVMUjU9FRN7MyM1QQKut+MWl0ST6JBX6mlHOmEmdMdCLd
Ib5p5BsITsxu+QbRtxbPVkUZNr4K2ZJU/sjtx1m3fKjyQBNNNQaJfiOcTpjv7Fji
JQCkwNKt8ie6RtKKp0arP4s5oMiInu3eyGjFJPF2oPszYnB2J1B6Jhkj/N+qrMz1
nMdFBoGzLq2ZnCjGmFMkNMm2pFEFZtj026oGtYnbwcjA3UmqoUrE6MNDn9NmSYKi
ezx32fmDEv4bep/wP1hwGWMl2XIp7u6dUKNEz9C6fvSvFAXX0pTrdV2zywGsulyZ
w/Vj2ty78aMhWtjkRkwSTvVm0JAD+ruRdKr3EyOW32zac9GvM5hjtYa/mCJDC3g1
B9bVlHdQUhrj8jMcslHA1s1laeWQveQqowhixmjQtXk+Em3EtDR7oopfwibuNJBo
dDd67FU8Ot9mqKvm9znxv6L8hO+0kMyawLX0Qc9hBfjSc23azrEetc7ntMvplHfu
z4ldD4mJgNtd3Ue90N80zoDEgZ21TFXp2PAHIibEfF1aKFVLRGq/KgtkSFebxSk4
rhrKtZiBwmGh67KF8gcxzuLuTwbEVaaNyRrib/Uw2F2UVQdqUVWEg5Sfa7veCeoq
cjfSEGzE4Q9SpH0gTJ8aDXtFaYLkyQ5NgKo3OWTFI1FB6Y8YBlIQxtu/zAGZbzDm
k9gtchZ78LUmU9uOOqisMLG7UyiO46YoHqVrWygJRBkVJhi3jKuuI2yBm0HOVGgk
YakcdUKN97aRO3Ll5QhbdvUCgO6LqJf5KPXOoPQEKGOiC5rg5aypQAq3GVAX+rGZ
ontVOF63fn4s1uqbUbjt6rYZE9F65L5+v8lmkUdS/p7nd7R+Au3zfp2rX9ccL0zA
FTbSoaO9XA2h0yOkMzny0Pk7eGzaL6z2NY88uFEcx27E7ZfQjDdqEYGphgcA2Pq8
Faf4wYZkVAmnrhOKhM4VUduE9wGA+c1sCo0U2MYfcgDH0Z6cyFKRzPsA1lXN0WMm
TgURfCcv/uLHnNzRMamPo3iW6Gv7hoShCoKg+YXsYaFIHjV+tGPLKBUklhjoH/n7
1ojEs7bsH/bWRnXfway0a1WCOr4knWcidwDSp/t32Wvr5zElbTTTG0XxbeaybsOF
zl7+IiN4GApaw6bvCRux2ksUVjdjC+OnIV9u/s15ffbaOQQyBjYalWGlZPXZyyh1
vRCOWF1s3h4LiW2st1QOWdWEVtdZduKfZh9OYxPcdehyXa6ezjow3x85JuFteBg3
O620LFJbUD8pxaFo5I7+3tka7f9q4qW+lOREpAAh3rBdgMr7VjrivctYV0h/kG4Q
c7Q6NWH57vPUo3b3fxM6PRYhngm1Gwko0eLAqS77nm41JFOKB3GccV7RK4w7Bts5
OLzorS/nrrMj48eFua1n3pdbToVk2gyN8Z95qhsMl001A0K1ERW1SnrI/21gRF+9
CAh+jdHb6/rMslsUPkVUTxaJ1B3r8S1Lwyhu+D9vSEK6ObiyGKQbpEoX8Y8tpmZ9
/z9TiuTHrZbT5kDIrbS66FMr4lPBNPfSZH6MIFw5Lbld9t0xYdhQseHlnXW7rmFR
FLVmwSD0MA6U5yg1xg9D1DqAfCGYju0kRK4Wk4+XBQghz8IbUnsAwMaN1NEn5JRM
1W3T8UNHD3rPO2c1zfgIeSVhkT4AZE+9eoIgFv/gQclAHFG3djeYjIzecTfGWazw
Q6aYq+IoE3ykddYbvlE67gcmIeBuitQJmxk8SCPvuF+vEkO+31xNujqsEsN2/tHJ
dqqV21vz2EK2txc9llWY8ofbSysSFq5ys6oK95XeJb62orbFQCtwbqZZoroufbDX
wdN0PDCgimSn6kUSjg9ZvYzsveMDNvtFXZyrUSUDeDBjbGGuNe0+liKXt2kvSHGn
SNX9n9zxKa3ZAUu4SBwaMuxuBejFQ/xgR5f0zENxc6LmS6jtCedbIy6iam/Eg/fd
eblPVJumr2vGjUzyoFHunL0QPRzqKTfQIFbssDi7PKW7ylm/mqG/GdxE4MilwjFg
TKbbu6WOoyuSOqMZKiLyopFQYNYFOBuRZFmk1DOpxpoZY4Ih3S+W9N9mvonCRz6Z
DQicJAKCCoWbsbapQzD4yoeE8KvOm16Thh2b1VR4dyNegSCcdBwuIBvgTqzeDqJo
7A0u91n0bxD9kMInPr37STRR1qFUm4+24KrHP4Z0bCQA7lnAkxh1M3zrPi+Hk+++
l/lOw/GhGr0+Qp0F7DLACPHi+lIZtmPXOb5Nt+DT4RLV8pEZc2VPwCtQolmOCqXS
/w8+6XBI+UTpJh6Bm5Fs9u5eRhtW5HaKwmAbfgQj9sWh6N0MeN9Wm6OYtyZeYdhr
Rqawu9wYrSJAcz+Hu+uTM+LAr/ob+bQZ1B/5Mq0ge/wCj1Q7XZuiV8SqMrVx0df9
enuizP4reqKf64F5JPd/85L8hYwRAr4lYsppF04yObwrWPtvT+HYPidsz0BEcXFP
Bw424i3x310XpdvG74JlGK5qNOiEXCb2RtQgjmxUk6OSW21PNQ5JH5ub59yR7g2Q
Jm5YPoaliS3P5VWYuwcgK8snZZkMj9H+ayQluKMo4sekaYpG3OPNi16vWByM3CpE
phKw8R2wVGlSDd3YDw3eRHkw5e/bwG8fzt+05NMrPf3cpDWK/OnpQGzIXvedjBgy
4/TkcrQ38L8BjIGDmKSpGSQiWY1cVvIEHQgO7oFqXBt52S+OjfzE8zzyqQTJ8FCf
4v+nyM6wsl31cs5nLfll3yxrgajbUdFJVFlSoPpVYYa1Gq7tWpnFZ2o3u1GtAEQH
uezClon/ERrAoDNVnDQCjx3xQQXMUEISEFqrvR9IwcPZiNB1SbaA3WiaOxyDhUz9
NKpXItCJAPL5iFU3FSw1uH2dgQbCUkVNo5DU0RNozebaIjj0L1C6E3+DrIeZlgcl
8cxRDYaOGdqWoy48AXKzXqljcSL4pKKUjViwMl67NiKRd6q0nMn2bxllSdBYVYVR
+dtClF2Lef9h5Fz+U0+DR9Sydou86fakvNqajKpa7HKzElM1LsgMYE/e7iQGRtNU
+ri+3cXkQhkjU6VgUTvtWbj8CpD7lec1otO6uqKbTdlhOi8RLNasrSz9M7hafHNT
beCaBud04VlHuyFc/XHXReXq9vejUqAq9Fj6tU9A8aeeJ6DR0TTSJJrKoSEpOHug
rhm9MJ8MJmGHmt3sCL5A+ya8UD4vp5KkA5H8hcZSPBT0JL3nBw0/ARWixBZ11C/y
8W/pE6lox6gMvB1hOj3lSmlzuBwlOwedQnTL2huCg0E+GmLc656E2JTJWDzN4Bm1
staC7a+eiBgxbbnnD/nCwGLRrhIaYgeAnCYjjEmwJWyN0Nc6yakqwqsO8016TIvV
KNl8K3qdb/vX+aE04wKRo2Pemqjl1LZnzzEO5q4SXSz1MTonduM+2iYL2BwPkWL0
BeFbQaDkdDoZfVczA1vHsZ7sbO2VCM/k+VEXpE2xEI1P77XS+nMxHpzWTyXQ1yD2
KBSg0bqW1/tkbIcZB++2IBXIr2Lg6dx8n+8rEm48S3Ewz718fgZtR9XQDB1wj6QA
rtROHTrd6G9CP9ULjonAC+VvglVvW6mFX2aMEbjwSsFVVXh/ADhmHgol8eHzLFvc
Ab7lLsrjLohtRyuXmN5UrXeTnAuKYpU4I4Q1MBSrMamBLlGz1eZRYucn5akmw3G1
eO4tzJDmeqqaKvSQr90zWGV16zxMpsCbm9PCgzIds+XjAAbYpl8/Ma7kEZUwyLzx
12nfQLsVr9qXFCGzJ4d7D6/eqb7Ao3nO0OCLgdgeI5sWM9Qy7vX5sWSXsD8XzLC2
NJa+FkXVdUflcAh3bM8PhqRGSe906o5ot7FdopVl/2NBDawcz3UnE5SjJs/Hjak8
Do0BJU3uTzaphOMnf8quAV5nYODPVOfdn7g4T2eGJoErjXPh4cTThDG2hVcNwWF9
ESkI3aTnklUR8XzYpUW5noUR3+wR0NYOQeT6uzO6EKuCJGMDaOkiEk+FkhS3lYZ4
1xeZENREXkqHmTJ6z8Ul2ElZIkXPLniRsklvvcDKNRuyrFcIAoXSeA23uuZm1cVu
D50NocMcpJmFqFSKBgWuwigapFkERcRDRPguyjJirfmpmFRyvrIg9oP7Fe7tB1ON
eP/rDY3lO/TRL3fq6WRptvwYF/syRYxr/iOjSM6gehzcyPjL4LBZodZarqlRiHOf
3Kg5BpTIx256JQNViRY69iKrgpaRDhMmeEG9prV1TRfOYOzINxTrqNZzgSOGM5jd
GPhltvPpzsVewSt71Wmij0+40tJJaC96PrdbeoRvF7A2IppxoO1YfZOV0sl4yAwt
nPm6xON1D9RAEZmqXjy1lQGoMiE/5YNKbfuY4qjWrg1tu4YPYsh3AylPh+cgiBpE
CyYbICFzl5V9DgzadXd8awDT8r2c/MrO03cORDhdFyWBPdPossTbW0Mv8uM/9jz8
cks8NWl+GY9BlMNcGvBemyKDhRDiOUzwUU/8Be+axmdU9dBzTfdGy1Eb6TYD22Z2
ekmmzqpfV86RncKMEJMehSOzqwpZUP6VPhLuHNpqjNQKNT8zIJFTKc35TzKlrCv1
7lXlljQBK4GRP9IkHqfP7Oxul659uUnBmZ4JiT1iZN1ywWA4Lz6CJX5ewaWUFqJx
gOpwCQdgUAVMMy9LXq0z8nDEphR0v9MNXytQPNuv8ZbJkcoKjA8g0kOA28GtMzDZ
ghbitQcZepckkY8i5gqdVmaFGC7WwjcdsElj6Ep2hfN4BzA41+3ebKnpDmXlf7CG
zDmeIVQ0ACawxpjFcOuuKSTEYUugt+mHqhrZqpmZWMpi2Yy3VKwPvsNmvcN2zRt9
Y2qXTJW30ePJokdN4aEn2zMYThHAcDuu8D/2db1ImnKjp95iL+2tSXCn5I5PsNDd
6K0O+dUm1XYeJpxel7rPaUCA2uckxMuvlW0fynddzPp6iVSnwDHBhtefMO0+BYCq
h4Tew/fbexi15tgxzW7owTtgOAOlLxqqGhfBzmQjW5TWMccn2ZKaGHUinOZFQOjj
6Pugl3cJTk0Tm9hDlAxjOHJNzav69Af6pTnErp+Yp7mnBWsiioQXygU92aRuQXrN
iwCqfUHPay4MPAaIcts7pc1Zuh4HaGLTEZ6G07C9Yan3JVn6e8r++5w8d047h8Yi
9dO7HkaE/ugaxqfG/axAtKwkaWmEEbNOHxaF89HGxTZeGKlK0/T8DzXykKpe+4Dp
TVEfjFqWLncogdZEsqYLTyiNuDrq7e/8DvOs4aqzI0RHWoMnw2Xsg5PYiajvtA7P
eNP/kDoRPkbgd88brpFmOgCgA5meU63+mon24bp2DmicMh5mBmknCKRRcuap4J02
g1Qusfk/y1Nu4xbdB3cUI1B57DJPT6vCrpIXsFENACK4iphtuL0oVAnEqNSd2aR/
90Y5Xc1yq1RjhmlhDkgPlyhuHK0YE9kv//QoztAd+6e8YuGw3pi7IiaBgzTR61dQ
BWBFWg5y1xP1jRwZE/lmWwnVfIu4GQ9z7BnDE2adfgEqghdK16pr5ceB00BJuXAk
eMUwvHsvo2HyyuBkekX4Q39cfx/7KKijhs4+OMGrJxRmGpzHGehktX8VfobkFzdo
CypNgn8GZvFB7vMSMbl6UT3Iofg1zsVjLHGxj06gnSrXOZ7pZtppivP2yCK8ImRs
RggcYW2lXZxMcNRRpgTEqVNAsYoeFWLrp+46sCdPQkUVm+OapxISL6E2boW+m8aR
xkY1j683GDLy7CJTULRvhd3MZY5p0ap9QR75pcBTDs3s5KK8FTSI7k3VITX6zLZ8
mGj/sJcBkfw0XfhH60EqOIkJOVX5vmdStDKsoGgJji0J2qw3doU0ziYDcU7NoCnd
99tP5ByCOPxT2b2rxPO1KWmfJDhq30htGiAiftQI2az21Fhu8ZD4vQdRj5PP5uG7
vWaL+eJhp+a9KBTWjqs1b+ZK4T8/HwMEosmNrgz4GUW/mT/hYyOrScjq4Tc1bpqB
b9jKiYjZW6So2fx+WzH2/E9v3qRqhypvHZ/4YN1p0r8yMVwQHcsRIPyAMGvEoEBy
b3ULIvr4PK9dCFHSmq6txfhZ2TWM+dZDeDkvHr1Gs/nBMpNbMvil0OlFXoj1k3Jh
UJmwdYSHxtoQha0rSaTZUE7wp2nC4bR9dtmRAKxFASsO2UCL0WC26/If1kONBatA
ojQqOXBuoggrsebpmdI6bdfOCxVxxfxLH3FJ0/5qqiyIgjWZB244Hp1Fyu7CduFk
Vwfz7NuGyJTRz4TEt95U+vrZeEw9YPWiNXIR6dsRwSCaX7ikvG+6Z96OX04jhNfL
07xRc6H0CGQMMJqz+Ut1/3BTqS6zkuccJfbp7mxHDLS5poXcruibzpNrxN8YPnzg
W4SPnpy+q/MXOVdUYJMtwIZa0gmFMp9fQ7wgVZBj1JzX4ZL+BzUGY29Eyzxmi07w
lnFBr1G3BHloFGIylKeJlXxIq+LO4TsmCNhJYYe1zEm8cXFU9rZbov4SXIMKMWZ+
TgVQozWpAamPtNP4cuJKAKjZEXNbgGNl6Bft/3Avz8170V0FPLe83BZA5/bXJ7QU
I88ex1F7cMO1RWtzErzb+vPmVFCgNbRc2oWE7VUT7iwYM6Paq9p/pXBl4vAUqi0Z
8q0M3sY2TjU9x9AW+p5XyOmKwa9wqIxpc4R7ftsb+IlRCwCbOlCySGxznhEJqEpV
X+O/4r15wNDywUphT9f1d+H1kBEhD4BaNUQUG3hwyEyhxkDVF+JbizddNV2qdvva
0yyofWLfFHygUzar2AyAUyomlXCUCNFCbqWfruK1B7Jt6KwGCuc7B3N3/8BNWyCi
9aepkGxBTlE355DgYTFMLpNY19j5OK6kN07JTHReogXYKogpzs4yUMfwRP6g+AF6
lNXra7WIGAhGUU6PmBFnFxiwXzfzbfHCsh7SBlZf4jJY9LCi7Gc9IcHlXyQ1Ua6Z
mvJ9MVjplFoiAq19wRFqGi9G6tYcSVV3/WQPI1V1CbHkWIxgRmESCsb2LGSCxvhV
IhdywxeBtcd63f1fTp7JX4jd2jDVYLkMX4m3yefq/hkgm0enwZZVhTacaIbQ7DG4
yiWE8EypICdqFVoh/zcxEpChipQV60NujOnmXUsXnkZU6dIbQ8Wo817fSk7kCzZY
n+G8RH8IwcqfJ1m1PDGQnblONbI5+oAYoNigtg1PGRVbFig9pWTFxDFmUEZxh/Yc
CAQPthO6Nz6ZD1JGsWrBUKHJlj3z/okgJRIi96dUknoVFyhxNOz912I8jJyHDNv+
K9TkGBmrCaW4TLDFf4mCQtqR3UNcO+r+fkXJqJoAiPXlmedSKfzOFCOSDCs4hPYA
S78lE8NUgp6DiTcFdBuHW7sKgYGUmvqxvnk+fIAEx/y//394lSQYrBuXHjssBGVV
m9iG4WTl9oqcf+8A37k0TrsM8PYdeam+y6ujcZV+/3wiauSDyCVH45T+OQNriekY
bUpeOwjp5XJiAG4R4LLuvAuJaw8Yy3wvG/el3ihCzUlXgrcYijfC4HOKiG01Xr1G
YcZTOvfPPG+xQ9x+PwqWnWyPL9vt2i08c7LPB5vR6qTO0zeEdOcd0cCv39Igw891
T3gzBdVschYacg4Vqfzy29Ne9uwwJBTZIFVXtOcs2xgGWBDrZ9j3AY6DarI0rlUw
5eLjG6p0jD3QItL6BCfm88XLMSuIT7FdsnCiQlRn29K9HuzIttI4FjIp+cM1zNl/
8xFee7nyfxRUyb5wZ6Rh4addEP7pkJK8vfm8EZJHZ6pG4y6iRaVk4gvFSxDH388N
9ycQ5Ym9XqM/71HMskJUNomk9gzHRt3RzA/A/iiKd8+8pu0fTVmVZyv1mIOtIXi3
6O9DSD7utVoHqXM3ECoTdQ5IRy9iqryEQx/YjR7zmTpwbiwih6VzGJnxywhWEy14
eEDeIomxp5otjNUq8cYxUJsJJyrDGeLETphm5ltmX28groVmvIxmaLh6j9ZM4Dpc
MXJjLAKy8k9TY1UbwR5wDpSzYVcOM3kOWcy2AmR9+4ibULHWNXtbUTeOgBmzYoTf
mLRzLwPdjU0nW7LDhtJWT4T5LO8idTx3U/6PqhgSBv5VopjTG46WZbxvMjTBkQuW
Warqf0aS3Khg3mZxgC3bhlEGDaNqxmi9NMd4/LnvxL1lNc12OL/zrAMIeeWatmnF
smZURn6IaFls7zCSK97TmOoaNDKmL2hOq/j2zH3ceu+rM8uwQ2luMlI4fF2WpYZF
PBt95ROkUjiJPZV5+ALLQAPYbVXf9zZH8OxiNKY4JwKhB7su3NAmDsPD1QfEUTVo
98whTmAkrb9Mg5atTC0yAqIJoUYIeTWiUO75hjMHLnKhg0C/952JX92P6nkVxWzl
rFjNGJuZ2GSqwhzNnNqUEBdBfwY3Ny0ofgjGdfTdQxvckPJEJhKlQB5En1pDvR9Q
FbvBEIm4+dS2j1fi6KvBuEc8pmAV3jGJm+1OQwej3l/H0SmgR+f2VwtC705NcRZl
M2Qcgtz3nCiZ3tBydFulxlxMPJTeLzlltVBsQDCn4e+C7jAiMY6HRDGT9Cjz/leh
VfrYBiZ5MiiS53p/vtKTobMiGJgSlEF6vfCGjARFWwjVxQpbyvNBOq5VdOthnfFI
yjtiwmtcvtBoWcGRVSEIJM9c6tzK2D7pK4gQZzExzX6X3VxeR23AWmH7FGknhqzh
J4xAVVcWCg/o8GbnZZ3NVJIZdQjlm97+wFJWhkRlahUEYSQhfLa17dQ8kcdnAc1l
YCCS5yjzv7QGCQ0aRP4H5erqGg9EFKac33KaW3VDMeeaCnbPes07W716bzY9erNR
6T6hD4SU+qBkK2FjHyyXPLlxWEeSvEoDAcBxOlKzC/YQXacDwgcxjCVGsoTScC8B
7R4b9PYbTn/XyoM4axg+rsR4ycb5n9wLsYbu7YIUWHg33blcnbfKZFxpzeloGtfw
LPn1UHoKmwPFWHS/3weUp8p069gmPiiz4PFqybjryvakfLoWb460vnv4sgNPOrEy
XhfmvnPmf0WFMy2ldfuLoUb4e8hS3KRCLF0Nn4fBQF/qyEfoKIP9ngybj04FjxYJ
JJ/ELVRvE1LcgrD5aLTXe7Xrh2tzkA8/XGYo5ctPUUCTX2uKgB1DTphGXduT9gfS
ozk/rYAdWFHgLxWKKXn2JdkQxPZWSuh94ELtM/iiso39Vu5+V7BWloCdyyrZjMbV
LUEhhaz2TwFq5PNo2B546lBjPF4l6+HulMeglk+4pPCkdkQlG5UDMzrQBhVZ7/tg
yU7K8povRdp+Q3Hx/1vWv0XYi+aPyh7PnXTcTORtVCPGWJsGQLOIpat4OrE8SapN
GOxZGDOS2cVtSDNZLZqDtjDTuuSAgea5oB3HhF8jxN7touH5f32npQxaKFQJ9Rt1
2j/1pTg/5b7TtIM+hpitjQZiHJxCy+5mi+RU1yck6IMDLwENTrdltZUKNsEf02dA
Ojs+b5ZnfXTKIvw/IACocMhYdFVZKkzqc+LOqYWukqC4Y3yLD1DTQFusj7ioBVRX
Rk+0iR0Yg/KSmywKnheZl2Mqy0zXuePe2es6symqvrWU+VuSG75h4S7A7XMe2oRK
HN5SpxpAJ2NMfSfbnqXko85D9s0s+vS3cC/xilqbAwoSIfMbYgZB4VjrqGXQXjy9
IKRuH1HatvYWxCaP0ngNru67pzVXT/WXNSG2LbT8H9Cb8OFoS4zYgEkENnwc/b8v
BS0RxEGDSqcRAOxJYqALDA1Qa1KOjqHRBlNeDOjM1Q2PzXjK2LMvIhj14Ruo2mf9
buq/tvKRJH8o29BmgvIzaWm8zJoxDMp0l04NXIiZz5yewmRX3LTcKt7D3TRbX4gi
+3qAxOnrod4dUAOSpTI4QRHuT/FO1B1/02XDcSOGFAVCMTHUFBbYvAt7fmLPmqD9
tTj8HVV+GNUpXNBPlyfEGycZquYUqoVcuPgkXb7iZyTrSLEZFbWCFY8VSBDnRHxM
R3dGBVEqZDbiIsjHeHbSYdd2mMJthEdS/Uorl7ugDi3k0zv5EpqONVtr2f1Nd1Co
iCfgfAk1ckrk6kzueWEyOPHpo/DjdZ8J2bqK5DefPc8Q4/YPutCb57kNgxv3FhsR
cdsDroZ5rrToEzBpdwrM0MV0TQ7XZoi76N6hUbySBV1W9zzvCTg2iH+UmZxWmhAR
aiNNpvWcKfsSe1Y/4b432DbwFdUps78s515ip3DLPEeyYnxuiykCikHcXN6swOE9
YMyiqDll0wp0HruhGnpeT1pOhWIGnsh/20E9zn9czY3k3S77qfakCQjY6EqRZifv
XTsWAySJfzOoCi81McE1/KZRnSydTrWtwd+pKvtzNoAInvcTaYXq+99FUMcnyvfI
vDG0FUL8m1a2FIRVTY0k8P+7wTWF/dmNpXofH7tI23bE+Cqunk2CV7W0JFBgajQO
A8l4GNkfUwtjd7Ysc7UCHDMFMAvVfpwZZ8VJ0TsNq28RgJluTxBcNC8/ICjlKwrY
+QLyMhudGS/l7NMF3xjKjoO5cM23njNH0LS8fM9rG1uxX98lMW5+9gqh4iGSKk4i
i4VoazgeMzqAJhgMHf4w15IobX1s1XHOxKdtX7h5pvKivQJtQlt/l3Sg98Rhjtsz
chg5Wt3T/4gRFBxkQHaLikQRQHrlnY0/DGtAuEr4dWhPa74dDZac7qhtf54y5s8y
1Z0NzIlVNOD1Tly4iPHodszRQnXkBxRrrOYKe69g/ZccadvrH0nNzh3SyM/d0Sol
0TqcBWID+gQv02SM69eWg5UvRL+nGWCKLl6i/ISMbzddEpy4PM8fcllyYNqbYoSh
Jem27+exBGRGoge3ZHetZ2/FacuMTlBrkSpsBDX5nDsi8wxCcGNMzjIPHik9oVr2
5gyU6a9wPKPPViz0TrB3/lTjEwQUYIk/B6G5JVKxaVHkrD8sDAR6PoqL+f7owNP8
90V1RIK3V4K7dscGlNIH7WpN9UY4IiGKEcT6NcTZ/AFCb9U9VnzFhNZj4Q/39z5l
Ab7d+JFKoIsZjxbS+CageDKJlL4iQTy+sXCbtukwa7mOMBrLRdxwMBPYlS3InDI4
iylzqxzgkOy1y9/rlERo1KY2L7IkENQaK9koo/R4PT/mx3KPOalbrTqtf8SK4XJ7
fDAcaEOlzLkKFj3z8bOYpKY53kOzSZbV3FqrTIJ42BbGbAnLh7JFR6zUv/nqeQV5
9N83MocGA+xER4bjuFJlJO4IoUBTqtBWw5FO8Bt51xRJzVoc2Epck5yWDzu0A/FY
aDic6yTINvcP4FZMfhAlokJ00/UGYPpAgBfgyeAjTxrOPhHRo/jLdHtYnMa8YeIu
xcpjwzw0U5uYneXLXKxX5V2aaAlSZ/o4sT38bAYVamhu4alRC/ZzIuOqY29ZxBqA
Ig5cCPRv6CwIl9JNBz9u9Ic7Dcox1z0DsKc4ZMzWEVW8KTiakizA1vx5tJWAmNw4
AvmR7DAD00o4MqJTardDo+kGJDf2YJkE18fN5NyJQ+bi1iysclOGTHVUFc4fHArJ
7ut2AePn6roecBBp+7/07lhQfxVSlgc2LRW0rX+uEYzcTN19FpG/TiUVqrMvYEPA
FxrYHaMzKoxCyWaqzlNb4hQkoshq4Df5TcvbJAhXGk8YNZRA3YKJZYbDeTyRqS4F
U/8szVVX/9PBMlqhNuKf1GVwc7OeitEHkAJj26VVpW5ETdMLhGZIG914KXPRv1Ny
nIoZN+8/yvGhLKntK2c9wIQ1B2WaNJntZl/gk5zNAmjC6eUfQ1DCyFTwDqq2HwlR
UG47O1Yh6EOulcU+uQBylnDZlhFSSvVjgYBLk4HoJtGtcgbHJZWgRsf/e2Cyl6fr
dijT4eo6YmGA+YBvS20chi4fDVF0+xjUwkTjH3jOIv1vRG69ZTghAKZ1047X4yPK
8zn/JONEYNP6vgs1rccT09I/WDTKIq/4SEiDICEW6xBfhKI+6TlyGsFfb6RzaNNB
0hV1pv7jYn3DtQZXrjNuVAhoVuc982Os5PC8KLnyoNQLRg5/vsaFXlR0Iete7fbi
htm1l4XqKr0jab2N+B850dLkmDqNEAW0U4SsZx6anf1F5vfLwAATxKBTOzvga2wF
twbsdRXX/wGQ28e1JOkev8duwHZVn4jd9vVW+j/X5M9Y1OQbzdhTwuarzFrrlRrI
+9njpaRuFdwjhKXhnEtPeJ56/Yrb6DvK3pLvLuK5IrreiLStfWmwiplL6pzCKrbP
9ny8h7HlhubZ5bzCQfihlMQixLN9VzV7mBRRunp+EeXDU+nc6wIlwxdcd75uuEjY
OjWTGc4ttvncIOrIKIawM7mN/oiX16/8eFKAOIUShsfagx3v70jqP0Aj6k2s+8hg
wPZaQYuzYeZKtNdjVmEUPUlMgVh4Ork8lHjB8eaMrZvCaF33hnCGAxxmki6++0UL
URmd2ws3uWvzkmFvqgC3RuSQjNyrdkIv4NMtqKUBso1+KWX9DQ8Rs2PlRP6u/J1k
UDUxbG+CoB5U8PM4uvsaAU5Yod/rBenoQdiCYV7QPfDRcguwtTUP5nSyfRQMjxF2
+kfGPYgBnwa/BV0t8ULlsw2j9U5PYyBIrPbmCJ/iiiBkvh0uYFWcevuk1jCJYss8
XV7tWt6y8Sfnv4mHXRSFdnRbJxhbmG2srTsMtAD+eyvPdzkTg8xRsdS1nexQFvBm
rj7PLjmtp5EpWD62gc9R7PjW7wOjKV5xUyIx//6owavSyqo37idFUUzp3XdnXzeX
Jxsr0EoVk2jPsx2yBpuDFUY+gaxQfku4jSq7gPiFQKuMx/ez3dM+VMW3MT8TstdT
ghzHDP9dXuf/Sl+QQUibbp5UWatmE0+AdwuDMXGeHhldOU0bh92VwmCcO7vwUPMh
WFSG3ElxonSF43ZoPrdE4ufzZzbWUpgbWLEKe+WJdwc1z6frHvIN3xcZybw5H01T
JgQSmlT+UA7PK/+KSxz/PJQP+anmVDMp324Mck30cSgdSB2eFt1ETZSIQsrsk3Ox
4GxL/IXRZIedf454NgQAsZcJi2cMYpfyIpDwoL3OHbV9zrZU/JPoezxyZt+bDAm/
Io0K0ehUWl7vlEcGb4Jws9zF9B7FYYY9uqjlepKcQr8KOtjzNorp8zLO4sNbFPL9
otOkp5dPZARjj9x1zxiPH/jZTUFOons5GjjUf1xcR7gJn9wwok5km452pbXlPtcK
pf65yxk4oqaEZMk3NKYvVfx4RGDQrL5BIfqPOKWhcV55QGCLMBI5K8VABisvQ+/U
5DQ0v74CWXCL4AUilRa8kcV2tvdCI1aTOhvrSwNlwBfFIO/1N4RtPtvm2MZunaE4
9W9rcRoZOWAJm8c5/q1lI0VQKlN5bI2l8XxQHWXKFbpOiutJn8NRchq/IturAcDq
ymcz7V3KemYFihS8rCqszvnxqw8GzZoK1Ng4xU/shplPnSQGvMflnN+adN6g3Hh4
NTocHOhOXJXxzbp8I431ZV0vGscGOpCXadvRHPdvH3DQCYMoH70LUzZPIsRs6H2N
coCSeC6kcvNCW3UQIshESSfRuzrwW3AaELnImSXfkpHWkyvkFcwswz2E8l4aCgYw
bhnrZ7UyNPfDwQxjPmWYO4yUaCO+NYZH8uy3iumal8rESwvCYanHSSatIbfIk1f4
QVCCDSSM6UDaFM7fOQReZXB9qBKPR745/OjZ0dDAAABGksQ7xuI5xD+NBWFyFUq9
ZX8DjuP+I+VAXnpR4U2TZYZpn3qqv7hialj4p+8LERFRbmgl2k8Twwq+zr1yGZWi
3nMVg8EbDWr4RJ4z3Qz3f1inweBgEn3meRqXNMi+JYpzLZ/QbESS05S5WEFiLWIv
TQ7no+BgCi5C2kxdeg7J6waLs0V1hosY1l3TVv9+4mm0/Ma5gl9LX4MljimSFSsd
dH52Ky/JqPcVXsHYJL3VXTLXW4xUNitJrVVUlpSt1YDha6ouXY5X36hLxN4aoC63
YUneeSTU4iBiuzEmCqPxipB0PLxbQWHQZ/KcUC7bLqaeyaHf/05w68VRC2PtGl8F
DP/akEuYgCj1TPg/yYk0mTJcy0PWRs5f4avrVShDmj+xVdB8zlLEZZV8S7Z4+g7w
yqSnai+psmL2iFTFbDXUFS3+nj60TTH8eVH+TffqDFTgtgwwiFLtcKBl8IB7T6+Q
TuLnKiG/NMN3JE9XUBCsC2yaFAMtQvrHosA4iZt+rRUJOTge6Qz8gh3d9B21Jp07
mSJmrzyE1ghObTd3UeHDMiHZP0LxMP836WC+pb1DHqxnhAZQ4zdj8DrtFJShbSzr
8jzRH4JWXKTQDTO7BPJEXhSc0cMgCg1GIW0akzxA73RR/ljYk2zXCmXbzXrjxLGz
dnif+pRSedKMpB04ahcNCzKCoh8SQnQBzilGnnOK/l07enUiJvaBue+VnD41vrBl
6dmOIs7JNBw9CNGf+Az/bJdz0mlBk6gGd5etqqZ4O+LlC3bPNtAUZkK1W/PIYCTp
mAkJL2F6aJzBRhXchd5hTSukz0vEVgw7qp4XLgwFv1wjFmvV/tdIqO/6kyRIDXa9
dvTN2zFr8Cu7vi95eomHLrRGWBo128EHDBF0zh4GDiQcqehnZgdB7ZVQ8V7uaCtk
FoJntY+/z9d5jSv9sZSVXJOw/13G28A9EwfGB7gfyqhTXyuiRsRnbb7bGnmBwAYs
ob2UxV+eD3/GyXWuXXHcdyUi8BGzb4QhtYjh7+RQ97/NWUogGbAxLTJByPjxS2W6
FCV5Nr0KBkUC/gqGIGYPDYAuMo62c+hGhbziNo6fCGt51LaO/7Ln00w3mfPmM+QN
SLJmiQI2ArZk0k2c/8rMzaJoxfMx+RAAzYIYmsA7O+2hvxvJmZMWpR3/wFFuZUm9
Ee12Nig9ksu7dke2aGPL618Id4oQBPbPh+P03wG6pXz0fc/Bu5WnvctcMrKyvFHw
yTjM3uutT5vtpBgFoR9HBQ9V2cyWelwJaYXV63yLWT+iuY0N7OZOIoSvJ9NCF+n4
ugqjVJUH6RFnODotiY+AGxF/NHeTLjw+OIiHD/ewptGhC8ntnVji2btbcnoSl1sZ
6K813CrhjsaUBL74WpiqnlgyjhZDIZkzredvStzksLjOjSF/YG7gUKU/mbyYn1/U
12lBt/lDIxhq2bTCN6bq/34+M3eeCy4MNY2PHObxwU4tS2G9Jvmm4kojh0Uksii9
C9VfHKlNw3BsNTQjMCROXTzkW1hc5JBfvPRi/S5vZoPQJKjfNoy1c1eHB3lB3gGK
IjTAF2/RA7KinUFQ9AyBJ/8zcGgIOGPucJKSknMjqmSmGGi7eHxkcpXKfquAJ0m5
YlFI8RfibRlV5xA07+1hy8c6Nw67pdKPwhRsQptewT4sG4TYZ+JdH+UYCD1TbLub
lSlr1haT0SDkgIs8bFVCvJ7u1CtQ0pV5aCxQMdfU/UfGNrZXK9VuxTNjenr1WlbV
p2vcZ0vAB8BZMA377h7R7EBCOww2J2bdpOpnY211u6YHIt1yuxDzbGlozBSYMK4s
WjjSTu86p+ioeIjpP0RHHWAROy6tTo9QnfQRwAsZMKbQbrjX8mAZu9T+Pr5+PBD6
KTZ93ovfN0OGf7h724CUvreKb5mfO9OOGqS2vP6ndzGZwAAegA3oXnpWvWJfwEka
qPR32WXtF0p9Ks6j9n1ZaMId4loVGjeQNXh/sdLrT2GPqttEODJuviydaqRTgMlV
bb+fxFFmFRm/rwD9Juj7OAnu8UVZHOaHfqGhvTTn1u1Le+uNC7FsAM9b9hHBwf00
lEzXg3sHKDUR0KCD/JfMWxjSRhmGFwG3D4eLJmpJhP8AS3abqTxlSuLIr81SdIrB
oxioGcQuOuovc3z6X8UHFs3EkR7I/AvAv7a6+wmImm5n/QlgFt8f+XgrezTPPpQh
Cuc5xEmDyuF4KXztHyxCDLwCI/czCn0biV0ECJK23STiZr1MW7sqtp8G8fkQZuhe
bvOfWRgPVwFZ4mZ4yVNYKinXbHu/6fwfLprcFioC35Qxvk/5Sd1Ca8bGDx6R18y+
+swBjXTMecnp3F+Pt+kpj3bdPuBPUR3HnmsZI5tHc3htPMhoQmBAfVl3yUvvvyTy
jpvXaC54iCAMeml/qLLdvgyEw8vbbm1Sjl3+eawE8MssAtGTFADwQDLhrJLvsSir
AY2QO1fa+xZpq+cID6rR3si1dkd4YV7dPL66WKzQnDgiUQtYG68kZZOjzbw+2tBU
o1COo/FLFCTATGsLXXTKmzvtroq/TMeoKRf+JkkSXzhcXkzhHZuc3V1s1lcP7l8v
JDteTkvtNcs5Yc7zmITwGo0udFXKIIRApCcYuQ8GCMBbE29wuUiOlntRmQ33va4e
FZmSHJ29YCXbH6tUYV66JPCzvnIvcCaMqjLFXgL7Qaj0KQdOqzVBnyjvakVu13B8
8Nt0XJWpvT3ri5jD0IrjH8Z/YAHtzvbsCuDWB3/auZCzvvBeoj/pUcqPQmNAko2+
mQjlLxm5O/QoMhUwtBZBjGWY7HdIcZGc1TuIFTfb8qGOMkJRKLaAFK3Zt0HieuGu
paCX+OJNiYzuD3dBdiVJBnocATKc4IDysNUFLUw/W8rD48k20vPFev25F8B0kBLN
uFkG4XQwHxQQ9NpTgg7Imvl9w4CBbZk7yE4DbZYmoDmFYi3psWIf7AwgXpdXAxYC
zS20El7VGLObaYttYk1r3lbwMYPzvVeCrRgubOrEZXsBWhnosCavgD1r9WVX97QN
CxyMVm/v71NFlshNsiwlJ5WDpGSHQrQkOTg232vv9SMl4kIllARVTEMX9v34fY6c
Jzw+YP/RGyHLf92WEcoAEH2zNbB3hBznzFIqh+CrjMw/w+Jf7xV6MaUXNEy7bsN/
H5l7EnSLMP7GIx73X0pbpV73I83nta8XtO7qEOLOYOXSiLFO4oYEEtgTLWpva6er
Mcki5wkwuDL4xOyCS4Up0VqIq2KxBFMvQXP55k/0OVuX/wT5AUMr8WIL2QRCQJH+
Q2R83wnE7dZaQvLI0r6Qvksvzc6w+up2y0XROMZjhzeeH0kDCStas2nkO913qmFH
GyQgZrkCyOfup+35/RjmUozq2hghdZR5miECQ6SOcut2H+fShzrgddX/4/qjetvQ
qMk0NyodhAq2ZZNY7Uz3QyXy6wD3+LtCQueUaoL+HlHAiVVhKyWIi5B3yEv+TnwV
DVKbrcANBC4+l/VmRyprMIzkWjAuTeDsHissAgrGHLyNdMxsc/z3Hf65TszCKpcg
jT+ugRsHzb9bFakg5TiVgTPLFW2mxxaC8y0XhsH5p9TNsy6QWrA8UY6u5tbidGB/
1FVziceknIVmHvvsbaFKG9e5Oxls4gsPwGVBHpZptWs7uzRBvCVwg6Eii7ZVvwLV
mczRne53ye5gW5QH9Wdu1m/ZsLSimru3R11kY3n4QAYH/Vk4R/T5a0FjDOu+K4jy
XUpOvh33698FJAhzn7ZLHozEQfOeP/NGE2FimtBSkSV2+PTppdnv1B5g4XLDv01B
v0CLakmPkOeFY8LfX9V9xBOkjAWZgLzJEdQ/Mo+wvn1VEDhiRO9KPKRqia+8FE7Q
nbAKeQ3W9Aqih6tu8Yqw/BrxbRzQ7Qi1C+i6OABrC1xODXjzOk7lagINIZdb590c
yIEjjsHYHm53owCnyIibHDPvIaxoCQ+wm+JIrYeKZMNcvzr8vq6H+HptS9cNlPTj
gQK9XAr3GcsD3UdA0fSaLQ8ojjGZLaHmCaEsKUjMVg4rTZafAEJefraCKlNSKSWU
32Rk1Lu/NVfqWJ6yFrU66uO02b/XhVOScxG2XGX13B+JCyK+3kwBVD6vyIMbDXvY
//0t93vfUJQTiNBe/Q4aTzHn5SDfuTdXHa5lyALZ0NZszywtybgUhSAkbmSMeB9Q
LnnQxMoPNXUFNvrqXSnEMt50YPYmOhJftgrEh8LGPqi2UGfsz8dcYCyXW2TYSxES
HxKP4utmu2OAWMIQuIkIHGJSoIP4sePH9+z/hAWmWt+De2fIiju5SqseViVJUWMm
mFrl9ZgL2twSgHf3IGoAcSL3zsGyoZe1nrswLoxApXajq07j9dr9m04XDSy29WmX
neu0WJLhUhSBWrKLMEZenNmBV0UV7z/ttie7jisNv9wIS2BcuNM0DW92XGSIMMzI
wcFAoGYbn9Ed1hv/Zy8o9zD17oU78dVOt+mwDVkCRwf1iibGPn7z92q7s8fzZ50e
y4OWJz6BkfmtTvlCBwvxKu0QpSN1bik+BiziHAtya4uvViw4CY6Pg/1k67l0iHRm
C+hYtDWrHUYyPBpAD6BoQa6a3zXlxMJCUADhNm0XW632/O4U3GXr8SlVrHR195p1
xJBZZtM3Kis7Ta/ZJ+uYm5zZIuY3Y3O/8Jfa3wYlNupZb1EEyro+6uVtPWpYD/8j
hrghKmigK8ALVCUN0njm33EvkSj5pg0/W/jY9+NUYHNts/tuRJxRBaP/6o41H9YC
PE4aV9TOyS+TLLi72x7SrR/pve8ct4parwcqmu6+pq+l1aQwr22iv4px40RRMTFY
hwh8NALmSyf/FfeIpjdATlrpT9sPcpgsh/0XX0KlmS6bMa+vGEYq3do+QCILj1A0
plHDAQZ8tYPntp7eDeEMliDP8PLxK8iHamj2aTpEVRm+Nt9kTASVpFUTsy8wk/lK
53b0lKdbxDVKU1Iti/VJcMdugQtPRSCFXkHvX8AlbYAwgYwB1Sg46WnrAK/xKQWj
gOhI4Tgwjwx7d+rE5wkwQ58Lie8uv6l+uDGZSkuqaRBDcm4RKM6R2zJ2WsdbSJ6C
WLW0kBOywZOTgztJ8TH9sTSDC0UzJHjDnRQr6jHNThksLnovaRAiCjjk6xqd6nUq
YuTTPoKYpgEM/FFue9nQjNm2I0ArgvBzA6irrSqEiUbSeGnZFlyEBw6u8jTx82Z1
+xoXwpnv74Q9UkMNvbbElMGqtpXn+ZowOnMfLNyocv70T08zDzpJkY7Lqox17LOQ
UCNMts5gdv5F8OnWFUP5as4zIjio6wBWemHbgnBAvlg2VJh3RzXhOvOOwdh0ZVJa
jqRDhjxoxFzInfT7dvnAkXv/oKQPSNIj//MLBVsBgAC310kHrn3LkgRoMDZnSBzo
XsxUZsSjGajT65rxdN5KEdZcfi2IzgFRNCFX4nmG6binfYTtriVONAqsQKtUOy62
zf7dIDwLYQpTfHx22WcDlht9XTiLORYnBfM+e11i/wEFRscA1J1Go2qJK1hUNnnC
lM5V9gEgOuBypAgHRVyGYvEYYamj1wvpORWWqdc61nBgstIrU1qiztS4bGjxoVWA
SE1MCwvK49pGOIPgLsAV2qzBzaTRVAghmcTMJOdy0gHJhHO+KfNp6Xh3kdgiIA+h
KKnVMoqQsOtY3YW34Xt/bIhelKmYPs3FpKPOsbLUjYQ9AykItSd5te5BnO3784Pr
QpZda9PixhfCMnqg01BBbpc/avsKw/Y7dQj9vOhxbuTkwrilg1ST8hcqf0vYYplh
Z2uneCsPxt0f4OIpngjernZ2+sK/bj5t0aA5IGc7Y55WTjLpc3+g4N63Dg04NEj+
YQKarSwaL89UYzj5pAm9GHIe8AvzVI+s9LTM7BY0RPE2VKM+d0FSgCG91MW3UhOG
cbZlNGyTSnsYou0gxTLaHTcLpOOmmLkX5eqdTZKyNNN18FQT30Rdy6Uzf4cyJBHJ
MQwOiEGeyQni6VmXeI8HelxJKB1CuR3VGiqh+13ioT+zcVCw0+qg90+6FXZJ9fIq
ZyPO4Cxv8ST6tYX25rzgCDFJHvJtUxN1Of8zl5RPmAJA6dnDYFJi2HaThT71Cn1X
1dKNJSvyOcHVf0rCFBrKRObVEDH7IXQXW7bLdE18312ZoyygCqpm04cYLTB095wB
lZvPzisTYhEntx4PkUKwKDwv59uhf+a6RRaBdttDEm0H33+4OPZz6ewNK0UEI+AV
M33NnCVZ9wy+ogRwww6ga+XHRCwPwUiVhJxIwbpkt9AzvbKGCgiJbxKMuW7jVugn
ZfdRKeXlRU9fzSax3qgdmmutIQ3bL+fbweRrrbn5+vLmD7vZEnrhk06IcdO+esLl
LryjcCN0PRXtBFKfcl7ChrAas5wBi6xN7Xuk1OnsdaZ67jw97I8gLDkquMmRbIXF
YSq+wn+Ese2dXL5hp7grBKhphlqkLByc0e7DZUHL+qxnnP2bcGI+ZovRyQ/aSnVw
I0qCt30yuMb3RwJFgMv2S3ZCMDY40Nmt+JHpIBa+p6VAGqOELlWafKLDQp28XpRz
FqxQUn2IK+Rhz0XxjqvoJTPsyz44wIMFURi4AI/AAVmXz42qJtFuQLXsoMHMTRd0
mSAAxHCIuj6Ta/ph820SRJyGnulIh1O/Hl9QFY4rJ0IWrVfbvFmmt5vTWx6oqr2I
hKzTt6eBa6m0lNHYvyqe3JQYEJq61HaeTXtxaNwGTftpub78Xdr7NiiAVRcxqrVM
JAKOYQGCRVabnf+jlhQfP95NrgerIOW7yoDUPlLIKH/MXsN/M2VPDLucSAbQYRjF
/Zcx0reDWAAmHAazQo9jc9/aVxBcSwUzlZ5e06BpBFNBBuWQlMvAj1yZ55NjQuSA
tA3gwFXs+JOEj5vXnJug9qNRhKgh+A2/14iAPLmlacrOABCQWpslct8QYO+yUUv4
ajajZFzXdFu8TW/QnD8GbPMTQHDBae2dW7pQBqHndt3WTMpgALn1wcYAdXKUsYbW
M2smCwkY72xFklBOJ3QuMrCWyarNHQ6wsSMBxHzfX6kVU2dPnXs+uCV/WaxAIMaI
9o/4bLxFPKt8YmgyoO1kiQleyJDgTLWub4+gOW6zm34wuxNgO45S2plnr0f9EHBc
ybEdhlaUCEnxRD9S8Q8cRnFh7lJ0xAWcoph3Xpn/tQ34+gSIbeObCqKtHqYhM3OE
qKck+Qv5q47FECZFsNDlMgtehBmwWxkafx7vT0EA6CbfY3gsHNMsUUJWyMBDIK5+
D4h1qTf9NKx8AUre4JiGaY1FeigsRIcABLlb5aTkF/W++atY+0lf37/dhX7Z+RGk
xiErk+26lWvpWNJMAqdv4FWsjum4iQHtrljxOWZbYF7koZm9eUMUuom77M3JKQ2N
gO5A/lH3VtluuM7p4RMChLPC9G/GPkcXRwtcn8pH8P7jJpIkdV+kM9B/QD+2Ribc
kLANlMBWDetZ0tvd4dsieiRcBGIsLRh8b6kXMhitrD/QzoegINfttQeLn0WEf/7h
e9xs5seF/XhRKFPKSa6v9jxlq/AXP7lLG46Qs+kHdHdXPwBYygcpH5cidAoSxj89
M6TX/9SokJsTd9IBdaStB5oT1JTxTtU/V1zC2XlyR06IaCj4xDPNq1f+7x6nKbh+
w0/bYgi8iwxrt8PytLPHz5PaGaNI3iupAGDgSvmbZ53JscPMoEcaZHuMJtrywKrY
STw7Y5lr4Zwrab1mAy/iu03iD/jW07fvDdEgB+Hz4Q+Knnpe8wHXwVjmHEbFTo/v
oc9E1aaVrFgLo1yY013yfchMVQP1vMU2TQL+cb0iyDpZIdd0kpFqITQLjUECAQlS
ms6dzDQ+srqoJbRMY1crJs8076pkiO+mQDynjHTJtEhLfbDoPj/GQ3/XXwXrjoE/
D1UdmtL1uMVVgOeu1zASQ0viNCC9eY7YOQxmUaXTqEULxEWS4dQ5BhWuBrSvpbL9
pei/HdJ28KqGepvE5WECRIlvXv1mxDSUPBVvHRhCWyB6/UOCkPtqOqvaa2qkRok1
pYUwiz0y0Wd/kHXpQu1hkF+THF4NT+Li0RR8DSDZkwbzQ+P0EzupHazJZX7C7wbe
lqwkR+Obwrj0AaZFXW+OOSB3Nnxuxi778jvt1IYcR3I8Taptt1gbGD57wLwrOfL+
la8Ej/YLovoCHji3BR4tkJYzaTFRFRIHag7NKgMb+idGPdGoWEj/c4pcddmBsz1K
OwXDcXcIQzxWXdsiioFzfNrrjvTAdWMmOPyT2wHN4pMW9lov0E5KzR8k6m7whHeL
Bx8jzVAcwp/pWRtf6CxVVPcNmXhprGCeIcCDQHrQjXR8Qck0UWddUX35ygpKmORk
rx9CnugAbrh1y/PwNyEJfMpKGD37qmrgBAF0YUGZ5WVsdxgeZWji9+7pqqP59xd+
xtU2Q76MUx8w6ds49iKa27SW36UdXxUMNCCbO0VO3PXy2cQJsSSoQMvITw3ljDmW
uaKvGwsDycP7NDU6+32iaGUNSBVBGfp32ek7ISUrwADp7hVGQGI5ReXqswcqYthg
OImyUjA5It3WjJQeGdv6Of/GZO11rN42JwRHWFw5rKIICZ8ob6eNUQB8v5BjFo7e
uSq/mwH+EWlGB0O7TBAH8R4SO507BA81tqG3SFCQtoo7s325cE8u9Sm/Cqh0zVPk
AnCLxjnkD/ovTD1L2mfrFEDGBUH9RMcDcD8+1rimqrE5h6W+j0Y9hS2V5Al0aMrp
h+I7MoAN+CtMXvzCQi6/jWYLkIMQ/Rhc88kmtUxDAcSkE1m6X7V2RHFL+tg9DlAg
BXguyMiw3Yl8xOV21eenR4dGJ9k7mJRtgsq+VN0S5sq2/BO5Cs3z+dJplAsTG0Kk
xVUCVhdpIMuCRhQMUTWkvtJRXQL6A9BOXSiVjyhfwMdH4URlgsBkrf2Did8bRSek
APV+qsl5k7vqrpuNh6BEItlgxR595s+0GLKEEftaT6oHsyq4wrW1gFipwF10nkL1
5jf1xjqbBB6Xjb/nU0C11JLrSzfmODJSL7PabTbosweGBVyTu9ijcOV7g/qIdruM
b7UIuBOempnW30ZwIC85DGydmdv531KbVOsknha8C0ywo5v/BblEOk06eM5i/W6t
IvqPH+OoOSICcZeeLn6ri/7mjxojt1153bWIkAT3X+dOmkxA2N3lHIT/550LcYig
MsTRg/Xeb/0jEEe2g20qYCPx2jzfOR3mfZsfQ7cz4yG364tDbPEe0Dvsal4JQ4fm
ZIrmOfxrl+pu78VVnIzl0FtkgsAJDNNrtG4hkExv7Klb3hPM27LjErsNkwf6EnHc
HsInNtpmtYwzETXl0VMPLbe3U4mpj1b/XmHcT9TbuwoE9+ZlFHjps6hXJhG1j4DB
7178fVQvtH0RKVBSW3Ps9DUEkxsQd/yU4D7QAWtmKAAX73n/STZ1mQft+UvMCynQ
QBfXCxigpRhaEXlXqmbicgf2ebiwTWh52nldh4rkBL5wVPpg3kjphTOdONuLsTmo
mRPMQf/qlNBmGylcbsBPsL/DhQ3If/bTjV4UsHOI2z3rSoX6TDECubIP2HR4xHeQ
xp0bUBn9CZzg1WLU3vXiM/+1e3XN4YGUGGkhrg6NbesCTSOZzIU2uVgobSyfq5SO
xL3yyfcuTmcBQhDBNGXbVsJPpOaNZlC6SVI02ZyHo/BlJ3FpsrY/0flNAq+hbIPB
bexNMogndz65WRfDwThxBcobB/qjoB1ZqjPQIxEKb86pjaULbUNiFGra5RIGh3jL
pjFJc9pp8z4IPQ/g0K5QVhoXjxmfZHmuL8wCp/UkYWaQMWmHK7bh8CjcaI/e2Z9j
NYadcsX9l1TXO2F02v25JJ//P1wgcfO4uVSU+aAvGE+KUL16CJJkFAjZ3qVjnrPK
PLI4f1uPvSeiVPASn5wGcIbvjORcLZU08Tzfj7GoxBNu3NHfr2p4pklU1v2U8Tai
qWNIrI5nR4cZDaX0clg07p/jaaubuOXHCK98fApzA4bq7asOn2fybX1Ja7lN1vvi
fjGank44xn8p0V1Dm/usNadRZOdI/Lj0nyS1cz9mgLbacQJiXAjIEXhdKiHI1ECK
xBLiAr2eK6nTm0n+zzq1b4XzDjG3kyPCJsXEomDZVq6opbMCI+fkPG+a8aMuagfn
n6UTLB9NXK2EDnlPy3Wv0whm9EP53a2AMUsv2emq2SiHiL37dJe+FKb4K9JWIvTo
BoTuI80ZzYzADLp2RzFXx+GvS98y1H+RHnQ6yjFvTpJ8lgAGmtXBOOo/3pjnV8Au
SkTCFKhXu17XMVsxOCOd055M7NeHJ+SlerkSwcCsOdNFZH/3S3DRe683iOO3J8op
20nmR8zhukfAfSByaQ8R/e5jh1QMFxzgZMkyfWrnwgDQUyY/ApLy3G750fDqlxC1
rIaN5+hnAdL+qWqxkcbM3DoekUaf4RDYH/XvHoUK8LkftfZLTKOXPWoETkQ+5lSF
edFcXCW8vM2udkbW4H0vI6eyrWfNPnLst4jFwZEjIz7Nnm0+Y0sCaSQwoTFRjuKY
TxeTvkjFJElk4W4u/j6kgRRsrmXGg5GgjW60wOYP48CEov34Oaqb6lLEMv0A83m0
HqW1dwngNH4Y1T1W2EkpoaiWgJJDKlZ3YwKG2HEEoa9khRaJZWuSjjXgUtdyhAbc
ABknub3D9enMeN7BJnNcbhWRUDoYtk4SGz1tUnHS3J3urNa0+XqPu4kujKgSuZMH
p2tRJPgNrxRTwpMwVImE+uwYvXetAQ5YSFfGnc4UIv6wmyEwoUEcD6fiY+ZCr4En
3cX/4tgoOHb0NloCP8Pw6yFt7Ht/x+VCuduNUZ9l6K6fPBPuORVypiFoDUnHvtpD
wvXRA69mIzSF7Wqw/ZF+Ar3XovCEq1uuXq0ZHkIAzGYHO0gp/BDdjiMFJzIINVAR
MaLEeQUag+2YpGJxIdWLB7tUZoEBM5eUKL1sIhyudcbOsTK9yoifp+Wtait5kpNh
UuPwz78hjgphNkoXeo7S0YRH/QJBRmeE2KGgqjp2d5NoHHDeXPJKSlrm8Lt/biHi
YwTP8fN0H1HaR7BTJybzByOJU8MhoXHLBRdUiBa/KObEHQgF3JI4L5u67jtzBn6c
E3oLsffQ8EUgqZpE8riqEhe5cul6r94hMVp1f2NWlGkJ4Ka4VQotbYkrO7IK4a1d
+MkAJmqQEGS3WoSLdY/Zctj3Lye9C3Xd2Q3HNNVmtjHq20bi7E9q6kSVdjHqDJDy
iDYoNonvnt3nH78m8tUYu74nBZEAIqSJtowcd3CuKgvZ2o71q6rYJdHB97HXNfkk
VsouQ+7rS1fZP8dmtL1hUioaPAyp+oA7cS4b9Ji0VoxKYyv2kNL++uomcsHG9hfA
2YaCZ4vEdYuWKl4VlbRpNPJb9vMusPH69LClhfzcwlUVB97tTZtLIhoojesVVmYA
aTWyPg7D2b0KKoS8gjpZfV6sPPHMe4VdpQ59qNFG4L7/Grf2gJ9Vp9wqOgimTXbm
j5YA4JWSxDivoQAEYgwD11fsnDmxZ83e1YgxBBYWQ99/e/5Yf4xCsBK7nf+V7/43
IGgb0HHo2SF+X37jKXSsZEj4XRSuSVWOGn4BNC7JsjiCCTW0IH5HoNQ07D+HmjX2
hYzGpDTxFcoUjSo+CxDud65MirAv25Ry6jL4S2hEc4aUgE6Q+sMMqfgSomSQP578
cGc0x/xVcnFw3M581F9Nup+i8ywqYx1rRzjN0RIIGylvpPQ+0ZoUG5ajvi/KoB0q
eWEzLgXrRmYYqSVV392q6+mX9+71NN9sGDVDbN23nqGM4M0XZDUtv2RFgYnpeem3
kZ4i+exnk5vtPc0PKtG/wOtdNbSbv02UD/CLSG0qpsat6vUXhqBRMyvsFBZb8XKj
8OYPo6gPCLQixq9w+tZyzbPdwPPsslo7rwwcNo6MWFZiYrW2XmXeQn9ef8o6njVn
uV4yIgS5rrF9wJpO+hdSOSF7NVYs08FCh+cA2QXE5Fwnc5cdu+8gy0UD5z/Zz8xj
lC6bDQAt6meM5I7ylQqNcGMd2BHujbXS7EYSWGN9Qwvz/kEwehbGU+TV2gRFRfFD
Y/zkCxip2rzgatFHY8AK6ylHGp/WlWOC/EBj6W4iRCjXmRbmVEQYZuWtNSOoiLWW
o/yFDZ0P22IQBZXR+E3CaIVfjJmmRdvfj9olYdYGEWUyzAF9uKJrzpueOef+lL9r
q9We8KATEX2EPfY7MOXH46l/XPiAPwQnij9/+/fivylYWN64fuJRTHgAKLbSY3iX
DOLWiEIxq3VWh5bkmQXE+IMy240n42oVuWgOT3hOUaK0kH9u00XCkjki6WVl77iD
LLphCJge7jvfMY+VPksIjcJxxkfMPXSFDes97nA93YDdFJHR6yu9UvJ/2EmPUkMX
hfTjevUcW32QArR8k2Awjbut8LkoVXT5I5siCSmWAgnFsM9zWjSWF9ygMJw9Mhef
7OaaOThSLCnGJ3NF6Dr0vXE0KQpawFFveESFGLy6QAzWm+qZGilvnvoojr5efSMH
HntvgW35FS68n/EHt/qILX+JmX7ReKcIkFuDFB5OIpvvUvcL48cOPopJEjCsXv9x
rO9da2zykj/EyXpDapAn6b5z+0TCOr/yGIl85/Y1QFvyQE4LUkEtb69IIygtUGkU
zBezdIxwdNl+DZoSF/oNBo4cTonZYYLRTeufmWQPerbr11jdm0y+CJcrrf87z92f
XiIcs1Z7X9nH9wrCq33LkGxD7zGBEMkD5t9XlI2NR+bkpJ2+9wSF547WjeNMKnVF
p1vM0hCYCfuWJ8QkhgVP+POGJInHjZYVyv4dr61sTkRy+GucfxmrTYvzDqkdh1Jz
nZ78fAWaNu+6g+UFvefnsn0Mz8/yfTDPed1VXISCI92+H3l0HnObPBGAZojdGEhb
NKr8zNRZiWL0h7UGVMA4Wiu4DZZbswEPlpXBXUrEjwJhAfqkZpLssVaofyODaOSP
Y5VmhNFfxlIArrqALnPee0m2P1hiv/Kw3AZBj9dNdqTiKf9lAVSeDm3JLVAjC24+
iozLBEsdQZ7UBSvOwGwYDTXZr/P73QQK7UrlpHLRxjbjZ3yJO5HtNDzhydD5Px9Y
p5GQjAvuNPZsKOc6gcbBoYvwJEKUPOjhYdfX5RUOqgm92XIyRoq5QANOu6CDRULd
3DiathJS5UdEaWwcyzsnGHpgrClvyxd8nK01GgLyjsLqjYA6s3CIJZtAwNWydYVG
3SsG9yrjj60b59hW5Y+n1GLo8Ma9oKjph/+sH4Ry4VY1y4dumi4SIsOWF1KoM6Pj
tNxDq1Bjr4tS6vB1QU6H/hnsKRKwivnmMmEO2E4ig/m8o8xA+YcQILPkTcNgN7jQ
erQpgcjECK4oWoTAdKjwW8TP8peZXUHMpn9hhbchpftxp03BlxelD/9Q8TfrbaFs
XwRpgFDLidUCLDH9mKunyOGGqyXUlWzs9+colV6bDHGi+Wt+ofRHrAAzNxSBKFSt
Dc6IIFoDuBbUlC9qLpIAS9qb7lizDAtuc2nYTLS/x6dkk00Ul0BTygylzHJwfY5V
zB0N5F7KX9XTXg55GJIFIaPXVJ9ucgV985yVD+yCyAZMg1QefPc23zmlv9DunTyf
nwhek3HOpNxAgEor/6LIJLncwBYKf0mGdy3cc2A2bNTdGxChzowGuk9olRQIPgOe
3LnBaUykXZnbnwgTWHqUXMvJHd+hXU28g2behh0zkuvFvqYg4q48zGLznjMai7x9
LoQPmx5omgsOzjxRUwiSnELxqxQMq7jZskfoLMidh8Jr9bdDYQGotLVhivyUQdhk
FYB8Rf5reFqgGqwFdt7qVUa4Hg32eqzMmyHBqa4G9R0PSEK7TGc5waTBxqy4pZSU
ZYm57OlbLDdWruQrR5EKmyesfpbCQVgVbxlqu3FPYNyuLPRzAgVZdArUwqsu5Ocq
FhHNGFyHz6xqlPbx4SpfD/6y2OlVQ6vqcdZYE5kGY2LdagLQ1arza0yQbWdcPGrf
LfMv1XOp1oTswwg/ANAo9xKQCvl0ugtpKZE4Z6bIzWnGYZdpFhyexdeG7v26LS6m
qfZU1ynH0arGyIqvaK2x2ukklJZimNoKNfiTYEn484kcBvtuUw1++4taaGuOVa8V
PGCuUaxuTIU5nE9HS6PcZKin/ObcmLEewnsrCPtZcvrkVgjv89u2No/uo2N7Qui9
229IDjHStlURmTbeH36nArIUXV5s8687tBzUGNXO2wkD5khVw1O02nUiv62yY3HR
F/lXjMYOz7daXDWZmKbKbO1QVm/lwrnIcboJMfgqqBeKTruHyzdTsDZ+0nCY7RbK
zyqT8MkbfZA0tXoRVPi49WTE91FFQtGLLI8hsK/gNmsROcC7zvlDNiUcwoV1tfxx
iqsxD9X7ALOpfJivqb6WC5ZGPcDMItLoJUCQWlQWxG7/+Dr03VDuc8guL0GkU0wo
qMCglZTNVs6+CI15nbdLwCFfl7bqJQgVzTXDf68VZ2QUZt1/QMZrhKz29BdI4MkV
niBttvplVoxl8YaCxX+XQRXZgkbCwaK7u8ll2JNt3bajJrUYNFohfl/lnjl0D2Zy
kGNIWUg0vKO/e/ByMsKjshPRE18jdUnqt8cgtrUWO5YUKdHkW4KNiqhYCKwbhmaG
EXEueIvs/xCn5tzR9yAEdjKEatRcfujDMbnsP8GAuL3Ole3sx5YqqnEPm2WbzQja
PWeJMJxP5VqeXEpvbLSPzOHwtD3ZCLpKRDE+kjbixuqvwOGK7fLiBc39tK1Ezulr
M48yd6Fp6oXEqvfvWbm4rcStjyb8qHBYa3ecn525GhxzUJ03ruXoNK8bsa1+ltEp
hHkyk6PRlVfnlogbGdauQwEBSPKkLsUom/v8pgmoQZt6ec9OzG3+liEV8oLPlLNw
ob3UbbAfEPZukSKL+PQMFt0llZiKQLD/JNGp07iHpb4hgjKiI4/bPZ6IvtDnEGVp
UtmAdE3ii92XIh4zSYi/+oD0fyclEdW3AK6WCEH879XmwZDE1e6ojM3LwMCSUQ8I
+iARJxwxvGEvuaPH4oANO+bwcqdv+PBni11SyblAehUEkinyZJu5oFLU/uCi11kV
ZLkAmbEpci4hAabTbfn7JqQHn6jPesEc4Whv5GOa1U0QQE4MNhNldnhMLpMAKpoU
UZiMnuG6n56rLBpvF+sA6IEavmDBBsjCd9k4FcKOBimzA93COEel4ext1XzQ0d0j
OFGT90KUBn5k3pBSJhR/GiktpX1rmzh5FAK4rwgDUr9d3Qt7upbfgTvtMveHB0uC
VYKQEixyzq5PmApNWTbmT0K/jcrZCkZRz9+wacvp4eZFopA1XyytLZkBP0bhKb9M
40MuOmPaH1hNUu14EdJ4mBJu9LAjkmcMno2D/clPPHyOimVm+9dCCx7vGlupacfR
PH95xuQ+/TCWAXhzDB2ywfperaFaVm1UQ0AulsNx0pMGoEjCL7YgyRVH509SORXB
vY5FDiKOHqUfouQRUhjynQbSADSr2GWX1tEJE+RTSvc+Z8PlejBes5zUQ731+7Qg
rvr+Z1vKgc5Y+LiPLIKf7z6mRoe3QBMH+V3zE9jMJrc21zMJ1Ib2E9YI3xtIYGOQ
Kt/z7e1a6wocWEIwvcqRLm8+tznVDzBWH07DldzGNFhJB+DM0Fq7VdeCCzD+6UX+
RLTRsglHcv+Yd6spriz9yDQ99nCBDBaK8Z5h8mAHbmsNyuxw1bGOsqtZJVvKUYn6
JgSJxUI0dAh1QoZkMwpmDH/p2QxJCcc9LBO/ZqFy4m1jY9mH4cRSbfJaL+L9Jft7
gli2PNyN+PKqU5Ngyl2gNmFZxrcMxaaruahxbCmFD6fg/y5MVStEMrkvcCwtVf+C
08y0rR7SWNExah2JnsuJpR5pWhe168GEzI6Vq9BT5mliypTMNuOgDuedcGY0avJc
N5bSMUlA1AgrbAXCTadoUHn26zOGOLfr32MQKr4dC0mLJwcfOfhv5PK3bjfiACya
wMrhUsGHZCss2YQy/qT4aZ9u+9faxOI48mj3jhnY02vvNeZJ3uxa2v2NA7Qg0AQV
A1YZANtjGuiQzLcwEDFKOPCJWef7YxWK/4NXc1ByyB15+SNKtXuz5YI98m83i5/1
vByVMPRRxmHUfWApLjx1Ve2gL0cCqBdn1n2+6YXzYU7Bvkb5vjB1eaP/S7UNpMxo
Y7oNgg2WeX6ny1GyDHySO8pVGKOyqBrmhJWlB5HliCVDfujUfwaumdIdM1ff30p/
oMlFgrdDr+9LDZNZxD0AWFlBJZqW1LLHRzJs2rSevVcqQ+Un2TO+1oc4fLZbDcNf
Z2WVb/cipyPHAGH6A+ZPL3ie/b33KMr6BgKXbIiTymzQYz1Zm56MV8DxnKwR5V5a
X73zrOTdLNGQg7VRhzeIhkswL7Uy27bv4ngSkFYuRlK87ax3BUVcWMjIWPT5cXZl
iLDTXUrdqXbpRXuzv5OFOcBcZpoJwdT/hE/pyAleoLpFhMNQErSBwb8nBmBg3+7l
KBW188016P8AbqVQvvbnWF1GY384ysrPVTHayqsIydFNymEMhTEAABu1nutK7S0A
/P0ozpRkq9ONRJ3lryhlXjbsy6eN1YrTV0ThEs9wnpNdkC6FjAKND6gBVxzF6f+g
GHo5mbaHHMJWIRD81MCYgm95FMqXw1oXSUmzf/S7yw3kKPeHRGO9ppSUWjKIdBTz
0UA3raYKiTBuvsSL83qvsvrELAk9mPX9E0wwWeMTGwBYiIJiu7X8ncbMS1Z0jV6k
hcvfNxjIsE5NjEh9wPMipVHO2jdc1/K1HycQCm+hEtBQ7E2S8iNPE2xGbWF8mDxl
sq9DUS+aPQ1MYEtJTDdWzW7CPl5FnJ9MW/Wus45/1f+qR8zoqITprYfU8spfso3v
3j3J5sr8eqfmv/YW3NQtr4PYunQYLZKz5mjhYI2cjMu7ilkNmtHm6d2Kdh7g5+iS
R3manOuE8hwO52+GDn8gsycGR6u1Tq46wuEiiCdp6fHBoc52d+gCkkhQS2cMmjFV
a1DGqjTCzX7JEiePFUy7JMWJHwIOs5idcrfHUkm4D7QkkCliqiy9YoKRUDVLBP/9
KoxR4uKe2mpBwdP4NawdPTlU4OA4R7PN+SfG/XX5cCsymv3oruxhyT9XhYMEX/5j
78J1PGIbuN5HJz5IBqp04uIGDkch9ttXT03kxb4kgW94yeITnopHvgOEAxU4TNsv
Lu7rRQcNx7bHISxqygnrTlIziyXhM538GGgiUlXwMS8PhpRTz2ad+k41J7yItrPJ
BaETjOeU18AWWplYUT0kpiPNC0r610GkwMIUWVEC+nzUv7E9IPqXCk54SANpP4y/
mqYaaoZl4DWICe1sc8lKd3sD5q1v9xT2YwmNItQRxKoE6AY+J8iSDpw0C1tdtlBP
Ys4XqrzRrOSHqxWu6DvK4pdlJHy7qjNb/fzlBIipOVe8kKzRtjk/I1ATkwTSTPk1
731rauatZF47JYcyh2bzxxOfmDgSqwC6YAw05e9s9yFmRXDpZXOQU9ATRSvjy5NU
G3O3IRNzqYZlFvCBGfymcXKJbrL6GgqEu8Rc4wKRaYS6LcNm5MGK07qyYVHsEVSF
CGd6olT9hP+GIAEj7BKoiC5Ia+zO213Ugs2VMrzKvmL3CKsB4AudbKfQBiPtVX3y
E6Ta3RRK6hekkmgs0t2dZSfHyjKuN4KWk9QvpTo+7albqSC/0+soweHEAkmQhh9I
pwdHgzKGapx+E0KdNkg0SJ6VVal2jbKmXCeE/OkPi/kQ59FJp0vaijUc90oxInQO
R4GQG1oeq6UTn5NvmzqwrKE8qWQCjGx3AS0k+beRJWkrVFfZQoo/SmiuQjC/8eoE
fWmq3+i1q6NE/R86QtjTubXVUsJ18YNLHCq0QuZJSqBh3iMM7frt0DeJm1/BK0VQ
CfE3U2LU3BjMCWLBloQbaTHg5640lnmzdYdvXi5azDdW5gYVtNgRpUc9DiY2fB96
lQrAX+xjvwwS4ibY3Fv0bsawEpkWJf90Nsw2s0w6M3QRzGuOJafAD2fy6ySeknTm
xOiaVPDad7dwe47yNzcjl/mR5XxmebgBmhHfdfLzq4sZhC6OQ/9lH0b+fCXT4w5M
cjuLx1dAexnUvxOJJd6yCW9mtASfHpVQSynNlO2/MI+cAUaJYm+tQuVJa7/kI7nn
0qV5x3hS3Wf6q6T6VLmFquTjGyewp9vrUAYab3GIfi45m6MRO/JmNKh7VrTwuyYs
pa0wn6bHsHvX606j11m8JT4koZgLMahr/Bk77AvI+eHAAvcMeHSUe+XYbvGV7iMN
30wgdFD70lQPBjXFreFNls9bFVucDAfKj/TVRHim9zDtDNtbnUm6ORMifh+f85xi
Qo4k8+be16SqxV1w1J5FPMwc+P1gPyrXO89ciJhwViueX/AmU6HrCGdVTBQZAhDr
1y6T7xIWTIyywR8wx4hpqugenlDK4vdvYPdNZhxkwRmnm070qwKrMmHS5ZdgYjr9
rgjoDfydEAv6W0z3cReDNRMXs1Sz4/85ovPwSu5Okd5YiBKin8GH8uvD23LDkQB+
FTTMFKUzi69YH8tQPT/HpNt/FjxkuAiDsWFM2CzHsr5GxU64QvJ1DbYzZYcCErTW
ZDB2cnZacAHpgZNSBMx7RvY+9pR8F+kjPYh3Te3XUTer48GH+8o6vH9RK32fz4TS
23V9Dsdye8ExqOTqNk6YXG4PKzxIgG/H32nc4S39mnXgoruNKYfUloz2+J7Zxucw
ykO1PrxMlsfxFnynEjp1lhBJJyHDrQXCG+5rTw+PTOpNX9DGAVLu9legkYPcZOdV
NNaeKvCddNuZbwqjjcZvxIVdVdLRlHDmHOZnG3KPmIcY1BxVIeCScivPEoYfpMUB
+WJmao/2EcXQsl/22/IQGFkYV2NuSqvDsLkbjY/UI/4SMi/pD4k43JNYnw/JYoj3
1dtMfjoWuenhdsxuPt8DdhlokvZl0xlaRdY/fMpi4KZLhFlPR2/fRumJmpbgzmvD
Z03Ruh+tclS8scwOZKPx2pnW/667z7fc5634FWAAqiw12u3CmizXikc/FQV1Un5g
pthe4clpuN9RZ89D3tRQVvS4fGw6fJduqYHQ5fIUxlyBAJNGtvC4hip/++GWkrBo
467VWW68bpz0jUQzAPPfPhgw5teX0u8CasCJm1JIob8T8k2tanEqmO3VaqSMY0pq
VE5Ey3g6aiC8Iqc1UDJ6PCH2WJrwkznSK+MSozxr0kld1GG8503hQuHnY1JzSURo
vS2JbDC6wbUcY0S6suXkQh6UL7oVKxAqWPqzTagLZ0+oD8C7dZ9VObMr6GWB/6WR
smgGd40pINsryz/WWo/pjteB44q/mhCBfB38XKGSMLd69Ji1OeQXADeqLQHSoKRl
FbQ+eofZED+EqlNi0E/SEThh+VhV2IPd5qeZGaApNQOXvZwQkwDYSbMnRvSQT7Ns
cRWtvG2XJjTp1tp5GxmnpUewkWLZGJpvex1BjMwImlEi19fCOR6zhMmkA82Je7KK
V+KXRbDK00lYXJNzLymJUJBgEmauswnBYak7FHuNQwQuvhbgXg1LJZrH9TuexL44
GMEVTlR652gYJj5riHcM5lFzJiwaLEqJ7+Zgy5Rdx0UMeF4QZDfmjCS7jKxFOop4
I5kYNWzRVVE2O7P48BdONRdJ/meT0q/HYoIBEDk8sW5xCtiBd8HXSgHkys4T5dmn
HeOHhH25Er9DHfujC21Hhkaplzj2cblxS7W47B+W6ZINC4BYHP/sLVZvwAikZZfZ
Jqjo98njJGv+1asR4ETpsoDkEFBPNXhHDbMvV3VnUkXGMaKZh54Jo19nS0IdKLm2
PbNMFrdx1WBXoCPH4EU2izx7JS5TKOc+WmhFUPVRyc/so594/telMqIPS4Y0W1aE
y/7lnjaEK77VmVOopmSxkBnACYhYJCEwoX4RfmIng9fdH0BUNJwbYim4UGu8FTmN
+hOkplE+BkPrv8C/M1e/r0bColZNfVF4G0g0VYEOOaqBUfaEkxB5nyGotFJqwDay
pot/6nnWVK12V2fE9TFvrUaUStReYCQZlwUg61DwJwvCI9T00DfogQAbnYTwdGqT
1KdeUyTU2jccy4irQMibFc4WqaDradFzqrUClGCmNaqOTNOOnXH4kkj3x/g1IeIQ
AYhX5dUnwWvSb0DHg8vRsgTVCQIrKohMIiZLahkmAm5ytJl6jrTa00rKbKb+OO5p
9YlEtkeQESUXznP8cJenWeVTdHACE+Ynei6mO1TWs3HnrUvYJg+0/Iu1j7U/1CPd
7TDgSUW29KRRMNXfeOpif1pROJUOSXP41MT9JLNpf2QaWaKlXnZYywwIWMlC8Nrd
+uPV0L13CtxRM8i/EYgP1zj1rADmFTFHWiJ1COXjYIIJSVsFG6eu71uK72JnmHxQ
3aNPrblto8pzG9BKRvAEqw0ycWuCNboTG3InYYce08bJrJ8+n8cKWHe1jHZ4K5Rk
KKUmuglvHwZp+L1Iaku0tdGa0UYc7ZKKuEuth7ivV/Yz1MKB39iDRVZeRtAuPhWj
NZw3Wtin+7SImtH1etRaYtXdxHivO/85c5dmKncJJkSaGwPFfwCl43YOF9AHSPnV
FKIq2D+BYVi2rNeuyhD5Y/iBxWFfPAlor4N8uyZb7hqpfeY5kcLZXiHCfW7bqkaP
zm1QsE64zsUOyMzdisufFF2vzBJVZYOAcSeRrwLM2hvZcs5jWcE8Xte/X/wQ2D3N
sXkz4z3AegrZ7WTTThf/GqVNY1EToSbdMxx/kCidur8kXpzYUVpdHpVfnY+CpCs+
q44C9q+6D57EbAHrQn+iEuZ99cmY8dfeq6DQZBJAjzUHQeBua2HwG6p/m1x23b4G
9skUsc7MdbI/YLIb/vwkeDWvsJRnqtOgf9RjNrqBUJ7iq1q1dH7J3uE0W5QZg1wz
zCA79+Vh9IIRr2jWkbC77jZVmm4HR+oCMp5b/Wxrasf8OlUVgsFzz+MPudqFwSTT
77Q2kNO1oZuDV854z7Umqt53GSrPy/02fFLAcVc83xEdgc5CRZ9a6ccw1iUJ7w4U
LEAmuvaEOakI2KvCsiiqwEso3HYiy8O5dM2J7eNUBwsf1R0hMV+ebiNUYdAQnk2c
YN7DDusZwDCWCfcbNwymAJCjhsveRGo1NyDgeSH8we77IvnZPSyxeajG/czLO9mg
Q6EvQ7hskWwACVDqevgm7pk8GZ92sjXbXxK0luAbpYEjrNe+zapA8amBglOHCkf2
gQEonhbY6LBkvSo7yMbMd9mDjazt2MenoevxZQfsGJJQin1epmnOk08COfa55EVQ
Sfr6qHe97XYj7rvs5X+QcoW/SCoV+BXFrn7G50ZIAIlCP83kg4MpKf5gEQ5VyiPq
L9OSnEEcy7MqD4NLiUYbEK294ex2t6wz0QNqX6yOdo6Ne84vCf3X0uLkW3kFoSuj
z0eqHrw6ZTY2YdJhlFotgSY1TFgn0Y1b0/DX9S+eiceO/u6SjzVEqJSPlto8yXzD
X9RdumXFoYK3/0EboKTpsJzJF6PU52wmusYmoe62kQc43zibc+6rb1uGFUlts0Kb
hiH05Hm3D95L2o22qwH0NO1oEpONZSN9zZ6xHtdgTewlLxhAUeTcyvfyuupyUh4a
QxRdycBOA1rs/EG41PZG3q5TUzUm9XMFi5vl1Ys23JnaDjUK0WLpXLrq0eKkZaUN
Dl2oY/OHfwdZ2gzkxddVqXbvnpO2PyWj0PTOQeBI1jyNPRDNE1lfRwtRVtZjABE9
DE2hRti/nDQWB1xmwC4kSEG4EeNTqFLe/EwcRsG3hyEkjvcU6/4BgkQFSRyIUVLB
++/e/ErHejNDJr2dNh9cX92f2fADISH+Yisem/yFUhyYvqECrRwhvLjXF14cJQ6w
ZHTeut4b7ZivHijGmY0lnonxzAgN15LY4076u65Ik19zuWNgf2XaAuy5pewY6ZwO
RVPD+Q1h4/lkq3J9I76+b9ts2PXaXjdV6raLjLvA2OdIAqqbR69qhj1WfNBrPwae
4ODWrbg1j7DccYOLWokKk3EkllHMNjAiw5BKOPW70fH74BooFkwNAhdU6FEtto2m
fEv579HdCL1wxIr8opHNfaze1OzVedpIrKuVlSlEplrCcB88iEoOmCpzBtm/d3VF
ebTqJ9tuHlG27vWv3kXw2upNCUWL2femZi3skRduLMjZNAjBOSr4Tf3FTSDcn37c
6H9VqoZICEFWqPQuY9Y+nwIkhr0yQnv6RlGGvb4+/nVdouA9NuEzlRXUSea5PvA4
K46Mi4PsXHQOd82QurT0/jsXP3hXsLqImHeKk0jQjJ7G0UvUr0DQAizllJr7bkYr
i0LxVh20K/BOpfMNobJ8sqmNAgAYArh6CptGCv/Zhkmcq/NRAWUOuAou7xp7SIPJ
uJrGdR8lNU+O3Ql1NWk4Xb727TLSGEs1OQsml0qx2p37he3EJ4mIRRP/ww7suVZl
Qyb+OBV68b1w09y0ptUJQeeaAnbYwf/6dovFOJnE1h6W3E/f4BRhk2Aq2dOSmZDR
EP9U5F1U9QKJrrzw9WBeuFc+pkyg38KVNEKBEM/IATA9+seLH5KBlDj3gVa6TJaL
CEuKnF+v0ELxxtcogNSkuxnE+KUYslpL3YHxbIUu5GVdBfZ/5J8xPFhVV61Td0Gk
80bL7vAqmLoptNt8xOOlurgsVCe9mG+B6yWc4wH9BCRMPZzHP5mV34RmBDNAkLI9
Nmgj4cIf8F1OXj8iOLuwX+1OxYN5Z7z6cQvEcdvtqoaQ1q+RmNJnfLmZjESrgc7x
M13SF7XohmrR1U+L3CT4BzvYRBQbHaT/8mMmHt4Y51dKV9rN4SZNaUeHQFudH2z5
7NVQQvOHE4O8dwySJ02ZyFK7P52oTesJrCp55TxEtC8jzO6PBAlfJWM8yjdsRKxF
BaDdN7XDwsNOoWvvtlMJZF+kiDgwukmVQZeCMLUDkigcuxo72Klmq0mQ60KthGF0
r8It7Q8P4wIXvOkITj5U/t/KdGLcHoDKndHsaCmvmKFHlEd5zPvusy7mR5AoeRj+
2dOG1lu5lUSZpZcNZf9xkBM4E+mLzy7Ce8vMREyngKEqkjvED4tftzQ4Fe+6oa7b
MJjiki36BeTrDQRb6l1mATaj2Lm7U7oWCK0WGEL74RwN3gwhb6S355M4nvWA4vF0
QtPboCkcxunGOldtxbPGe2nD2op2Mxc/H56gsYrjodZYXORDMj0XtxvFDjoqZEl0
ub9WMxBG//HaxewL39Wri5RwD2Ny1XM39s8FaQT0ETopLzsU8hP0Aq+nOUAwVxtd
tYDVWBac+P5y2N7d+XjK/7Qt0hO16lyIhj823w/6fmT0msXSefMSKP6g0EHTsJtP
3DBKDak0GEJi+jFwJiFuaRACy6VaISsTk1PivzdbAHKTPM4WaBEpigWlLskdLGQ+
QpJ3CIDmFRfovrmwHP2N5rppCe7fCLi7mq/VjNs6TQV0alOg0E19JFp3VL/1uTJL
qHSbWmtNABsDnRO54qy44AVAKdbUtZC5j7Jleb7pMQigY48X34FgfuO44heMVqaS
dxik6ahJ1XOlahJqixeQk5+SuRoLb2ljWdSVECaAj+P2cHnwy3iNnKjmS4Xvqj9y
3rdaBGNEdFaq+bZQiYOVPYH7X4KUAq9LuOTtOK9xsf2bGkAzB9B2z2cyufLAPXP5
KxsNWtB9R9mZyAYeGM5SOZIJ/fMjQ3DA1qOwwMa6/PJavIg5QM1SS7vuFJ/mH0Gn
2WlUMzaQMO7V6GY3O8lkHT6svonLQwFubpTFIaSuFP3aMrgUw8IwXacHJGiKjD+W
5/US6IlKDtOsSET7bdXwHdshtBWvbo3oyXYeI59rIQAj8umiYhVTLWrUNtlISVA+
pg1+Twr32xZPZAoXmllScHkKqVwTAkLdUSqLRxwNfjhduSB76Kcu3TCGnmGEE3Ja
IIdp53YOSUeSNfh7YioB7hVO8qJZOqPIaE07t8u8WgPPqUoaZ+NTCi8t3+RR1wgD
ID/aUv54obvRDjpwezxp8j08woRa5tgS6Alt2KUabKFWrIcKuRjy8HCsiaq7I949
7dxpx8Pf7tkwaCz6TCCr5drR1PSWKTNHbqo7wh8fVwSUumkAtUxeTjiBzIq/a5iI
CUjd8bQHt15yfjqHn9fuQnUgZTupKFU0agfUBUuugSK4mmBKohxImWzeT0G666n3
EZA6SNmqyhcwThnaQUGQsNNUN9nrumXIoHyTK4ksb6uNaJzWDfmJk4mkbTvijDEu
6xSyazE3s2NPfNSdgq1He+TSPVf7PtRnV0mBTI/EhD5FpLFIX19aWrB5f46Xk7D/
eLt2jlDJPCZiSdqqOIvz15GyJtaTyrlAfOcUdjkdnV/ENKz64LoHq0LIqCeKtkCX
WKl2x1r88D2hGnejY7daw95zkRBkoxFQf8ds1xmHyFRFP+SUiSV/nQybbGsfZxv2
s4BQvoHvjInvtGlfvdxR5ERaM13nqM8Pe7R3NZdpaLY60d/wi4k05MPrAgM4fp8m
am2nVrWAmrdHeU9zeO61SS4YE+bA8+4fpg345LW4Xm7T/1SIgB1B9th2wRz8LF8F
1pAOkyTh/nXkq8WeVy5V2zzGMhF3ZC60jO2U6JJCljONnXP4wNlnlz+RHXl90fl4
RTpmwqB+BQb8I7/dhvSyWNXG5tKOCqW6fA8fG5S28/F0QwS9sT+7eqSPG1oQV7qI
EEnPDQoE+eE8oaPzF5HLMwgk//5Df4FqI11uQQaEIjzKXStJItFi34FlJ83NhX27
YD3Xnbb+QKvkPkfHiw79mFQC7UyjM3CD2UUm7h3IulgKrX5ki9PIKGhKWwiZc4Om
RiZmDqsycc8UzlRrxTZJjI8plv4/s64rbtowddpqlTqeKpk3rwshKDwJ/+dSMg9C
TYwBnxG9XTojWHGVZcrlq0zTtUxJ3RQfAGrekjQS+zz9Z+4BPsCXjaqUCkAPNw+V
oXS+B0miyAs/WZSRplpGm+j7SXUjTbyVHFM8PIkzo7AkhDOfYOBZieOCPkllnaKF
xP9pzXMTU0E5xD9qDMOUhrBwC8fOw8IQYqtU0GBkZHfp0hpNy8BpLTQmhFv1f3LP
r2Cz7+cVeU4dZJOXrPdMYLxCSymsKl4wZD62K8HneRWrhgeJgAVF3Jl7esYwD4PX
K2752/3uxtcFvlbYhxD1WDjvV39rdPCQHUhpUmDmP4tqVY/PyZEfMylcwTPFNMVv
j1CIpxW2KmWgFQPQfNPcpAsPjjKUzccnkVEx61j7EsWQcglSZB6CJv+iKZp78QEd
Rfxwt3KvztVctLwZuVlThHmkJh6jxdCE+Vt8Qwe74a0BXjEmmXiyx2IsllyHSuki
Q1dIhTiMBMfa7c94RAPPB68b4kZJRfnAJum4Q4vK4cljF+1phFDgn7D8ezwFkDpH
JeqPNg1LNkcqco9lAYsHEoZE5hL8CwZXp7iiKEAG04U3UmNcIELHTRkC4xgzECMu
uVN8cjpVimXmyNaHLACA1YWqeMLFzGwzQaTnCRcD4W+Vp3rlpUQwOAW5LS8TtxnW
9KtdypPgpsmhvBOdK7BpwLuHz0VyOfv+JrFPJ7UvX2jWwQOdI4WK0qxvOyM5vJCc
501LpSbqomil1mPX7Q5/MODGtVi7w4ElEAhAZwyGA9tkTfRylqrRxOHF5dagCPzN
nzEeuV66aDXVvw+uJPAtJTlHpoljC517AvdBv6Pn0WPdw8F3jvmbtGQ/1uAfbWf2
QaMDd0Di3T51y2EOMRIAxMAq1qbrigjieigkr0YCNBGYTVYGnP6cvdbmS6T2mfkn
wmvsBzpOaDCHorkYMXuf4Ybe/6TQD2URaubvGZMsNeMdmpQkQ0T+KG82F1Cv/p3y
NynhXggb2evaCOgja8d395xgUv7AR3/PWvCdXbFq5baRelBTlyJfup8Plyu2dW9C
j49IHem4gAMQQSDE617VWOK0ut6GZc4RA16tLcu8TGezR7xGMSECMJFckykyYfHN
WoHT+KhFxgvXlItkQvdCyOrF/hxxzShXRZxFD+LLrZuiFuq8n10b4cPjGNcQWIw2
66O4mHAGPWcHB0V99vtpM1YtLpI0lYLkSfgrx1lISp7jvSrBKqBBAq2mQYBmCBH2
xEJC8cVu6K8eeV5RAiyTlFq261xWMno8FGD41+5y8xn09YgysDK+W1QVC0JjTA+N
QeZcsWg8RkhF8pkZjuvoRXz63USG3pv6xEFnoDADMIxssHntmSr0tseoB2DfxQGX
HI9qznhJsAx49APotWYq49GFaycv9497KkSKWTVI2+BKGCn8/9+uZiO69taxfByH
bI7VZE5RHFLBeMxVlAXoo0GGhRsZIVe4OTkbDQD5U/aY6aJv7g3Ua/CoJkyB6sA6
IRkv1fgQ8dyq0taswd+6O7Pm2ItnhScFi1kmMTRBq2i2ZkobV1sqMfsaUKr+3MvR
81XYLb0vH3fuYdoFB/ku6APX67HmilwYKCT4BlsFeDIzyh7+s4Lws8xPTEHutkXd
b5dIgQR/wVvg5gtsZFIkq293RevPAOHXXFkqJsk3dG8mRrUlccA2RsqimLiFwIQD
1vi3YfeKK6qN9xY8Doo3i4wM+Bkvw3OVzAeQWeau6Plxzwmt981jEJBOl9JEUbRt
6PDiwrKZGDAUzxcpuIlGUBdxPE/E0lUSo9KammmdDy6JmCCH3GP5vH+9jqRz2Mvd
rQD75llWPyMAmPaUZqgPocd2vEuagjLw907IDb0jwdsNWW0f8Jbdf87gON7VSGER
i1K/xq0A6guBPplBXbR/q/1ZqDt2atUOfSeRUxKsS0JA0+L2wEJd7SQDnWrqu8bR
4k5Azu3C21VWYO1FNdC1EMFBIO+a7F1FpgkxYgbQZE4Pn9rwtzabENhjliq2n29C
xQtU6htpNRGMb5H3JMw68MKGLjKW8i1wW5sUPCV7EZe0xFu5al4jG59S03TDVbSE
PiXUG75UDu9jRO3YSlDoy3xN5E0k2J9Wt1pUjsOk3iVOyJZXipBqiyU/n2yQjwcB
pbUwm8MniyRNO9fAK0OiooZM7F5PeCvovMRhY2uFcEI/dkC4lnWDz362MtAOeZ5H
vXigpu5Q8349o83vtyqhsAM0W/JJqZ3D1eplBb3d2wIDUP/xpTtlRDyiIXUaan7i
iPXHMxTYd2NKfRXBqtPpclz/NulxAqeOZY0baSQCDOOGSx0G91sZpXD+ZjNh983q
cqlpMPhG+5GA1ja+xWFn/EtgtsezdnRpnImSIdUK/VPO3lTD/YE2nZ4Q0iQOGmMR
G3XRo9l1Y2aPJn5EPibnoETxilV2dwjadu+1SUjGMXMjFihCIbiIePiZAuk3go+z
y6sgN6dK8K+JfQxnk66RlNFUOX5vg7RnvJ1mXK9JdtTUMPb7xhFt7lfOuQbVesJk
D2NHvrMd2j/0qq+skNwsMrVO5Ay0D5aLXvl/RzBmqjEYutTSVast0/HIf5dm6V0J
QNoMF804GwS9ltYRaC2xXoPlsdugY/QDMBsW1ULcvF61kXN8Irj8oecSRP+6nqlD
ROVWMzhvay5S4y0RTNCZFTJzPEvhw9Kp4K0HOqA2dmLuwbbJZUgtioTzrvG3mNwT
nv3fyY5mXFfr2jpw+2EswGt3hlRXhZGx/ZOMSAQ3jqytaWmA/gEgo1srCSNoAF+i
qlM6hw3DUc29/rHid0HndX0gsUsX6MY4CD3dqy/aq1fzLyb/8PYwZTHhGbZlWFQq
LSyQPFAStnNoLoOjwKyPeOu9WbK6QftS/4vpdmVcTVBU8XRFnkjokqypeqOI5V1b
1N/WIsz0zgVrNRFGLbG09ns/0rbh93OHasSQPanWdmTi1aFtJadhkL+1wtGTMfys
Yxlq6dP2oU7q/QwYBAIhscaLvbOKi2nO789BlEPyEJXITqlB+lAJ9DyCZJyiLSCa
xH7stTjHqJRNC2LsggPSUT9zrTawAu9XyGSWCE5r5hgnE1m2fW99eSXCytk2KU1z
G6+iGDtrUjopstKuu6nJTkd48MtKXTGvkywlGxg1Zkw9bY0BT/PZSqO3XHNdNIy0
vbjANDQvWVA++3qgjDk05G4w4s7vqpBb2erpOoHhiBr5TY5NMXxRCwUI53Bfup9Y
NpgiBWeoN5yqHuSdfvB67Aq88mmDibFnOJT+iXmXKa9yutAppcQR7+1BrOQeqSzb
z+seP+pdLsqAHty8tnu+fyJEkGPRGg/rkY+S9Qeze/KzwgXOK/u3dM0R+8/2febk
5cjh/Qt+wI2WIHXXjfqaMYE9QY4EiCLHLHnRy0X54vzu7ICmt+H9TuyWAS9G9aDl
SDx5K41Trl7vr9+3Mqw3k18A1bIthAP2okZ1moqKkIyeiikcmJKSmcA4qAyTVbb8
79bfGVvbBo9NjOXu/fY7JrBXXjr2c/0RJBJ8izMAt3NuZIX6zmWxYFuYcnw8HVSQ
HPdiwm4ayV2I8UhARJ4l4Jy6s6EugqD1XpXb/R3MwiZWQwUfmG6ZY6r4qbpg873H
Vo6AJl84UNcFGp3eKyzDO3uvNs3EyzxVcAce1CWf/9MmzHk1F6IJlAxAPdigSqvI
0gA5nJvKKTKGAOVVbKJBCR3aK9bTBOLzVF6cWdeV0V/kblTgIvWM8Td1viPaCfyF
SNEAYcc9VZ1KuvbrK/5J2zCAcJOqrMK/54sZ4GMzPGk1Iz7EVwIeQCOF5Ay0RT2O
NAHc3mRljCgWjttbOY++VNKBBAm86SizsVw9fwXlnhGUSdHq1ocC1NlOncNPBZB4
AkX6ctYJ/IQfySx0Y9XfIpxLncxLtVKCYyh0E3MTMnLIFmp2qi1XNk3QcgCbSnly
BV3nQJUGCuTJbGxfWzeunvEAaUMa3/Ge0cACOcviqb/QG0Pbx350QoFXBE86GBGE
h9a5U40lDVqxK84FqJFhxk4umrAgaTmCb5D6zGMOupxqJ8PfYKCb1FZMaV/Gpa9R
FT+vfUf89iApEOC9Bbo8hdLN0t/hyXgtOjajQYjynAoomr9ZE/AltBGRgC/x5kEo
faiWi0UPW1numexai8PEkmcfONLyJF1RCTZgFnjSS0bdkZoZcZFAUe20v+ix/GTz
5lMtaZ0KL0ZQVc7z1DhULaSZLGzwVbNIWPxXXuSFqW4YM2u03HCe9Jdky93RbBAY
qMWuEvhUOsxOFONJFtr/fScIr+qs0Ee6mna+SsutaMaSPeBlpgT4cdyopPa0bTw1
LJyQn87aq4yydwR3QRwtY+wOlD3br0X7dIqTQwVSVA/0SdFmaTo7IroIHoFxt7+G
EFxc4ry4p3+38cQy7B+zAyRg3igdGMUJN9uVO6sHKYZ3HDVqqJdgZpkHmUnqWLAG
iH/fmY/Jjvhl8vrKRU55crf9+4hrj5/SQd+LhyguWob3lRgp2nnkOWHY366Kw5FR
AH02C5Mw8Mr55tJPD3fnsnhEzBW35R/uwfmeiUzoJyehSQqZQVy/5+l4PeBp3rqM
33CUWRXr3BkMcJd7LC+TBHshk7h5D43NVRFMFkVqjy0CG7fRG3koSB0xnPkZwfgc
xd6Xzn2BQYDbUsBoGgPPvqtSAyWg+3cy+7e1n/UCHeT0oYwt1l9hdP/dewTITBIv
+1SFyHps+NZLvjLAUAF7QRewdf5Sk1Rf0pBB0M4nzb5nEeK9qXUUy42TozX5Fa35
f6LqBWPR33XdLGVoyPi516AtdxHkuXgF57TkcTWukGmHEcJUsNwsRFS6RY78azMx
c7HU7SUBfaFqYpIiwGZ9yodK/qsc7iYqUz8aLFONbben/cozqoWGq4EBGQri071m
PeZpwiMIy4PhjQwiz8feMXbfkFCq7Z3XKhjjED8OD/WajTHsv0KqhZYyrlJtps5m
xK+Q8yH06MX5Rqg1WDObdbPk32JTsc91yiA+5n9VHY9M0hR/9WsJJ0dv1vUqdT9m
nisBOP4h8BgucM0TI+Jrv/YQxf4rbnfpWdQVEiYt1Gg5RtOmgTs3FfWzu50JuerH
/8a0PqMqDxgO6Om3ymjqZAhfNz6zHahIt5SeVbWM3h0fLkvfAlexA+psTnJJd1qZ
ODpLR/ucmeb4+NS2zvnegK2BaalMTT2Vm7ku3IIL+V5v2GjTG0QTEUKEA9JxXEKf
X5rC7mJVVTQv34i5F8lddcbuahF5gGvDgCph0wfN7hxobIy3WUS0PTvne6Dvy678
I/1LiEJdulNlPQehSn2bMhFtE4X/vmKIDGdGNkdDJVT1URTCa5GNAwtHqRbn2Us1
MYF5+4ps/R+kCrQn9iI3OUuP0PzTaFlkET/5z/Jgqle6jqS5IiBPa+qJnHIDyHSC
rKNpvFzMKiKmGj0f4a7Ua4fMQ3j3mh5h+r59OJ6lY+gICYFsn3EDthcUk91Dlu2X
3Kl04NT08wN6KMYp1IIR+Ooy0uQNTGS4tOtMt7usvJNyEysFt0Btt1CXOqHKB3hb
rF8J9cGHyrMUdq1ATfN+KTdRjaUqct6zNEeZQxHlwek6bGlgQqQtoitupt1ds5nE
pbnAYmZ1N9+pDnOL85jB2vlW2Mp8qA+iMjo/Su8k7JM/j0SlqrBQqvAnPy5XbVJb
z6HJEG5pI6nHvYJJYuuJgzcKIou7oQ/GTdPLBwD8os2niY9Y867AQQc0Pbv0T9XN
+pSnOCeBSI1V7qnrTTEAIaUSDIA4gMJytvq8iPVtbKpC7XUxg9t9RuAGJjL6h98v
M7mI9wiMQznfEvJ5+zORscQ6WnpperDmo5c9ZXhOsU+SAorscROCoSoBdwk4ubY6
v9wB3NgNnKXGdIxeFEOfbVnL869ONZ2+ZmPVMPx/TDS3DQ02P6M32+aAsWV0PstU
ULny3Vi2ruOI18kd3W3k2MjXSiHpC2CyUo/C43DHRyU3mGFzVlqK3atJekIQK/0/
zGyXXNIDEmJC3IDznlOFBM4TlBFc8IRCVJDWae2omJ26+DVoT+//baBBVThVKhky
maI4+qfolL1L3zQRLg5NCt/YXGd7nfr2wkJHDpcxc/jlo3WDBcTPEf2uy3f+Zsev
hMjwlV+GolvwPEOCpqioT1xFEVmo1VjuJR03CsSOwN2sS2fKApVWoXI7uTYmTJ4E
ryLKl8/dQzC4+EKuxSXlG60UxYyprYLl9qnLsiakJn+mvkh5Z9jk+Htz9/8jMRuw
ECKmYg4iwMQIM8onKIeDkUAm1ExUJRX3I62fRCCQDlt3fCdZtuB6sBG9x4IXgUXw
QN7vXbGk91PtslCJ5FAIyLpFKmxmFc6eLjphI4q1wJosxUmi+knQBwv0ZFOFGxrM
9C+Smj6cFDi9JemkZgu2zD4R+HK1LH/Flc/ubrqFUKrH2/LxK0yt5OIkAeNT7vH+
78sWZhQnTiKmxl1NYaX3Ifo67fALsZDiyCNM/wEgNIsxydkPqxCbsHWaDhBC4WzA
rigROXFJA5ky0rB4znATYxO3KXAblifwgMsv5SI9ax3/xd55obGAVhxGeb51H47P
mVgniDcFANrsJ0NDvVQ5A9HqbNBVC314VnKA0izCrGr8Ske4/j6LW2Sx+agJ7swY
l1glXSMKzyskfdowFAAPX3WagNondRyx0C70vEWL/dtip2Vh46ct+tQeWIA9/Mlk
HuLc/YqKulQNP/A7R0BwLKo100pzTEkCGr1Rq1diOrZ+h5rOosVEeeO14hPj56Zo
nk4NYR8KGryyEGGNisu6TH2gniE6J9iuZFuHBi95hzEHkEP6Xc15F9qdaxJibmFM
jgiJ4m+G8OguKwt+oqC5Y++bsSktCEqC0aA9ks+/QYXpp5yO1hSSXjCu8SE5IGpW
aejHmTnV3fXqSn2h3oH+TtLcPAFIMVUBekeV1/U6pgGlSRUk55XO3w71x/Q/t0Op
p4oIwEB+a/vehQRMFR6xZuFXTkDWU8c/LiK7c/023dsHKv0w6f1bqY7ZP3VF3oL8
lZotrlEF2rXxkoSErCbzpQ/SidjdnYi7MbPeneRYr8lN3hV/qEn/vxItDBMGddPL
lFn+mguT0Uj5d16NG+8DvcXHGDtZKbZoqLiOVaBgPvgCRJ7+1dHbEEXjc8efG7jP
VLnt5EVg3vBfsC5KjGmuuH0ukzEsPtrDdhH8cm93OirvZGydT3UNVgcQoJtWXFRz
3RGkikPoSMtuDDxugfFPleIxN5uc2RR5xN4Lo4Xq2hUCHXnlkRm9ToLJ59j16F+p
z5bG7Vevv0Llo88G7Jc/K5DihpkL/2VO+kyX6emLGz9/1a3WK3qWu05Y1cBFYQU7
qaFxeFDtuQALvn9qYE2nfmJ3Lkw8bOoYO3eKa3T5t0hjDOqIwXhxC/yJGKIEwVDF
f6UoxOcsRJj7TWM5IC27ikq0em1TNMLUyiTPBUmgOLelzfIrOdrfNUmNRXLuuMhA
He5BpLbtBN2qSXO0Gs6RDJHiHZjTKiks3U5qgRNJBNldRBQe0pHCXElYj0g5dBI9
M+DkBIeUynZbEpa8ynYefXMsTyEApLJW8PPO+jZeSueLDphJ0Oz2IozaqmEGvxqp
COB3YBAt1sDxmGL9WXR0SWwylCnHyyFyzputlMm0n9hfk+ryfMba4XCLa93qZQTA
QT56DoveP2DnfGDbcHwXIJDh/t4Ma4fsHlXBVZGXnF/rbDcvYKOJ8vtHYuduOqzS
scFae79qikc29sLwlt8xQIMOL+3mj4AtOZZlr78K1/tszOhHto8IpXZRVq2b6qyy
ntytQleAhbD106MYGkM0iruHOZqjuc1SBuX7t/BKyh9pRl1+PzI8AtU/OR8XMLi/
aU58faceHPbWrxHkVXvQWVE2p65nKF+ZWITWhoxG4wcKfB0QfL2wY6V0MZ065zZT
v4TJSE5gpDT+odMIAgVPQ5ZXQikDTajFjSSwPKGAHGROnjeNUpdA5i4+H2UEDZVd
U92fC9saRPfJM9L+zPpB7CBXH1QqHdG+SEy++784pPNQNvuHSePjJX5Fq/OzYh8h
a5T5uxwvsVZaiFDtKeXqLsGmUVBLJwJgPT0dExnJ4z1nFaeKmDLh/hm0xlVI++1h
aM4kYkSxHrYzXgG9gJHmMkbHw1WcCJSwbX/EAXDx4cWqpijFGQkJa6lsanJzweSB
u1IjgBAZSkh42SvcnCZIRhfqdLa2yGVJyk21cV1qnD1RKPK5GMQxPxuT5Kpjhtef
GNSxK0XOBWTZeu2UH4EsZkg5BvGwDGix694MgsU6pzKNgWGQ71j2B90t9Dd8M0MS
clEIdjrcYbrFLEtIJAsLfUZ7HvzlVQq/Ot4jERoz1yU7QcxFhnPHLZDpA4TASUnN
QaUNcHo2EXvu4+brV2oUuRnCXVxQuAf93hDW1PZ6mGm0OeKHrRD9wDNc4Wu+L3RM
7aIjgwyzlsT+i94uTibCAwagR9xwaFFzsGBqC+kTXYYCm7m7wdhQU1JP80wgHGxH
OR3pkN2eUYI8QHBLFw33VezQC5fPg/l2054kXFtUt4OyNh5hM00iW+RJ8fJVTXtk
WLFCFzp0Kjlyqew8GFUNRmuZzPcbbLIq2N0Kc2nEt3dFSJm5+csmBHyK6XZ9oG7a
zMIo7Aoytp8Of7I+5xaCV5j2zbLdY10DYSdsFIT1ERhyxkR1/G2/q7+LfpalybwU
l1MWMjND+LNc5URstOUDEP9V0CHRww8uSBw4tobLIx6HqSqIP9P8fUy44gPWNBdV
rTTdDwsq5YqPXaNn8z7wFsDfCAduH48ujAYI4gljatEXPPUOCQhYlfctqhqu56jA
EpEw6Z78N6z5B7mJHboRCaxdfoAgEc/SuAoRtN33UmMBovUaGgyVPDcCVrQL4z07
zvfaerHAXfn9fxssfnznToU0agfWld55KcDYGS0MtS37JIlMmFaDfv0zXWG7MzXj
zolh2h/56cA5rLxRHePpuS5dGIl/N8FULVJ7qHNQCTJrjVuLLviBCL8DpywlptHO
Gs5Ms9E9cAlt39XNYFwGT8+65rIqCicHXflB5+EauYg8Kr4uL84n5LsBeb5W6c4c
1sJsRbbOc+sIi14/5YJPNp3xaAxBYp2dKn2QeGfteELDxVWp4DNRm2PObaF3Dhxm
bFdtIBNwX/jUxzzy+CgBJewnIyBUl3EUfyD+XgmSbHHYm2v6SuSh1Aitj+WrYCYG
qL4beYEBY8JejHRPdudPLNT84bG1xt5qfvEe256lapir+/7X4Zxu8unG55RXziNC
C9+7DhaGRnCyC0+Y4G1Tq7wesIfBILdfoTpy84tlmCZ7sZUQ0CqkJcgTJ5Uk7PUm
0wsp8Gf/dOcVIR3fJCxNINKkTKwsC1jVx1NzaIQEG1BAZxyRJwZyeIcUfL1pnQVC
mrobAAJblpmrqb665yYOjuH2TppECcHb/xx4KC8xH7mOJUqISCihSjFuKonvRK9t
uy4noBN7Qy77DNWml1VZRA0QynGh3O5sP3dR1xrx5ocOOemcEhS3zFV3/iSPi67A
zABeBFpV5244CdCWI4SL1wbBo7dFwGA3Y6fw8ck9G6wasyGP9A7mFJbiJEXUBBVE
hRYhMAHzV2h0DrBOXEBGCn3zZhF/t/9YinbPZ9rqm4sd30/hkIaDRrI3pAV0k+dM
NnZlUcMt4o5TbFi0hi/dHkHRmSTUo41SmKehLdaoBN3m0mkelqcGcNjpNlHC01zE
n6AdwPEGyiPFD4OEqx9LuUM/Ko79BRJyhnvGSMcwHsxA86Mq0DlNsLO/OhmFIQg8
cm2ZhayYn5djkj4y6Z/wxKCp5hXNkue8lRj6u7+Ig04AKyllf1qhJS1Yz0GIhRXO
8oBv1VCToij9NygFvfhTco/hT109Y7O3TSz045P7kd7cvAacuIEM90U4y9O94VnI
YAqi2fkP4KkS2u8c/Okb1XjWeUfsq8zEQoebgzqokQQwMGfPR9WxWurSn3qtC3NB
n9sJInLN3le6wVv1jslQY6T5jpXLK1oxj7QkQUcng0T4ju2ddcEoxqxTI8KPqI2J
6WubPcN/RpMOIEq3u3NoV6U6P84BkfEBTCJEcZmf3yW/yYPBcykJ7yLNAJ2FnjKX
zsqL1JHTZ0/30OEiSUYnBol5N54MQhAl4o1tDCxyvfdKJ5M+b0EyhkVAidvvRhHW
7yBlW1QF62IJpKnNH/GOIpfRLppS0UZL+hz4PCXsxSQ7OwgjbsJNI3hl5lsJN7Ri
fcH1mCIXD+FLEHfZAzekP3ckN7hzSSkITA5dgr7xUoguIDH71CbXT+gBN5l6b+jN
CaRM8D1fr90f0A3/zd20tYHAWm7e4VdjTLYrUMQ469Q3PaShLsCFuMrgRFv/bAUK
Nchz9rEIuoVCuuoVt9q42qYwrAgRLe43ruUiyy8ZjG5iUpqXbLAFwtEnQ4R8hsTx
I2+NyHFaLQexdF0uqUtjtF6PMQDuBo54CKlEjsIzpc1BiBLI7gJus8Eb7s+O0/Zy
Juu8BiUAmxjKs/JUIsgbXshsQhZkv61fpupjCuIgNmRuhcbP2xbUbIPQE35FUuCa
IG6WTUBhEFPSt+MCsbivM+ZLkBhuK0PPOzAWd1KFe3kx8kZNyPCOlPzb1JLv/QQH
e49jsmR5wtta/YS8932ZMd30hHhnXw3NfGx2CnkMp5APnYxV4kSIEEsavmdSpyL6
nH8JYR3YGxHV5iFESUJ/OxnGB1df/cv98UaVDKDEsdtNtwhAYLhDZriXEOPUaroV
crsVK9mSrvLE19EwSnOZc1rYA1VP5AWIZUrYoKW7ob3OHOvjqLzBHUgnJO6dRCUU
KdLAo/8P0TR3C5SZX15Fh67IIXfOWY871ofdwG9m8yI8Tt7cTFEE9Y1j/fk2wpz7
gTfyXDjeCZDp0ctSoFv8q/oiCE+3Nd6BXgRxUxSRyqI6aEn5poZBAWYK3G1VH+d8
99OBvFdyqXiRIBx7xWpCjzRQTSG6kJ9jUZNKL5r4aL9ZsP8ECbAf4rc3Mzc0xcbN
F27BtelRK47ZT7yzrekkLD59V4xLc98bVOd+5cm4It6EaIotzsXcWScDXaXXpKtM
wu5nlNTvQaaJe9VfWcjRYPHoAlgrBNjzS+/9hL+40QIR6Q3l7ZSfIHh664Z3F2cH
85qY/qHyJJ6b/Q8lXi1+44MCt2o9zbcMPVVJynnv5CFr2kue8jgMnlVyRk0J1EJo
1gJMgg5Q6QI6ElDJmdCZZi7WWyDmKMIcaI2Iwoh9s4lly0ddauO2r4q8UTDyueOw
BI+Hys2cRsRC4/QuOKYdatjgmXfOZBmHKr5wLKwLe13KxezcF+eAZvPZ54Qw3v/R
A3YfjuUqM9QaYsnnxdQDftqpup8rz9yFdeCRgcg+zRhljXdk4+SOS+wz/hkN+w67
8m9SmGtgYp+84fLfPkULIDkOxworK7no/XxRnbo+o+ghD8N3fZYzf0bkRpxLdwaQ
hbW8mayLBB6w6dqgKrXLpHBRWqe+jHUFn9F/Wh9G+76lz5/iNCLa+9o7OSKdlXOt
joo5Ja3wU50PHJrjqcz/d6KZ+bfp1R+ridoE7wcOaSzhiz+WVaETFNcm4lM/ici5
h2ApVsZ78+LrvDIFwZDnnpgTa16R7vKyElgU5qZUGLcY+LqaJmFtkKLNuZbFruwj
D0arA91Zq57KN2VU5bK/j++W9JtUo8HFWA9rntc2scRH3silEz29kwQ+2drGj2f8
o7Uxob4vRIJ3J8kzAwnAcLLEibf6ssdGP7w4VWqedLF/F4V25UD1B3+8b4SJo/oh
U2SbQIwTKaSovKO7MZGjtlNooXGOP6nrTPFHuX9UX5R6ELQ8A479rgeqM0Hiheot
QFt1t/qNcHrA0mT2YzouVKdrlE5P64rXkkviHT/gMApWQ6dJ6hqgu+VzE/0OGvW5
2IaThurcZS7bmRcJtcnmCKGcs0fBESw45U5v/8bFLYb103B+7JOLs3QyixHImC9l
41KuuJt6zjXwMkDRje8QftySyOKcbYICHEiYo9EQtRRWJxD4CRIRo2kk0j76ZdP1
FBS81mtvWfjsKjPB7ox7TGExl1uUN8Ft77jDfwYofOYK8dtHCqau59TmxUsFSAEC
iAZXE5ejzb32a7Ld8gfLT+rCIIvGWoDzMoj9BjKk4J9z5bisN1ln5Q2LWSCFt2zW
6wb8rwQymwvwOZe2fXbl/bjh1vskqpAT4FU2/EWZa4p0G9ugr3rM+Vtm+51Uy69r
7dgrcAPa5GN74O3yiT/JLiIOxydTylApvw6eiMiizvKCX2VWT4f9uUbaq5sW2Ds0
uklq5HTZ8fIZ8EHLE4dupJDh8R2pN0JPh+qLUBEqxI/6xibljG5tD4JsUf2z9LUb
nftooDzOR5ShRMPvT+jpY5FpMuU/NXLHYizNFnHdJQ6M31nFmZ8ME51oF4SS7RFh
DyQIdnQ8nfh/WHPSRaOePRne+i7AHc4BXG+kloM6ggfE/V5w4b2ix7hR9G0dJk43
5HrpoMHtlqRS014jR9nAiZp10nroZRyY+XNoOg5MWGRsYfzALFqg6et8G803X2XW
SFPtGDZvyiMZgWIe7evpJwEbu2AQhLJmUx//w359k7LCiBKmroNNpi8LogBAjpp9
K6q/RKDVDyB4pWLnptkDqkMfMLcryqgyl9K1QLmcKr4qNq2TN1OInopAu8wXVWmb
OjyPyltw6oo58V6+z+RYk0iW21AMCIcOPi2vLF2n0yZYnz9FwSlJyc7zXsnZiJLz
gX8SQKhICqN3Oxx4+MBwUdBdOMPEvk/xl0wUMw1TkReiURmsAD7JSMzLFolsDK1L
SDJQ8GAjUkwheJQZPqp29Q5BjMi8EdGX+gOi3dmDOURwDlMu0CEnD8EdfIczC6Fz
woaU+c89/fa6bR085ORtq3HRS9DLLT+Q+MZWpUq1gBPApjPJqo74x47WV7eKBf6T
yz3J/7ikHCmwRo0xzsr20yg0LPMXrDTxMyvMsPgCqmBhicpx3HVb1ifJiioJWv5w
H64ucLlOMQX3Z2Rot8w+C+G1eeO3Mqx78dh8VeviztCk7FqpAFyu1Lkd/nU+yKbw
M+e9xPg7Dh+2NKJ/jb9JeTfoqodwKQulN0pej2gtmyn2PUfgewltZL8UfhgAicR7
9ROYnRXqF6IVVcwcBrwOHYb3O5H6q+ysPuSV2uJRK24qZRInYBmn7QvV/NOc3LCv
whDPex5dOXsp7ynin9T2h2hIREh0YqOgXeeKnblrLEdAaOgakaMLXOUpvTv30zJ6
Ob+sl9hBuUtEFD997wLaGmUDkcJ1Jd3V3qp9/oe030Juiw6LyFlh/wtVtjYXCqbw
2Rg4Epqr7Ynaafw3gGNL4g3ja8Evxyi8J+pOMGxQQi0+t3qiuwyU8GBktQbk8aBp
kk6NX6aNzH6pAMkalWC6rN/d0RnHeqQ0Ivr46f7RtrhFgRW3x6QarJUmhoojJUgg
HO/F3+5y1UWSXdzIE5xtP9jVnRqdpCthTu+iFA6hSNSC3zoy9VVrjcq1eLJy1aEB
IKxhQtEXBzQYWI02lbfQJd/nEro5eO9GS0Nvk8yR88eoULUZ28NcvL2HilsPmvM2
fQ6zUhQthevdszIbpD9zMVjpj+xsr3D6JL/BBf5jMweYM7FS5zD4yA22iFO5rePZ
MOUuH6CH14FmIRU+QWj+rno3wZRVa52j/hRapH8/3BcOIf8PVCbGj6exNWroNOHU
x7Fv4s2T+8I7nTX0gxjMMyQekdcP0SntUneMOa2BLjOXjz4ZD1YifgWZjgGId54Y
SPpKplrQgYtOIjroZw962AUgd5jP5SAKBUeR7hlnjnqnFefQ9/p4nLAP+WKQG+UU
G3hERnV9AMIYzmz015lB//zEOqkuv8mxk3Rdowb/q6wOc1wyEMj298xxI7aKR3V3
SgRg6JhD5sXsPRlh945c+hshxaGtZV3w5/Ozs1n7EZIPIi1v7m/onyV5rnhzOixz
QvykwipIWZ2ZSY/FyVw8SaLKe3YYkEQZ4kpXuJeufJejIPOroNqLiryf2q7QYtOk
k52DHezwbSAS9pKlziDNF/zdbZq6hDveOJMnIXZ5sXxKCIjFOw7xAYrWmsDuMKhO
0rte/YXxxOB1NURfzZwRqVOgamuN6bC2osMMzXfhGrzz1ZFiF0B0IQz1Tbkq4jo8
YCd+FRFfnF2YsdujiMaaDoLk3/yMdaS7EdsNjgFmdd20kNDGXHXLF9DXXcPc8ni4
G/3/eURstd3kAYsVbR+FSSSG74ZM+DKHcEQmx7WdGNksQIQ0ZZwUPuji7SKZfX6C
30VM5GNBnkkMlTB/wA1S5BojngtP2yve99X4GBoTgyxqZm+jwLffnvlZArfGaCiF
t7M8XYwUIbvujs9W+2ny010puolvfMbKdZfbTlZGiMi97/Eg4hRGiKdyhwz9dJ20
CzFLFxFEmblLyaYYH38SohJFhjl6EYZs9ZS7eFTk9Qvb35u/ydAvHr46QFUVbBuH
QAdvTSDbwG4wegLRPd/wUspsGTiBsz88W45A6MgTFTtRsJ3HzrfDGLvEyTs4TtY2
asYXHas9XPz5nTPVb8q+r70Dyvg4RVhRN6mUH5RTugOv8K3+AfntCoaMtgx0WRSA
AyAC0rFjU6DW4/PzKDDihUOYPpPzO1P9a4yucE8pFd3/E/FGDgUEeHnj6cCa3DzV
Tf3nmk2w7+YHMOJ1jNN+/JiqktpGHXE97ZDoN4QCBkDDfw4U5Bz/c8hL/dGN5Vf3
Umwvaw6XXhvdR5nILWonJje1/Xw8laF5zbH00Cl26v88q7KMsVH56mzzSuAzftST
dRc5FJ8LGEbLCc6cw2yGLYqXNUq3GJy2ZBcFmyX3bbeyl19+a4O5ud293Wz4iZ9h
+ltLLiMQcbYaH5dnRpsVsSBmuGod77+hnZgkR1DZiZ1NsngLtmb2SZmWajCpEsM2
w+QWV0Omi5dcRhXjvDnTNBNQzydYgTWHQ4Y/dVmoxnyKCzb//y6zc9Frp+m6Jk9J
eKrMjESdbQP1qB6jS9HfsvL4qkApvgaSfPB6RYHDUXGtdkQNqSHpQKiULsqr/o3r
B/sHdv/BHWC/gyI2rgIwzNl23THIS839G3yw+CiwyA2eSbkjSAykXU9dMEcJxhqc
YBdJmal6HxuzbIJqRv/NCEzPKHKjvew8rXTgoqnH++HSSNLDVbFUr8qTpOVXZFqK
UItAbp+TMq9FUdZXtAorEHHsUhVU+yWlBFkhyxmXLDX0iLb/PFq17mq/f/AXvOwZ
IFrYidXfAjjowO4l/ObdefsyojIJI2WRadBdZ/LNAPiz18mxj5HHfmp0Tc95Y/6x
ecqE6s+6+IIY+YHG+SXMtJq9jxmmVIMITxN896pE5Dld13ajPL7RlE+dEO9R5WCW
JI7mjTyFblBL20zbmQ+9ZoIHSSaWLclUwn13H7MxCh1fj3rEqOqlmBBGRtsc08bD
pnzKMs6avKIXp0fz73yZeMJKoivI22LV+MZlksmiwfVkgCL1VKuUN/7ApfQmAKD3
ajC6TUwMBHYB8mWjua12tctE7nql4ecL3cIvgiI7QopNxoOu8jD6jjx/2i8nf9t0
Y7rFeuIYatjnH6YlvcPV0czUSZTreLXQdMsiyST+8Rk5Bt42zRtoKKCvDsHXQjvV
fpmsZO4/K9T+Y/rpYyj3xJ6LJiYErn7E2ynj08KxNnKSkwxmuIxK8B3mL4lJub9H
0ODa6w0G+1k+PuyUQToFC/3KJmPjR4tCvzf3ZnLRTzgnIRDUHsWcVMme3bEk+Jos
EP74B0d9KwlTqwlTOraqhwx5aX9R/qQghzYefhCGWH9HtG7I6uxFeaQf7tbA3Xkf
oH7RUT74CR82x9Kjgq8OwHiQmeL8u/W9hV98aSagwc4e57IHWJDxCUqNmrzBDlPF
WVMDV31dTB40EgyyI/fJuAobt4UwbBfanV6D1TzgGHGLFPcJmEhBTDRSCkhapIkK
R7ZL2Q9ve/RRESnCdKlePQuX1Qkq6IqB+AdnJbMA/Z4KqFFwgo7Tp6vDfQHkqS34
SVuugY/7xpZMczWpKWaA49PrTiXzhmISud44KcKxb9H3uxPTt3SlBIZ1QJXq4uVZ
QSF6VV7dH/JSJT0023WKxc6sTalIVIlNUskm84Q6t7kILadIBR2pkJJPMZBGUSK0
bjfG6jUa9lQ5Hs4QuT7Pk+d8sH8WvIY1DjOS2kP/p+ABAf0BomOwtzirmycKBsi6
wn5mBmQ8hoFv9PdoWdf6TamnSBgQGMjta1hoDvuBZR6w1c91/A/9ednfTbAMIRp6
rkMNk/Hm86N5FEtpd2ifocjRDLdm/biimeYYFn+yqh8CjA2JEDHhYFVZKsr1fDXz
cFugtvnEqHDsdr/IhxFhdpGM0GZMqkoc2OXDzTG82pCDLOZN8hOr1TtNcn6tAEKA
zA2e2XRbrcvnn47i6dE/zmEd4uftoKVZY4IEXduXGOHBt+TTHaCwS2G1pkkr6mGK
dZYZajFFxHw8UnBexKhrDWdEeK3p5B68KhiHTm3Ifgm/UIPAPj7opa+mE547Il3E
Drc+BbKpW+HNG88y6mf+Hdcr3wzDsrHRPzZ82ZTnq2L4vS0IQF9A9k0cb8aSi+/q
c7Gr6lfguoU2Wu6e7xzwwszydGR/5mCHLnSjqe9XbPvfnEmL+SpT0H80pWntzqns
g6uEl1BwmY35AdU8X5YCq8C2WkI/oNSUgxnQlNdJ3kBL/rfbJabPkVrX1YiYKCgJ
luVZztRw9MXoLPFIW12Ij2o7GkEKdx+CZsLqbh+BcBzJdt6SqS/Ho7Lg9MtTv+Ez
rwcQIxZG9Zkr+ndY50fkxnZzvvgHfXJsICDIZePJEZkRoxR7F1DKK+vnKZ8th3+g
iuMaR81JKS67ananJUg5m0/1JQpIjF+tKThqH7aThAcpKZQhApLpUm9LL7O9XZT+
Or2cpdoKFN437cXmNZ8FzarThXpmrNjaghteLYmBYQiKw970t1l9RV5MXRRL1syr
8r1ga1cex2BD1FkNmbwBxvbSRgdCC7n2Dv5PTQdgRYHgaoKb5KRxHSMTBMN1P1X4
l4fdPZ7q1bz68hwvWWfsPSXDK1+aoV+8amdZg8AyR4wt3A2MD6wyIeuskfWYXc92
QLJuF+RTU5NhpNpVOsRkmrM+msktJiBlRILKQBguZQqcK/W4uCE/fyy+JXbyNNGH
eJXEd11exz+Lm3Z+RL1HT8QiI/at+PMqXz1dW39xryuLugsXWoe/RbUHbWB3MaQ1
vktXqqNlpuDnrf0iJsMj0Bqd4aOBo7rgF5AvjAQundt4aWHI1f77cjvI55Sgz1xV
v4Jr7pkg3rbti136paiVV425ODpOJxQyu4CGDb9f1zZQYUKzUSxnAQ89R1jtkayB
75GthvtknEce67Ek99ZQN7PtViZg/2qsfVIbv94PMgdGrtJ/21kq3rtl2CeVOXIs
iCnW3MBLsHIxpr2VlSdXMYX7Lwsl8ddXhC2Nn59aJv7amfrNJGQv0pgjjj/Gxxoq
w4Bcx5sKLcbuiyoOJaLz3d6tAxp94J3oqv0R3YRmiLVlJw6mKl10eh/DVqukIvBa
A/AwmVkEf3OP0naau3DZiO9MhuXI46P6i9SGSKva9zq9AhYLF+JuN7B/sDyOOmoG
Sz0MnUHNIKhBVcrMnEGqesCHONHU7yLe/oH59i9WczUdVKGd1CNFHR0tswdXXzQe
ojnr1UVPcRZ2g7ohDT1YRn35kYU7EoCV4UnYrCIK6aXtsV9tyjxDxsx/RrZV+nOa
bWAfDYkvIT9ITwaxU5wBTqDCW8VeYYpDl8VPTbwscI3bdT1188s8i6AGnX7ujD5/
wPfE2LMDSK1Wkq1iPKDTjUjHa5IpU6HLrpf+48C93PUc8Nc61olvzlURi+0CnHUh
694QNohexboGJdbLThhSQzp/55ADnBhI55pqfi4glrirnM7IePjekz+7uaA3DHMq
aGCV8dgCECvx7HjAyEtfwHkBaqRNYYlGAVibpvXR+8beCKkztagEYNIbgH5qwqIu
sYZY6r583e2SUyKDi9HHkhRGrlrwGxEzCRDtWHrLsPIjTs3t+tmujU2y9CU2bCB2
/K/2jYaTLiXK2irWzkNQEBId0cgjs09KaroEPiQxAGplr1w8NAzLQQkZteczdslS
xAU+8qib1IDvHG08+roeLkYfQwyxQ/S0DHUNHZ2R7+c8BbAoy68yJExYMAyKJixg
LySPgAiL2LmCasxAIFZdLdQVTWjX5AqxmvLyAb3vmDpKrZ+g435Mk1uGVdCWTtOp
2puCugP8wb6gou/77/FlODF9339oiIpsp75mzp/spuqWPAyBOEsmRU0tLOu3RRm0
OHkFiWgV0f/EqYTZYgsHdby8SnLDJnOQ+6pG5RSzisCkkezZQF0I+SFxCUg5VJX2
XGymBrOKLKxTokOC1JEcl/MbWCqYsQD7Tk0UgShb1JalFBgS0M0+kmGN/Ec/UiPl
x7XFoAK0lOBNBoNlydZ+ffTvWnVDXTBdgPVBSHVD4sUXjmXiWpVw89hyL8JhbC74
bV0egLn6j9yRAXpigeEKLCBS78pRWnVxjGb0RctYreVIfXbz/7yTB9qyjX1dc0js
5We5wHomKB3FVHWazAadv6xsh6wILB6n5DTYSnjGqAg7Sm2uj6Ne07aaA2AByybC
hQ9dKHGl2GpVUhua37fpGjDT6ut1nsBKwJ141aK0WMdvZDA2j/CpaCRY13VdWv6j
OzCf0Z/aQd4zqH5gxbZEhr2STvZzlOnqdOA2WfILnAq4WZxp7zaaoZdgEfhSORfm
tV0RG18FgkXDG+T6W8SLmAtRypjspBLS0ILK2B12b0JNq/eicv8Yp1WCVGCUbmo4
lNRCL/ju8nVoU+mrs6GxD42eJCeBzVCWi3FI0i3PCtwC3YSn+N+4UdnpQa3YdaSi
youAH5qJieggygIrOrJjmOkrTCMunFlkCkeljt4j4jXrGsKvMUgcgPRKV2asuZf+
7+GRjDzKXrzJu5pEbzXDkxTDYWjP+knaW6DcdLg2/BzmKiVf/BoqjeeYG3Bm2/B/
wpsKrid0Sa3P+0xQB5S8LMiRQB5eOlY7NA4IJpOD0fpuWkg/JuVzKpWJi5e0Dmwk
j+IbaH4O1vlLmyHrO92A8Kic65QXgH4E+dVLDLf5SDPOoPbsy2YvLbrlP31RS92s
LS57rSIvsY2LYYfXfH3Xve/46a3o3Erll6tKRJbowi8r3ybRsPuHY9A16OhXvmrI
ji9ydpjp1VR7DDs1i8H0u0Bz9FuYGV+TdSPqi/xxsJSsRIa7C3pnAycP83LzWM5u
pyoPB5jBN1PJNWr+FxB/umm3hyljn0yx8RSELpBzXTBvwiQpjLbEBKFIK5bhgmmd
PB+AKNWWF4ARVqNlx4z4h+dtoppVnyq7r6zMiD9rBfaSP79KhWjvXJUN1jBTdJmN
9OsOE4pjhOs0c5bDaPbh0IV/ozf8HLsFCIFZ4q2fEJNVR5o1/NM0bVyWfSF6YkeM
800Kymkw/IW80kCJ/Q3rGO9TTVccInSTnJCyDpw5fqErjwr2/iHpuDsUbTyu7KO1
pVGU5+9+GNhUNJ5MwwefF0a/3Nc3IQ+2h+Qj++ocC8YVxVmeiujV7EozBvr6vLqE
+WXvmNEj5JCyD8ZgDwM1VNEcd4QMbVrbILBGzv0+dOZ7TgXtB9yfOsDQg9Hxy7Yi
5QDNjzr3yrBvTAl/iN6uUEDQkzAOQELEIIJIorwMeAZfINqiEWHTnAjbyVPDyAAF
fy6ThuhZvbWofsv52JGDMqCQP5EVIua0TLg6JJ3zPwS5IEZFNLhZyUv57nKpXDu5
h4KGZ556NpvCEVuOmtwRKwk4RQ/vf55wqyIg/HuGnIjepYNIcImWu/fxfwydW6SD
E+J9IDszkivfEah2uXo48K18niQ3L5+mASEv8rBZOCJaEzVadWJpCDPio0HHXEmn
H9p7N8DUs/KOKlOApO8cC6L2I/TPZBTSnFGocdkAr58a1MWXMmgyaituQgaXnQBv
UqOvmZ8Cisze2Fh7KORsA5JWMPsN36ACmWC8JRJ3EhIqI/F7bXOQj3PoAXV7fkw1
S4MONXH9g+Wsxb/72pbcrjGJE0157m2Agb/dtUeoJH1rtXPQjTb2omxhLrljtC4O
EZ0XFWWBnUsHVo4Va9Kjb9/p7YxqI0CJBx+7B0oGgvuKQ48pCxMz1LUCJi3IlrLT
TPkvfy+uVcMeLhQoZZVKBleB8G9+ZtiNpCZ/z3WI30g2vm86ByGyrSitYvIcQwMm
dB8cxlQwLBuRTJEkWSq4OCIno9ueJT1jqmzF7AEMXP5dBMwa3ILOnJRWrtz5QakV
0rhZvfv8LQCVWlNeak6F0WeRLbCUOvDMZWbd16tuPCWC8W0PSbjD1ktjlJjG6L6h
xrR6o6jWrLJ4v8+x6vnwmieZ1yyEO5KzXDXMV16ogWxO57mypfZncaum/ENgYK73
ZWyOg4VxoV+8AbQDloTR86aesq4m0aD4jKgXnzjLyXEI05Yz9skIEZ9WQT+kLp/O
0zfb2nMU6q47hcdPvPpByTjVStfPkwZ8Hq/xSJeGs1H/mt5p0cXKIkQCNuowAh+a
ZLFovjqPMpFtRr+mGu27QRnnfp5yFKdQmkZIHcpiu0fAN6CdWdY8Ywsu3o7SsTZK
mpukprjvIqBV3Q3R9YoJrn+8ekGx5INOQVHlO4PoVYBBTgpY0+GhkCnXmitbwTao
0+fwpcYhrHufdecfC2/jyV7qUpFDQDOtbEqVMzM6YElhc4gOWC6dQWxwtnFPfrrE
lg6SzugZH+qLrAYkmSuL1Q/c6BUsF4KxafcEKGnzC3TgxzUQ8DINcNpNeXGT/aEy
uxuusTOKIE24ftar3Hy1tYY/5kQrCps9wgl20X9IVOt879a6SLQUl+Nbr2l2UWWM
A6+KuxjVqlzkHCmoGrP4p/MN0dxdrnXK+l54KMKuIqJSvwoSgODrC8WUX5RhwKu6
zF04a4mcB0tShvsmJFWaCKo5QtbKOJol4krcCSkJUy1qtVFMbKyUsOZPAkFpYLAP
xbV5nngGLlhXtm3VqdXi77spk5C6PdkarB4HLv5DUlQwusTEVnrFYSakSTvQeg3O
8fZIcuRJhlttptxjK0AxltJoiXTHZIJDt0/6kg+f5ee/YN24vz/wQ0p4HJDvil8Y
TQDdyStbhuiD+pHMPbuKEzkyOxu/m0AMyWv+Z8qkWZYWHTmO4T+Yg+qyh6GQXVGz
HpI+uK3iQFrUZHXOqHruqLORFP8/CHjD3GtsSB9XZbpTSbxJ7WOGQyf25i2pPpc9
bCRQAgzlaEsvLT3HkBPwigNTp+SlgPLYcU8EsEC7PM1+qe0WdtGDvSuJqvgVB4EK
yTaiYB8Emm94QQrHdu9XAByYlpsC9LhMlei2hX1bA1MabtjzKKBAvln22yxSxf0A
5wqvy54PlX32XtUawZU/20s0PkhZfJfMlmMqxu8BdKDGyMpe5J+1NPcTXgs1JDVq
LeYw6R3otPjQyX2bgHR7npYDce/VVuyggKVueViSEaFIOCKbVtjHQ0Tm0H2TA3th
vNLP8svk3ItTynH4SyE7JX3pn5RSutU8iLu22EaFZPh/7FFWZFeD6F9hSG8ddD/p
Sb93QB1o4Bd8g5Y06U/bg04InsSJ/PZwCW0Tmzxw1RBY57+6Q8z5v9WRbGnKoSRZ
nbjKjL2CotfqDdQOD4id7mqdz5YQAaCcTYy4mbGEIL3bwX/CzO4fTVEZHKsBs8/+
MaWS7u62tI3gKISDKm6sz02ZEa18GYtdypRJ6KDwSSl4hxJGxyvs8LVn4MSlP1Z3
4IM4aDJB5cToSPEEnUPNpib0E2QE9ZBGfGBdHFpEdeTEsV8ZrNsq/u4xJLUeqjoC
Me1fQDK6ye8KNt2euZ25RstZ8vcI4JtcF6jG94LjHiz96l8KTTc3WPANoTt1X1+l
M/2NtMtj84gN6BX4UEpad+rI6hMhoRFInjLFXf3aT9PUadfQEjUobMrQAFOOj+ji
vjYWhjMAVUFgb0+tvh8YhRBsHf6oq8in3zMUBhzApSkJBkxuQbjjU8Y7sPHSE+q8
i6UXh/scjNy1SDPa22yKw0KFPAnoOVO19d1FHaqYUzkS5eHU4VTsf8mjU40u9Um+
CSiyrqwtSEArteCSGXqKxWE3TIm3b/gUbBOrUs0TWzARRSjHSfNf98XSBItpkiFZ
SXenJc4Ilxl4gtODCFt1RkqQxDmF0WskoklFIi1F93Pi8ZkgXX/qKAwDMHFizNV2
kqvFN25UozWepwIU1xmR59BN6rFmr+GxZL+ChMEfBQz/4XI6S4mNFV8dkxlp+pCR
XqRJeSjxPXMI0i/9xCTNoOJgXJ7DzhGpJLxfQ7RY1cyJaeLQT8VZrQ6DCQlmue42
jASbJTqUhuL0n9gumJqCH3eZZ0P8smOFGAlrWE5J+lbrEuRCkjd8iWj5ad68Zl44
7drFPN1ZDf95QUf6tM15X1mzm3fYfahHH2GRjzVKu0rTLAP26a/nKuwIXIal4ho+
13ED7S0WGQPzmLJJNegXtZ2PoNlCcoVlvaT9w7FKDvr0InYQocypK1mMjh/6590X
/xWp1Xmhz/ghNNWuq2c9CUFYobEkcx6I21YbEbliFqhiFx1QDaqYf9ySjSHdEkQT
Qdbt+tXbW9nFXYAvw5C9S8L7GsTv/cTGDXZEo9I4zOgI0YahjufhvtGVCTI4IHDp
bKrLJFMeHabsq8eY1zzTqkC/VXOQTA3yQxbmmmtzCo7SV2+IAk78uEe6sZSrk4p5
0H6KtM5kkVdYJNKrjD1j1yeO3BDzLHthzjtq79T/WO2iJorBW7f/Whppror9W2oO
YRlkmFF0VwUPQ1PlDPTnItpmDlCyOBnX6881Ceb2Cg8dtwFyVCY7d26OaB8S/6di
1tWs4VJIaYoTxYJWtYhGELUfkTpACc2qAR7sP4YEaV3Pw9xpT6+6CXk3KhoTTOcq
zrYRjSmZrNGTfA6P9Tq2iYku0JQ6fQhSDx4q5Qaizr0pigPk5S45vC9vsPb9IOog
p0NalK3BzAmHB46H2y9+vWhsy9S/Y9z9z2S5Oc92Ne2epgFyTFwjf5WIYB6mJc9B
xporctd8figtg0UOh5ltZGdAgLK4A9KDA8fkkAhp43Uc57rqP+huaDjS429LludR
JNP2vbMkIiztNswVzzAUyzBMaZvhJKOJHkj6SWHZ8kBHdF3y1/jW9E7XYF2Pqu16
eoEO8MR5S2oLlcck+49buCzVxebjlRoDVe8FL61Btk8uaxVf1i9gQBomxwZsGGVE
8RqkSowlAOAjFGRr7ymhP/zhxGQgj1uUK6ia9O007saoJ6G4ke7SszeRMj51zLfJ
pnp96UlWy6CnjXlh2lyNtjmpSyfieREXsr3hTisLiWR+CoRPwauPWntyIcTkHcwQ
k1oGjhQO8733ua0TsiTY56ETPK6bMj8lHI2swjJgF0TXcSOztwyteXkER/W3adk2
pSTJEuguWxzjPLAMbPH/WehTkWgj5vO28cPSc42YCfbj68RwzsdNteodClKYbXuh
q8NV7HLM/rQJ3FB6LIGoybE+JGRsD8ZCHeFz5D7AO0mVFZKtJh/IqycbJQEbf5no
ty01UzRKj7h6QnWdfXwo6McEaIdud2eU66nEOGRNTTIkpS7DsCXWDR7lppkkOoEU
jE4UYMMIjedFV0/m6Fo2JZXRCoELiSUDlLZR7QvsBpdSIaS9sk0Tg1BPQceqHwKy
8HCyQL2Z/JGDi+XaO5Pj5coo8tsIRFPQN4Hf+3uCekBlDrkmMmdh8uvcyJJxzh6X
jZs0CKe8/HFOb0Go4Hp5hiWEe+xmfuKpzGRqGpwJC2FJPkF4KaPKotMWteSZJ3uO
LwjH9QMV5LYjqKghpCkJ4uN6MTmLMsFntJgbRNd/uOygro+f3eVu8LfFYX06XZTJ
qrFCAc/Gis6JUTx1LAREzrew96R0HblQF98nSc/J3IgwkczQpLwHfhkb4u69NUWz
4pe7Fnk+AN/kmmow4LXY2grfy1NgW7Xz8kIMOzLEKXwDkgHgnmXTPrXqtDfuMSLv
gxhjPZ2EU+NZjbyoHxrmWUNZMy8LefmwSOKhMeF+I+UonHjtxfzGhdElalOkcG68
tAMmw0toTuhAenPq+A/zy2b+ewdo60EjU+QwwJuk7MYy8un2JkakUa6r2ZYJeOwm
R1UqJMA7eah809BhxKsPrHH6/0NXlpVC/AAVMxbDD+cERsltSaLIFy4RQDSlJkRy
+rjjvmobNFhX3ArdN0651Yy3nCWkfzXcrgCQR10d3uTuhI5rWy3C4TgY+4dNhFUX
XTOKO6yR2LfVMiBBvm5iYg6s3EkzZPuNt3W10Jyv/GjXVcmHhnhFb/VYGx4Wl2TR
UvdWF+wcfKSaTbKaaZ9d6VPZNaFVi+ixG1hdivrZDIWnhmctkpCkoTCg/wVhsk7G
k6Dlioqkkl0vQeTmhEKO0Nap286H2/8hgn40Y9UTZI/YuiKG8rLnoQ3ZxDmmbuBI
pFgDAl9ld5drs0u43UvFht9SBRApqMZiOHwHhF+Y4rz/S+jXmmiabcgNxjaxTlaO
j/WpQEwoO5ccEKeNdG49ZFjbpxXP7lckVl39PUYiyw3ATQ3s9ozmFgwhaVSlRMBv
10v8qyzmrSDCmesuLbPTTu9afIa0X/2jp+gr+n7Xz4Jm66ICfZoSJMHUa4VZb2FC
a0P2Up+lN23el3OwDyfodThhtxpCRlKjshcNJYKuHaGJKhqQpAq22Xqh8MQeO/K6
yPVzhN9zs6GjHKOzsFmU8ghEoqDc2kvdxIkVBd0mR/AAGET8l4n8ARPdxXtNQnWc
EqvetVPi73SQHVOt3YApVHGuxBpHo8nR+GJ9kJoEBS79TLFFIn8Fqr35keVqg0a/
q17UXTS8RwDbrq0mPp/5/OJl2rDnT9wQDrVCzko1kEmASXEOBsq4PEX8x85DgRhP
wWscm3IiTas8UgZr19P0odSl1JlOd2pc7CVNuoWEI4mP+nuSjzbvtzrxNO4ec0bC
KEQYGuffq55qwHEyKmZfCht9uxQdYOWs3HJPAZrIIqD9fboOqdU9KgEH5S7fY+0Q
fNfIyXQeq0o2lXPSI6bF3RqwJyuH9i8DgwOmqgF4wfu8xej0ImFlCOzBqlvskpw8
qU9Cc2KOuD5C1/hPpQXL+puXzqlcfEIuWQ/tpyDHq+DmhYGBEMT1Y5RwegkCRhri
XyGw28+LNzjv56QD2uxHrcQspWZse1SDRjvlDqRLdZ2Ld6e9rDMY/FpQkADIJXZc
cRPA1v92FsTIZxMkFpyG+OvAMAFZz3hRxHVJZ0DM43wOqm3IviEHCrNK8xrP6UCM
2KuFiED/J5z/U4/OpZFdHmghGVu333pJdwcfvSdlWk9hAeEXQBYVvpCrEA556jH4
g+oZpza5dZXrX2G7+WeJhmISn0KWvT2gzVut74DKePeMStkuMQNgclF0hdw4zVoc
MxIJfNk0L1Qms+XxYutH/KrU35cCn9AmIdsUbrN2ExmFPWgk2uC17Yww7MzKwGEa
Xd5kPQQWv3819/lYcn/BZD1vlgIiylBSllHcOh6Sz06wxhN+AOqFmiUkDeKMcE9W
kzK/jeEt2+n6NrD7qa9E0fZAhXBCA67mf1Ww9ql32TmpgrSqY4MK70xVwm0AMG8y
Z6hdu7XPE1mmE2MycE4YS5e40qeSqZlk8owusxEkEv30TiNiIa6HzklhyHzC/MEu
WqUYwXikHha3FlkdafM9wtzdDGnz3rdT+AIX9DeGmFIAWZNAVVaqfyiQ+mEgp7Ul
DPbOlgFHYGmjoFq6sFEMPeidnwTbBolXFDrBJXlRJB3DsTWLP6jCBpAN9D4zThiY
3pQMEkwWnRV3ByXGlzRjmVdrY3j0OL4bUb6ruf6TzwhwYPcGAtYL2uVOIOjEndJS
dnq5rYzzVODes0C9FIKCo3ynMsNtFxbqAkSqKTS279aI5kCSHjfJDvPqwog8Jsw5
NDWHCIq5kr40L//8PlG/39aA0l6deGm8JoqnT/hxeVwOyvCk4QsSV18S7gMh3yip
UJOcv721mXmf5DNxf0ws0d4B1fh+k/0oqXgSfCTiIfUs5ht6MOkO5BN4bQY/3SFk
9JN+/eM8ZUr+Gys26u1BiOxb7692OFlRiQx0g6Jcf+fnDWQlVmxsaEHwFbwTxl3l
1GDr23FGSm2BPRSYzuGmxO5f+qRnW8q5SeRT8fJYCtKlhvXVxC3VR10Iebk7yhNH
e/BFkx4fb6eb+Pjtnzpla2tHrQ7RdJQlffijx/Tj0tAQUIvcdYwlvQIdpV1QvzRI
BcfyBH2m8PfFRIsCeaTRWtPr8cFsLe+YATnJO1x50iXtQUq3I/eQ7miy2qBA1h0F
2vZNlg2l2ALEHFjsYK8xwm2xSWJIpH6IaDUhnfu+YoimPRt4jtON0vqXvRiOx+yY
9aDqsc2JCtuOMCj89IN7RtW/GXWU+C4Ic6+ztcGNHgmuNKUxrz98B6RsG7AXPxm0
ocpzXwxNINmjinqLLif44j9tKSJ57QnUFk+Ue14IXuU8Ixd/n3oKWUJNfUTrwxsD
Va0C5w/O9fkB1HM+YvAdeVsnhBPPwTS967QA9hqPxPjyykjOf8gacd3ob9uyQPGQ
26rAsXP05MaQ86POFrvF4IxS8DfJ6+fnjSeC6bxH7VztqfYrK35Hc9RavRpnyd4c
oRjD249noL1J+yVDoJRXS6syjEra6lrGXvBO4TNLxSHQsZp5Qb+A++WbsigkQklD
mg3usYN8jAChv5/ILs7Nv80bthA/IG9arxWHFzHN2EWkZWocKEn7PIAhtU67h9Qw
c0USyog3AIzTzxLV2+JL5VeIOhM49TaspuYroGu5iCpQTMc/dZ8EJqfF5wVHVM5t
mFORmJgyUXwD4tamzHgrdMSZ4/oLGT2GTzLWRVEzj9+UwZmpQq9ciDlCHHnJrUM1
IPd1/tBMtSrDT9PCYlIP2Rn84rcNrl4mGEcWFHvZmMc9LNUQ6zdHqXr5KmbTv+4c
FSyLLtXetQ8wv6UyyKY2OL5WseJde5+L4SKskWJSZ8a+j3n3nRThgj/heLcVmWHh
V27AGBol4SpypoATx/EXdJtBRRTz+jrEdsUdHvR6U9RvVXG6NGSadzYcJZbTtlMz
odhYdgz/op1iWYQ9rqigdO4h9IVSacmJBKQuYE98fvlaVhlw/APWn/wiLBlmZ9NN
fQ7Dw98BomvlL1g97B7FbVH1xmBQCiySFJgmwt1i8M0Zg3r1QxKcmBSJlEdgApY7
OGU2bT4ZK5uQcT+INDF41sWkGyKbdOhdQA1OJn4uVg+Mr/s2qYJMke9PcQNR7Akh
FPMm1Nbv9L2cDpxukgxO+5DDF809Jp4XhI5RnHHYTA+5VSi63YH85FhAk0c7oeIG
+6SSDAspmFhsU+xybG5pQ1kRcnCr/xAyFzHIrZPuMqrrkwfj0Usd7ePlepysXTQg
e9r+r+pqBFrjC38jBNTF46Y+KD6kOEIv3ampf1EvOeNSYm3nmFrUoYfCthPzL9It
zr3O/vhzLJtt0uS7YQtCK+vNW3KfiqHLEkuw1DeXzhLKBeBs1jQPPsnbyM9lwZ3b
lj3/owkyrmJUMucEt/2PojmgpyXHAqtStbgVcQcGIoKkdwD4zkDByLdj+JB9E8nm
x0RDQiHC7JOU1s9jrINHKkiDC9C4xGn3nW+EIojFYljT6kAXzAQhqLzrXOMbkrCj
kS0Vtmrdr3nmdTMtp0Gbt5giNPiZvWl4WEGG+FSEarogl6v/sFH4iDa7Tyw6GOl/
ZK/s5XqnoWDQqKxxALAHBt5CxkUuhdAyn3oQBWZ/tkiD62FNTT4WJJg8wR4WYPzm
2QHjO0wT+1rfceQDQthwW6OZWbw4MbfZLyRcVf4FEGg7CcBzetLc92CFk0KfU+/g
wXra877VUsn+2k3YFG103SBKHZOdLSkGmpIHWGz3Nsa0lZu2FrJSgaPbkEBhwoZA
hRl38BGZ4w1plkZ5J7gn0DmSoHD6Hi8zT+wbGWYUKEsFVS1VjHfXcFUHn6ARDg82
ykT+EvsnMJ82kw5V8Zz1d2STQBel+aBDG2HZwUTdoEHJ95Sz7A3r+q8XP+jLVfL0
neohw9qEfKByOw7D17WxzCS3IrrrVHk+q4zvyM0zfnv2124UFK1kIlZPvGYOilF7
yLkPPMzYwg/twvROzkB7IZYyOpv1N+8RzS7Z6DMF4P7k0hQSsfrG0sJD4npbEUko
M60TASg4R/U38c+QE2ckQx+7E1Dkr6rS8JIv1ZlRPQTtRUZd9zrn58WiIgHS+qUo
K4UmsEXFouT88uJnEB590PKjzVIBJ1TvMWcoXNXgBwSMCOAWOVaGLY+wzIV1s1I7
S6y1bnnLWQvH+fXZKe0u+hdv23XB38s4niNU0CbUHSugh8P7Q2g2InDDffEGt3ly
cJ63ZQLaBzdRV3HmMDFmpSrfn665vFqfmV/g8bl7JjK631/+1PbknbOSvVwWKOSC
2eaJg27IZoV95WYSKmLAhx7mV9rxNMdbsnMGNMlHbCSrBiPkx4bKWAhp2fsNduQR
qmc9ZFTVqjRATG1L3zpl+Ga+8c2tqqsLIBCL6UvqU70xWJQtAb6nCzUiC6LKlUSj
lO/Lmj5uYqd0s3ykAdQK9xrcBZc4a9LDK1NT+ax/RgtVkVf9jgkgAbO9VUS+dhHE
rAmlW1zc8QGuRV1dtdq2TdMmsTDPDp2FRgmda1T/HJH3hbjFlgQrCa2pOIBkzVIU
aRwaQEyvHLCyPRN4qN1ZmLAlL8NF2Dol1O9G4YwQQOKp/HQ5TFVNKwTdFUIZDiCk
uOqkN4fhovmuHvVmwns8NB6RZV8jPe6mJmE4NGHopND134+4QTOXSDhJ8XhuBWXO
FNN3GfCRNMmV64sqSabAiPdSYXuMRLutjXlFkcx9uAEr04U7o7dHZ0VZjVISo4Bv
o0bdVqLK1OQ9JAvA0cXP761JDr5bUzuwhDedPdDCh29DTkPvp/0ends0TSh7ECZM
fhDaOk1xGD2Wtcm1N1jrEiQUQ9QbflFdc8fAZgLDNwGjOJExCOH8EprjN+oY77lZ
iT7BcNqu+bLvFVgQLvwPNY62rAITuQQyl7Dk4Pp/dqAAXNYiTFMPlUJLa870dTPm
nUH6JNysRn9sTvCqcVebcQHS5flmtsg4X2fEqkbVgKN3kTTdoCMnJT0Ic0W/8Aq2
1hbArNa17/caOYNq2TuOgpeGwZxuP4KrKv+eHgl2/IMUwrLl5B3wjcI9/r1LTUYD
xOwfLdZBW7/a9fSbwPiG8VEL9q3FoXErnuZv9HTO4fTR9cn5e/8HoAM6LdvdIokO
yVGcNFx+r+vUeogcMdxSvvcHBEHaRAqqRG1JKYG6a70tO8wx/2vOsMPzVpAQigCJ
p4jB0e7rLdPqaGN60uMX3rtSwHXSn+ENgYmeAdhWGd5nxH1a3VBfYKNkEVGF936a
IXcSRNalmYI81m3Ji1pExlHO5aeuCTVwu480aiesElK3oL1Ite5zM3PoshEECzh8
0iI6fpwkDlnESqgm9fTbwsemqwC+Zev9al+1bBBQnmNVSxEKsr/vYAWmSPQLGN4m
hx54GVotK6PPVie2L3O4h3dpTW3zDFmeHGcYMSrI0QzMDUzGvt7Rf3I4frr2TE8t
z5+6NVhUkt66f8K+eqgvd/XeNfRpcOY92/0HPvLDKwv372fi5RB2Wf8sgvie5X2+
H2G0Ggl2NaSnA0zAAlgwHTziYDbpSwJ7UkHKzmKWRYyh6xynbqbigBdf317yq092
neqdWpFhNsrTemyBO43X4895pEpfSaBJ7+6UUP6/Ttc5d0+HPBfn13476lCrDL+8
A3iRAYMonShMojfrzDaX3X44TJy235jDiaxN47Wv8KMvFWZNPe5xA3lmNoIT6sDw
5wpuYssu0pWw7agHNVlFfS4IaQdZlbIQYOFEjxZez7ifTS8kUzGv0AsWh0cWq9G1
oxtZIcWqykhmJd77yxV4D19ptkN9q8ZxinsOmgAC5E9Sa02QUS74Tdr5eBbxFPLd
V+W/EM1sqMoJXgSfPoA2PTxmDO/n10w41lJn9pF5e/Cldd2jMKxylj3PkAU2riRA
PAR5Q3HdALe11JbPdI92XkYr445xXzpuAr08Ip3k9z2orVRUTQNWeSwtHiKDQApN
zDf1IuEp/m3yDYxtTlLlIGWUXEyPDr74zNbeSueiCZ1Hh4wQtl8F6Pf3X1uIo1W4
+zXCyCOB+JJU2KPDOXzdDcggbsAv3ef7AEvifmTW+I4LGywPSh0h0hxxnMjZniEQ
0LuhAEdFbVc+9VTGX+/5/bq8QmX+yejMjavBNG4kIGu4N0nwl+QxBtfY88TLgagT
WmLcMig2JAiahgBrKF9UU1jxXAHH2+3f8Aau3l4Rb2tBFGmm/kz9SkWucSTjnsGU
wn1m93byy/CfbAwO/zQml6tDk3Z0T9qQWYfHyoEYL0fZdMPuksCnQLXGfzWlH0Rr
JSO1QQgYyg0xFo0OXimathm9eyL13oZNisKuM7WwggCkGrmYLfoZrtkpQ6nAnAew
khYIqOSR05AD6b47Ra9o1TKDPV3apKW+GurJSTNHyaEr/0tVXo54fxY6utNC/zH1
bdltqinEhy1wrLnyFGzwSkuOs4wdqRxxnS8F6MC00mfNec5KXCrssEjbtaQd97wG
RaY7przaromahUPkMguxBwOKpb4LUoIhQaGbCGzhD0qAMyMf6iEzXY/UVTjiTm9y
piOvgnJPdyfrBeGxwf0Y2GmvKQzo5koV+tzbxNss44tEGsXeB4+vOVwr642wiQ0/
ibxwFf35wJOhfEdSH/vOrFAGFcfY/l7ldGG83LaqqofB1cfrjuMAqb0NGWDzP/zq
rFBQhg7KLRQQtg2mU+ksHNukE2MKxmyVXXg7ab7gg/2U4SCFHtsxTugS5Kk8zwww
xUtuNNy5sAY2Nsicl5UMOHt8eBpI8pZ9h48bg5bWfs7NM4TOqfkcnkuMcHBitDXo
DtZMulxMikS7ZO+AIsPu9ypu5oSOnfY9yJTEvAr0S314B6R3lK/VLxH8I8R+tqPa
BqnGsdIkV0ayqkQ0sHwE4Gq9KrKj2gJzNSXz7FNL/oTgVn2iQk6DrzysPnpE5sdX
76XrEQMBYp3mMdPrhvBbLJhp3qOWFlO27REX0+2qNR+m3AaA30PDG+HE82UBIF8y
53m2zG7Apuxiy9tyt7ARghB8hkr+iNuQY0cRKkKf8N7HEBArTYd7VjFSbiMzZ1O6
hfO9Nb5hMOI4vaMNetX1WM1NunES6gKn787VKfnukk9S5+n3W4rn6q2WVTdt2OiC
BwKRozluqTEYsmBUJ38X1SX+ZBe+4ccxzFN6hB1wkvAUphHFPnIGfJUO0bOvXklM
yq7zqlYVC5/NmaPUbi9rnTTkQy/919picsXx4QrnbBjyQ/Gh0F8LtusjQaAhmwWc
gzyUep1TMPDFyMCek3SzA7dASc/DYOuTLjgcjEIu4JgcTrwPmtnyqHurlPZ0B2Wc
RZCXHil6JyEwkXBVpqgfTTKcbxkKqsZ0iYhASMdCDrn/caw7DKJ7ArwkD/m3CSCq
Nm5WYY/Ifk1QJChsrwjT6NBsQXvZgNIOzyllojPU7Fxk0egfpg6KVfOOR6kQw8oX
DVKWCCxcwKHEa2uPI6DK8KpJMmKrDE+RyPWwqsjhD/n8YkJMF/VVA5a3mc2Dngjl
yYZRz25lpbR8GA6NmjeOZJ0ae7G7GYoc4c5niXyZCDXbnuX6wy0p1qrpVt9Y/OGB
NYCssyXpaTnnN91mC76bzMxC4EEhti9IP3NdJ+6RPt0wt4QZFcbYk5SBS7GqaeCO
GYPrTM+AsKKYtORfu9O4vEGSzZXpM3yVFSdF292/XWot4zXWHm/y1pPHI/ZqGTcS
0NJqj7oRQD1YxIKz731PwnC1RiyQsWOfxA3e2y7UEeIwDWjsbHORwIs8L/rVw9zA
0gcnZMOfx1qGiy9S+YJbaVh7lIYQO3ojXDkplDt3i1jhiM0JfRmlhQXDCEpPyU8K
ri+EYnYM4+CYN+8ZRUzBgCforaJzNxXvQpRVJ/0sFDdY0rssxX/wxnqLebugfO3a
djbAFN8gexrO66BssmkF0nQUBopqHXj6WCUVqt4jcMUfNU2ZA02bikOiV3JSVByU
v9eMfVo+BHk6IALopZOoHycAO6JzMCa1HlZcdQwx8IX2q9kPgbAvxIqJxn8PBGTB
qgh25aKs/l2u/tDjrSv7K5iWqQY7XtEUSwBD8qemEmTLthmBPg36XH0FW1WEeuDV
4weuw4XmlzXmCM7RWRjWbK72ZDV3c1L8EicVXqL3D8Eyp0UD0VcjtzW/Jn4HH/0A
EIY6PO329h9TdoyzocwZOA5kbF5377XLBef0ga7V8vS/ssp8I1m8QfCTSK41n5fM
46eoQDQ90EmYkOtJrFSFDo6ZmYHQO/mqnzeG6E9CutWOj74yu2hVw2kik3+JmsFA
giRLFRXAXn3Hml4T38HANcO6HD/X0RYWuoxmfJOp77l4UKCI8jBcKv3QSU+Os/Ip
N7HAaEz3y0rpKNOdofZ3PIInsbduHbA7phXsnKNtLkH4U8aFw3dgcBJFBmaTz3HE
PZTUesztNkczR88GvHb30/kjv8czUJrBd5LkKWaj1ndYO+8rpgmwQ1AERg3ldjtH
jK76tlnAFPLQinASLQqhcn7I07kKs69BlOAB3RlsuMdcFHRA8kgZCzyNCKAj0bS1
KexTegaMHWAYSyZT6I8pgRbgzogtx1IXXG0NfZ1f4huyrmGi/Ys4ww7lmjOCGm86
+n1xnQ6dC6mQ+hkHcDv5G4nlU5TrCNbj4VKltbPF2c0jOtJghqCpv6cCRIuPaPvU
vBgktyCwsgzUD3JEQo+ibCziBZyRNnXLNdz3NoaHFln5VLSgSHgXEMJaPEZ9JRTI
aEnW2cMe8GtachvXyBuMRoiRxg99xCNIS4KnzulK50pt+G/VXF+SYbxJX7ur7pht
K1A0A57vuVJXAeOxNpND9XZh0zkn08N//008YlnhXTNcVmjHnu1tSLrlls2FUANc
xi6/xo707iQDxJvKUr428xp24vvwMHg2pIIYdopZPXPLpIZFXKO0c+/qQwPh13Yb
V0wX2g9ETgB7aWo30j2CWn65Wio1WIWSad2EK7/3m3OruS+xvmXBg/HEdkJ49y87
xqOvDiWxuRU/dbPdL59SiWlvOfYODhGGrPslGpV0xg4pvFeNQFrmdn9yoo9lf22e
OSb2xL7CYpWRSx8Iw/JxyOt12jUPDOxSdkZsCoo+AoKsYoMF6gq7zEEX4gkAxdVX
i7FMf5wVCiG4+Te8S5z5iP5XnzMwXuXlRTe1OL/aRRseCMuOaSEoPPwYoS6JWbGD
4goebz0b5arWXBcSjyVT7Rs9zQhJHJ9Jlu4peYY0Os+4WXx897bb2ly0hIj/yB2m
KpJnZyD/8cHcAfgYiBFysx5tn2AOIraPNDscJMWaOhZtQ2H8ec8Ik0Q4aVT3EJ2q
HK9R6CfJKp+mnKRBs6FWHXHOrl+QotfANZFK+PyVqQ9AAPgc60qTajL3K/UC70Mv
ICZ3oHTkujnF4GCNHvmQEvTOcm0sqkw+UZWrXBCvKut4Q9syHWxmamFhMUqsMlwG
tt05ZWH4p3FDs7bggSgXm9vb1OtErfF0RLlXcXAxSZE/jAuLGtkqjzomZEmVMuGJ
OjjrKZDPN/QfdzQzLZ7FJE8c27fy2vNDCQdpPferk/AJV8udnAFw75WL+LW6YMt6
87Hn0OTVugJM6ZKL6l5H5xbSrbv0YYgl29oIdsBhkhdY6Vog+D7yIfJn95bCGXrH
40r1y+f5Oa7yVJnEnvvav4kWpgolkQnBAjqZH2MXJCYHuIpew+3+YDeGorskmYf4
7UvSPpm2YaR0UxZIvgCQC8JWS98BDz9gp/utfjLPED3yo5+WiBEqez2xRz2HEpwa
vcIqK+2wiKwe5gRc0+51lI2mz45lkx4jWYu8PEDkqzS+GRgVzn4Sue3z2bIO0z3S
HG6YQddDoOtlFknXwJuf0E/GUD2kY3HA+7dyaA6Bf5wUTvx8RpLB5r7VFh5dpcU5
7QwXNJ42JQon1cjWsnLR7LUsDbqlnwbxppGlZmtNTTzBO7bHX2KrwL3+AuPxXw12
ieJxNqBTEkZVNYQ1bKaCOOzpup5PxzLGOhgfyrvNoNmyLbkL76UTa0ql/fe1QHeu
hJwPXkWiQRzbj95h6c58vgJWGoW9T4pqLk9MYVqdpAqiI/cbCF8y4G5D4CyVXblg
onkh/GjFet8F5wmr50ZgesCVIXbDP9e4tpqgZdamv6R+ZP2byWa7VBFjo+joVJ9b
hVVVIq/mCSIx5mzNhHP3YL4ps6yrOv++9yc0G5K/1R+uEMoWtegqJ456HBqKXIqJ
5Lf2GxmL28k1kTLH4896Ck3ie3bW7VzNX0W6IXby/IfBxsXck6i7VWZWfylbRVSQ
zl0A8bZD5cqDaBG9lER/obLL3SP/f1Q+OzVFzQiAjS02+0tMd65QT1o0ojCzaQqw
8JTUTAN8Cl8X/nrF9WPUJOYO5G9yNPc4B130yK0kQBl0Nd6V6JArQtLw47HjP438
Z1RcoG/+q74OnQNOdcyaeumTTTvecynD8+ERfOTsILafAm5pKaI8tkVNzjNww8VL
sWxZXfW12iRpc5py2ea/AhU/qaZBYEhJBd2zlgYF5TzQ7ZrupEMQNov/oJnkJjVP
w2bF9HmrEQvOEjhHy8DymyuT/UWDA+YMwE/y1hGsV+rMd8q+hfkTrrhvM0XE4phC
MojL6+7qwilSwThfIfbBgUCKC+yZP2+75I2RnSPfbm5rZhaaLZi7Pcishk7LdRkX
ISSQEJevSSH8XD6P3dDSdV7G0Hx3yiU30pB5iWhstPYMwJvqWqSkirVf4lMmJ109
iHe4G+sytT8Enj+y0d9ZmB+u3fJ9QCs9c2KFTE0EIsvD+MURzQOcHn1ugT3Tgu7l
IiqB2XYWdv5bPln0RP86fg3HwMa2i8DbjS9SJxM7haDPU8stKqlz5IiH2Sa286Ij
/bVYoqAJVe5C4bSqsodc2JM9ZZ3dK33xeXxN3oe1/qK8p1u29xvVNvDVKKPBkFXh
JB6gYMK6zORSgDXWk9DvSHciS3geQznP2Rv+5pXSuqXE00JZUP7SVFxt6fXJXwo3
a0icUb1ghgLRKV41skaXtXchHcgp+fOjeUNn3cSw16AXhljbcSqYIPB9Itp6huFl
2tYxyvtVobSufZkw6wdoYOeKgrFbwlrtBeDGjzJ3DrRKTDnooUhf3tHhlIQ6Jpgv
4SI+fAho4XPiDZYJXbmLMXWeqHX4kPMk+7XSuLJTACLkJ1XRKA2hJqjxXbt1G+II
QTLR8eu5tLY2zcbxabwvzS0Rq6zbG2yODRxFOSapNwzfM97iakBZxDJimI+hOiO1
VoVrNltiTDyR5hHpJaVLAEn9L7NZAPYdSkz2aFizBDulBc7ylG7pFTvQMGrLXcZ3
Xee7hlvz5SLgGaTYkbqiNkJw2ZCVGm4YAWIQOC6ekXqRq5lMquT+FE5SzCFidb6/
x6eZA9juc9h4rRqPkanFlNS82ZnOa9KMuX0sG13P/j6aWiW5uu5QH1B60dwA3g5q
eQUiw6KNNSqIZYw5AHgqo2XrZvJs8RdR7QiXySNXJ0WzVgxCEJCWXhcaWGIoPqg6
GcKCcCPiVMBqQI1M31N7fWULM9pppjJ7t8jY11HPhtwNDps5oEtT88jHKU/NR7df
3gcIjaMW3a5+fKTwr02wb02vfm9KXYdwh0pqgC7MpuBypM47na4U+oSbTKXnlyT1
pld19tixadPofv4AHV+uVWl1QmP34K3a1lGXUCKQyU75MSBLw+vK6awezODJxQ6Z
EfhI/EMaBBBigfRJ1zqRysc8ewJwHhLKqCSx/S3LGNDyjh8zYeIQU4iH30i5RMZf
pu7QRJ2pUiMQHc8VTiYosoqEs0zN7OaZGfqYjJj3ZvFq6oYu4umEcStQWJNpKYIN
t8T9KM9uuGd+xK1F69wmf2Diaexz2p3ilpzGp+oRwPFLV484ADM+FY7NHCzPy/of
NY/EgldMVYvwwXpiDDO+w8zaNhvU2kuAchUJnjzdgirFJBjOgFdVo9Q0cpR7m4Au
SJYHIo1uDhdH89gb+zBkrGWiA5sJptr4kWqcKdPtE/vtbC9PudZqNLSL1zzAlfNh
GHuUrhDIdemMdAmqG9T4P6CIzQA2AZQq4RsEMaRsACfAA9wq8+susMGyNbDgzXPX
UvzE5j9klZep76GoPv6B3ofDD9h6tCGwpSwl6GJV3HSZ1Nt2+ETLr7Rtx9AQhGXM
ryBVvmoNEbaAq06zf2Rvz+mJteW86Tp/Z60lcey97InzAwypoh3ySOc36e/TRrD1
cjTkh/hLMKhmIpEEU1G8o6Y4lf7tyZ71u9ARxPFCNq+0ts9WCvruGvmuo4t/TUSV
XYEM1oBmTKItMXSkSTxVSHqZB65C89Jfqax6lzMTuvwjZttSHJlPlwvkNxw+Hsbx
kJs8D9JHqrJ0On61/54UzAxPgZx06a+7Nnc0qtMnmUWOr8f/vHkrA4HPfMsiQydz
PfvrIw6P8qRsusN/gLSXQyY//Yl1cvmf2DMt+BoX1Qvgs3SpXsZWnjk+8G7oni17
VaXidI7hNngUsRotEuHo92MueS4Zw1a93KIW4aHskcOpXTeWws518R7U5AjecCNC
4oEBdDj+ylQukJcKYdKuHClYlSbO+jN8U/4Z/RZHkJC6EFOCVPMWqWVjwmqM6p+L
IJ15q9U9S2VP7IPxVT+l96rEhnQ629nb5t/I761OwfTPl1Velj6Cc0VM8jV9umkk
FniBtvrvwm0WwYSEwEK0kpxOZw32XgnehYCFKMRbgdySKj1YnG0TnCEmTbfR4mEL
vlOcQ46Cfr9c39qMvWrrjSZzqeKantZodIUu8tEZXIDQREN6I1p4dLUs3oUa4ekM
3Ny6EBAAMII4O1Mh/TlMVL5Q+XDfkeHs0xdbLVYxWn7naWEbnpzykYqFU9FdbQ8x
EL8BsuOOTgPrNrWJ1OAWoxNVW7eOlasEHDgtl/SpjGHPYqyiQd/QoERZaTUW40J5
205MYEOyVHhudtCb7YXzoc93+w+yTgDXGmlJeZ6+ZXFBJmak47tVQrfT1BYVow0f
H8+HVsrx5KassPW9lTPQ+tLFilkEcS5ybBlT5vLkcM6fWKc5Y6iXzb7/bkwtKgaJ
rOJ3zXWVG1iN8innV7eZqhcwmXxZeFopN6b4WCWiY107HaQgwh8HRE9iBKK41tnX
meoLOTSXJVTL/aaKQLxtovNRfUzZjRB0uU1COjeHkrGguScudum/16T9NKnLh+KA
oiP+xkjdE1HUiH6siE1PuaAFhduU25eXJ8LiYOGdiuHdSoQDzzdn9RY0PWle4s3r
ENmSvYjrW9kVWiE60v3n4oj7c8SxykW0v3+XbzuEy9WKrRPwqjzR3jKVkeXvKr8L
3+l+pLATGF/47CKF5fODT2W53vnWLNhPjw8nS/9tCyALaUg5Im+AEsgzj1nohDP6
eFnROA6BDJy4kQYUD7XDbZJyco/ruGC1/4qT3l0iYMLkfwzFaA3Swsb4AAM1x/H2
41PpWtPqx0exA1a5YqP3wteXjujLvqxWqOUj2jv8zaKVWFXKd0QvB6CM7tLEesre
nkpmsUaz9huYCp7CTaGhzTTD0s2A7QZiiiaGLD1nY8keVg94Ps2QMIuRZBTE9dSK
M3X6vr/Sgmj8kwwfyZD0MBHtL1jEuF40FzBoKxJ9Tqju0H3IoW/f8GHCFYbn0W2K
Ybf7RVzCuufvuaM+hnKRsSsr15JcfYaOVbLx9LMpYIYAFzK5mMkfL4HfwCCiqXOM
AZNQfQZ3G7wfYpnB3mcCpQKswU/9tYlvv3+bFrVQcTDfHfh/+xl/QEzgxctho6t3
pvsS1VXKXXiYPpJfDV6ejgrkgO+jX2B58/hicFGCoVwbK0cyYGjp08TW4AqUeOZj
T6TmR/ZqXHy+OMnoQFaJi3d2doFavOsemMYQGl7INrHa7iRXmaFwNB8XKriB8Kj8
z9NXUTwsLNnfFr8PeKWO0V8AkBb/7WIbWa57x+QGt+gZ4xNvOyVn6Hv0l1WgkBlW
0exdrnnI2uR/BlQrjkDcOB8E98gNjrcB64+za1Iy9bgVFioIg9ToFWaG10E4Py/1
5sxYLIjdUByjIbo0AhsWEZpR41M4ggt/iYd6uMeVUYEF+UCjJWp2eOlwmEaxB760
JjtL0afEjAMhiw0mMtNnmul0ukz+uvP2IOL5/Id4+EEElYp2a2dm4wKGGj1nBnq7
fkt51YEpzHGNMtv5HfAcplPkEnelk4H9ZnsmevWGOPRKBXZrilf4+PMv4NP2d8PQ
L/MYQQn642NVPQ/tbdFHboqpaCETnYYtf0zIIgpXQFBXTqfv3/kasCxraWC0V8yp
Ulm69rIQ45ysGzc54r9TAoTQ/Kwebew2mwRrswGZfeBXazJBG9bwnIKz79uTUGZe
b7k1bhimW13Y7S2Ahi/5N0drXOTz/m6ZYF3qoKpsG9jDdv7sDkyWTc6vG8rN8XkR
mAf0dffpSEC10Deh+Cr3fOrHu7KbX2ifGHmiXg1KarmkxaTBIZUZpWBIsHonS8r2
zSUdNnOznVueEKX20n8ZNAZn8Mcjc7knjBUYLrh8bqvIM+nv7Eb35hTyjKuQStrv
v6szDpUeSID8y8Tp4f8d+8FG3e/CZfpQpAkuQC257TESeW0tx3iwYShWQluWTYGx
H3S+IL5yaQxY7CKCQZ6uN0wJGWjdGyJyDFUr11p9tssX7rcMOq8befAd0k3erani
+DSKlzjqXPLmX2dYr/ZPTBuwFg4FtNVProshxymAj/nxHBSX+9j21Q7gUR/NMJoE
SFGgbPFq34r1KZ7KqPCPHmpSG7IHn+rGlT+DWemvlNYXl6uwuHXlW1X0fsuP03oh
pAc+Kof3TXjqDdYKHSeq5VYBDfL+KWKzms13IRQCOhRrfkqJnKEwfzYBUQfBseP+
oodgMtPEr96pF8neMHHxnnGmKZE54MSRhXaY4kM/y1qeSFS1or8S/ofEL6R7bbmV
IdPCVMJslzPzYlRfVURtxAMVAXXnzSAWsAUauvD00xwpbL1d7GCWD7RfK6gUsuRB
1N84u5MWgIouRaijWwSfMFcgbTBbhTzEOGiJEKwWsf5oT4QE/62cj0tCaixWoVcu
chC2lSj6+I0kzxv2+4FrS29fRYyiad/it0m6V7gYni8QqIvdWq8yHh2VhS0DfTSk
F6TNO7sy6mi26lmalKm7cdqmTSP4XNFl3gIA4AA6U2K1koFLKCNfutOtpWUoAn6U
gWeAu8hHC8dh4UgrUoCkZnz5Mzg8GDX3oiEs4g9h6Nt3eRlwYy6A25tY5Msl21h+
qoKIsX4tC3pi39PSsXPQi4dnIYxdxSPcySws7nZtvr6O64iySGOjlg7qVBKjsLOI
H1NV9DIMtcXB+vm1Zr4HKh8WuxDAqQvhkva1kGxsRocH4HGZyD0z8kSRYkiJIfSz
FbfhBHgaIX2pP5gYAExIm9u4vp9WAkeJTrlEJ34oF0cZcygkaBUoDtl64JEh2ToM
qfdhcXm3Kh3cmH+Mgo2at37F/coXVNApoAvWquk+q7OWuKQgHDgbFN3QKPC3ZeJh
ROnJAmwoOwk2wCoYaZRwgV3os2lB99YDC4HM5HQH57fWX1M+Kwyacx3TecQHdSWQ
7eLgKngZTPhl5LEom02eWB5cuK/oJgmaFffm87c7jZ4TNwTI4jdeRJ1z1rbjVE7f
Mqtrn81c9ObwJ7W2gcjePvbHJ4hE3AIS4eyqfv2N5K1BlbKm1LMEm/15y+81WPeA
womTmlWKntF7NEB3xhvNb1OdUZyqV0Lpp63WqKFWmXE4NOv1lvwLzSCNttGMmxB3
zi4iZiDb2h5BnK6hBAJ60n11A0NmfJpEXpCkT0g7KSmJlaFeRxXgx7xG0R6m6gbc
QS4JxULhrqqU4jRRdEM0vqRaqb6gGDeM9oCcNYtraY91bHShPij7yesv5tHjCZda
QlL9O9lid0hSCUQwf30zaT/+oS5h1y/4OCWdr38spRrXqYMbXNNKTRoFIya3f80D
RO3Bm7MsaAnsUCb5pHd4nJhaaR+37Bf7xd4wZwZ+Q69aQvJxsDTmNTQ6ofuOZVcC
FqN5PA7gSILT0PUvhmipFhZ0V+0BXi3L09B8DeoDIUQl37LcGhdOqT3kgS9J1b5e
ivlMsc7QnMZiy4YJDVtYY8HClw5ZPlsZoX3wmh6snExjmjpScPrLCYxf8YHTYFYp
H1J2Bv6seQIQ2pVRvSq85vfYusvBnSakOV1ncIGfvKs1GvU5Ric7dmOp13dB/8zt
DON2m8Mfd6QOSB3TUiggvriEF6BuLA0BiI5dT+MXMMAmwtvOL+ThSbCZbELQ2GQD
sySDGHRvyDM88XqIXH79yXS6PV4K3xrM1bM8EXiO4gFMLESSc40BL7lNv7R5Qg6i
4TU9PzllnfewtIfimfoucIZkLkkfC6Q5R9tjWqjR0qu6DOctoEfInzgnU08TZ9va
JGjeh7M4uErQajA5B+oqj1PwPZDaUL7/Xneucd+B0azzaZqLqylmYgt8fAkW/BTR
QySwGVNxwfs+2/dOfHo/IQTbTwMTzYFsjy5VQOba5Ym5OvgncY5CrNW6+By+iA2Z
pqNLThzAkbit8gQPAa5rQ9oGhohV1kMGb6TNYqF96I4FtA1Y0Jw1z/QJ1o4B8i3T
9q1hMcEPCIvoai8wl+2keO9CeCsOeKAU6m15Yz3iMVEiG+cMMDn52/zSgiIrhyH7
kTZXcJpBLlzjVPtqJEzPqvpFIim4JQyoMKx2+egHHY9aZqwGnps7fw9DBA8eN8uy
ystpyqfQDhwsZtIbhEm5E5T6973CzPBrCoEf5xJ64vbeiaNyoc0cqC7lS7iiTqLD
pnLfLRqTKtAdEfShIesFQUFSRMw/lMeNMGUrI3w08946O2/YnfdJSl3n9BkbeGwx
zmxfvXRmvqzFrrg2soiZbwi4CvFNJVhjcEfSNr1COy34eAFaY+OI0mg9vjlByGVa
4XsXvVwrTOtlhj0FJPF1yUQYQ6mjsilMNfBPNA+yRK6e0KWxx/WwjadDKquxwKm1
3kHnt1WLlY2Ve7sI94ZqDeqv0Iyg7zfDFd0cYdqXOeJub6P1Czwp5tjQtOhjNIvi
LffHG8dHmbjsOYZ7Z1cPxk7VCCdMv6NHleiY0J2R6cbtn+v5stai8A/peKUm7EiQ
tfaQS51B30wxPZgpdGQ9gcAbhMpVjm9+HGtHrcfXFAjgwdS1LuUdwYF1RRIxqo3k
+O8GUPD4finOJVShnAeLFgfdDNQOtmmiK0BQylrfEyPfuG/nvcdtNj5xuXeRSXvI
YRFogEvnjKlAZNJiMtrx1tTOdZEtI5MUayjbMSSoM9QjdcHK1aCk5+xr5+0dnmNA
DZ9BrA4iDOkHP15mqNecmpehVsf56ZMRTbtmKNf/sIKOeoHUc1rhRWg8V5H1ZHKg
un0poYv4kWBVvkPuAGut8GCrHca0Fh9SdP1I/YffjynyTcxFGbehzuMhs+Y6SulF
go79VN+/t1vj7M2jnPXbxxhOCuo0neDGQ7KCQ8Lipge0JtSZyJmGD5kUZi6CnJdX
27gFZFYs8OW9phsbgA9NUxHl0hs6uZA7dGR+XVSVaSf3ZR++ZbL/+lesebW4lh5w
E5Uxz4P7V7hJqn1wuQlERGbPnQg3xtpiJvDquHt6RaWrfnCH39APUCtAKovVU/ro
TwMB70t45JgkDsZA8N6C+iJNs0h8qCIOWaESgEieZOPsJr7ipvH90rmZYxdQaPhF
IvZi9V13pQIcZfdSc5U7LGHk9gnRNg9LEsUi9fmNb+tECEz2Dz/9/2lu4q5y/OOW
JbHg6CtYFtos5pmQsuLzR+nmMNvdrPgPZ/6NuFsw/lRM5j2mBskc57+6Ef4NnAVM
LKX2HRS6gosGbRLyZjF4UW2nvz/Li9sJ+SdES3QKHiax00olx4hERMxvfEnoiSCQ
5v3V5lly8m2djYas1OD+LIVf2KBaoZCWiVVjfgCSBAgL1UllOIIzN59MG1NoNs8K
0OR7vmWhqttL48EYVMpmKearzbZSLnSM6nuwVHW+msDrha5cQjRtzrXN4QckYidm
81g8LUWxA9p1HMCiH7latJ5W/r04bjkgjjdMFuKbCGYy/q0HUIeiGqf/HsbI2ljX
uk9H8zdNJuK/jlhRvKLtpFFC+b1/AiT5ZMBFRmobUfd8DcVAvy82pLn/opK6ZWBc
5oxDZPgQphQVyV2LixZULJ6q7h4mlXPkzfw0yqLf6GujRD8ymmwrCMaW58q21xhd
df5T5V4Mo8OvakLauTMFh8OqkDsxw2LibklNsk4vJ3mZ7rz6J8eC1SqgwKTbn3rj
Fd6JhrlR150Kdi0+g3lWt0MCd73edD8e6m7z7sYiSe8A1I9qGSiiRi/Lzry1h5Ng
dGsWsFFvgKruUQ5n/a8ym2rmQnM1dSHCKyDNvGApraA/cISMlkQM3HgPodMJiBL8
18NWzRwgA9v1K7hwrJ8K8mCq0My0DF+uEhnXyoFND7cFfw3o/aoF07cJCapxBq+V
M5Jh17dFl4KlPsJz3rpmYZ6FK1/iBoI+zee4t5Od14rIyf40wyx1pAJyJryY+HE7
GG+20JwYYClT5mLwyol9EZ0y+jVtiWo8TMl8jAbdVX2E51YGHn5l5RtxBIWH6ZnO
h45uDGt6/m+54OKYJWWf6Cr6UEWd8CCOpx04VPG3q0ubrHBQKJwESTw7HVQ3Rg4o
a6pWZwqqzcXp3A4gVS1Cyoh+1Wqnq2+mViUgeRiOwJ19T2uyon1aeHQc4ZxvBGRG
oYuW5rXDwAVMresbP6RT0N1fUBFJQWHoSD7FWxvrAmf3iFgV1lCCJPw4OjS8xnW6
Pe5WlBJnqPxzIVdWOZe/o2dsMvn05F2WeNgjjw7JP1u065v/mJ5qCExTuddgG7X1
e1GkLAATC4hkru9o6TWHjbcfMF1oIeGNgEMidluyQcxkAVBihQwwdM0pb3/bqglH
wOfUGoh9mI2NP9u5GekQmwokIgo7+xMi1vwa7Fa8YywOvhKNjpRbIaTbrrxurQpn
I0ayYZMZ4ZPSQFnNPyj0MEekus6yT4RAiwtEh7Bts86/pPXOSUwbrDQ9/d0eHzt5
RyWgLZDOUaXwwEOZrmpTgZBASA+SOlhM42ANSo3tdPbImaIbHW5vEnKgLI0h0Ivm
za4rigmxOL+tPuLqhUD3skpNxKt9amY5y8Hq3KLQfenBCjWnhs3tXliNlaHRlfNQ
Q7hy6FwujVQsON/GkQ45T+P6k00Jg9LJ5060MamKoXxrPg38AvzV0yTTpYZ+cgLf
huirYA1NS87JHJjhLEaF8Nk8bNR3xX/UPsFujNFtRd+MMZiBSNZRX9zqKLBMQSRZ
iUlZ3c5sR/RgKNYNj18KbARTfGoDLmy6hySp0aTCutjHO5L7gmemEdrqLF7HbVt/
wxZ8KfnQylEf/Zyvpjlf9fzL9VUDocdoxy1WAl8kfGjGzuKgIku3X8OpwIqkkzOy
Y6pGX/xirKFdhA6loq7ZPJuyBsgO6yZ4aIMLARgy/KJGhdQCgbj7qnJB51CrGd7q
Zy3mYRTD0nHtxA6mclJaHDDdQFnBv/M7yGHp9DVS4cAm4MMkIE62BvGXAVRH0Fe3
u5tev8vwm98J7Rph0w65YLktRe4sAVSMwazPWAq0FvPkAxK/EFoIKmvWxvyB53ky
nwe5FMBt4xHPrywkxlnvUuuvl88yKDkwm17Y7zshM0J1TVi7eXV9/FBFwVZS8cHd
bpst5mTzZHrIbMAH6Y1BHwlPhwxfkzPslqYJR/rg1lmQ2Ok1jERh/bJ4NiouP4IP
JEEtBTp8reEpmZ1PkBcj4BndbtRqdxUaQVBgbaPnOiEIoegf384WQ2ZRC9A+j+DU
85CdCYdbrfMFESuGhKIjS6iuCrbTjcaLP2R/tmfx3ws169vJE1ayfJ6HMrPppwW4
0kn4mA4bW+4YiZuL4wdHVfct2Y/zw0TLn7bxGNICfmnaJYjlGdHTo+oBjOlWOqw/
Ow0g0o7lxpUjn1Tpy34L3dF/XNdKejjLfOaQMxJrNuzXRJ47TV+X9bBN8Z1B+ONQ
DK4DEpks6H0TJWg67sGFrBSAD7ty01O7uqj/FbUaN1AhB5KqwQNd5ZrM1gMsuWSi
Zyg0EV/2oPGHnElrB4q+ECdUaB209IxxVSu0vz5XjF/lNRhdeo/WEV0jz/40Rfbg
e0TBleZYvkhKJJ5yVE+PtBGdSQNjG2YoN+0gFcnHADj3OwbbaTL0pK4qeYAgqFlN
4JjaToOJpbxP3Q+AutruhgO7utnU93iYSIgXagsOUwooiikg0kkXv4Gt/1P00Cz7
dYfYBQE7lcHlQ8MPqxp8Gaz54a4INfoMuLi1rRNZjGThzLXheZ7aLV0qGusnaWP5
aHkgoIYr7d9DvIYsuIJDsJu0Y4H7+aZ4yKOhtZgWB5koFWJ09KWeNH1u1cnVXs8B
lirFFgHz9YD9GjsSYLgrnWKanmcyudyEb0p/BKzwYNGYUK0lpbG6TgBgCjlfChFj
vi4DBVdF190wUH9RFLeEgYwTklhuBqGBZbOpWSWjV+vKGkI5PsYBD1jDHLtBGyWq
hvMf93M1s96KGJeQbh36PVSE0aWTkDM0SoJoOPaAGpYcUDzW1ii2RBKNoMQsADVO
akn52pNyIu2TIwWY+0iyTUk6NGMqiXxVkFPcQL+zFyp78DY4yAzx9F2gNrJ3cRk8
nOXh6F+OEmxSm3JBVUI/EoQaWiYUjU73bFm/pRfijox2O1f2X3kxyrkmmPTVRo8R
HlhUjHEl4RlcOU3mqy1UiR7auek5JcvC7HlsQllQkOuRt1wj/oYzIMgMeXFnih56
2n+/bv6My+hFAWuY7Q8oEYfBGaCnEdE8pmRb1ztqsXMBFyYf0NuPU60yVb24MqeL
IcOO3d1q+eS34fG2xdggiTvXjY1zW9oe/B5B983E3DgqzPaXpQR048XIv6tNoFA0
A82Uj/L7uhXK3Ilpt5CLWgxG4xmmzDXdlmNeEGRJpbXlPX88UzPsKNeFmMa/u58l
A4LJam4d/uZ3l2+d7q8OPSSmP5d6q4ZPZ9BNCVXqm191rZWXUhFSP4RwJHDafnLu
Arj5RftIljFZUbC6CeokoOniHs4rruUF5BQNw0ie+cUvvsEOgX32saABbCDOIqUH
bbrYOGWbQWjw+Iwv8RAGFg/LKsoLt2icSWLwenl3hGypflyzXtztLG0Z5FFa6AwP
u70IcvVqie5r6pTeKAIIkVdFWxfgiYb4YVKjJDV4cjpJZNOUugdUZ6SaIh3EbTVp
bJYKdwHcF8Wx0qUnAuVWSDajU+StAzD1iOy1AjYh1Vv5qkEqHFFXNEX6VEIEbifl
WIU7WFOse3xpD2LQLgd9n1WYcSvLRwBjZey4XWvbp5AhXF3Y0s3iicgp3AfMyzse
xRw845QghRT+xk/0r45VbxMBfLAlhzjLtM3bBsCzMQnfvd6bBIyW3L2jt1MSdPkW
UkPRecyb4kNIdGd1r3dICU15Gol50OeCkMndGXHRjySVRH3rUFlkLulqtxvHIUD5
QKSZENvEZWLqBAOs4t7+OBmUTTmOWp0Rxc7a21suQYJP77i0/M80jIeV/XiPFQ9c
T4wH5xQsbO/jZgU6pTErNtrJxGxseK7pFefd5LaWawAR69BUsyo5O6iaNSkJMhEB
5hm2WhxaKRHmsuvymCPZAkezjpzHlVz9ZyUN5OqJXwpFwgcno7jhDJO8K842FQiJ
xVDlSm7Bd9vBoYE2luJa1Nbua0AHvHIS/htGs4tRkr/Kw6NOoBMw/ORVFCb37Cxd
kuqJmbY8A4MiRPxSWSKzaPlhsqjkLpqY9LVeximGmkrXn7ISp+Eu+GKATiGXjSJ8
Mi+3HeXkwd+FlY+zB7837mntNhBN27abX99L9kx0tllwJjhRVwOlyUA5EHTF2P/t
Ign3p++2B5kFRuS80LW6le9ILHN310nzldq3mzXyrdqNkIDBgJLpskLQMmsV3I6R
EBT6jNpSXBlRfSzwWzDm6SWlOie/4xEzneji071SWtldvhlKsWMbYOo+Hu/5Dk6Z
UV/MpZouzeqYLyjZa8HJDLnT8E+2AFoRnG7J6iennvWMhNPMysKHDlg17R7zCzMK
qhZaXisQe80x7uoDRxIIPXFvtYtiQ8GkytBmWcu79BkhFRmkpt0ZXrmdQ2XLWkU5
x91BviDlX8jTF0DRmLHnY/D6pM/KQcLzZ4YQuIYHNf/+fxyz2/OmhPtTcJFSr3yc
q9R5lblnJ/mblVwOW3E5FDuoFz7FkKksHIHQd94F4GkQrd4aAiwIDviw/qKn/E8W
Fau8Yt/1Xt4GEd1lupUFELWdllNfWH/C0kPv9ms0DUTl/yt5RhxkEV1EDUV+fM3M
0vdZg/iKm4vDNgc6Z9C/0vq7dl2+dixV4Q9s6yNOMxhkyTtIZXOrn5r3poeWqMt9
PeLJk2/pkJ5S3rUQEhgbE5jTmXndjany7NJX5fwQzNEicDwfaN9vOlIOWkqE9yyC
4JpycwQUVVcLnk1V7M0ADQVMt2fUpOmGxvBQO+m8Mf2eZSWcNM6FQpTao42gVCfc
mzN2cbAvG2n85+0NIh21ACaJr2tKNyesCByiBFCIFJGtPOjEiOTLDjSZNzj6Yj1b
GLZvdM5FZtFLQTuKFOURbljibKUJ/33ZeGFJ2IlvYyN6z6xeP2Is+w7wst+d+rNA
JlWdofvqvnA3wHt0yFkPYIpWJQvNsZtiU8+veXMN+J8g4fyClQMXH42KC0uLw8Md
+/j4/I0BRyoNuhGCpFyigNs89X1JSlIdUWgcCUkmZl3wcHwIAaesO8XIONfYDnae
L323iWY0bEHilNegxfTVpk7xD1KooxbWMDjQZuBxsfmI2+epzALa5hyTv2HberaB
0gJF/s2zTXjnz/OsTpJcsStMRT3OD+NcCpP88NYx77FjmX+qKhIOOdp/cdO1Rrn5
gG9R/ssC/LLYRkEvb4Q32/LQ2XIbABTMeSJyqDvK7JiIAUVfmRUo21y2bQ1SdRx1
WdA1tk9E9y9JIkmKWZxpIumS5TgXdrP5gNfuhOOdZNGORdU0MJh75Bs76uVXQRCX
Cx4ZrgWfjlpqi6DdCvStZ/7JPBZf7+BfxYNbcXsBZnuyTuxlTKG8Mh8TiA3greN1
YPM1nWRyQwQJh7gTBEarB7n5YI70MR+XbHvZNW+mwBN/UxXfEgQLbBB8OjiX782o
8ibmkuyXiD/+BgzpS+zqv9iuCeJp4YE9YFU5EGopMX3N0FYMbqOXl02W1kP1QLJL
7lqPkeXlTH8N3njUU0t0sga0fy5MjiV6i09nALh4SPO28hhJ4dXwwmgTYm8WItWU
PC6vUchfDAEZx75cw4Qs2eR9SOtuq2XdqGaPXM2mgHFrlHos8x5fRQM0ly//IcAw
1bDu30V4nlkwo582HRl1ex6Olg8lqXzMOM0mHkYfXGk6bGcWN212hvoXYTcHKiBh
W/SkI6ZDG04Vsg6mdX97E7mNYKdgTY1+iaLtNLlcIRwdQUOqRK3MAA2Emq4FWUcU
cUcjzokrDYd80Uc6M/b8OPcwuJmYdL7qzAIR5myhWr7AlMn69+OdjNQSBmmBFuBB
cKRRPWCB1kGjXZEjbOaYVUOY8/AvwMX3TnS+svmOjXPDgbqSQzWw85D7RA++7FC6
88oX7K+LALI5lNO27tTDQFB8G/dlWhIXmwrbvTNRBtDw1bgS41TmQ/ZtNEADFF6C
bhKt18ykkjjdaOMgdHnJv7IsTgEJLUIn2xP9Ip9E7QmTy6Dh1qu9+12S2oi4TFrr
gBwhAN/jQiF8+LxHEMe7ubz3u+8B9Et+mCdVIMUdk6r2lOMyp91H3pCnXhDyIpRH
g2m4PgDlXF6B7MJ4m9xwW+sXMmXJSrBYrm8wooTIa0GZOWLcl7+IlX5XRv0CohDp
BIwLoKKa/8vSTiBlnCMxjRiH/QG4OTzZMWN8cNd4HbQ0hQCRgTs1lSCokkbu5tzP
3Bv7onYzppq4kJSDttcdCkUl2hBso1aXDBVYLRrSDG+c5MiACMMRnV0cE/4GB946
BPDGzdLYLbVoDLkO0unfSAU7MBavD2LUq+6qaYN/Ov4Yi0Ju1LaDKF0Lk8mzXozX
3NzTamPjlqpBQYRv0ujC9cpbp67la+ApirzCAUJsi0EnaUxfz3581dm82eEqiQ+2
P4sMJCdJBmbxlRGs4tKPxzqY1qCamZCQCtOUybDIQzLd0K9HOSVwhO8XvwaEXYQq
A+apLKxjjUnCp81idKC05thgS7TOfzec6/5OGlCCmG76cTUokb+NX9+Sqd+50RGU
iz4H9rcKAyGPrpb/8sfLPdx5QmdEjj11klKkYGiEQuU96q1nJmG7xiT5JtLVcKuf
AlvU+DUd/kAmqdv+pp/Cwvif49uDlSLwCT8/qh3wML5cr4a2iit3yvOyV/ZAyWwZ
mKrIuuUYPVjG8sJD8pEK4i2iahdzSppnBZeYxXxo3xz6MVxkH7AUEQn9hmPGSEPb
OMVZPekkw0y5jOSGcslO4uSAPGSCGZ9DF7X73n8TW0y8xSH4H2JOa8wzxjT1Rpvk
lxHCsODJ++ZE+xY6O2TCZiQRtTtuSDJmv0lx68LqTMjlUN6/MKT3dAlVmfAi1jbI
Eh1dRPyzJfNSCDMh2V8Zs6xiHWW1ecA3eY11UvJNDpFLKg2haib9tvqopwGGyQ6/
su6GchGGSUKQzmPtyULJe3W04hpJIMMHGiV1XrNd7C3zzyLEa+PLzGJZZJWQYk7h
qXB7HNxPxUaMyshxNv5LmHzGeIQeg61Oi0fzLwNbxxCnyxOqGEcgXcjJ0GYwzbTo
cxG0uqWtquNPf6cKLpcZ3X1Gm8GRugpSSWTnqXAu2rPL8Fxskf/UwfadgEmrMMuN
DaztueRTdIc/ZiNgP65eaTaXW+W215WHGguL8aUvyUAEXUi4ITP4V0cXJJYMuRLO
BOs4YjKs2BDT075JcxoyW9qz3az6zkK5JOxF+TQOJ1uyEUZColear3TeXBSzMtvq
I44T+8uqrxv+4oyc4QWbrs7NJ/Sb+SjU8vOL3aMmcIYyjBIpalm6qUHsQUjj/z/p
zRVDn9ig340wTd//uXXUdQ6CrW7iGQ0Aia1akhZT5QsbB/5bEIuQccY88nevSjZL
PTb0JWEt6OFVvC5QIW6AXfOELhmKD89Pa38v7nLgrlKdm0FRMK30oeANQorTETug
Wh/NwWZCgXS5paIOdlKPb+2UG68LN36qOXWP3IcrEkvb3He1ItIZ3FfzqzYajsbY
MEjqiJMPLbR+WvDH/qldkospjoYfNEO3GqIXrDbPN2E7mOfgo9VIqG4FkYVwlOIE
rRbAtKK8Gtq/7OYIIZ45+T+yFg4iddkE7+HKEYw+DPzQZiQ3FEKWL1ICweyphXwd
qfo/SjBuz5PYE2ZMT33+MtzcGnlIALP2UQ6TqejY5bTw70AhNNN6Dg+9cKZz6fav
7eTn9M+Maanm6EVLxgBCx/zRW7AZaruJ/u0HNAkkTx1/5/sQOjyncf6fsSoIvYJS
j8bYSaJf+imYwHDEQ191fhnkK5EDLaVu/UjtjkYxyVdciRN3NoAB3j/7e2m9wGLy
Rs20V2EudcxKWGrCoFVZWcHLTq1tIJZNGHgGzNXL4RoXDrQ5oRQ4uvfmFRNvqb7h
uiek/4Ta2R1ohLyo427abmoZgsjVZhFPIEXc63xHomfxmEpG3xVtDitMTxR6qqnh
ED/m5ZtV5G28OwYfkVyGLJci+zEiXKSDSP/O2S4qL8YBGU+dby4ugDuwbE4N1qaU
Xgk5QnZP2xf9W08860GWEeCd4SMl3ncY2dERp1tMDd1PSTuJdvUyK5eqHMwOQBRV
VohTob2neA6qevWc8fBAcKcmPVDBw2QofS5zPsKVs2Kl/O57+ZAjtBOtGguqMNln
Go4yWMXmVQBR4CToti8eFdBpztRDhXtYKOuqZ1cYR+MMVzaOScwriSMf26r/mcJZ
DwuYfhokvXNIiAnrWzjbVTW3yPg/uscFHkrZuea7yugPUQ7FMH8v2+EXHLDqevoH
jlw4mJ+F0dXqFrfKb7NTT/A5Zm9ixt0hu3iNpiTRBikgu5uUMaFYFPNq0LN8sqjR
j0Yl2zAAoAPYGotzciWWMdbidC7K3BavLyb68zjI8r1gqZzFfUYoov8+fI/ikgDF
+9Et1uQNT2fjOMthHeTMoptmTIvIJ9IDeKXcypXzAtEjU319GlTyG119ZOWrBj+D
q9fqoQoHoESRQ5AiEUzcQDO0k0qtID4xZzDD3EedRMO9aR00enUthV02Upg7hXpu
TpBDzqExr+Rezqtls1uWz6ZMmkgO+Am/cpFNrnf3WppC2RX8nT9TYptwNit+2M6c
IY8c4nCqfFF59O1dYY/uLqnWTM4VxNdZAnWxungOMb9M6+0UBCpA6IRdKTHwVbtm
/u3T7SdKB+iF5v04ypdxpfTdAMpTujIKsHTIFW3aQi6BVDNsZUN5nhSFNf+aea5o
sZgpOy22J6jUYIUFkXOeKfDmybFFriqonYsiVJrvgzpoC4rMIioOLCoColAaIPjt
FvZTENVwGa6iNPgD9TkqzvAM835q2SCE5atitKpYv7I4ITnJ3LxrMHZd2MuSx2VG
DzhySVNhGaC+3msPTLcgXtEEsmdvh/l9RqSJCYFFL+kv59APrC7p9xINVmDAra4S
YOVBjMYUpnFWW799XE73fjJmRPJDj9gBGgnWRLFQlkO/uoJL2iE5eoQcVZICfdi6
JPzwI0vPjS78QlXHTqgyKEAnBNcFvmPLuO6gVFDZyeGz7remZtqNeolqOFg5TQHj
ZFeW9D19p5j/aHgVn4Jfj8Z8LUlfdmgkwCqJA4tdT04SZZWmcDd4BiajtvsKOqKU
nSoq9SsnC8yknDpNtJJx5OhkrAj0vosHIygk2icoODvgHFTOMKH0h7QJVWj/nWeD
tJgnV4p3Qaq5XnOJJ+OwCiLfjyOtLnjEoyhUF0udzfbxBohQj9sDY0fQnn7lxi1v
91oVxDfW9UhL1MEUfBxFUdzy4TRoWTOCE2JT1cRBLPvT3Tdl5uvIVkLQNvI6F6ow
519hV5Yqj5xn2fCaPdOphebK+jkPp3GxEqke+J82vNt6Hjmu4DudIpeKsatGQonv
BCgQQ6QcNXaTyGv1+B3ljtOSwwJbAs9dRyt0yQs2OcWwbNgpy/ONCnAg+kE8ry3x
n6GSPUmjg4IoUxqiL7Qw1IO8WkMG621f/xWau1XUcVDZAr375TQ0eVqQNCOJDhxy
qSj1MNxwxFGX8uTqDV9r5cBWTbB7voHvAJLWPt5yTxebrxuSZLC8S7/nzLp9dY4P
fX8LxujfypV62HoMjhGGbuEPCoz4lvf2oDIN9z4DQjHMq6SttW6i/hGasNkagzBV
ETB/yyl/EVctAWmlvJYTOABuyceckwnj/2U9+NTeW+vwqzpWHHU+GNjFORumdlQq
eyIc6w/BprQYUws9xqgwu1Hl95YjV2MGSAaUcqJSqCYlMmwTqKKuQZPnJDsXJDl8
QW7KD+IDS82IF6GCk+kaTcBQA9FXbG8hyXnGhRISOo6JaWlpJC2IjrWIifqREVu8
dAgqyDdPOWxJvCd+JI+4qCL13Meb+2xQ9Jk6gbzMbnZ2KWiWUnvA/+SpGIwa4HL+
gnYf5ZRm1NuIfiwbT0ihQ6X2pO4GaYhl7bzUtIN501B0pinEQQMpJDJ2W/NwxPRb
4UHi1W0MCqNOQsf29/yYX8FFIcSIJe6rJ5aHgZrj3GeChWUk7Ntv+fEyvW/MXOON
7T8y0mxQ+Hgq+WsBf0yKGib2z4HB5kmKU9fsuRs1JeUmvbO+n8gwVC+xwtgcCeiC
mEpP7pSw2b0ZdeI5h9bDuLyE+58omijMYrpzpdn4cjn1Y3RB3JVdYZKS8Wd8YkqP
mfR+Hfygd0Og+XVC8h06MH2hdIyIsvYFQFbtBDT28JR2QdED1h358sU0d5DVFnRy
t2vx8lCTlWd/wI//RNLuern9F9LQUG05owfS3vTdv29VZh3XfLjoOsa6YDlXuzTj
e0h7fbZ3nBAP4Pokg7/ielemtFGF8+uhNCmOdMuSUUDFidzWttOueZB67gYPF/r7
kOiJnI340KNGs1lqK18nfCtik+pUQ0Z0PMUDhsXGd1f1wvuKI4C7K53tRtm6Oiew
IfJJPFSgomfjOVlocOMQtufnfGeDYcVfpqB3YlkDF9uFvXnfKLUtvGd8xm189x7S
OhCM0JE0kOIII7b9Y8bJEK4nA3WFSQQeM/af0aKtPqq7IkmjOJf89h8Kcf4MwsTw
vQm3Ame0xG6x4p55vg8cRtSealoX7ysEhYVB3cYj9weADsBTV7z/AauobkdvjZOM
ppVrtIwAKrYOCCoTB0QzQF1bNsrzU20NVvR4XtbjhU9APdq+QoRSQ7xuR+0UbBu4
plzqhTCATk5jCshFdGkytXsmwBu5ga7BuJasNs5vgDcSP6lS6/3KJFIH+JTdfqmk
deA05i5i3coZEMymRxj3oN/uYRAOv8g+MygR/g4v/ch0j7WCZ8SmQQFgLbqCysGU
pdZ7awS1aOuQNNgaJYjm6AJOCKRt0R/5V5cClXxmQ0ZF1tHFWI+oEDMQrQqDlzG1
Y10FskJb91TOgzFQ37w+qbVuBrJfoWaTNIvelTKTfn2XSifq0oF4Y8SNkIwIJprF
/tpOeO/GWdHjK9RQtQtTLwavCSn2446K9EkdBr+KdwOLAktWcBb1/1LTvyOK2mzE
fBMKTCl5uwuHMO5YuccOxzd5IyctX76DlUhh40Kdp30cdz8+GypVMgvG3lm0kJKO
JWua7bsXwxM3FMdkFIgsptmRNvJqnVZlF92jU74/4C8kT3Y8vvIUMKJqFGK6CVeV
ADQt0F3afcurpsc8MPYUa/3yDi+8d8VhglrWIK/HI7wie7oqYToCXDhX294znW4t
z6mn3E9SVKybotCWhjjavh7qCPnYRT2SjltqdvoJkM8Gew2kEMOTVu/V/Cn+t+hJ
/W8mtb5LypIRM9aWNerKgGmUwE+1LndDOGeLxFMOYgK7rKbg3gnSP8vOmORhfDdC
YlC3lYyjiQcUNsfS7kwwwjmXqNrX00Gr68bGycRVxAjtuJ60e5Fuq3xoVTdo86dy
8/pq62bLJpIXbBQknGPh/BAc31/FhVn20Mz2ZHwS4CYL6ep+fsi5q8MKEQPLosbs
bGoOCFvyq5dU3zdKMDLsZsaJbm/T6lBXBdPImyMFDnk/1oW93x5WML7e9tG7Cm2w
9t/J9tdGfwYFgHK0lNdwJn1u9AfPVG7Jtrm0vnbTqZ/2DN1fHLx5Sl5P5jWXT5JN
zASbRPVI/8poKHXItnTrOOt1gbag20GojyOv5KKjWxN7ywXeV4lxYCSwnFpHR3MI
ui5yZspeJH5iElzupjYULI+vzLxknNQVQNbIupUxqiAPR84z/mEKs/I9L4BfYHAj
OKh3197XGPIG33JsMp3RX9TiEm8POUFlXWJwIYlQW+dqFwclnVTSOMqsZG5I0k06
X+HyDhuZUZ8uu0eW7rLDTfXqhtd9weAM/WeYaNmuQd+cTj780iZXzFgOzGgpq/vf
XN3qdMIqjWWpDmZomEybJmX+4wwG4kkt4NzrBdogGZwAvujFp8QHP6OQZdG8b8k7
hfPSpoYOrH5Fq22jHupQEW1WB5uX+5g2GBJp8qd3Htygw1KwM0phF3lRlXq52P8B
IYu9PzjeyIu86+REg/sRxcgxZjyXwfQFiX2QbbkbzF3ZqP9M9pae3xD23bKqrOui
GtFYWOih4ornTGS2Q+QEuGS5Nnh8XbCVpGCnqCXlifKVZL3JuS0s1p8TjSl+rwKi
EJspieAOf8uM2RG631CyXmghUu4lqnIv5NST/HcqjhBjYvMOpYLKRakFgfO57jsn
UYJ7eFaxB3dxGnPOSmPyR5e7u1Y21O6blPATO2MOsosLV76Ba7QZkrfOKaT5Ukmz
ZpbMNMG/EUSiF8y3OjK7cvpWIDIJwc+hcQKZXcZM2iZZhOWaTqrnEz6cHX5jT93B
u9Nz13GQcHIxH0vJ54naMIfVsAW2SzpACzxiWQ3ZwVKBiJ57+qCDzV9TQBTikfZH
L1EHElh8yzkYLVJrauNPZ2+Q/1xsLlOrKhoZIYn/cdXD/s5AFSzhHWJxtzidboky
YYi0VSWhNK8ulbEdY8sDE1x9cEPqo9ayszMLLv6uBofZF8w/001hGr+1kzrWM/j9
j45vnl6SzumVnhDNsagd6s4N6mnyFiK2iKOBazQxKOjJY64F9O83oRDNIE0fwtGB
cJA/G4nLvM6pf8UfraJwhVrtY57CKk9hdzyA32QCVc1yL57zEW/vfvpELARbBrU9
7nB+p4Gnft/ms+WVu7ocCEF9SdEw4zIhAUQyXEtRAiOgR3gpCxdndXFQbsDjFvug
pM7PWhburGtuvfUoltxlz+FfFCfOYm3jTj8v7jHZl8Wpq+2oGkKpr40azJxpsTKV
Go/ZjKx5HQWEaV9ZDzsc4RqxrTU8hwIweXXz8CUTMbv1foTmW9dgaHs+lldIfT9q
DvjWe0s1v4Gcg4ZW75KJbCaSQXwqjX/7odIEKTVnrXk1mIlctGsflTeaNHq9kKKs
5HRSVm+tACcpN+iSPZvPaoSQC/58/2i0f/9pWaujyaE2EJqstsTvY+XGJ0gZsxHv
CUvvMIo9rzWZQQaHezfs4TrpPq3ePOtY7AiBAEbxvN30mJcXftsaZ1w1OvV5dh4C
yfQbO8U8Dcd+0jjKWvtIjWyNb1PlAjHsdsgoDH2MhZjpKBY9hz8atUOrrBnne8QW
wwNSJF8cqfAlRpe3ak+TBRTzHThP0gIZ5ZsK3GeK36FcFsW44QlxWoQTSJypgcKT
cfqmXWXndk6OeeLWbr73yuZmkL5FXfEurdUxPPia6DTPWvQ1nqs8K3DUJQ/CpUi9
WXHfzxMc8hJea44lRWjnP0ChNUAaEbDvzcTPn1pzmKKpck61pdwYxL2aOEUVZou8
46gW2+by6Rf5NNx7BmlUqLaIjFTGvqReAVOIB7kvJ3jWPxIvcdYpQSWSFXlcXs6j
jane3oJw3+H5Cqmo+xLQuD5k3AvgG27f8Y3P5jYfv1FGMsd81S3H87dKi/I4Rki0
Jf8y0uQp9H5uazd32t20GBpvk3FGfELivWGJrT1alBFqHccKQPpVrzdaETagVg4L
/50TRQPQQ1TEJjAItt6uVEJGK+kdNnOYdygr5SxEUrIWhXfkoK+CYVxoWfaD0z/L
UUE7npWZKfcH8BUqK6qFwe6c3UkHrzPmhECxM1daMIj+d61E+P78f6+UOynSyi5Q
4IFtUHW8wtv0KNzyV0dCh4FNEJlIQQJPQbSptSsJUNGLD9lS9dD8X4HO7SwpbfzL
qmatYxdB2gqr7JUxio4EypvGfUXJ9KgyIiL2dwA9s9J9T5+XYY+SbQse1fBt8tgN
drrdtzZj2NwdRC5l10BYnr5tfQF1Yb1uA6+nY/FqZ9tQi/n2Qk+fGyJtOUwASs9J
mwNGr4qW2Vn80xVsrfFme9/1QcIzpcTlKpTA5IVgsqMgUAN6P5FsYR6ZXbkEEzUu
LnO04bCcEPkSSAtvpPGr0JD13CqY7/yZK6ati86h17t9yRxnsi7ys02uDTZOcVf7
XN5aDLZRw/j5ppeXZ9kEzHytzg1uJn0OxJllwAYnJ/9BBw+SHEHzn0XsgkeepXUq
4YnY4gbf/0VtRhnu4rvCdvRvmWDzPDw9r3UF73IblV6LOj9SllGAX52utcETyG9R
OrkKFcH+sCQs1Bqa5z6IQdiRuSUHD86OYhkHTDADZzQ7J6BOgQKLP9PJoCxzR6Wl
gUBiURvMpbUfMHfs/awMkzVpPeYJFOm+uqTnJ52SK91tUsF57tUcyxOUwAZN1MVT
1FTfoT/kVHKIVgfE4s0sf541cCp45hxVJek6tgj1RkBhm5CceRXtMHsx2uAJeJ4N
df3ygdcIqCKN3+heXXtslWJDRNke2Pws71gmN9RZ936+Nl8LpIg5e986YeBtzL0O
PPXYzzcO6CnZkekEyrF0D4aKx/1bt9vNdg4Wz7StM09D7Nhg0SZHrNCSJ5u3mvt4
hecPfR5Q2HukUWV4PIaiP515nY2rs8J+l07rhpak6Zco0qDEfb7LtfCHbTNzBt0/
lUEurgt26hKK/iqpxlS3S5crFoXHRDNcGBzku6IH3992Ce+6v0GAMuym/DYzGEXD
N9QEErFJfjYJL0gSZeXq85BCtiDJztezifNQW9rEi/VaFgVk6qP8I3KYcR2esRwJ
aQeznQrkpLQt29OM+RYo0IscNKgVCb+NHPINDbFVerVaG4Nc/dQ0Kr22CypbcAMn
3x14DISI+wz3URpX/QlwZAKjgeq70mBHphJASxKHqxHFB13P8qLyW3qM0rCTCmLC
bj89vfRooUT+xxdX4kncSVE307JBT0sYYFcxTOkITXPsb5iCIqngzUEoNh/D9Yt9
sllHgfew8sp/GtapBSP+2TWe5xCey2gZQjsQLGA0NZ8ZngNXDAI6FJ4YewyGRJSM
DL9NPQsZjQp9LJx0VufAmP4zQXH0Ri1bVT+ODMufTkRcancSWeVheOYT6FbTmixe
PWVVeZKasps1A3L3vv9UKIOPNiijy9qJYNj2zhgZA688qGE9H107jYfIN1aKz/tR
8AzqSpz8uqb7H8qO/PpZX5ITgnP/PJoh6u94u2gLdStk+qGPX8fcAy0m9HZ7Eahv
l5Rv2U+nQFvQh4U53P6Jgq/jCzgx2GXPoHMaaUkhNsX27w8j7Eswnb/s0wQbIzh2
sxJQsDAJFqoaRwlFRBLkh6FkxU8bYtW+cQWLOuhV9RhOMVe1UiTioqsmoeMkgs5E
Nlu1hbRmkEa+g9YWuSNp3yjh+Rr4FIJzKm3nVAdU5Kg10GC8/fDlsYntVvjNz3U1
SjbXns6QGkuVlK066xfIHGu31h/IRur/p3DjFmiIVj3rPuzxSAk+kMqcO4aoloOu
ACol5XqI7O8Xpa+pnMipxUvpfc2CCqYQnteWLZuJ9BCBG20UvOs4kmtkA6Xg+0Xv
IIU8xWLeZIWgOSOssRbup+JuJbHV0kpITeXtZ+kE8WNCb9smEHPnY/LfmgJjb2uS
YC/ItxyueO4WKB1f1ekibbZNdr2+hI+uPhqvGR4g4KB0iLauIl89zvPheY7nS3zR
lZIM/tpASkP2qN+p/O8rzvkRujePBvspcQwFI7klxvkNyiaTAoZQxruPgMsu1Z6W
S9KcQ+qqrr73iZit5798IUsAPqwIKD4FSBoCRrDeFzY27WfvTodD1Cc3g5jC1lPx
oK8ezle+nai40MbK8+tkyTJZ89zg5KP9tnBb5FZTFv2JHvWQIcSyKEkhBCDHAc5S
KI2GZ0P/WEFk/tFFBWFO46aNECJguBNywyLcvLzvQWdg61QTxcNFQy8sQCjc9U22
YSs2N0I4IZSWXd1Jh4moNr/y03broOIMzCE4yh48zDwWupn187d1Og6c2Hpu7y32
oc9BzANJcOAkd5+RDDgB4WJCXBWHTLZHqWpHx7R4MhNud6JZnvMEo4Qc2QSfK0ob
EQjgL0Ex+JmqZKZ49+cpqFAwcxxB3HvoBrfhlU9Py/0s/DY4fTmF+m+5AjOUrTn9
GNSvsx4PvuSJd17egCIh4VY1YqrLOhXI8Xe9TScRjKk80rSWprR/bpdFxMm+Og3u
k7rO/69darICpCU1vf8ZT2OyBdTdGusM4SXyAZ9kgdLGSkWssXQf0X88QjdwOpx5
muiwA/P8iQXJKqgIPmd3O8rNIIJt5i7a3n5qQNCbuBHUQEJXv9wo1SZuToCi3dsw
EHS8YOK7ALqf5H4kI0aAEfoPhy8p8/LRirja9BNcF8bQXDsnyaVcPjL1esmq5m+0
a+MhYLExvPnv3XflCDImUHO00vKO3QctCjDPhNRi4HRd3pEcEEPLM4LG5kWZo0+P
8n1Vos50VDP2wlfg0WNnx8qAvSwtqiquNw/L3ESx92gNleiwpplVuehLOAW8yAVh
up8v26R77iT6iVbOJa7MlH/aLQt+Z8AjTDmGEfWutoMi+pBrcsQ532U7TZt3U85h
JTi8FBbcczCZ+70s5fU1AnLEcIDsoVa8SDOJk9fM0bwTxmuOo7FnxWkZsaVCY2t/
+Ls+QVtHnHWtshIUZ+QljIMmCQvH9fdt4vkeL0IRGAeeBReKuf99E+9uYYB/HlwA
R9GuFDvpCZ/Ny2JriTNPinwpSLw1mTRrtOyOPf1AExF0mqJPqseCzIrLNemraDDG
yJu2ZrUErocn4CUJb33HC3ClDw7NpWfgxgCRM61HPQCJ+ySSo1BnOvpukll/trbb
m85W8JqwyoGRutccYuVQXI9Q6T4NgpUawHZugvs88eviD9E8fs/spJ4Kbc2eoAso
+r1fVsTjvKSs4HzqKDK+PZAXWmqVXPiAoNNrLXweBUP0TdhoZUxdI4w4DalgSoCb
V9ItPp6WPCGEmsHgDF/aR4zx6wrE1V5ED/FX2nD+MLRIagcQ25bNC/G9ps6x7p6V
S2YqvjTPtuGMHWNZC5kU+4rcEKsMyZHe3YG88N4D9JjVAECc++85lFbKcUY/81vO
YcZdZJpqMp3JMlnKtzGqbWq7pHM0PFYEgPZzdXGpscq/WSdOQGVnbefs3DeGSyuf
pl09BuWaneR0hhA/6WGpe0E2u7umLym64LS4Is6nqW9iO2PWUW5uNTeXXpjDponQ
z+oSVh+glj3n8+8i2GJyub9X1C0TrXYc+oEEAXSfKryetiSH4Hgiab9fyeHauuzi
MuQyKl/x5oST9/eY5IKRfLUPypaj6SDwP8PGduDue1Veyo1bGMo2TYwPpcUavmBJ
lncvFub5oEUzkcB+lfDsOR6jwqe8vz+0foKS29VNv2G0vvV3Bjr6e6SNpT+rzzH5
+xBD5axw44qsTc1y+5kEm2NAnweYq5hdXbQVF1EVnan2D/yLw+JVharbiI2RtjyC
WQ6GFGYEDt32YBBuyhY9Yr4kyqDAeoBIvMA4NKtSp2j9pxoD+Hj1Y/nKM7WJaLdp
THY18ZElySlJ2LgQpyiY1UlMMJMi+YzwMy7yG5T7Qktfyzsnc9gDzc43OZh98Xwm
qT43jLL4mporPz4tEtBx+5U4B2kG/Eb670q1sQ79Zy7A78zYXgMSB8uuhT2ySbAV
cGo1Jef2fbx3Fm8zTAQ+IWSXxpKw2hJgMM0u7YWKCf8pzkJDW6VC9YROfbtbIVmj
LqzORvLe19vukAZMTNXDKL15SR11Xf7SR2v23S/H7Srz0+7fzDTSz9kE8ZJfKaB7
GTFd5Kvo1WRJP1KhktjVVxiWxCOY0ZhGgeuOHuMYuLjAgDuUf6W24IFtVZJcON6M
WAh+MSWfLho8zUc4N/8Z/JKz8dF8BUxCZPrJ4SeLkYTtTcHnKXSH1oubi8GadetP
4C1gKTUTuvCf5Rju975KjWIRlbt4py9AXsC5A1/NtXvZzrLc+Z0Os1hUUQ4RsfJI
s2IHXFCei0SxEvfdsTYt2hNUESEa4Hskpun7fT0DV9HIUPiAmXHTXxBD0UdCeym0
3AUKJHWBoMe6p25zW+UZKclmNjkLQ5ALyha8DeDP/tEily2FznEYv85OwPJnEXnL
Yq+uwLBmHD6z7aNIgmnpFyl4IU2KBQHnYgKeP1qaiWtUBbNfxqAFrlFEHlBKCRPZ
rqf4hUTZMKpUnWO4Q3bwWuGE4aoRn/2PTMdhMbPy4uj8dXSNmW426DG+d4ly7/3Y
6zTpz/iRACssVRw3j+nef/hqOHSvv3iHLP+yJT62O5OyXNYVWzyntDa5kKBXZ0K1
htvZDcIP8UE3EBz8egAq0B1J+wLbwVe5Pd4GW6rAkIviaPLOms+308N9tPrpXOGM
/rXi/zX3dzn26nSL3YaGGLSq7Ksj6VmmzdeGh1lFoAH2fkCFhNxL5Xqe0/HTRTnH
lxK4ZXGjTSGLmQGAIh6kOOyQdE0BpQiBBqz47sxFAr7FUEm7yxAc/+KlZygNRtuS
5yDdiXHX0WCFf5BVIOR2qavyAJIxUkDM5ynUMIIbGJOMyojWwuNdOSEBImeh3xZi
kadomvcnWyBAjgD4Fs7cC3qP9bPcvYivqavEEBkp6uYMXhUcwlPzgS1ISJtIm+v2
HhNOQGji5wePUmtZiQWovuwOdLXCHrkBhU4NHOnL9hIvpUvDpLIaxBDUiJGkBZg/
y7SPqWzmzPLqbhUP5yNLiolUXAZdzR7dNyG0vU7dyBu3wlwWOUkx0E8yuqe3PSS5
9VQCwpYjr0XTJJA2y4aaxZ1ZDYP71xNT/MWeqk5qn40bwBT7kQlHx/YQ0H5LxMUl
BcdMSCp3yXbfAoFCKtCYXV3DrgEa3ihhcnTqh99J8GOWxlkeInH7JslOQgyszarH
/wHN7XwZ/qnejbnohaH6NpX8ZOkEiUlyOOUgFSAe3bwCgW2RC1Dd/DiAyo7idPBl
k2K9AsPkLHzGaa50m1mYv2seAs5xJjIdP54pxfNkpWIHsvxsm36TuekdDf89Lnue
DcacmtaTaZ+pT8vArrJs6r7g0kuhNz/Q5HDRCT+VJNKdehZEi6D6VLmKSOeL1WqV
OWObGgg4PvRLV56Tmoen2oaJbT8dOkFyNlnNjyGOd+/dI6HR34ke4jzCuA8m9kNx
1kulhsSsbKnTrOK6/TzYSKTFv0xUUxIaOozGiowA+lPif/glDDmle7lrRZ8jke3I
MCR1gAxpg6GimwP9axspdnFp/7hXYkwt3VUAcpSaMud+IKZYQQ6yEEUXhoOevpA7
eFPInbeToJzX1cqSEIMfk6a93+HhxnhqIdTwJvPFDt+7PBNbYbhcFCpmQ3J9NxFh
bg633a15lHlkCBEwFyG1Hxo1RTnucPYZRyMiB8ykHGjA+W/600JwomGk9C3y68Kr
wIlAg7xPo2Bq+S3sswGEkKePWxAQcaQCLXJ6XG7la3fe5defZldt3W0B4yj1ut7x
TbizuVogAQAFp0zBbhfceVdVUkjy6/ZVjdv/36ziFoXusTHjuPvzXc+mpVLyeOao
Iy1vB59j2vv9iDig9tKIniOJ5pQUiwlyrQxginHMda1qm7RzxMYM/AyXTQ4hnJEV
qohAfX+U9V4Qn+qKtgjv0K0WBlea2f88xbfFWwy9LyOu6GeyvIPuVEvVmsym5Y4q
brJeWummVwgbLtI+aiMxrP4/r6pvEMp3lMjnSZWJpNID58JYKmzIrnyfPs2nEeIy
3J/3wyU3GAZTLmhCM7uJ3yYa1D2Z+FzCTokRs56dwDpKTMhEC3+pUCAQunwh7u5I
Fc2SURHck1AWSZbuHB/eEV/mytBx+8szIhTpX2/PkuvHmXoKVwgfTsUTu1/x9Nhl
CDYtNB/tBfwjgAtiqbv7utWt0CS8Ze9d64zCJC+dYmNpySa41fFs4pSwxgCQzPlg
j6nwMi9FVkGqDNS7KCb3epct2GmTCCy21AYtSPiT8Mm/y2rCnSQxSwiCGIRQ8XY/
uPMCGy0nbTfCIWgT1piwIncFPHWPeyV8jXxXX86LIb3lpXHUxbhTNGyg92YrlrfI
M70cz1FoyQXmiIbfoD7cbgktD44MMcmBDI6hd2akXlAXU80rnnn8TeKL0h4IuY3b
4UFN871mRSGU4JsvbksCz17GuvjY+HH38lP/Gr6GwsNq6uV1kRbkhNOmTwmd5+dD
OaxW0CGUjG1g03quzf+UgPpe+gRY0IPGrQvUpGCdW1G0egeurf8DgmFAH248kRwI
wFq0/Kq00Vv/2h0Qr4EumOlpLU1VSdoMD8v1PC4Gj1jHs0ledw4SO0ueqPsaq94f
6TPTyWVaVBiU4EVqTZmZIg2qNGATAYmEZUxFh8eylWimsFV5owk14aZixx6tO/ds
MVo+BfUtqz2xb03RFbc0OvcFEhYDA9nOWHF1gaKsVEOqFXIuyKoEdld68Ga3rix0
R2R+wEYmyNUIRagqQZshbTfaEKyzw2WlKYL5xv+aQLb5fAU+SkX9pA5ko7x7gDUr
/U9KLb6xMwxbvsJ3d9LFRqJBxYmi6WqAZeBGRJlwb4wzAxegD18p3BKjttoDEn4G
kRmXF98HnzOWeoczk/tJp3Pn8FEntnzplJ3zIB/wnQ/ZZAVFdeC/5LYx2JsRa/cs
uqxYMGuaPz42/AueUgG4AxZdJrMJ78ARIpO8gQ80lAJIUJKdRIpk87h3XPzG8+zn
QiIXRJJPfvREHk+JBua1yXmwisrsvvV51ojKIB+wPQf5BD1yslyPrTFjPKBCKaNI
vQOqbaGOLQhBWJ3ixPr6bumKL8LTxMDjvWIT7PPWBsKUHBWQuvwOJOnsK/XeaTZN
RmZxiFDLefD6Sqk4t98pIoGlQczMiZI2mvUFcFUWCzd6Hbfk8hkHDL75e+HVdqtH
92nn/EHTc1NFUJeXZU31cwWnEV5umQinM0diX2xJwSxO9ptjinAj8V2Vw5MMtIlb
FHKd+Ny5ZPZCWSM70jZwFboiEMNHt40PWk4JklkC4XG3OtvcaD7g/49U9OZnX6Me
00zU60WONpztfhsYLj62wA2f+TIaWugHdJPoXSWwRee91QUKuCT9KB6foIorLil+
RGuG4NiJzr+cqnzG776VedqOl74gWxoNjSHitR/n7Wg+kPP+LydjJ+sE0JSzNoMl
txxAFji8IwbxjgT5eoAYa15KQS+idw8zngYwvWobja5bYg9odTG16q0FpbKJnQdd
e76XFA/H6e5WSnn4pujD0TqR41qrqdzZI8+gSI44G3gvU6CWp/dEwMxdPLbgHnPt
fwD4Qr1i9DK42cCIjGXzD+yHvP1C00juRuP0utoFjGtAssDYaaPQ4z4ls5IeFAc6
GhrCKAE+AvWBvS4yndxLJv//PggaE7FYphUwWWIBnwModJR+mHZ/bZeLM+DYGm7S
AHdhLZuBBCNqyYU4vDJ2x++m8Fg24QCCW0ydhm9GorAZVG9X+MQbARlQmI6n+1xL
ut4Q5b/qrOwYqKR7x3zBTJqzHpDqCQl+psjtVd9csQzAMC4XCRUPUb+77itBtynx
2x7PVTzN7EjlA+rmwbC3++mPdhiI5/iJ0nkCgjaA0N0Y5qDsezIuTipkdSmZ1nX6
LLqokqu0dXDYCEMhJdpE54rDdP5Dw+JTskxExABQwkINyVy49g+q+Ek3IW6vsd+n
+qWes37ES2+DZuVWaMEZrPiBC/4PgHs83Esw/CbezvuuxT/Nldwt96SXrrh2P2wk
fyisG93DNqhIJNmQWxCQmevBDbV2XOcm5HXeRflNWjxtio+GrXLHmiTBv8ibvAny
rgHfO4GZB9/maoRlFG14mzZX8b2TSqmrmPbeJLTEtoZcjBV4MWH89la2jk4FQtAF
B50eRcPGCXT+hlo/2fA6CfioPIaadmmvrgRnE0TdRK8e9ACvv9q3Mws0/wqU+w5K
XkJkxwGiXs+B8ci0PTD/koQLEwc8MKia3aByhbRGXUhACJQBza34SJM7309sviXV
fqNPIMt0k/JR1/Ng1T/Sua88zvreMLst9TYNeS3Bw+tED7OOzP/rTcJBblyLH/ce
vsEM6vCwuBjs3WH07AIG8ZlxsWGPePTHYZPIaI+7/WTeed7+2Axozk0qpniLxraf
3R8Wf8f/GfLPvOOUpMRXa1CHlEgPrVMlHu7842O1aHND7TuKEbZ7S7yhJ4nCGYI4
hkB0Ms5fQNAWk1+UjEoqWTvSA7FHrB+oHXR7LpJascEdHaRVQEmpRu4QTZttmlxL
e5fvM5fACUY1H9/tcWHJj8k1BsHy+RaaxnJVpLxUj4XkOYy21VEhEZWfdQsVGed0
5egKHBFvRxExjGnZ9n7Cjq1K9lXUO15tyQN8lV5wyPCzbrhmDBNpcIUIcg05Axuj
IFncONDj+IZIIHhsGLCKNorumNNLY6ZLL1bbNV1t+GskF9UclOpaqjVQfCBpbe5f
Owh+V/FAHOG3lSEfgIacVG/ZRlST1D81PR5sYYEG+sxCyNGD5AfKk6kYFO89qLEw
3khnuTvboeuQkYpxyO7IWQdcTWLXWbKXuNraRtcrohtZLfp42OKUoD5bf9qCwm88
ObsJxCqtiqzZ3d3yk5/Q9yQpXcNr58QApMLD/Wl5EQA0pkYhk2G+BorCJJsgjxbV
UtInLkL8DQEIXCsELXUEPQMVEJL61LBIzZdoteZjy3V9wBJ9TvaJZob1rod8wkHy
svzMco6gMD6xNlJft/+nw7ouAQ6Q3Hw5mGNPsbGOpAnXv/zjNodIfln/D2jzMdaq
v6AlndRd6QUSzYjG60ePmR9bj7+0L7elJCdq0NwvZcl271AgTnPhYrja7AbYH4K9
tSFnZE0AcDwF2gkvcfqkYxzjOTGG6a1sranXVawbucaNhY1a5mucyfVE9y6FdX/d
G8ij0rKLZNfOsLWCHyMg+KFlKM7ByQ6yJzOpy612pG3kYVJfkolePeqx/0lcS1G6
jXZ0oJ7gAcXX+MgDiqmgRXMSZwuVCKfRWtiyA3mDf5eMwuDG2fFBopf9PRsoG+ue
3ces1iDB1ZV06MPfDn4W6MglQQ1sTXGIo1ye9g0bB5hgmRtmhUgpVYmPj1mQbf3v
kEYGQlu0LtifA/09xt9FUmYTUsEHSOKwGpoTSmlrE+3dz8pWZVryH+C7kOxW4NK5
4MFYgF1Sdp+dd9dy7xc7jcI/lgv5fBfpH5Y5MvUebfJRCP/zb1vvqj/7gEaQhkgC
BpGfBLGXGxnvMYZobKYsOjxqumJYEOKbfq3uCCnDshFrW3YCunHHTeVho/miSmh4
wUMyhJHtVDcD2efxA2aqYM731c+rbJ7ONVGIh0NJc0KO3ChQsFzOdIfTfEQzRAIK
HZSbjTNGoND12G1Lwgw5fp0zS8hseLzCKf8w2YUGiLNsJz/C079J8g1m+xEu3Xxz
0E9iiyeGaKAlkW8P49pVrGENtosaIj/dfz7qeqoOoCmY024RWzZEzvOGRXLQRSS3
51zMpLJ7i5oGT19MO1O+LcXU7NfKEwaEcJKqStU01+i54SKN4OHwsEBkWo6wWkyR
1gbNHngC70ztvrZmrPYR3Y5TtJzgdLqlhkWfuDBCCi06H7ck5+j4sxKRRvzkSS50
YphDjwTF5HChksvCWEc7PBUAi8lFcuXSVpbjyzNd8eM5ftPgv5NZbnvmbJ4slqYW
bzemM/Zt0CEynwq6oUb2y8x4tamX8GxoQBxaPG/zJPViYu4FCTcU/pE+ZsqJRb2s
NEkaP1+hNnG5KewNdRE5GMEvQfeiPOwPx5rLQ+ynQi8d1Wyub9HRTxd+W8HUmBzY
WuUh6Xv66sZoE5TH1D6aNCkTTYjwuUiPcU179YsM0xOA47WGa3hlm5im+1KpM8Vf
E1wK64BAMO+NZeN+hAz6pxtlfwMKSW5mlZNdjWNzGiLMobnyKnYzNKgRH0IZS2LH
ZN+Tylcd3Bo0p/FAGigM2IK/vx1N5hz8b7p8XitbGvmPInDbeFiRGRTEiWwtM77C
nihIEst9aN8j7ekTlQGKKSDF5uepK4OfwVMUobcRijsKiUz7YFaCcfqf8YoIdQ9j
SjvF8puO4DFZoVrd3rP5bBrqh7DnEgPMVBvjitF/N3ho2vbDQf/+lKg8HxA7CVMw
kLDUEZnVYkj9S8mp469Xp57fP5yQxNeWVSkY6yxQjPMqR/7bTSwUXz3hwjn953eO
EHvmY3V8Dur9lLuE1bccaSsgwMlLbyJLMgCD5oFZ4frnFkCq0yNQ6AQ8Hb5TF2nF
gRuB6aRJDWDIvT9tI3+rcb1dGpW8v6VL0ygtgvYch9tSJmwuOdDHOarxCYau8EPG
foXZa30cZMauSoy3sJGH4sWiuR57rLhvUS+VUBCgUHYujBX0YXI390pUhNFLJc/T
W6Nx/X9FG0shL396nGSAYAWQpSQZ6K59sjIppSDTnObFi93Y8vl8I2yJTEGUief+
ED2bp08i8FXwoyq+zFGlggD89fnLULINppln51e81qyTXgKud9PAN3nwJVa/7fK7
hwA6ikSP++zOZ5WQblQV7e8hc1U4rw8GMlhIX+0zBN332miFgap8koi+nhw75ZYY
ppX7/XSUbw2erh5HlzC68tPWG3vGWmPnQ00QHhMMJuqjzSdx+G14IBTVY1FSqI6S
JFkuim6EdvTZtI8QxnHgk9Rq+i3bnUhHxe+huqXy10rRO3NiwYznd199OhLbep8V
EWxJ3m7Fkt9E4BDP8Ek0Rk0UdEQZ46lhZJSdxcp3vW1YxMWIXOiDdi+Kual0/tXr
xekQOwqyGREog9Sbm2txZIyGvFKj7L3ht+mYK+6XTB6bZ3F7c+u96j9AgG9Tf2Zy
ms7o6hYgMO5X/jHuILvml6WrZKLHzp717AxutwrqAuZ8afqe0Ch1/ncXiIgvF0J2
aEvNPcz7/8BySv+VjuLNGph9p1WULv+H/fBJXt9rUE6YdmVc2oNDGA3NKaEPnKJv
dr0YdvHM6pnghoonuU7zHp2cwIgNn6fDAh19me6aOuidChzmC5Js6nK6pWC0LgLc
gSrp0eBTBgtv4mR2iYoyf3bgiAf1+cfkYAe9p87UmW9MecxM9hVGKRCt2kuHK3KG
eTRKihr5l5DgK5N3WOrj5SOKpze9n+WHJ06sGVO78pPFg4kG3TFCtbHNCKKJs5Lo
smy+YUK+3nYz65Ow3Mni8Sa6BC+XHg8r4S44822aG+hCt5KG3FzJv97ooKuwjI8e
VZ9Wvvzz87mGysq8ttkl3VIswSEl1RhzkUrZ+xUrMbPRtjww2r/5YycjJMi7xHu8
oPDFRh6UWCr8JMdjotfWX3TyUgt9yd+0C1LKQy6q2ZWBWudLXJBC8UeBxWzO9izy
hfWusH3hQgnYFroRgsXx2ONhXTqnX1FqNRTRAp1604pXOCYvmsZLc+1qtareIaBV
VzAUN/hqmCnG/xXTmjUkqDWRIyF4mIa5JFEGEQ6sg80cScQrMR1riLhjlwlks813
jkd+h3KdjVdY71nofPsmMCqe5iq3/sIxFnVvpMdQbhS1KliRIZM+peHOIkFpKqlr
DEjpzrK96QbOLvGFHcHx4InsVbgidwF+umP0as4mj5dNpHGhYKlY0CWBX5TmLezi
JS45WX9N9KXFYii5wzu8ZtdTM2TmMm1sDqZ8W8SWAS+vjZ8mpHqllrfsg5xYwFIS
LjMjIN/ZF6BlyVHFbhAblh9XJ8Pt2uU4JYtoMkeoui3GRAZ2AWeizfGnjIV5vYu6
sdeOI4deWfUHTstXJYkm8TA5aygE2yoIWqS8Sq7hSGX02EaQuiFVM+oLcQEN820c
gyHGKcDGka1agDHbr94jfvXg/nq+1f8Aa9pWfS8qk1HJPhoaJ0H/pwMpSKXAxYVK
K3fSCx169vipmPO3VAKqR5CsVao0SHI+bG/WjvdbpS60frvkFK9l4kgrIlIVoMRt
ccG3lwfgGdmmgcTflN8LZshG3KmsDQA0D1HnH4l5ytPqlVdMS4mC8sT9TBG0vg7Z
c92rYh0GY4c+ByqeCAFkbRlhnI+IP9PyZtt/h+x+iTs80u59h+EiA22USgsDGQBW
h8838OK044al0bpHN+UYcOTv06ewa3Ua1qCx+gi7RfkwJHwPID4rQLnpu1c2GSHH
B92ndwd3dHlZn+KLJquXLjrXsC9rih4MSCe5/p3dQM4O6JJUUsrw4Bt9criUIkKW
vMXGw+EwimPcj8A5EPXTcspNn8+5bNE/cVhljobURd3Qb05fuZW3+797v1nqPAMZ
PHyOU4XcHS8ntNOzc46mjM3+FwGSvAHDLs+niGSswJIC+yAIzGsTu6uvOxEGS4wo
ha7l5+LqrswYUkb74oVSdrT1VBPjD1J/RC9glGMuC62z2s7M2DgQd7R8fAIKc/eJ
3jIfPdGgka6Va37AC+fJ6jiyFyVFnpongy8EpBnAU0T1u5Mr1TTf8RFhvkEVDnMu
ou5lJrL8MLCpV3Sj+HcJPjSwObR3cbedacpu4lrdVVblc39kydviZN6Ohkerg4UZ
Mu/sfrSHRWdKKvacgDNP9rTNu+pBTfT8GXLcdCMATEELlWjX+TaDcImAJxn1QBfm
a2OPDtM3fMXzhQStu5GtaN10AcIetl0Ak58jhS/flO+WZtuI33HGGueig882VT1G

--pragma protect end_data_block
--pragma protect digest_block
rz50bVLXZAkS+GciPq/OG30BqSA=
--pragma protect end_digest_block
--pragma protect end_protected
