-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KnPy3yYTo1SvFHpcdsaQy7k0sq3UYY20OPuLqT/tkIQAUxuilS3XJY7zqTTrss4CXTZp51e529GT
8JvOi51bzRZ5i9PDmvkQ1XPm+3AOTzeRed+tQel4mMKr4xj6h2xEarfW1ajHwblyDTDItjkM5XJS
WiHnlKQShrpzIqGHsRK5eFETHma8MGE6RZMcZ1E07q2XUsFU8hUPflRXgubo+PqFDX8h2O9rNeXs
xy6jUqgnuhHP4ncqAFws/HluJfEKGif9t/AyoowtduvXScjaW6JT8P5FDIaoQoI71w0uUSHQsMWv
fSbxeoXbnsoj21gPqaj/ivIjirj/kmZXnQEUjQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9664)
`protect data_block
Qh86CVCE/mJ2xslxdGmKqHdGohGL1aCfE/ZcPcgJQujSPwe1Z+fluMq2MfvnsZj0U7dwJG9mENfd
asgnlRAiFs8iZdtIBHxC4Ed5Z/cMwNe26U80iBZf2Y1hiiG5ugiyS+7m2EhkFUK0oUOD9w+0Pa16
sYtpducXb14H7v5IvMrtpQg1aeE88EW8AUVB2GRCoQQP8+eceOfuUjGIs3EtXyOm8zhMRHA86OHA
FEHTGke/Oq2kL93Meb5cJMiVb0SRfXldK3kt+ybRahh8vd+j5HMt3I4kLFEtu4CmizXoMJlG4Oyk
6FAUl7BM2lWXZ8mGDbau/6JIaoG+1Z/p0w23xEoSByy6uuCvjQYNGhQsiG4KJblwNWRGRn302uYj
ZdqE1SdwkGpKfuUvfsrjp3owAFjSnBa5ca2wn8vhYE8h+aes7qrLiyGV42mHyI4jH2ojQQ9iPPxH
BAu0eRBFp9pIXQlKFr5/3cJHb1RHIjUnL+6EbHiMlatekR5OF3u55l0YXGTJzr1k6SYLeQnujQBP
1VaiKJOlRlZl22S+AtC0B19e7XAbZjz1ZTOmzFlwdYpIcTWayHJ8r7xBU+S9IkIRYQioI8OLs1VB
U7dLBd0MoNShKW2Gi7rb6jd7b2WkhVa24m91PfDM1QM6cg2lEgike5QPS1O3uNiL4aWGmaLHQiND
LhOeQ/xOxpcXdYg8h22Z1sXnM6YIqHEUxx5Kiv7PmjoW5K16z9/1qK9i6cSCVLLqsydoUNArS09w
V0s0DRN99m0jEundZdW1++wc1FG0Je65LMKO/ajwAqM24KFPzO5FEIz9Y+2R1uCsFdRMFAVqqZmU
0E2kHgyAHVH0Z+9RnqaHWa7Gbm7pN0PV808xF5BbgFjQip7bXY6D2hbCwMXfDcdHBGc1FlYCq/cN
Oa/4uhrBO1SCTBdC57gX7q/Kiz/w72MntMVAuiu9xQ26nNbRo8MqIrokF6uUayvXLtgm6JSLQEmr
dkanZZV7rtSJOwCuVCLAXAJockpAcq6VszzUicveGralE82sLn6Cj2QlqS3N8FQQVogF5MZmtR43
kLTTjVMSqn3OFm35kS7AXfAOu8YD6je5yZMQnmUTabWO8w2tbgC7JxRJvD0jK1RnTFbuq6bjvKj8
8xwma98QB/DSob9Com5wEqR9eus67atfenP6jjDctg2JOfgIXUfsqbA6+V6lp3DB5DAjBgPKDPKw
iB9/aPc7I5OmRvu1z3YLFgyqBvbyS1QCI36vElBf9+d3z4ZFgKM99hrbg9bCuiFL1Foc3l7S8/Rj
ljlXP2/VBmT7lL/V9i/5hYDqMXy09bFJSDz/JZ5EnWLFvR1JZWPrVKpNUxan4cus98CcF0JOBUyP
zU3PHUecMdCfrWsICl3REkeA+Hk8XAh/1X9qYIcv2BUHDoVa+9tavKH1GjgMM3xIAjpkdfNufEC4
mtX5OlfORzSts6JoXP4/YNx80YLnnC0vJpp7DBRSe9k/suAg2JjYTg+7elttQ6I8+HgW0l8ISmU5
R3fTuzOMGqSj34OwusMQWt+2cOVG3lvKO/ZfclARerLdLGiZobrtfginKqa77+iH6YIVA07eZEN8
jnw/UfWZMLnLQrrPqnZ7t3SJQZgIfrfyFsmqdzRT8XEX/RR+dkQ10o1AcLlttMc8nwGXLy8ljbTy
4+3B89TwYDjmZ1Vrt97j+ZhY74glKrKGIb4btvhvBnK2X0Jlq1+J9zUgQBCn2ISNckL/Wls2m6k3
RxxctVFGEvou18/+N0qpDrzQ3q//WvAjRzao7TiCfn9vIxgePxOtlYuTuG3gBDP9u+yufg3biDsS
1hqQrLfthBkg29pcrSY9eKvMjKldvC4UuAdHID5vukxcr0zfxtEQRoFpkAICh+aO+WxlxDt9ztD3
H01WUMRHMEKWvmJgCsd8leZ32bbFV7FYPMZ+2Q0Mu2BylxtHcLqCVtKLa9mmxihcoM2N6lxjAw1m
Y7IwFkVbXMMduZLB+nH3CGl6AZfsOo8CtqMVpnDRFgEIxBqRPljK1VUvAwWd2J8nfq7uyTqjU79V
KPoDMTU6Ncp7/MczMyvKYKNYtx1fTf3WTZZBdt9d0xSjOHh56a6cB2uE5X7n1IAus5DQ4Vsls9Kq
h3Cfbi+VAW3vNHOKGlrypOoAY3z9x+y5yxN4CFRgufi3kc+OC9cUsjgiqdezIH5FQsCbN8s1UKMB
c4MkbCq+UG3v8onSvPGwYqFeHYjYL+TAGOUXQccSoKtdwg4P16vZNenPiQ7DlYqZbx4BdUONoutG
qlsZEE0Ns0faUBS8bsJFbSOb9oge8wNOZyefA8VOIhEEo1KiTROFoJYOPfRAczGcBnrgifj1V1pA
34Cdx3nYneYnTq2TjwGucDj/HhBgVD+mcr6x+xilh7kgeMjQvBWlYTnOd6HrzEdvEGU7/CeqGyBx
G/qUTdRrAgSNcEXdFr9tTC0T5FbK3jcEk6bwbmvnWSNf6wMimqhY5Btj3Z8Pky132DuG6tjijenR
FF97Lee3R0W6sK1Q5FeCQm4mQkeKRlXove+TmYz1vsF9ij+8QiCTKIAnei66cqqiMScZR4ObOigt
xwfhAIjGGhpcRJTcBcQ706KXS4x9J6MtE+7s6Cg6/Q8o8nMxGdVd24Xt0n4Kf19DkIC8Wl3SnRH7
1nEe4YiNwMKKTPgcJHm8q+7amWfAbnRrTTAuXDXfnJOQ95/C5YBvKn/1Iw/AKElfXYUb2/D0lbl4
LwyYeczj0yiMGvVBpOG9f2rf7GPgKoY/j/FJMlKM7byxjJSUqQrwFURUSEbxtMEuOaHMQeP1GKyd
HIZnp2kWliFdtaIft8Y/VPgQ+Ve94RA4NmIEIC6/jWJPCKw7o6QayXYpdZeHRAvcyhNfUQPtlJrB
dRtr10NeljlFzRTImQeMFKSkOGnbCd57Y2hizKI7MHWFOFjjXGsAVJFajWvseUfxAjDK4PsDcfFY
ZxSyVpXIxONI6bRSotov+2lMfBrONcEKv74ehPfD0bLldnvLaVjA6RH2Kh8r8KSHYJPCxjVYY24V
s4hy+drn3Z29VndmWQc8s8Dqtw6CKYIZm7/nuCGVDTXuLMTbpwyqJPUuHNaYDgLp63a1tHasFFzQ
FinYJyjDZs0ZfmEc81keleIM6uDd8cgXfHAQRAr+R8JICb1oC6+jdy/iWeZZdc26j/a8wzaVenmR
KP+k5m4/gWHU7B+dkHCMeKXVk8zxbkE1Id+VzIpRLghxAgi/HAdtp6qYFi43RilWVHEedkn5aIi0
Nvtic5EDEsu+tvG6uR5Au/kKJXqX5bMYD9MdUogee5OtLUYXt3PcdQABaDvtV/9whqqeEkbBBLis
M3bfmvLJq4Ps7XwWq0T8W8X0ZTRJJKe8ENUXLXQB85MGwvBD4VF4WNCBYRwNh6rw/FH/+DMZhWCT
WkpZL5vdr7g262zbwjFk4/QlW6xtqE8L1Ad6uYuMIKsIDNU9xrqfg0wicT3eu6PgZdCU1hCwpqit
Zc6X3nOG6r2vzq0zg+XK/AZdH3T1AEMNSmjmN3AgeFWZDm1KhbS9Z0ljGuKmN4eus5wl3uf7fMzK
94+YSeqMwx+hWJrrU6ISOm0V+BpPYRnnhrcrJ4HlyLB70iLSK+zC5tmbOKgML5bvitE1JSUqHo/Z
rDc+miXCNtAOT9aT+kYwHUQrhYEswkqXL75/7/Jukqo3DHUfJizPkibdlelQ9sJZjIOEqnGbiQjn
TkRYzpTUaI1giI/K/6P1nZjSGakRjuxEcLBKJHIerePlDAQYYAON8Z2VM5e5n05vWXrxQFCTa5IO
wwvmcCQMnVh7P1mOzY0kSsS1O70MjSBgdkT2o2oLwQLTxC1jHezSEMb8dn4tNPS519jVSZkq4o+A
GZ+U3K/x1kpQWHlvBHbN0kGdpdPJ/RLExX2piVTwTIZwcoaH73L8TjNOr0/XWz9TmliezT7cG8bZ
/ulqgU/f9WuejI3sWM6n5bgGI0/e2tQYEs8FLCV0mBCrasgJXwrvMLZEQrojZBwH2eE+7re3NuRv
hje6SPTO3NUkL3xocjYlVbPFcDCy+5nG/h81RS9PuYYqyWMagqG/XML6MChhxXSOEw3Jb3lczFl5
YTgRXncISAiaCMFr865JeH5FvIvApmBRXDBYWR0X5tD/royT14AoYosLLCXNHMPcPaTqemHnVju+
klSqW6cjcov37a3qgy9KURdyBjBbYRVmdvd/vAV1oCimyPueRuYahJl+sqBHw9qvifQrmdI+jjdY
T8G4eBrWbP6MC4NNIHBRiF12o5JfQZ6gNk6TEhNQnf4BT6GbikQ6M+7cMVX7NJhdXVAXJuF7nTj5
4b5PtrqjkcudH2AV2x7l2NGtwrAdIsWEtPIwh2T4f/VB1E269xp/l0H3nGTw9v/p7pJg7Rvco2Bf
rQ0RMKDTr3JIG9S/uTbixC+K1yFAVX1fX8+9nokQptzbXoGtIRCqkCR78Zckb8V498dNVTzwPbYR
XmoXLCCenD+ECmAWa4LSnYBABGo76kV0Sw79ctNrxDJN9exWFVolIbop+t3nhn/kjoOzGPhmRUw+
x9m61VDG3kqqYmjSY6Y/OX9uJN8M8Ro4u4/VyVhOj4AO7Oz1A7SaJa20a172Kr32ybkIZfzLuyPR
jr4YE09BUeg9od2IJYG00usBtttoaA28ansWGv5piHfrMXeDPL0efF08msPF9m2Z6YVJYQqbCbMR
or/BblYaldHxyZKRU18CuwVe8gWdwPKevpZtomAYnkfppOWnkpSXnzt+z/tE3i7vXKra7LNxH/lw
lkD1LCp1UTmMzeVDkF9qG+IpZP7lr8DusPuTnzdbjnkLrWNkIUYqwQFTUnZVCryjpXnTCH008p4t
7/NijsXhia0av1EGYQp+/iOVjg4nc4lU12MAOk5QRWF5/bneqKOa2K6QPjFkayn13SYMTrbFfdVN
JjAf6HmGKo0MgMgL6QMPhDxltx+owqtaHbeerT85WNdF9nvhMmamsGi4s/q5ypcbSBp9Ah6PMZF+
wKpHd9ajmPcVoBhPcDqgVqEbs+zXH+Og/lVPOhrZkVn0H/dQvYs++PhlpdjhOMtTQFAfXsfqptmp
LDyQ5ekxW9TkUzqqyTVvDZFNyIRc9n0PmKt9q2O+2OVtlUa+LgMAsOp9LqGZ2R2KlgwfG2+gaoVy
b+h+21XSPEum+hNh4/lhfZ6/1W+/yldCx5OKL/zZl13a1c5v/ROi/DWqUgZe1qYDuCHmsJSewHoi
zG4+5uKRd6FeXQw9J5ZKtiaTMaoQRCLaGvTj+mudgeY7eSRHxR8oHDAZDVtdDZdZhKGCycbRBP07
/Yhz18uFEGKSnDOAzLNJ80oyc3dR2NY8LMSCUcr43yDmzyqDPPscWygcSYTyNefqZbmckucPnH47
TAmwwBVsD4z6IjCFWra94vL32KJF9dVrADQriMFXCcmUFiaAHHlTPeI20K7Lb94J8e0K8TDN8628
9+J703KjhZLdRhGAn+BdGql8cJq3g2Ljk/+oM9X09+6CmPdKsbNcTyLR/dmk7RDsLyw5KA6FOe++
qvRTaeFCS1PVi4o9ZVTpgQAlbwc7CF6hOzq7mR80794AAFxnttyjcRvsOdui87pfcA7BnZjSIc4k
b4cRsztqwqBVLPIB/UutxOyKb8vyJtUu53sNHlRMnS1/pwrCJUz2z+/1tgGlScGWooxB0GeQDNn0
YbOClrIOjfBscTKxMg8qjGnBSNaFCCgKMtMqzIJYp7a4NMkxzKJB8ENwbrxCRMz8mTYNrvjAtwgO
p8EKJn1/QsfmCRvEjDMXax3aK6kyevjMZg6Cd8Y5aqRZ8kTdxy/v8Q8faxyP3sWkVUy0dNyvqcbI
V6ENsVvKSkxAsDQhU1arQ+DpdHWN8dZ6KkItfL7/sJOj5mkIflLikjsA0gly97ccnw59+zX2h7Eh
Lwc2N6Eynl9pJknx+ayqMviAmo7TXbKQ0DKO41kVf0nJp8b92ob9l8i3WLp7tAiQ1BiBONOHIwvl
88j352YxxyK39mgYWdggbEi52SBEcPaySpidNWCiP84k3YbpwdPpF5mO4RlGQ6TbF+GLpUI2lyC1
MFcxVsVWWJxBprbLZ0m3Dshh8lPc6TpJEz0e2aonJulemZwph76cJJy1OSY40n2kjRmKGlIEMoRz
6ZduufqoXHLDu2lNqgJgR6vYVk0Es1TTSbJDc0JZxCPD2DyjwSRhcZf9uAcQJOJJMpt5fEk6XKal
B7RC7sZ9Ix80bWKUvpK8Ef+Wq+kAN35VDKNzE8NzYpFCNkqMeq0olh64zB7sfSgtNm7u77HxU2KJ
IoUqXn9DR3b4xO58gKnGBvW0d1bxztg+K8MS0hKRJjSAGH5+KDFyDaQ9bL7EtFTlFgxcorOsdW8T
z4grMXHzARAYPQBhkuWceD9WX93850IscdmiZL+z+4x5ApABD1AlKlPjsqUPLkmbe38nN0m86A7U
HmNwolofQxS0dbmGTlU7TUJntRfSga3NAfKmYn0Wpp15nN4lCzF0ds6PC2pmljpkx0LLErfOctsU
dDFoq6xi/Lw2p2ZpfUi1I+OPXKwzSTvanMLGfypqVf1tHTvNBpvGKUKJzbY7jAHciSPbEUgAUtpm
FVRMYK9KSINouhLYFdrorSahhrNmqubVC5JOsRSZIFWzGnD5cmpex0Mc6yaP0ZoQ76KNh5aggC7y
iR8GF2QQaatItM1Oq34lFoWgkCYN8++mTYUrCjJ1hKWdS+QRoCOs7w34eii9arZH5kd8Y5YJXbP+
rtaKRa4V6/ScXMKig76stwM/b1zdy/EipffSr2fvcL70m4T2ZgpITn09lfU7PerJsmx4Yjwb8JMv
RknxkrmsFZ7R8RN4xDTL4ZiylzkL2obHHQMJ/mV/eF5tPPJcZydPoOyxNk8wNyMSF8SslZMu7rTF
jzviK2Z2ax3FNklkWKO7mAqBVX/viYQDN8l5klVo3zUM/t3PEACnkCusZsnVROjOIPbZ4gaJlsLO
NAGv2LMLGvA4SV4Efh/KilufM3Ta4sXW7IkGjqnAs+f0Q0dy68xCmVul0FBHg3sRxGpxzPCyqdnK
mFN1+hIy10jEP70hu7GWwIoqDX9ctWYTgLDwfFaSiFjC8lzPKJXbW2kGkgjlR4G6QMplcxn/FS4G
5F64rdmfQsuf1zgTm/LMDoI42WVgt2zHPwVuoBpnZ+EsvXvJaV0+4r42PJK0zhGnyNaKYTdQVO0W
J74335ojYVVjj44+5KvY5LlZfo93kGKjp4Jj3NyKxGjkHPgQShlo3lAN8g0qGUMGZQZcU5NRxMjS
ncRSAjBGcjtvWFbyAIirDjdEUz0QF3kTvC9rmQi5a/3//4eYEp7mKHK3aEXbE53YnyG3HdczO3MX
UxYTcNHulvVJK25UahkOKATn+rDh+win70YBDZJuR6oF5jphjbL64YSw6T+8mX0Cwu0xvjVpzTsu
/WUBHX2cfNIFjqDb3R33kDtiWUZgJHv9Cj6P30/AOse9f6l2VZE0jwwFH7I1JSG7JiCmNwweROQh
uJEpj4TSzLUq+L9ULIIDXqFRTx1GGv44VaXtJb7RG2BWsR5xACn3EOjY7S80Wm6YtdwBg0KF4QI8
yrx6EqX+n7tiJwwk8gjZzcGNHOd5JQpF/uaTsbxhU1chMFC8XlAUNIvKhnwGyJ7EhYqphS6+N9zb
WLSmvoskyBfELtZzx5PElX+cdYMz75HwvPaBvGtt07Qocq6CPktVaIOz0mh8/daB7z7uun0Ur+95
TG5I3DxcORidnzhcEZEzmrc5iS3zFzxMHUZcXF3FdLj4T5uAZxJUNq6LKvzntTbvc18+la4gBkKG
CtQnhIW5GQYE2HoLKNGTswnrXChSxwyQTtiad8xDrKS43kwZWaY5M7wBKwnRtM2Bp9zExmT+m2pO
acY5PAKPOK5MMqNwoCnoj1t6ZMxHbYMJAukCY26x5zEK0/MfXAQDXPC4x3yEq+0FDb/p6UnKq89O
D14l4ArYjgzL1irxrlj6Ik3JCGQJI/M9apJ3k5NEu2G/DQkEUq+fcA5cZFxh3LnlE5+XMTXyehAr
ZnmAcFovWcxtmPh707WrJ3Q6Rwamc1p0sKKjfFfQ4ib+rcHspEo9p3shE5DW4fK3t+rs6AonN7RE
/Bw06jEqb2ui74pulG4zXe91xYFVvths8ATu4tgvh66+CeHkxl9/MA8g8voQ3lsEsoQDO8HoXw3l
kv/M9KxunhmSiN5BUbufy28oYPpl7zurC5RtJVOxkVpbgGqbvqsDUmWGnm3IYDRgyd1X3gTkqJPo
DHG71dzKRJa9uhj8FMcRpv4V2KulNWVls4FMxg+impotNErtrT3AzSTDUSCPd/d4SwjNWex7tZCI
TtYRO7CAcwKZ2C7y73g2YZqPMdYJOzBhEGw0/k8vKrioo84n5UAPhjPuAj3UsNNWmyS+l+UsumTw
mGgoh0lEoczJ+qpAJB3WGl8VrAXZxGlX3VEumAdSOoq24yxp6arvi5vTNdhIzeJhy+ce8JE/yViF
JmtBeU7Rxj6PXr/nTlu+rjG6/Rq8T941o0/N1sxzI6rpOot8kmXJ+Awe/NNyIt1rX0BIXC7ui7F9
n/LQKEmEnbtv/tpmueQTJTsMDhLr4Mmo7SbypQDV2avioI5fzsBpR2Qcl0lZW+70OGqvgPVebcYA
69fEaq62+PCVW4Vzt/BWMHiC9Rt5SPpvemixctz66sRpjSIrE1yJ5ntu5mkZO1BSVrU7PHVw9c1M
RYLTI8jGNAY3B0TiIK0IRVAx7+YrpN0hXUg5dUO6Nb9pJm5CXeZxkDL4lJWgQnwP6VOBe3lQOy7H
modlo1Jxt98Snz7pVp/UNYJhK8J5ED8Qxrvd+W16Wnbs8aiYKMJzybVn8AROzsuH4T6gRpV6Kspu
dtXKAiZJzr7BNr1xAO6Y2tK5tX4PibgeSB42LsIl39HCgNmTugXOBUcTY1/e5QF4xazi3FGoghIg
09d3KvMNob9scXYO/eGSzFVea7vVb/B7FDMyk5vilote4E1k54w/nu1pwTZTgV9Q0ewV0jfaAOkH
pm8duulyQEelnwcUvU0K4lpJneWjFeJPcWUTMMWZMYdhAI5/yVdLhnMmctXoGp+WxfW43QxRHatW
EgMz+vxN0dXHFZqydig7RtlfkstWC85PU1O0fKrG1+G6uvcjsNC+Wa80h5M3bOgmLlRfdX9S+dCa
uxOJe2Ytn/k0JxhnoQJdKXQzlQ2QVa2nPQr7shYyGcAk3YG1GUTZ9SY1X1HXEEqMzkJHudCFk7wy
Yi8FJcQakrZMrGGLHEYygO95cTCRhD4LKrbSKyUuNdNXUar6fHxPvCq701l6V8IFStho28JPHc+u
7P5TQRQQtbgVJmjbaHd3S9cWziepz+uoo3MATORpRBKycdSDpIROj4XXtKFHO1WJM/jofd0ojUrP
4dCkPFh7N4rNebQFG/vk5NhViB8Xs/h1snM3S6L//ucjeOXxFMRs1XYZfur2ASKriZJ+WH+cynzf
4ls81/GQThWSXlOxUtFbgzoOGBiOmRHrfKxrTL69RJEWLfHSWiaim4Smq7zFpT1OyvQgetsQ/384
y7nbKh5pcJOiLd63QI5+5o4ZndRb5yuuhqymSjawcMWbw7sVhHCc1WELMww4bdRsd/zcwcR3ajj+
M2COpcqyXjqkibAi3JjVNl+vsFJ6BpPpX1qHDP9Sv6B/OUkmasTWOfTfFAcgJNAyQBloiMFjqvsc
cE4bd9C2+4urkSOqWF7PtmejpbFzse4LabOcD85P2s2e3yOWWM9Atm8JRAA4Q4oCfemL9FtSx1B7
Y+ONQ78zpb42RHBbmVrUGj4N5NFsYML2mavZeGR3B3TUEhDqg3Y91SEwAhYS2vjn8E6vQjISpbHP
uzBePGb9i5VD3j16HBsMBt2g9ufUBkib1+UozL1FZHGuOXEwOn59g64A/L+74iuLsn2GP7r4C3pM
faVxIdD+SAITbWY7ekPpbt6Ys72tR0miEOplhED1J8v2GMOqP1LUwQf9fFiWTu4j8jeJUjsOpjKv
1g/iDBxM7RIw7FM/7kr+PioPGJD8YbO2F4uXgc5x304FMdjmajhWuNU0GwrFWL6Yl6SahHrQuXpf
eA54MbuVoxaY9UTV760wDLH1GBlwxCx25fWXAh/vpLtflMwI4K9XDj8UbI0/ktbOI1LhBOipCLmf
WPotChCW+EKe3clZeK6a0iC/dyz5zzKtyRSGLxKmU0Xb86bQLDT1kuZs7PNBqMCSPeIYU5Rw+UpC
hLanWg0NTVEKCL0r5Vr35bcb2lwhuzJH+t/fX55dle8mwb8taRYWFbLOe1kfVeQtkY7PkcYWiLWd
FpwseZbPA16SeygZFiv53inTCk0disHgxjXMleDrlxDy/luyj/lL4Oew8XaMB9XwCpLCGikQLFaz
ocA56uu1bVjgyAdbLbAONQhcKdMVG24g4qEcgrlvd+IC/fIGKnJp+oktf0+2Cr/EdIlRiRSaJdqB
y370V+fe7HfrnXslL22wH9h4N+uw053CCbrWFQ98DqApBC2G973LpgaPfrotjSTsUOedIC6f3b5d
YrN5FdeiL5WhfT0+i0GkKZwHEHZePbvkt+hdufyb2jyzFRkUNFquFQSyEE17Ca01e3lltt/kPXIZ
bm1umTF1U6bRcV0xY6u8lSqjOA9MWmEbyY62nBBRxg742HGI8Z8PbE11vt0+LTo8aDOuCjAEzuk7
G7A9RWeXct10W21PVk85C+7wOJzXeSjgZjI9hWcj6ZDUGDB6pVMhmwFcCJMmYv7qfW0PYAyJ38JG
SJ4YOBA3ubDgHyFVqnemqP03D5ZFLBLtjzSbwv6SV97PB6MX8UMrAk3LJL4qsbJkA38QG1SuGT5c
OvypBAvA/RQlUYa83s9NyrEqhHsy7GlRFrCtoOPYAg1JHGQgWC14rHsA7+7CS5xbA4ONoCjiyUgz
f2+qoSladJzeEPgveLPAoI/fhXIa3mvv7g6yBv7aOsK4PcI+SUxCiI2rkLUJQ/b+QocJVGHpco1O
OVxqbiImuu/yNRu3suNhgm+OzCcU0kkmVsenxQjKXlqrQM6mbADSi5tLc24+2FW9DNokukY/JxkA
okkHKIYKxH7lQ7bWf6iesgw1VfsuTGAeEF9kxN8yup0e+WjwFvqJ6XL8Cer1d7YuGuQkZB4EUCYi
vEeAczI1N+nX+OIkzt+gMj/uMIwbXx+5jtBOjdc5OFwr8yaZp9fgHvITYj7WtduQiQgr1txvxveI
RoEkufALPcLITLAbBkttBDHIwpoge4k29iKT87TWaeJJE8eYWjkNAtn/C3nUQ3+SddUyfxuWqCaV
AXHbhQfOrcALVD9LCMLz/SAAaV/qYsWWqvVFC0lypWsxY9iXQqHl9wiGDRXvuh6Ggywn6OOVdHHf
K3aFf0bRVIc9EyG6oTf0o0ZxqZ9knCrAk+y91d9pDmcTS2hZv4V19741sIpIFtYrPWijdb1ge79U
8/q1SkVAPkVE129RZYzGFUdHf+i21ENMVNuMTaP/QOaquZh4J6WxCxejES94O/SL2Q/fYFFWwxEf
UlBLqgcDL4tPXE0b5MyJtfirftMLAxV/6dH1kzECNyGBveitFautL9nCQtStJtwuaDXxi4JptyY9
uQzXgpWhvtUP7nBN+897pArPPguK1bYB6f5CdpVh7Sr4NQvTf0aiCKgViYlZPLmyLxxpBtA/RokJ
v5pfJCmeFzU9NLs62jFzuXHmwuzA0aaoP0hD2iqAPm6UqyNILpDQb53i6P6pyQtisfh/YefdP4U+
GJozWipt0o/x+5jJNWVRdEZRb4PSS9LgqvO/zsB9zVO5XXs5u0ofhzwo4/QUtL9iQG1N55rhAdEe
enRMLgcomnK6t9mHaYoXg9YPBQ/fvnvK/haLIO7TIYG+NNW26jpx+frtTgqYi7yNtqGkAix45TLs
tFSOhb14jPKUEj3tUssl/TaAGkZ/zK40u4yIRkTKlXvjrq5Cgan8Dpi4H3I7zsf8tAEgzXwmnC6h
A3Cz4+M7dlY9rcLOZPmGcDUitxAHAN0Byu0291JpeGrVS5zHoLx9e/LbHL2AionAPXYKhAVE9FVG
aolcgFkYzKN7K9FrDYVaaB43V6+VCtXXDqSRZ4pkzC70f+YSxo+/A09b7Lig2L8x0nQb9jUXiMz0
Bx83TjwauM5N+PGMKOzF7uhcQo/mPn1syi//Qu4bvQeJJWMX0KkZswhxiMoO8iukcvDI/CTgjand
SL4sDEyf0URe0tspXXFDTxUuKV0s+PKZwWAFkIwOOqjvv3usggRerPOXJAPsozeybFwXQIfpb4ot
GN0WBUBUitayAjHiznuFGTCvFdLTkQNabpjGBTVIWgskF4aZY7VeV0Q4djiRmmxf5+scUnYIzchM
KC10rSD6AA8YIQPMNOp10LfCymsfQFrhyb5pniXWoduBpi/b4fNAnvoMPHXm16fcKNQkEpfAoJFl
NOiyGwqo/qn4dQsAfQ6tw8jiC91xhn0KVqXKOzI8mXyFByKZG8tQvkWPkIIN6k4dl5xYtYghCcah
f8qp8eKtUMTlnYKrvdlKLzwwWAEFDtHoXvhcU3dtei28YG6BLLoLtkuH4fXp4iW1jQe2yjR5pE8x
f6DSnbxLUa9UCWQAdrNZ1d3p1pMl0YNyQ6GaSeBPjtJIu2KhnYCvA8h1ZzAlMrfH/ZIVCrMJw20A
NxGmhk6mlNpdRWVehN5lwJLuVb2MCup5PvLaceDmDQlfAkhYCOViwzv4GWFW+IJpvTyba4PDvByr
2iX2htb7+3j5zR6mI9Nq5u7MmZ/28DvBszlzsSWcoV4qIoxfZQV86WDQAy0LK2feGR1tvsMl3/6c
rjjT1joxFe3XO2PAmHc4jsER5FkU5Z2ugH95srzTew==
`protect end_protected
