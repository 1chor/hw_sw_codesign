-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
WbCn9Arxdoln0Utlw3l+8nkMAhKxAuoYZ4UtkzgZ67SCjn5zSdMdjuODrNAJv0Hn
RGYl/wHvUSz6r5CJnv1LZIK5M9cbjGXejrMbnKl04aqLxtL/um9k/7CnX8fPm7eJ
XhnOcj9bszDGGzWH2NSvl0YNPhcj9+kXkcZHTf+0wmA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9808)
`protect data_block
h7weKEgO1bIy8tnzKvmAnfnupCRjvdpzDPDb6hiaeRvTqJDD+twlpptGvpWT/YHu
zG+tMl00XRSjg9r563x4oESY8lu0vkwYHnyMRwQgOSB/L0n1Jie02nh2pR6i20UZ
lW0abCVSgUlKsb5ZJ8DA4/2+p7Gf88zQiyNOlRXJtCagfMcv3Z2JBweX29/xfB5b
lzaovzuCVNCsSUutTnH2JBfPsGzwTKj7uNf8zqDVD7/AdAW1O8yyL756K/Cfi4oT
Z5g/JcmQaA+fgZda1tlBiSx8J4Ljdc0jVc3YyYbPmOvDajuibqw+MhA3XqYAoLWc
+Gxg54pRgcmotgMMavZMMeeAocQbcLJf1hKZ6425rYaELv67HIvZnlidsjNINYGz
rXMa+Eh3tvKBVZunk+30ySy/jepQeAR5E85vCUEQ3/36haB1Tz00p0yCl1i7sSg/
EZbI+KlF1sd2uQI72EY9uZqwiM8cke/0/umXOzMunNASThFUDhANFBQslCDYsW0O
5vUWNoAYGFTP8HSnIjM7Z04aCQaRM2EqCEsP3XczykpxYZAhgoHdtyKs5G4q14BB
dUVl6r/ubjI4vRUHEPv5rE3MUWcDTkPlQkjh7oEHUfba26mYqB/9Iq+KyUgf+Du1
qVQKZP8U4W/VaTSR8cFkENnZo9BTCv+P9skzNMioLgDF3sifC4a4Y7gYUXDJPXCe
TN9XicfvmD8uMg+lxOjW64hSShGx8fn07DPLsJL/ZlC/b8JKvbnRI26+jyrPLEkG
nIi1IaxVrFzSjjU9uP91Hlm9QcDL3IKaL6bsaSExXelV36Mz3KteU2izAgk1ZUFR
Wt0TBVVcELnjh3f0aZyM27qPgTuP0b2nwF238R2cjYr6oYyu5/YBzc7prQ0iJqBc
GKgiRiuDhAjAm230TacFp3DX4biELaIMNHbHM3QfOVD7m6ZOQS463EWE1+mTBpC7
KpSVi/USZ9y6co1Dq26R6BrJmKVTZzEhkO+XF/n4YbQ1LYPZ93IefHTs5Q5QqsNz
Iw6XIsmbcG0p8z3Cg1lNeHrSlJ6TMHryRjbrHMz8AWfzC7ak0cnOoVCqDt0OxQ4A
4nmjkQh7KgaA+dme2PlQfzupN5XP5ul4HjKvjQsMzWBpk3hWGZBQLkT+qKgeK9jC
uRGiQqIzj2ihm5p/c7ofkCVV20KBbVPPpLK3VhpFjHR+LTZcHgtC1iqakeE/TUup
as5EVCfPhlNnZaH/rSg5pKRz7n3amUskRNtbukpPlkgMqcT+rR9+HCO8d/wsA098
Xm37aQg17qAjDEqy28/bGHzxetXpu82ZX6rjKzdlQwWgi8BBQsPXv0P/mIPLNsT6
U/FbDTHc8Ef+KhSCT0h5f5Sa7SifsVsCJ9Y2FNiKobq6NWWwj8wK1U+e/vgxJppy
Rn0h0fAnVc8P0wLjb1NuNNTjpDVxRR6LAsrAzWerD4MyrF7xiWoOgs+lK9MZLcXk
1OCXV/+ZT+gM2of2hhw0phMF/madKNw3PzpTrbluTBDN3rv9Yyy/GwXQEvBBfy/c
ISlrWDgz6od/QiF7tMHsIRDuPER6TJ23r/ZWgwiJajhG54aHcun0EqlGq2i+ZCvX
xyn00+e8ay3gIMKr3R/VcMxAsNVqJDhuB7SQCn34/TOUJXpnOovlF8wkcBDdabtM
5nvAELTaUYejoKP7SfIwnyyJwdChwhsFPx8zMpbY2f1yROSFk3G/HMwDe99SVjzy
giy+8mRVjo30oq5e7dmowBCqQIH/ERnQxeA8umA3vsJFr28Cv5Z9NN9+9GYcHhT5
HQ5p1rwLb1LqPu/NwStVdA4/Yb1e5aHFhHDoJTQoHNz7qaTt2ut2QHS511PNHr00
qZyWfgVbGdeqV53rP+UqiUb9pKSuGWt84tRwd/+Ih0AvkXmo5b3zuJp5L5xm7xEk
bnNmSwK2AgzOIEwIKEAt7k960HS873htwm2IkSi2oFyJDp7H2FMI23T4yDb3ObvX
lzn3M3AQndJ/AwCMPLLdXWsLrmGVNPuDCPwG5OfrAsoOg79jbbJaPLTqVvaYCz34
2iMDrXYWSImaUh6KmMiM6e6cOPHDNF+MuW5lHc1CDjXjBVhaEJAk+bo93MzCILPi
OosgR0o84yn00Rg5tm3LrAqf+MxFlMTT8HBMRtuUL4q+NJ7a5hQ+oxFTMq9CJOLH
B5BH75/zhnGSSS1yUqFS6rRBaRdocez9zHBV83uj/KltK5CFS3pPLV9jnvAy3EYJ
iiAuraQMDVBAnwrEAcTkeJ/3ZmVn7GqoDS5xqmq+/63gU7ZaJktsiZCis+v9Kaye
ImM48JpoYyFjwwnm3l805GlAiRvw8wQy4Mtdl7icThIYznclzKo8gXyUHtvrP67r
HZO+D/TlWSJ+4YEisBj3TnAzl6YAmwAnuB8AwOg36iQCEC90pniZHAAPVhK7vc2J
+xYG/QNUBLx5DGot3i4+nCCmkX9FVaair93a35zMAvzpJb+IPN0uVchrvRtFnPGJ
uU3S2tPmNdVtUV7bB6qQT1PcITgDOHHS1myEuitB+NYgONMsInpKYV4oyyb2Sv8X
cAL/KG3rLjJsISsB704tWpF7d4NeE7CpNINaEeIy56JO5B8SrJahwDzVt0R3QMkB
10W+9VW/3Ozo7McBWOkNV9BzlLZ7YTe881IF/FUCSnRYPwpHzQ7cagPs+YmroNHl
4YQAzPEv9/zLv80xCsTIXu3pGmcJiIjLEKxUgLiVZoUya5hXvhJ/PY0BzlXb18+A
/GKEhxPj1wpLb9Ujzjl+kt1QVyRrPoFsEz3ycgU/smkeZfZx1mF2VJt9iXrj7kg4
LP10rwPkYqyNveV7wk1eEAMMjFlOjAfeyW9aUtNUyIpdFbY07onLe1ShXiXou6hq
MUa5d0YlidinJXDDh7un388nPcRd+0wHnkkgp2PVYcZVntXE8eK8z7WxzEpIIkTj
iSnCXy4PZ34MjtdLMAF3wMSTmH7d2JMTRAlicqalrTmwZFJtImmjeZL2XUbZ8pP9
xmPmnIvs+472YCGKC0SAVQkl/dVZQ1LZ6tFQAwX9dVB/SEQ6QqzAH4n5VfNlQx4y
xxUYGuTUvGADoalYiwItU6lm2UfXd81saF+XOCmYVLd+losz6+BdysjrkQqgnY63
n58q7MhqjFdgXCG18U9Bxd45LmKQWNN+gDgS1fdhRoZDhZi5u3DikHaIIWMsqltF
811vAf/xBef4HCjsxIgD6cq4gPNBkW37iV6fzo8BCTstilCVyoT2iL5WORVQ1vuM
1BxgtrmtjrrRQyurQgrpl8i8f7JuzPKtEvETyikAwTTfuZ7J2LdoMPfiiIrFud3r
afN3enx3o1EUUQ+uUDmIOjcriPNlMmtI/bTWrX2mO2VY9rCb4//ztyJBz2hRJlaA
87Nz9TzUz26wmQI0PSL+CeaGkTS3zrFfIBO29n0Zln0qI7xDT/XIBPNlCldgOo+Q
YNBbj4tsaKPQpVbFJ3JWRhl3tvtEq2EZZQ/X/PZl4OssPNXdwKmeG7jtRSpUAVG+
96KfZdBxa1MLHKE6qBD/wCtv6Tlg3WL1NkLdG/5Fav71U2/qEF+XWK3DoEfFg2H+
TAnHujEbFKwI5FZ/EURirgz5z2cHV6c/Fh8ies93jiI9z3eZTneBp3rKBDho7uDK
gt75mFcRK51ukHCLKNgc3ZppZDwHpTEUIvw/znwqcB3JO8AtfaOLD63HyA4YCgyr
EH+9wWjwgDuNtQP/+sgMMqHg6fThr5RJq9PHyU+GE/oUurfdi0psysb2cj6GVIIu
WNhum5GtC2J33G5j1vWRKilPWzuHQ5UqTkdbOyKzB4Yc9nwpzU8zXuM0r8Odcb/B
k2AWWIca0MecoPovoKPMd06HA1J+O8w8x7tzIrhdt0NXH7BsjcKBr+BLNuguuQ5/
VwE4QpI9/1NVz/kqeQycjA6saC12zvBJWsKwPe0+FtMaISlmXJ67YiGwLXCGcEN8
lVVotGPM6xYLEMJMTgLwObw0T+Dq1V+fL0Zop8w11RnkAAYt09OtEjsC7XJ62siS
OcWZuyZqoPFtFgiFB4nuF2SCe2Y5JVl4Mo4hwrjbrLtAgv/nlYK16OoTktiFN4Px
xzfjwfzB0wWq5oDkVTnbHytvt5QtOJZN0tkT7rCHU9QmDhO+iW/Wn5svmkNw91+i
n8ykaoCWFyivmGVnNhAUAMWx2/kr5TdGFtE1TPhaWRhSB/RVj4go2KjeWuugxje6
WUP8cfrhQLd7NbEDCqsHytl7/SV0mmn20UjMeHr7OiMLJwxAqbN78wI4KsvYMWG8
XBbVG3w99436UvQ161Hf3kWD9U5B/0TK3nQjt096HH8XCUiDF/xCHTuPd+1BZ7yJ
dspHtI/Y+hfvIcY2PAalt5ae7jZTgmN9F7J5nEQG4kmv1Xv/pFxDtRL0t5K/3Ipl
rS38yzggkOke/Ekz9/MHPbB3aKN6AjDo0FfhoEmwj0N/n/xoc/D3072kXYOBtoiR
ILPCe0NuRVYtUWJTuPa6fJp6UTfal5nsgJuLyFufvQbcZAFc1MYEuVSvxtUgjlH4
BVhbDRypAztK9/uyPjSlRAsa+GtmExqWu5b6oYktcm44m0Hiy8chDJkPpr2nDpNR
pGxng1c7DWaw4LEzgmHbSL9lHvGVGbY07dzEGLXEjNbTMCLqQkoEQRSNJt+Udjxv
ug5yJOUg8ZIhaJemkNOsEmh0HMOOOXkLEdGAYNj8xRZVS+xPebsfYinGCK8Lhj1D
aK31cRjDfj7LQBmacrnsVLHoAVrkv27ZcpkfDVO6qRoPL8uEQ5F8msiYRcXq/Jp3
gxIYAF6MR1+ls0Fx5WDjG9xh19MMCcQ+/EXoIpqamA5xM5pVf2vhsyYxCaYmGHrD
zBaQXyMgEzhH/7ynC89pd3mvy7/YDE8u2cO79xD2vLKzyBLkEEfn0wuW6f0/cozM
MxtJh9xMoOXEcC4o7Nepz89Bf5sQvOKyl0lueX2OHJpOaz4nKfQfrIDuhTvZUAoi
Lb7kjv3oSPVJRv13M4tQSWqXE+nkQJwuuiMNwcXYJFxIn9vaxWRGno/29jd1n12A
huZrGYJ8vNdcGpsv2c5ACNbi3Vc3L5+761TuSQ8QDAJu6qTCLz4aOfUtteyMrfrB
ueRormTkY3kp9mCVlruwiEDqgJSxIVj4jwFfFe60RZl9iemj0bDRou6LnDA1Oygt
gWqpZivFtRprp01RletyPp356AAymGWkY4UClFdT/bWOd1ko4VMXDgHrVL43+Sxh
C9MQ9P2U+/hUEBD+pzmrZx3We0OeRJga870wYm5U4g5i2VIXkMG1oSuOVYp9gSIx
KlXuf41wJJUwtGhpzjPvkfQ1ZXX93b1wZt6KIAvLtvIF8+Wgkprf1LyrK+0vUlaP
Ff8o6frDbCCCv1FXvKeeydmM+mP3w5ewEumAXiUbgzVbVodZStlWytKb/PgrRCYA
Xibcp21I/VOcndNXp1XhRcEQ17SIm7M6mcdp7pHLsRSBoNd9rMplIrGsFkVHupPg
xFVstfoTBUCllyCN4irW/AKoQh4EzMkQSiC8JjVdGk8cANk9klajYStxqxKOyKRl
M9O3mdsV56qYUlTHlCfe0xaq9B+x+6kBHPgzfabQ1PgGvMxL9pCa34dUILgvDj0J
QBNMRjMFuy0u2F3cvreA5b3qeAKG94fZOD+BSXDg2nGIQmh6S0zLB/Fs82MmxfaB
yzTbubLgBaRwL8wZaUCJxJH94ovdwEK6n6jM+RSGUnSVC/wP21XwOcbu/kua946y
NFRnvv5sXp1pEMvzcgM+ItbalIT5nGNQmQLTEZpL9YB8mF3kbKppxd8cOLI/kLnd
Q2T7s3GBTolcN/dILaHjEmxUVOx8r6i1zEyLLp2uASFkkkq+X0o6uL1vCtp8+LDj
JkxN5PHPEi8ojO+hO1DtQ5nstCbFnU5iWwO0gWlnDfvUBIIQec+AXWEK8H2NvOcw
q2HocpeqpCQYGjCKGp8UHdyi67g09yeRL6OCgTPuPgAaG8giC0KbpaEqrOv69voP
h2hf+n7QN9pRltOhKyBb4CuMqXBVbzs2ioTBrS2rq7ejMoeLXi+QaE75TGQL305p
R8UWafvqhOMLm4EeL0qvoR0v+Jk77+rUokHz0Y+u7LSgRy1qX0fK8d1ApLe5+0Q1
lCnMI634FhAb+Qkc/NDPxuf8+yOcG0k5FSZQ3wdhKxRRx9k8Rm/D9arjBVj14XPz
V0/Q5vvwUvzk0kyEEVkHpMOmM0O7A8XPmzHaaO+myJuXeS5lbrBc2eDettrCru3X
2bzaz3skri245m1a/RyUgy1fzMM9bOEktStEccOaO3+GT3RmmQRFYwKFfzx5RIfG
WBxN0Ey/JM3CTOxuQrgeZCCUPIQ8l6DzLhL1HMnPWBDyEqLpulNyKFaf3MSdzuon
v0MMLB8cW+JwftyzF8kJ9RdDLvhEc2nVVN1OmFLF06RWTjZE5eoW+j0u2eoPTEq2
n6f5kI7rMVP1vhmerSSayqDeW2Icitsr+mANN2Y89Lfr1onFlTIw1peLlREVKvz0
/WUbgoep2OAwaH8gX1vp6pbRmfChJ0szDdHMI6cVdyKPNXgqi7MaDpAQuOWMB5hV
xs+7WTYa0xYMZPGhygMG3Ki05xvPfS7IWvgY8rwAz7h3zCsjvBnZK0GmU7lYQhPg
tLuI/qcAc9Bnv83wZuO+5MiUg+ckTUcAD6old+dwUcJvUR8yhgYHP3E1nG6ubSB5
Vic/jCsfbip/y1ZleO4/c/lyGviMQrXJ6m15MhYh9GWrT2zqWk02FUxbPxxcD3WL
XuMuEgf+Z6Sxwzf8qQhH6b3zs9IVypZNAt9ovXWSTqymVSu8lAwiVugqJNyfIDU9
BbDUzZS7tZLKkzE8MVODU6IqsYhrJUfP9THZVZgl9RUfW33dvptiT1xAUbFWCvA9
0HQ2ayV4nQoOXFOnMts+G3uJfIVz4kLZIHQhCopRmOY+Gweqx4vzYzPPKqSR2pit
VC/sbVWCdwjKz0wmnkCFyi8BcUQHa072K3fEhQp2QRNJKjUmGSPCA2sF24Kb/j9N
m5dWVOZN66F36JlBPRD5MhbDTOD2Ina/3VX6eecH2HwXKbK2R/R0PEZrQmqbEMga
OUt9DdzszDOK3i43dihW3KKbqAFehjEcxj6cozyorzHNcS1weNyhqMyK1IYl19GI
hSZ9OZroYLY0s6Vae9IwtFPpSf9hmF+odxVy2wx5PG98GP+8eOuGrSxZ8T1xLnFr
lkTgPpHe5qBwXR29NSaFFbpuqh4zVp3lmhWsYQNqadG41iLqG6v37L9vUW8c8zNQ
ivfRuYks60Jh6MFUSmTFxYF0Li3+21ynGrC9BiYLjPLOtakVZvIJDwU4plY8LAyO
OLB39sbfhvsee4/s3bNBTsFMIyXaHuMzBejCxb18LAmLKJOZiJScee7XCS5GtMD8
iKbSfiIopCJThx7mvDxzKUIg67KHF3CVif3Q2U3Huz1TEi2Q+19DHEuLQoVydy2x
Uq9AALd80qf5Wh8BV11Z36f2fqDDTq831wFzw2+uSPmuyW8Y08cTeqH0e18NVaCg
HwOOekhkds9OkFs0DPFHw2nnN99AU+mHRqhLyJsLL+eheh02g7gkoHPN7vxMx/rV
uIXFYqql4PVnIhbnqT/CTWYTqN3/MsPYfjNE1283CkE9GKDqR3NE4B+EtjHCfnqF
yPdhvydkUl2I5I7W2dXCdRNkAxKiY+iob0D+q3YQudZLfN/4bnIEbO5ECsCpVGnV
Rqbz4zQlL+2+ZV/mhTuHO7A0a+9xA/AMprHZ/dvHo5lpzKB5zFcrspIJ7QORRqRW
jNvNvmK6Cj8dtFmLq/Ig3OiSuxiO1f1Ow3zY7nVcrzQwm35ueVyKAfi0v+xJ31Nd
pRv0cRrD/IHZlEmEDCr4cWre6L/moZ6T6FQF8W/MuL8BzugGEtnZ46s2oWmZbz8s
uG8lIu83KSyz/Ska7uq9IuY8b6HiSO5nc8fsdAoYKQ4rvntSHhCBSWFzWb+SNvyG
SyUMYf2TBEi9HuWy/ojEm2ffvkSdP4nlEF+4kOZx4iU2kTjEHEYCyDypqnx9CZy5
ScJP3oyeV+H0IezWoYG2Qty8wJTfHsxRTp8sOPekn4kaUcCCxu47/gu7OdNezn2F
nMxpAKiWl+VXmovvG6uLOL+UAcFrgtCRPR90MlhO4Two5MA74RbiF+Hv5vLXjuBt
knCk389Pf26GtfTxT97g6JyJiNOERVDZ8cSjb7C9egCunxhqJEiYPT9ffr8U2H5o
6JPZ8+lCOf7QtUii44bQ0J4dT3w59rP0Sxn0H3+hCuOFzkXAsa86fNO5b5xw2FrJ
tSEI/o2WX/ISRuem+sWJrCxtS/WqOdkHdz2l5goiS8n5Tkvl24uFyrCry/2oTSLc
4PcrigHORGuXBw32YSz6Tgkc/i22rZHA2P3fpI9fjk3aMiFRiEdg2XWQVT+frTZP
5hr23cJFKf4m40o9Z+vkeYtkqy4QItZU3qpCJ23BEawrQbHvPRpL29jUDKqjV0oh
8gxsUNKXNhH2h7gDgfXzxnhaqYqwTte8dG1Ri4UK6HwOmzF4ZwrxuhjdSDP0rlUM
3QmeVt2utAsiqyar4529tFyo4zwm9JvP1xdcWBYupUH/qNgr+2tuBvQ46V1ufrDI
3IKfPaCUWSyjhf9ANJF2Lfa3r31MAHqpKu1xoODzKiuJhwQMDFWpMm3oyngbnI40
7v6ZZd5NHaVna6yzR118NEK5K6VWkV2XD3xSn9FEaJa07osh0VF3Znrynvx/gLv6
oXIrwUtPX96sBqvrj64Gv2C4bcpPzefTjSWEQ0ZMMtqdmKqxgG1dvH0O5vjsBzUR
2ynQsc/89BWxD3dT/rLl7BmXsMEjBci4RDccucfHaM8IBrxDnGc1qbyxr80NPPuS
qQxfswuZKMO+BW4b80IP22+FFREqQEfawji4bjzi/RPDkgX6OWUkpbmEsiaaDeLR
ItO68LFieK2xgiSdRfPc/cgaD9Egt2EX2XsVKr3qkim/lKyPJCDdg1S17D9Vn2Dm
OtZL8zMAikgLksp00TyKfh3br1SqKsLvtX1dIdqbx1HbX88CLS/JI30grCMHLv2O
28wyLDGpr5GymKfSvDHPFB8VS8pUO/SOI1BaRZxcXLGQScI1xYgHAWquXRC2jpCu
VpY2YqplA5Cxi8aaaF/oeBg/SqXiS+zjjC63FgonyvA/Pv5IEKSUYn7L/hdy6Xrt
+wXdN2+VUFoGNbINLCv2vMmQDws7Z0lxGuXMuXJxvhx2rVeHkq40oEqxMVUTA66l
yLBv+nWxOn1T+ASRoRZWvuRiSomBspcPerYJQNBL+Dq7C4uJ+2DgOUPp4N0eC2Gj
wonrq4G+1tP26JCvn/MbSK8lyl+HKv1HFfdrL/f9rLLNvQvjJXYYJ+VwOao2GI7o
QI1uWYbYveOpWOEtB0+OmHU8MY2kqbrcSqRfZKfXX5QU1a+zdldLl5e2V2zbCclj
dAHKYWWGIEfuZ/l3YOe9fr7ZpBs9m0ZdEe0BHaDq99ZFtiHPSumWH0a4u3t5hT2U
hKclZjIWZBR/M3Lnfd0pM133SbQZhCfqAsQ+UXSyVO/r1Bg3rhhUsrU3QJ8f8Q2T
d94s6DARKdxWVpjazNQad2gGKMG4oOG1SxbVcWSd4J7/fxM1eQC9keMDQ0w34kSC
mgcHkKETeSHjncVkBhVvD8WXKBFhq+Q/wa9XyKVbDTHXfMVSlbNl49/cGyxopTOh
p3NNzPk3ipDv1yINJSLt7bFWe1sNU8S60M99AFQ8b62yVySCHiIhmux2RhESkrCE
PnlCGaxBmCRCWRgyDXe95B5vmGxmUTJjd2A2Ym0RY0aID02VZBzVoiQBgagHTTbE
U31pcR34QTfUY38bg8a3mJKxsDfBStoIgfKOYj7/1I+NiPhWmYdETnNalLdKmFIO
dvLXSaNDWzXSiJfjoelArev6Sbbh+nrmh09wvahZGjiVC48Zew9wDClOmVFycsuk
GSMRE7vlMFiggs5wE44uwo2ThtDiF1y4Wp6AcVY8og1HjfxpjgXNJTn70niDG0zH
MgnCWD+nKEIcJO7QmcszyCXFpN9JoQEw0Sa5TvXIns6DNI21etiS8wi5wT/bQI6p
yjsO7Yim1qAcznIQK9b9ffcYrKZOQE1XdAswRXQ70hKtNRxCqX9S9dgfNfMJJlgK
fHChW46gjOTVC7X20IBiu5DpxCNG+jkOA+OqIrOYk0agpK+YoF8oMwMDyKoZzuhV
KAagZZTK5Aj/2hagNM/a91DnUMTath91/O1C8f/EV8YE/bcvuH3mmQJP4baf+vjZ
ioD3J8PeBsiC/vL85Z2pnq4dofM4IoytrQHdfssSTh34wQxtF8vcSJv6hQcpluaG
AhVRh5OR4YLut3y5Pj8ZU68EfTG8stTLrul0O/RdHQTd0RcCvkIjqWrPgJ+Me5oT
SxoPy3JUQjIWDMeEV8EMNVT3TmWjj4nDGSCSRGgbxMLo48qunrnb2/f4xK8WA3FL
sJtWHwTbpasiF9P9wcu9Cs4GXQ4Exlfb9wzXNBaBxrGRje3zAZHfxZSPwGwWPktb
/sYhD9NuPaYe6qQ/AgpCSkN9Ejj3h9Z8ZaxKpYcbMDvvn+duPRzuUi+i6J0RYaZ3
jo9EGvuWsW0qK/LKVTZtVYEP8mLOBJoNB/4uTlE+UtJxv2UniNVoYspabYF8Xsl8
V2VlvwouC+Nox6HFO4UbGe4GXnL6A5cLX016KtboDNzm046YDMdNq0UTbg2rGKBs
0up9LM2WbztCmBdgLOjaeXmEpetuvDXduGWBdMB5EfZDeobh/KZew7zb1EeTZmZn
93pSf4nQFAI1oLcIZCrkDUpW2pd9zYRTclqtqvqd8XKVaJm5YMPWDI1JTq/ZUuZz
vxbNCPshPEs7CptaBmU2TmO3cYrDkGeLibPguZ/VfGK0llQmFNVdrLb4zar+ziaV
1FHTPFlZKstt1bvJWyB4FwbQUgntkIOcngoch36lyITZj+N9CnyymhL34NR5RnCE
43gZrwyYVRM1VakcYQvVziQPhymYBK2MoCeeidLdyxYPdOfcJFrFhWBQG0vWp6yy
XmZCstq6He/M7UrYtKLdP3bZ9zQBbdgiH7GdEVfzsuL2ACiUJ1cUz7qUZg7llWSv
JyaZRDIT3syVkjSIyt8fLkxbcOSApog900pmAteCziN3eDlgrPm1vCyYQFa9AV7d
3X3xwpeUhei2hLzWirW59+kn2+ZVIMDHKiLyQkwG9wDH1kVHvsZK6GpTS8ODyYgz
iy/OQgIluKk3eSecfQ2VAmJ7XutOZf4OFvHoXd0/+rgycSPhlvthfU//PwuMA17V
3Of8VegMV3fZrH57PzOHaO6BcPbCyw8KkbkMivui+RNgx1a67M2GyeXkvONiM2tZ
wYOXBjHosm3Cfn0PHD649eFUExC7uyUEDY10pQ65peBcJfZ2P8SIkPSGBu3sjeqk
iq8duUlpMsuzjFmaxuTLkS++p0Hy71oe+CEK5zyscsBdVCmaESoRvPysclhqFa+6
P1EQRN4NG0ZwIm2PvQXfAiDqHbuOWmAzqX+97SkB9SxPwjlHvy3J5MNRCPsRXI5f
jI9VmS0K4BN5PwOjyWHIdCnV6XsYvKieD3YLBPVOBe0VYUtptL6mBPbDGtM+soyT
90VE6c0JamKtroNmuhT8xLDrKRuTv0UgoA0BPSaH182McksvAzzJTrBD/Zw1BrPk
7BHtgWMFvB987EELepgpM8mVXjafMrTqnKDfvkfGDZUEGxMCNownCzB4YQkcZt+h
rGA3Rir4nRCLNftdo7jJxHY8DRXW2CCgLo35AttNLWetZwPWiZj4z6y3ZBg+RBKR
6eTzf35ozdU3AoFFb0fYi3f54W9ZwpwEW5uK7ZN35B+G4NsHGpXrj9wms7qLLXK3
t0tYLwRya63uipVBYS/dGd3oFQtbqKEN6oYaHDQC/UEcp1tHHqX/L4RgElmRehDy
ZDj+VfHi4kkfpXi8N4+MJ2w6GqWLSivYjf8oPE0SZmVVF2oyS4X9XD05Yo3amUCJ
+5muU5QfsDVcmF3K6j7HVfPzRs672psm/zQ6gV7h29+Kv9HiJXukZDaqqzP0WVVP
kHM8CgdS6sTO/Le+ozvtCnUK7Ge5rfncE37qMQ+yE2ymSOxw7J15YkWd1APH4DRi
7yUGBs2Nw4BsihHhihoG8jVGkMkrfkT1ZQjzHTtf5OTzJoApZCZ9UJG+KvMVFlH8
qGQ1ufBJZO+YJxL1FsjQnHnC1P9H3vVto6Y80h3oh3py8y7W+S7bKfTSR+Xt8gNo
e0PDMtLwTIoJMNGUtMfsPigyi8yrlhTgNK6vwHS7GoNZIV6xY6q99DhN+DatXmvw
/VHErHJFM79pY80yqgdOp+2/XUfXOHozehllsjWUJWiK8k8KJ9OBOYXm6qzRJ7bj
BEaSqZ9sfZI0HImPngt/TTz8pEKqUFEsTXJzC9vK8s58+5jB/rGcc1XJC0TWxMbO
Bsg8j5Df8KiDMf5+a0E2VkWzzmgjJPT0ubbUzEubE7VZe9hE8teZyC19RCggV7U0
jx8fom5NPWI0bjK4rvP9wtwG8GmNCN7wAE88L9mT1JGVWYdo0sYrW1Ke9+7Hj008
2/330JVz1QJd/iiRpQrdoOPZP4TC/69ADiViEelWtXG/6Ca/2/L5MUDUv8E6eDbV
SBHePV58+p1/8XVM4wtMV+A8pM9uEDHFa1DE9BW1uSBh9EIzFxoh67Q73lOlC2kQ
b/BdxfGTmL8OWjJzMLLbBQmdTE3z48tw+yekUBRP+gjNcarQY9/JdyaVSeMVOx8I
m712MozGx65pmD2iPbzPcPDHQV3rq529N7P9gUgjwGJsy9q/2MUMTOpoNT7ACfZf
K4KujrcGAJ6BswsQO7I45DpwWCkpxW1yI1gKwcjjq7FIQKsedwnHQFC05ZVgV5WR
RK3YDKzK5ElNQeMNylxDuZC5M9bYL9LecEjC4j/vEB3kA7zjy1Wt9nk6vCtV4xsg
5dHIuj+cawYqfEZmB/EiUgM/GiM+KGpNzKd+kuLhVizYHlEAhEqn6hrFkzLg8DSK
tHIv6IHNIwljRNTUuoYFfQ==
`protect end_protected
