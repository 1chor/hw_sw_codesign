-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
jYM89tSgpEtjiZQV3aPgt34/WxYoc0TJEImSOinsq5MjTvQNE5HpMq5Kqn5sFNuahdkw/GxlzRSl
Af89SsarvXM5Sr1dJtPnfBdxhQ3GdTjzkBdLO54KziICJ4QxMvdo9pAxkumc2+gKd2tpuK+XxDQ5
jPas5DRSMwng4kamoebPT2Z5OnvOzq2KnaeuqsY9UjlbfmC85lcX76+i4LKnbp412+gwoL3exhCz
kSuH2plcAkxWipM19kz/Elh0PBpDC9X2l6V5kBdyXF0B9hqF1gaW9jf89bdJGlibjov9bmYYQ7GS
3uAz1gCXeH9RLfDc3jdfg2haIGE+ouZJ/FOOZw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14240)
`protect data_block
uGP8m6Idg6wL6T/JfQ6N31kCiP5aJUeiqPIlyTLBK4bZDUScziC7WRfDAgKSlvRjUCwaZ2BN5cLJ
SFaF1vrgP2MNbG47CbmqHA2Vk4XCiWoMsaAWUn/x/Vj0W3DBCQBgNV/6LsxhNFfpV50OUQ4CLBc9
R816EYNbsU1cOpyC6bJ09B3lIPDzEI2D9IMwBMUMNbVAj0XfmLK1nIRRy9TU9wcbKuTCvLC9da2s
nZLOJwPvG2mBhEGQy3QBcWb031IafJp5Xw1xbkHOjEi6oOYNkFkxYh3I01SUsmsYx9AIn15H1Ku5
am52qhMQmZQOhCOcAcWeouAKF4Key+BfRO/fosqh/qCkwANVlgUBELId9Eu5/E6iW3ct+t4eRxkx
8/qfJpsnO+zp3bFRxrc17VmmisvbmpSaeVQw3PDtm9ppTKNrDKIEpkdypH0wcJCTwtwXwyze/Rmx
SxaTIN97n8xPR1x1kRdKJwdPD5HcgZO/Cb5T7IjaKHOz8Q7iv78W48gaA7M/Cb1LNAapUfMjzpl1
IeneWYHvBg1N8BL4dAGnQiuNp4tvF9ugEZvwormKA2qcoounfRw1LIoQMShL5Sa82RwS7iqJiaMe
JvKE5pEaWAz0yvE0r47VsE+vjeOon5xJSZvdPIJDiJYjG2gUDcqUHc0GHGWyAcEGKxeXxoTwE0iV
cfPdZpA5BOSeFJRqM6QUKeIaus5angvMU4LFWT3hv+lpfBkUY7TpG1inUfLu+0Kqb77bm0gFj5+n
P+0ZZF50ZFcv96i0mtfiCk58D861z6dDvIgmtgtVVmDJz4rReNSQjVsa0X1vPZQvtulWZjV+oiIu
8wb8klKC/2ZvOZc8TQWo2pjQXUI7C+6DWgnfCoH8tlxfD0ektdlLN4DdLxKdhIRq2dGgAXgq3K+9
BwGGxQt10RzG/w/OVmpgLybDAAzFZru+nhJfy80ZhUy3LmGZfCqZnOCxYDSfk3MQavfDwugibqRD
6XKcQ98aM27htLsefmIDYLPZ3smt8hCe1d9o0OG2/Zh+++Nu8ISSo/tXvalSFvPwaUgXdYugXXfo
MdxCHCjkHvyVLuVE4kcM3IfIbVUQ6SEftEIZiQh6ulNOXl3HpLdIfcZrKt2Q6Qm33UmL52qhEKmF
pV+PyUaYwkYsKn7YU0THGlkGidUeO/HRdqNJPpg7juBDuMPC++aWcYLDLAsS8DEjSMPECBHNQyD/
aIkRYxEM0nn67pScFQ09KODh//r5kwbzXoBDgGXlq39Me1qkHsIYrUJBp5NZSK2amKw7JpXPSM2i
oQ4tTGPG59enFmg8vS+UyvYLhmS1AQSNUZ+P5vOLmsYdlJfw/J9o2XPeScWW9/0KLsFxY47QPMi/
W2okhULhKJRV7I3gxxfGZJHKFDGTzY0KxYOOzyD2t5cAdG44mNrJ0rwQdtsBLMXK42wJv8R4nXo9
ex3JO3/zz0wqkOg7x7694FKLN+UC1Egbc94FynjgmGwwy7WXl61915Ya1+nQCehu35q8An7zou3x
7P9uc0YLnx4VTpVV3GYBKyEGAREbDPHMMWyI5qtTw0NZa1s8yEeGp8srPUkbXXOr+BmWIKYr/eLu
3jNhJS2MBfuXJOaDYT1EImq1YHQRZefvfetktP6UDihBd51fZa8cnCaZAM3i21e2d1N6bkFdRxhu
RVl84MsY9Afrv/4Gx5NqOLHv+zyBrjItjl2xe4Hm26d6SoL9KEeTjCgfHy1qZ00tT8qkYRLKMcDb
H1tKmctNwHT3Rb72oXQ/SzkE0gsw0qGSZq3vhyMej8EWQn3JQflZll0bonDzYUp1EEpYkFsVayDr
X7vZWueLUDCydqMWXYk2CdMJFr6XKCUfU4AQKBNoor7s3BkrEg/936bbX7CUHuftSs0lGf4yCMLh
yYSSdOcTbYA0WKqsr0jf9rFosfOsRBVPhGXOL/AJ5hIOjdEfNB3PUm1DiFQb/gq9BGOcbYAbXJND
9mnDCz07XBa/Ph2xr60f9qBv2jxvCSHYntheVBqShkoQ2Jq717WSVynfYIfUe1RinTni1Zerf4Q5
Dlqh3LicO7COU5AqeUeqciDcOlIM+FmyaBiU3Yg5AgY+zGYwy3XOdYAb+/zPLqjqRtFRUdSMod34
Y2juiaJL+gUUJgHhTrV6FDLuW7iesMRl9JQWchfMVFwxjn85tg7o45SCegmJlIyOeC45CpVnvxjd
4MtK9otU4PjPGa8wsT58IFli9KyXKcvJhOCyqUIlTeTw4SjPHDl9+C4KJ5S6t95muhaf2LhjSgY+
21xLaYtb1PEpG+LManukKnD1vJ9ZJDOeKPQ5UsL7GOA4T/BPoINiWJUMc7oVcaWgBvJSfeP1i3+r
I7+E/s1WeYPVaNjY+BvzQm+vmL0TRSMuDtRJ045UQeJOVDbNEvImc/6nkDbTy/mAIQxz5wNvM081
Ldwzbzxm+eLxJ4EwWXLTnlDS0Jsr26KLJ+5DIl/WZVxFgSqWsxmHPHZRAHfnTLsC5CJHnssRXBw9
Jx08x9VyRMH5YqdroERqrLGELdU2rdaAPCGq+vehZotNMu3f0vCfhYm+vPjlcERJtSp/icKfsWAs
nXbFeLdDOJJiGCyJnmwhIXN2fS4NKR/9f6cWjQHX4s2oKsQcxPtAa7OysOEiWLXjSwDDbKGIRy/A
0uyCnbETxD7iulNA0xzL3kWU9kdN3IgQQFBGHj6K7ShpR1v8R/Bwg6IA+p+xki2V05bl5uspe5xA
31Srps1UzVqBZu+uiukUzNr0m2mn2ehgr7DHGdRlR7h+qKNf53+evjtkUwzqWO26mZzTEriCZKEk
YBkLE3XHqmEsm5IcDZpw01rpncI8PhYUnyh6vqDIcgJ8vDaW5Gw6DToT8BdxLvSNjJEehRRSYOaR
hYEPcb1elbXy5zRw8lgBmoG3mGmPHrWsEJ2SKLQvNYWXjN6zJUbRfjUwmqdv8cO9czUASx5wmq3j
6c6HK7Mo9fJgLsLmDvLz/HjUjYFglqhkdm6URjCpqZZDh8YSgptSZNyoDkh2ifgGksiuQmkmbYkn
UfHYxbPfS8/1tcbWs1RMuG0EnoWC6014G0bKxlpV3xY4EmLnkELPKHxySA0OebK8qw/twWeWqX/s
8LWmOU7ZupOIgeaGHbiGkFC4Iqafl8TMHRtSBAZNfiz7KzQIX8lEJkrNikqREGEhsbVKbqUCzOpj
nb/h+cPwLfxhuuEfyfBNaOZaqGHrI5NSIATMYK5wH518oVCbu6t6086bXeZ5qVEJ7R7zyECebzHX
UpxQJ9FYQNXB4P/ptSpfdxXQzb1C2mqy8OMYxUBOPcfVeDN0e/GYxcrY4TTFrStXZpu1Qy/FmLZ4
ZSAYoPgOFjEzb9SYTrinoGV+scjpGrqIMqrzzHeMHwd95b1rfCvU38pt2n0+ghbQLhYqB8Hj4NF0
vLLeHxKq/t5sBOOt9AHDIlyuw3o+d6Zm+Hk92QhjPehMCjr+xkTWidrLV2O2sMJ2N54z9W767wxJ
vZ54h+FEjYmCvJPvsbiMJvtfAvea/abmpZcuTAelzzAHZk1ExYSd/w6rsRsceeH6KJkZadvwJcSJ
h6taB8qe+SuC4t0UNZS+8O2WFzouwMDZSUU5kBbZEOJN0tVRrzHKGExjQVe3Y0g1ySnHmXhJmCiO
tlBrp+AIe5JE41MCXwxmpBimFMDq/oyx9AU/Q2JvDySwcHGZPUUP66zM6psbg6TwiSkxD4JjEeH7
SuDJ8dFhhEsfWPZW7vq8EkzolpFnTfUg6LSoH8zKjJ2/5sepQqrogRHZ24lhLaGiJrpp4vq+9nV3
K3SBTSsak9ECOX54TV9/GenCU0w2ORqGhLMxBeOVDovgcnojb66vKH268CkxttV0ePqOI97+HCp/
/qVVqqlSHFA56KKY1xlOoSRdPW5cXd3O6bcure/2qSHD3LkzXMJ0bpMl61kUDIEf5kX1nTMlVHOi
pyHQ6Z1Qmt7nnDgtXvpJ3dCkDB8Li3U9TPaXX3pxWPNogfOSmUk2VL7YjnqJTDFJQVLYoBnfRE0J
XLSW1LDgZwfacjK1HmCOuPziQJR8Rdaua4TPL0ENk+V5Dq+JvKMpTkm5U98lRjlm0zfTmyk/F/U4
lwK4NjIsOTPKDT7LVpYPjcVD8z3gkEyWGa2eSRAvPQMyYGuQxQ+X1iVlTzKgXUK8yUY4qzBchWGn
u1gI4pfwJwgn2tNKi45a0X6iHaRKo21PH8G01HU31GWL9KXsMTaB6Fq11wrPjRAgcMd434mO2vZm
ABFRYDWgXnpvB4Cf8lVJFTaFHUWh5zUtRBaVZehBIl74A1L31H1sITonSwwBLKffkzUkZIR57zmZ
d74950XGUEmAl9jNvPNESdO5KV9Y54GRpInqmPszcUBQNX+Cib1YC8FshSltJiqIvg4vkG57COZX
U9j7knSC3DpMlsJXXF3FdGj1MNVgzI+x0fWdwV0SRJu8bdjTldtjMtfcoWsKIFIYuSJ/yF8J2cM5
h/Y96+Es0bFA3a0w8WhCZ9VfeVsW1Fg7cB3dQUOp1vwcIn4NAr9JT2O9MFbyxDeP2HA+d0CCXR1I
c8rhlT1AKeAjPDIFsgrjvTb48txErTBOMiUhEyG06bTq1j6R+7Ju9KdJdVwkmsDkObAT0XT2RxlN
u5c1waxp8o2Zy0R9EGIqxiPm+J2oMQRd9Wc/UaSTBHNNYGiyzK26bEeZp3jcAtUNCIWj2Xlw6shT
QytXrtIWAeNnG+zCaC7hqyD1LK+p499AVRnoRWoawXDIcHcKXZkh5vq0hG0cjaZl5NTM7SncPB0Y
h0qUXfCzWWik61nMnVL22RkchdswKAyTkveySh+4r9w9qTE69ZFY9Zk4aP28tgL5NpuDGtbSgJoc
XNBzCnxlQKlYatQAnUaQpdOWF8fEOWkDgXZ33mCHHjELIYdEbmRwpPZeTzxU4TLsIj/BCGCBm9B4
xnNLgHEzUgiu+fYxtXfg3uOuMTXdScKF14spD6QgBiTmVviDPNH7rrLIVC+aM/Ql0LyWYpswf/BE
z3i2YWrliuHc70PxKbI+91WpkqbvmKoNpBvHoIx+Bm48uDZ9Kr9hUZedln312PmINQFULh2PXDob
YkKGxVrOqEvStXZGa0hFey8v1wGtNMFB5Nu8O8mINfkqFCHjG9Sdm1gn/IPhP5Es+pvQhdpreUH2
XIPPfNoXunp6skbo2932kJyk8zoF7lMEtIQeMYny63IVLM7spbMVVz2OS+p8vvUuxfGQFkFMiFxk
ZoPWjoKHsr21zbm3sTMbvm7BMLtWgSKjUj4+8z/MGKZhoNtQ2wrHBAxo43tf31G9Zk4v64On4ueS
Z1a9azfgx7obB7oPHuU9cFqb1J8UjFsHHn7Yk5bQn0OA4tqnHx1rvUSvFUgT+rdoqGZnfJvg5UYN
oqxCW3JYCPms/d7smiTqdtA9G+JZg/ve/4QGrM9S/IZD0cKYTcHi6bVK9uC8qnZOXdjuNCI9wQz/
8c/vullflp63JqkZAodjnQRi66AZktJcpeD1PoXB3KM4WYFyHFb0ild+2KvgbakDZopnn7d4Nlmc
tumkgTDfexajuLO0QamadeYemqD+lVWj10rKCTRsuCodNGMz2MhlH5PEiZzOLnFCMREAFzoTioXZ
IMKo/1yNQxGu8DJD/VBnruAxBQTFEduoRKCFFfbh6BwZ3VaRq9I1GJ9DhNMFb+j8BkRzgQWS3oUl
lsvZitmEiNyLr1M8I8jJzeS2HM8YXkxzmlE91dO0a9An7TfWuI7YptUFjUrcGln4WYKvJ03x3akO
4mYfmZ5kOkf75yP7lC8n4lafrZLcFawgjiD9fSnCM2Qczw+IDwqYP9tNONO6aBODPVl5WCyI5MwF
wA3ARt7Z+vV1x2eiHFBk4YIxFTzsdWQuJwyy10zLkfUIKBueAtoFWwAMqJli4Cx1bkCQugtj6oKP
JO1B9wx4dG3062ggk3DWyTJxBPFhb4E/lxjrLh9rHaq0xsusdQ1BXFFh8RxpuK+PmTJGPGOX28Ag
eFiBLR3sjxlDgLQonSV72ywTWbyPIYiXGH6v+j3IvmIFKict7i7gLYr/Vz1Fkte3Rfgff4RGU0Du
rQEG0XnSk6GcMOn9CzJe+BWuxC00oTwpOcbWr2EeKjAPooIvfzWkZYvB0ZTXmapn3uGejHK9yrj3
cuQ3/cj/0BzjzLmbjlBl9uZE24eGvOsqA3xr741wSZjN+u7CKfzE9wuQSmm0jYkfKLjf9IAA6zAZ
jAqNv7vLDHT7ypJ+0ITxEa3sqdbOR8oTuTSbxLS9u8ZnwdFwwVecKxvmuxEMv7tGyyHDaEGBPMkF
HmYcAlJaqkL7nqLQPbkCdBJRt3Ow4+Kcrx60v4LG+j/0/AF03BBMNyGONloKn5p/4u1CskTJAnTv
4XV9RTXkW8cLizvcuv0/0G/nljy4EHe6gUvvM4tx6DCnc4cuDYAshn50E2pwc1YKQv5i3mA/P7R1
Zp/TNtlH2yoeDCextqGGQipz1xCcxYsAnymBS9XlkBbaeHDFWSyXWFmz4qaAOMoPj0TrmvJQVkO9
m2v3BesgfRPPf+Pulj87Y2hOZuxnRUTQLHjCgDsBl79sEEmF3PhpgKDjudsiPFd44huLjDicsZ8t
N1Vj0Y++Pc8s7ysazCQnST+zccGFEKV0g0/FLu8G+MBtEsBnTWl1BVXU2AAjCg9WQAaL4+unsa7Z
8QObn8ehsy6xUZt1AdywN+H3uOX11SOargV1AzOqbqqayY55iE9zZSFmX1zjAHdYxIWAL1kaquRl
ZHMEqL2SqteM9yUDbDcQsBhnRYR6Z79Y+pGwh6zmTlAAbusYaaW6f3SpG+UfrFkcLQz+3Yr2cEnf
OaVEOggIv7rzYI4YnTSg6cS1GIN0doK2SGk5xh8q894zY1wVGCyTW+yPESSP48QCX7yYDYiNHKdV
F7gBG8KGyftQA7Gk2GD0pJX6zcuwooVqC0vSzcWPhEf26zUyf5Ais9xr3cdz/tRO37zV+ePLWYio
6JU218vaECN71HgmOjsbfEsggSp1i2Ax5JYGRuiZRqYd1zQsUXWihEZoVHhMCdLCKkAtsfWLXNDx
KO8wFEo86zCnKvCCEYxbkanfeD6vtWPmx034mCdmSoxtOR7pma5P8EL5RlRT53bqwaLGausgbDGA
mGXpxCGqW04oqHE7j1foOcdU+T7kiY05Sur2MOH1a3MBxpzcx2g6IWp9ZBRBjKBceBMGjZ2Cc0ph
i+EffCWNSWA6MLcpBwDh+1azSR4P0CsMOJyMaRcw6WES2LLmcm9C/pHJ6eAe9+oREP7y9K7426tC
RN7u4g3sLXU6xYhEpn1iumckKxrhAGUpsMVyT1f1tQqMJRlkeC329G5q0mkuLjxkQ5/v4VXPiB/r
PLmSKtIDq111hJo/JygkjBvCJczHOsIdnsSMDwVoR3mpAR9fdupV8I1QOiJlveR6xLeGj0Kxj+4I
hirQTjB/INbiEy/UxdpMBLVOnaMexj8pKjPWB9zy7fKfShg5TKFg+WhMoCSOBbBjc5480voDvcfE
vGAqzLVOfPZYyjtwsiTFPnZaAsqmb2D2wAa2nDIQjD327aEAdCYaq8iTAW2nYL3wyQblV43ixl2r
48O1j55w5fRRHBjZG2zgo7l6G8e2t1gcfUBL1Dn4+QDdOqi4QkcjQ5KNiBGX5HPK8ZGQiJ1K5mPn
I7ZigSIL9o7+7s+tPpev7EyOuq/AJTy0fZWh/uE4HY30EfHrsBzaFknGLaX7v/mfxdwW/E4SaTuT
UTZe8rkLUuRhcu6xk5xY49yz7pZywNtjKzak32ooBc81m9zMp2BT1Td7Ne83PJiWkvLXvo9oc1rp
sloQiTl7q2/L3UBmOCk19h65NceFk0oYPEeEgIapJbBdF0PuI2mhahlz4P2YBtaAaMQ4e4jDPdKk
RHbuKGv61umIJAsTwDK5HisMQnU1rhqSHPjbbZT92klN28s7QiLSabsz/37tn/AK1ZwBFFCh7sce
ajPh0MOmUpJTbRwh+TshLJ0VMuWwS6D23Kw3SX+OSqW+s61q9pzGBl5nCU16m5nZXh48El2rC+YO
WO2zZsyIO4M4GDEjPp2+Gc8mw+t58ey9AhtiUexcxrVsdv+HrCSy3ygE07ZNbXEzDdLZSCSctuWB
fRpSxnX3XEYp9i7fTDGZwZeZvwIRVrvsbXCLlaSlAlWKYy/LkcKDGshC3xvOxuxKEXfR+XSIKb9Z
5BIwbEV4uZ4niinEEPnlN7mJ3v6bUSxGGmbaNnxE1C7C0zqzsMKiZbw++DLofxUnzGHA/EHsfYoH
/KtTSq1udkg/sjAo6m70xiTrjFRjmh41Xkls+CnAOSnWec1ysTdWeVwTnm8lwhdj/6VB9STkdCjE
XEfio/FSEbycGOGRhGnvLGSTEQJ4oSKpn+TwzPCDCh0xYs56n/ncgYVSdP3X9Wyn/ZeJHl7sAsSF
tbD9dSmwBiQmHIi8erPcvGBFP+mcBV8/Cyc0juUg+wAY77O6IKH1QCNx6ecm0L6HFQsT2JKOmrl9
pYAwwuzEL5GDvVtQwKKZ3IbWkcLLmKe9b6RnNpilVa4hjxtMB0e8HVsGuS16JVZ2sBeaGJ+9RQ+r
TUXjpYcnyDe0WPC+mGmsz2AC1xfJTdwSfpchVs+WKVcncvRP07erb5KyfCDulOIQJ3/2w1l2EvBT
HwjCfSgna/6U8Bw8Prwihkma9jHsIkb0nYfcq1WDGFhcdSg/qQSKvcRoOFXFF0R1Z4p5z2txO0mU
3mgjjzRJzekANDgw4PmEFk9LbDHNF5RnmHzcfKn6gpqZyjutA3QekpCiTCHh9Gly6MB2UNSsYZfT
KTJQraSiTHl+5u51WQE45MTD7UbQkjeUhLg3epXN+ohS1UXpNQbUsCQ39nj+YBxjKmaGr7r8qrht
U3VvuRC6+CNjV4kWaNHqGonCqK6kAiHoemjkamCYvkwb0NbY7W+Pcw4ZJrhGHSia8dEWAkR71JS8
Qxmxh9X+yIYXSBe3d9mTkgsgsqxpyLzavd7t6emCHJn3KRY2tqcTqurFoeOuMCchtcQDvqfkuzld
1hwz0UYffQ5G72qgYdnG29CP29OLquncaWMYshCyX2TsQRqJPRj9xaT6CIEoDZxXIShhWj9AZ+O/
vqsF8P7QOs622lTTVYGzfE8Un/MMcKlxXURX6GyzOqbXPiO5EeKQxNPybpb3n8Mx+rFed1/aBlRj
kOgc1Tv+CB8oOdalu2ekalXOXPxtnxVNueT/m5FuZLAghrlCQTeUM0DtnpccCd3lxRKqPzBBIJwB
9BhVYWk9JSr3ynxvjGBntj/BB8Fj5br4YHpl4YjlDD74KuAcfmJcDjDJ8Pic78QUNbHn/gJL9gJ2
GruBm6dwi2fiMzjyRVaF2vmur92/hSxnRic3dVJy4AELpgIPkpEDSfWh5qqkcHhcOBEtIYaSqYvt
IFlt9peDTbu+A1UqOClm9LgNAgjitTQHCtfI9CRwe7iBA5UMaMF+skrqMPbSnx3l6/mBD6IyNWB8
mLZBY1txrNxDd7T4TZIDu5KMVjpA5wkwsl28TQ5eGAipacAgXtX1bZ/H1U8Hp0X0biyX3ya+QXYW
jEwoDkMiZQyXFmOizcbIrq/DGv6k0pihuPmtt//yPFoXDyRJj6+S1IDcVTCC+mwA+G3Fg4+lHbU+
6DsiOISl1ydXEnJjAgvk0t2xAynvtqBLmN4EDXsTRjKdFM5dyij8cfQzdmwzifProy9xKU7H2ELu
34JPrfDioAK1/V/Sg3z/pfXTXT7ynI2twxciIFgOjmLeNRJ2YHJDbzmj4d3D9jdhsj5CNkkav6kP
m+T4USZGrjg1bLsgUHCZDqnJajU1VWH4Hyga5WiBfvUfacaWKmc+ZTq8CT9ZJKQ4Zolnp0+DDxwb
6ZDsx5dEW38Wo5Z1b5EFtLa8I9sme4/gsmxZEjhLupbWhA4e0Nv+JKyn4BgCpzWgkIVFFBtWgK6+
xNNnDb+TnqT6qMWp7TRFMdik+ch5/2YkMW94sPpuMQ93biAyr/J55tqV+zXCiUC+l0d7wn1m5uWE
ItYkfH8s90MMOto8gcQiJnzzv+gK/yi5WK6OaCUaZf1YN58KnkGaVJuykXtF5A8g7UCKjgS/Gq2+
zvotDUOc0A+OhxdooFEPQTsmv0XC1YgZiMBrMIDQBhzVvv1AudDi79pgdES+SJlmxBDAlAUYxZaU
XID1uNlDH6p6hme4ZKJ9HrF8s2wVRUT+hTOXkJ7xLz1jfqnWs8xeXmuoj5+zCY6KYEWtCcm7YQrq
vX2oryMacvCwsxdTBDPpjTbHY0XLmN+7JYFl2iOrPQngsx2XvaFDnSBKPAmaQUyTgLSkw3qhkT+H
AcY8uYVM32gdisqrpEMLWPtOatW//9K4EwuwVnEJU+H3z4LdOQlor6xMbOxIWNseZku86ZcF0sOe
yVQSA3V96WISDl7K1l9v4kCIYc8BwV2kVJsW4J1TyJQBYKEKr4P4wda8gyR66mAKdbye21/Hkelw
j0pGiC5u5Dtesxk4+gLzYLKL7S+kdbViAvLZxMEUgttKdBiuSwHAGOHMqVpYFrdObLtSMbOyj6Lj
9QCyj3J1Nnjgs8nWqZV0jRwGek1JqXsa1UmaIX2r8akxr0sRuWZwl7KnWsmOjkW7eDk6FT/cx6l4
RSlOhyo6fnfRjxb0EW1jA2JaP+Rj4HudPCu4XJadUx5UWGM40mWAXimaZAuHVYeYVScGtxQSCeei
lPoyvO0Ivd3fCNnLYpQADxw9MGVV3D1W4xht0I+NXgrEacEXOU/ZNtTqR3/GuCb/8nAa6iYW/+3r
1rU1hTQuz2MVt3s9/4bFydAgESNn1KjD5RM/DB6FfcsbPvDVZ6TkRfmImdi8mdc7OdBBvvXgnxeF
N9Xo6hB+Q36yQ1JlLfatoGoQfJoUdBEZanVvGnx1Ew0Dj9101KG5vCrFWLn0lDvznaO7qkwTECi7
1nhop52HvMMlwfvc9yLpC84KEiCRi0YGCGGcigGvswVaM8gCrjVRe88TzuWKAbUVpE1btt1JLGwT
HNCCtQAO8xzj3qY/MYDsJSEK6s18Sm6yBhr/WyP/CUcBccwUywM9rwxo6gxPWNpNOD/apucn7GF2
YSWJczIM3NVzXaSXicAvR6EP2zP0gDI7QIgeEMpwqxx1rPYms7BsewPjB08GUF6X+zTRnt5w4Xsu
/xPYU/TyCY16+cZg/X6zPkNqyMjafscQIfFmtJXnmgaz3CHcrSpZikmqDlHNFgQ+PEPxVPvFhn5v
ngc80tJPudiWr/kWrh6oKw+GO8h3r/5L728vS75qENF8cYqTW0IcihVsnK1RP2HJLWiGxIdbS8EH
GK/7NReo+qrjA8a0ng7P+VbUGD4AEWbQdab6u+Ny5xLMaLGB4jKYouxtOuqRfhwQK5KWHNeUOYRV
TiKQFyuZlZY+qSm3BHptNI7Zdxs2MlZZRHYhDayS/9ZpI9Psw81S0UkrjS+hSX72giaFDxvZGH0W
cuzGc/hhxxUOY5qkKrRg1qgUNd8jhZOwL7oj5K9nonoSXQm1Eqs4XciMwe+z1HwbSK/vlkNLcAdl
rJvDJOd9ptTl3Li+nyXWadWkg8/edCFXsMzDIBRl2tMdvjeZ9nASN/5nkd86OGmwTXqSpZmVtV4V
8/v5at33nJ4yJRZO/LFVc//ffn58e3+gD+FXf8PYN2dJQ9YG9mc4H7mSoqgcpvExVLsP6vEtWNjx
9UxAXbV+t0YBhVhA7f1hCC4gYWC4SWzVjRtxor/EFqYl0JbiOjJzxsDzqu3gkTvaPFgO0jnU5mZw
5117D5DyHKsfWKlW3asVt2hiiDfn4o5+a5tXMA+C05sJlUGoJn+t9xvgeYeV8T5V7vvGWGlwG/Pi
C5mjzI4HN4peuCnuZtLVyY3atUvR+n4W8cfDEiK3InhoCrfMp0NHCXTAJASPQdW1PvE98jnWGV4p
+BfYpHFaAK330Rq/U6McbYw61MjtJTQAhAzxYZXFCnh0FdoosFeHq1uxOZA/AcZ8dHHxliecSBJ6
TDR3MxeBScR3Gmcq7/qnN7AvVe+G6x/+ynkAAap62tswZV88QXWPsKoUN1csBsAPudzEPUUUiNJ6
/FTCAqDu4u+wH/9HpJ+N9/bXhULz92xpSc3OhyjtqgdKfCRKrogjn2VaeHvIBHY2c0Cmgdh7rO9e
r6xYVbBdWMW64rukW7QhmAZ1ObpHSlzTZbtQcr8eD64j5pAr0d3yvGbRTHgQJcEVktjwB3FNuyWo
t/UgSYwcZi1KaDWFyBCqL8foMIEHNv+m7mFBDeM3BqDmVkCVzwNi7CBGg8e8tV2X2g6yqwUCfILJ
u6wvLXIGYSf6F91ru/chdzlHSUXB/cf9/B2bSGIFRACi+z4izgTOtXl70/MWLFNz7+XeVrRAJn8B
7QakLUWMDolOVxozZLqMR0gZWpULOWznRGMVj/kpU4oHBoFps4dQg59sOQqZ260vPX9VyHMzIXwE
K3+rrCGOhX7+i+52LDd1Ef4o3JRiiPQjcvQVTBSX/9xKBoMaIsQw1oxbyTIbiIImJRT65t9YXSiV
L5M4k6J0QeS+PC/q+e9wqmBJGPZOodxd6hfmOd1Xbt/r9OMM7r2t0Hg1p+LkOj63PYrzh6Lpwkrl
nE8qPrIuOcgQdgP4nbvDDcv9EL4r9NND3yNk6ps3MP2aA7UUDcppaBSiDRN+C6vPFCB9tP8KVB4o
sbwyv68HXnfBZXGEvzZyi2sToP45+30Qgy6RNv1FUFr1zXvIOYRnFFv85MOxpkdLlF3oWgbSHR7W
OJIOOJ5sYbaxPLxbTI4v8zd5SaMrkBqC2+LS7QyQyR9wdU+us0LsYOHHjSFK27O6F8jxFfchjiY1
Axqmo3AWetQ3f0Om1QFZItA5JqXwFSossQaxLNR3vLPjxj0qXtOJgD5hSG9j8rrTyHIX7HTnxANI
9pKtkvN5Ux5pWbaPpkQj6Epwv0+CWYiMg8fOvJlYWdntNULuw8+1cz24gW86S6lynr4BFdRAcKlE
nVSXzdsSbTp1HqWdSt/VkLSFzayleGxVYK0g7ZJPEYpPngLdf3Jnib5u9i8EFlKRFsCvEd8MobRx
mgmsV90V4GO0Y+PZx2j0FzJSVYVC0/UjTnxySj+GEeuzmp6DdyuIRpDV+/BPNGfKIZ9ubd0rJy6b
gApr7YMmgrI4ZyIaFS8ckftYrPrP4HlOuCahEdDk2jjwr/tL94OuFViUAVRB70Id4U4/iEwRDk0B
CLbMYRYbpPVJCsHRFs29xlzZth2/RIECWzIO9gJY8ufGhvM0drnRFBlW1DUuTjwnwMdnUqcHPsPP
dmTHzzMTf1SpuSL0nVzU/hWf/emKiosSj5/aBEjcuo8FIS4RPTzytBFNX/SyjM2D1qhRApMNeHT2
ok0kMvYLEiHqFKc08LyfK/K1SdWJ8c/6sz2VUakfZsUEuzTxfaX7z0scaAJas4Vls+1E0rcDrZLu
lj0o1zuqqXlpI6eAUlFsx3A7R3CGl+ijYIE0HBeDNVoBB50oO2wEXhkECSvQnr5THt+0GUce8J4T
+4T7EsF8sWPGjc+a7hB5VQqv/+ppfJ3AYberyYrzF9B5IGIhd9XUMwy9M/hxX1j12DShPavcZdLU
VNvWrJASTHI/ilkznObYxY7Yb50s4RnqNDGT+XGwQ8ApC+fb8k2od2nHrIYQOpNlQR8Le5+JrWaN
+zPYUL2U3e6i1WISozPO53zLIK4oZAfub4V/bv6RTBkR6gWoYD9XCMuUYI0YUcg4aKgXo+pO2MzE
66nlC7BS3qmObVJUFRCn21kraPaNa/cohhYSfJyrtaMD/VfouWFkfEX2n4U1Yxg8ZoWu8tsGt0X5
K0jTVsP16Dhy8A0HVPJTFBZvzH9IRQebuuaZLgiyz9OzmJkavC5msO3a94NQUOpNmgEPGjDRcTEF
Rqk/zHd27zxdLTlWaY01z7Wj7tbnyZyEluHbWy+I4QFFveXbWSzDXqtT2hBIqEfwnALX7TlHEaZY
if0y/BhY/K0nSronFtzNFXfGvI8+JZgmTBotmvRXMZ/Q2GyVrviCGueDAl9LGueYeiHVap1KkeuH
1GWvnNnwaDhricpU/JBh37ZwXpn+gx1sAbfvHhqYR3F/7Q/7mm/v1IqoUY7SQEFl5+mIxTDNLjHv
+pJ/nQcts7/mKIt798AEObJJ1wUo2fWUM1X68Lf+v3hh/JlxbcZH55gvfwJwGjESN4fuP+79VDpR
yJrBbhGCxXn0RKZuHcxWQF5NTZgKsaP8bFNt0vyVNSsgmP0ZMyPTnrOo8+OfGiezWAe3c/lFFzCH
IKpe2kqxJNm1RRWD1zQRag2gA7w5gXwJ5rgnre/r0S19tSpI2OuRxv6Ry0N8V2/WHxn8M3XzA8p/
4+uU+Rk3FusFN097zkzfKT1aaxAt8/5wlFbgbvIfd5+azdqVXyc7GzLgTXOc8DqYQ6HQkbgTzKGI
L3oWqjuwtPfSe+xMP1ItpPGBrmSHcVvuWDZbABI49zo6qQ/1EixHuGUUVqDXmhaah/aGMw4XlzZj
KKPhnr5XT43SEgV+RTVKPskDZJPS6SvMwFBlEzDMO4x7xqHx64OU77PQpUeA4FxLVINxaZCdM0nb
bW4TBaPVvE+FXlaX50saKMyre/oAfe7GyuCZcwWEFQHGQm7FfTS8esCHdSekYQCsIGnHKuQtW8uR
9KrXkCy4aPVhptZZe3dD3PTV035XcFQsVYH4bjvjIESM4111mA2Tp4uZIKpfAsU4bTF7mKCAattL
bB+1TDX/fZTYnQ9Deh7B4d74L/0JJ5+ASLI50ny/+3oJGa3AVpAp3TkE69q+1G6shaVUVYglsEMP
ZT45pSkdZga1nKdrQBVrkKffYg0rUzdzhW618gJeWAuNzYNK8t2Fd9A46VLJLE6Ftx7kdxFq3M6Z
zGMDvGSeBX+FTcblTpFTf8sYYBLA1aDQfVLHcFtiagEGw3EY0E6RidFh5+cxFPpKYvGOfZUHTBON
eXGAk+yYSSFvQKWMdewrhNyqytBz/Lq0anR/g0C4AGIFjHg3Y77BzT4vm5CqKQ8+r7FuLhGtjXTd
c1YEXd0EaNEVVoHUJLzWJvzLC33YNlZA8fa1UkLuoPshqoG/aP/dv+BQsjSNq6lFcmkhwkXHjQbw
ElCOD0SCDPcuZ9esMNrvLJn7dY+sVhInBeosU4GKz6DZIG2hy1F8Oj7T5Kis7PLIMUj4bnnNUZOJ
3MU1U98m/kjoPUF8zwv/LEsoP6Z6fq1lllIVaymjNGCizfE+4myDtnkyeXQSLBYkKO0hoUA1pGkZ
Aeid2t4sE2faOtinfGGAotURfSjJP9xrt1MY/PIxenolNERXjJG5T9W3QjJSt3/zPGG8P8AIWE+v
KtIowSBzX6AkrSMrbHf868VAnllG0HAVkLd5yORtwy+EF3usOQqiUvBJQriiV8zfgjFYT71nM/xo
AuZqnCn4KP2evT5LeS5ATD/lDRGT7RiA4+zBsd1MdZIBiQrxMwNL6Nc0FIjq7cCg01GwnxfWBj4n
yscPn8gQRWkaDz+lMlwHUo+81AZSrcX+SaeeyiNtfqgMMCz6MbVXYPhnU1zEBQW+CvFF2tTvlUEE
1KrNyPrydwipmy55VRpgaxdQWqM/ST/CDXqrs241b9NCFNXqWBTy4nsU81fs0CtVaGT73QASZVgA
SK6mmO7QtPBU3ZkAEY32fdFF0giDCYxNhVVOTR6Rf4DrkZ61rNonYnza5/mleO4jY5MM7qlCpFAw
kI0ZohOVfYTusAW7jL+310hEj49PfWdhDm5EiGbuoRempqh+f3ceo56EMNNbohz5WPIHQBTMSGNO
kljYv3T0oe3/G0Qk2YXHr8Krg7xLsMtXOir6OTo++72XgC+a/sb37CFmvvFKs4Tra/EV/dI1LWw3
ssdFX+TyrfFA5MykFqAYNn1+s2cn5UyZ6e2e9jhV1qxhXwKR678S7se3xorYtjtHyO8ILb7tKEBC
mHPqU6/Bap8vM7S+l37NokJVc/rvoZvDVTuLCGehYOsXev39vO8jhzXmbhSIUsfefxsPLEIBNd3T
tKz5N/civBD7PNPW2dGCYdCPhUgd8v9maAWW045waxtN0kUajWhnhPc9a0zSABUyyEUYELUtScE1
IiE5OhxaERJb+Xp17zTSgXsWLrOCmB8mLmF3fUcQANOIJldykPBrW1qjG6Ws6dLceKK1OU31R3tn
eToMEfnYrBQs0XuxrKbnkQPxINioISqVvU+jEDlfYgiH0xZiWm1h69+X8HtZYJ7DVSKXMdNECDO1
Qo1LqKc6qkaPsylzz8pTz2Q26KpE/ZEZLn4bPox1YMOSSjmJNsYIoX0t6lbecdeOIYnt+S8bXU/Z
rjJd23pF9xjuCDH2QDwmWaNKiW72BxhLKercaZSKQy9708p3bfYl3Ga+hApoMcPGcr479p9FoNQz
h16P97YrFDMu3sQoa3kEqzHugPH2ScurMHZ7Dkx7c03QzoopyaC9DXXfkxwzOI6nqOYr3smgsews
Gg1aiLUzORqskLXMfPNxBLWk+xFsd0KO539X18U4Fc0hfrPldKn3QXq+EJj2E9Spbd1D7IWaH/zO
RlSojmEyZgim43IZeJrN8zICR2CqSicFWrTuFYHx4dQV6a+PFa/+ErFF8ecUjp7QMzzh5liT1ph+
mCT+vV86tZ05t/6mWeNXaE+8ezAFbQCs9i6m3Cqgd3+uRt7blR079DbExZ3YGuN84fb1EH23YDLb
wnUANeZLv9VOM5Uc/kvbdqDW9HX9OLeM8ED7Mu85wDJPZvsBpvdeJP3C/3hdGv0NNjXajg8Z3t61
DR/HDMQrcAysTu4LVlURjVrDZ+vXftiNvR6Mba6rWI3ybI+EODqOJTk+0GwoZ4SrafCZxiW6kCF8
poUF1t7uMN/1ydG1fA3OZuWxbV40J4+7sjmzZeT5f7w9wV3mQClO7YlhULRxT7KIE5AfnkHnWY3m
XlklumlK9mo0qqXJuxsVYREX8L2n6w0ZeLPnfAiWt2qK2CVWCjRIqHv3m+wFh7BE/qC2kBpcHAGD
12DVHfXYg82/W/gMATiFbcquLhIAvC2jRxFRS9ZtZQ/7EVhvHt6UrCaxlTXN8h53wZqUVnTmYSst
LikbEKiVnGJiZ7iTuQXIIKytr10Rmd+p2eNqABUn9Y39Uc5pr3VWMDw4cSrwagIOY1GCsVzcQHEB
8sB7qHRqjHSs8Vu5pX+ZFXpro5o0bIgR9u1XKEBqbsuCr+BM2kEuZ/gV9En46MPamtK3jJISYELx
L+PxeHLwb3hChqrXHm3TPM+mG6s9a5g/5TPzhGcE+oHrVyWdEfuCttz/0kF/bHt6y4miVCTrIguD
g/ufm0mpvrjUggMLQyeYrpgv0By37XKruBPwxsV/7lB1YwSg4NBq1fkISxW0blnT0rtxctV0FyAW
q3OFpxS3UbyjqS6NsIqPRb+aAq35yWvnxylNWWyfoeF0xgduad7Pt8E6BRArg9mQAo3r3vvCWzZ7
PnKw9ywPEsQp32GifLf9JuB9WQE49gNgU+4BmxLwqCVmZmAcYGBDgWxWK8Fb1AJhMDqC2CDMvUKr
Y88YvP8j+jhOfNikcRunTSMDbxccYcEv98NnGW++65b9p8rE1w/vuwcHcSNOj9j8ANBTMD28zpXY
r9GVwmFExDip7pw8Vq2rapZVsqpfYaa+A72V/yZbxI1dEl5deAh4KRU/z6RXbXnbweySAonqbXK6
0ZEXvOeu9qU94vHqShnL1RmzL6MgDj1DHcEZffwTKiFnoMAGR7vvG0nLqqGFgpGZKCSFa3OhApeW
mihlX4ToLzWJhZ6yTSV8IqBCCQXMtP5ClBHcPvO0TTRqQFEzncjNeZywF2z2PIywLYNeGeHIInoB
5cqQcAr4maHJ/zTYPFfwZ9iR+tsHRZR8LOClXysOj8UUVS4shJ8pN2rtccCCwcl5lczoQso/SLdT
96U+iXjBOLyXN5KEGwXPsGwDlhhQkLelQNUAjynS0YXnhJY3vKWbs+OMShIFH6f8hdmNonFJNJFH
IHW0OCtLi08QNIlGNbladUlMMjjufEpChnnUtTYcncXOU55PAMzAFUroODyFtKQhkB85zHvumQSV
myrCaNUk+LJM06jk35t6a6QZFxyyOpBaycnGEkOSlvY+pKqF5Dev/kqXWty/Wz3hBmJZM7/TkDen
tqq48DebyevB0+Ioap/Up4Y8Pil4lg+ZbcJUcs8O4nSEw171QekLhrmoxDUrt30NCgElzeJYtfLt
Reozt49wqRZhrOZ1Z/x7P+OdIcvewmBVcUuYOowzCU3WL9Da9qTJCBRU1A4dzGOPiyR4/zODJ0W5
ZhstUbQ4aANfy/pZJGVouMFhV6bMmQnDYBIlNtPB6n5pxf6sUmVz3HDH1pvXVVydZPzmywjhRBo6
5lElbCpsWqMAB9Uqwc+igQVyMW/eD9gLLN7ULzPJwO4xIC1uHwm7clHzva6eriTP4OK6aHTj2b0A
0j0Q3S7P24VO0iNgI96/r1kLZr9DFgPrfBgwbmwZZv6IOyZ92YxpU7kNVhI1BHvQ3HKkBeklETym
a17+jypufw/pCRWQuh+9Z/J1W22OE5hpD2ruaBmXHwH9dCL0ju7DjqXKPnSn++chm+aUictPJ6iR
p/OTYoWtCs6qpB2+kJDe3qqis1zrRuVS3PDRfJW7qvGrS7tudsNng/rMEDzETkjY+aUNoBnND5/6
gAv8ejhO2Pb+VmuwkFTuM7SvBGO1QUS1JZ9dP16kjJBv2/s9vF8RLR9QoRvrLkd5Nb1cIowVKNrk
ALjHmSE4fMB2GXtLGcQXv1ch7y8R/1Jr7fDCM0n3CEsdgZAejNKEBvsC7IVSkKuWB3g7xPt3g8aT
HfBhCKXuhqicncKrBtgy05FUHfagXBhuvJ/AWJaRKmFMAVdUwqN+34SXa6N3A4YD9w+G5zMLrWzY
tA9TYow9bJru3EZH2U8SSPWPoMwaxDhukuv/UUdMRsDmLnuNMTUTJldo7xYJzBk=
`protect end_protected
