-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
9mOoSIVLFj7c43BhI0BPAfawtk0nzRWr5bmrOEWBD5/82wt5rNzq09w9w/gIrWBM
0yTdBq5P8q4PWaAObwbfImwedOHJuTSu/3rRgkGTPH5LS01pxMJU8zdcOxFWBVOk
/guJNcs50yZK32U3Q+BczvwhYArdZOxh1bdOVDg9MD0l9iGWtmTnBA==
--pragma protect end_key_block
--pragma protect digest_block
hIrxp7KkzW+FlmQPMelQ1SGJbds=
--pragma protect end_digest_block
--pragma protect data_block
tBUKly3r4spCTBC9qeWf0XWewqSc9aKqeOJrogITIVsW7NROebCf+K3YS323E+PI
l3a7IqrZlNn4FOrtrsgNiGpa9vcbJwu8te8Fcw9K+GNoQDW6EusHJJLhz4wN1e9k
/v1kBTlnSeVi1UcL1qWiJtn8xcl+I45yI+/I52HbWi/Co1GRYeFWx35Ri6Gw+ymg
auCXYbycj+eGDB94iC9cjURDlEp9p2eO9YilFZ/sPfX7Htsa79BEecQqa2JA2EFL
zjmIM9XMD88kxGiYQs/Zs4c4cUBBomgM09zoqokLNLTNlr28FWOTR/WGBCxpP1JQ
RiZT8JFujlyKiIKcaZr7fLW/hcLIGdeThBg0tzlPbsVxnynkzSh0Un61jtLGKidv
XTXmaeuoM9iFnwuUl3+b5CU9EcdIhwElm5H5Lgl5MIqyO3PyE1k/KGR5/eIO40sp
u8kuJ007g14BCTWwsgPNi/asTAXPZuNzDRnaBiG/YUbn6qjwK5NzSInZH1m8sZiT
dVA5Qas/MH6RoIcQQGCV75OvPfj6R/df7Rsl9LujaRZPSosUJSYTYuWLJzYo+kLL
zIu2gmY5lHYyC2jWAoE6gL0dSB9BAnFLTbWZ6vRzv4ikgH9LIuN5Pi6nTHp9x4NV
bVhbhX5OmLU1e5KOhj7udYJdtZA7ZVluT1tqd2gmqKKaHBYvs32lCrpQSWQVmH3D
nhZlk7hqdFsrvTs/IB93/EK9vv4ylpKlYqprgogylYb5PFC2jTH4/ESzJNlTier1
kX627K77NIza4r/710HZmVXfCo/zZTEtkAdUyo9RYKE0UB0VJ3fHY7Ob3ZAOLBz+
TKrfvwunS9ni7bFVSZvFN8u2dNOAFgh/hDDwBqa6bHOk52ijFhunra8xGeT9SSbv
oLK8lId7U4asH6r9ctPJHWkv8Yc33NdaZjzFHcJ5u5jWr9KpJ6dSiowTmzZq13z1
I0HJk9pQfoHDS2fc4e5/GxfjNvk1RK7YSGSSC5ky2YrWll8XiW3k/R9gWrxnwBIc
A3KmAHLxr1mqRg76/UTwJoJKk1XR412c4XeCh8Uftwkr6RzW983iXBNUOVIUr7w/
E0beImV/YrpI9NG0TUojCZRQwmFcLtSX/xX9zkEams67OWfNbQ98cp8a1FOTCPT1
IIrkt5oFh7cfQPlhFcyJyxc7NUXP0QpjtLVl0INpmY2nhWF3FpC0ORirY41Ygi1i
0hsCNzh6Uo7GcsiJAUPyEMcvqefJF97YX3gedwh0XgeOeQTj5+fed53OccpERfFL
bDEUzNwapjwmBdWjgYZKjPe7x6wSlUhm7SnP1OfR0SelQ4elem7souiUKmpXpXYp
A0t0/knIJt81cF+YH0xWFQ8F7PPOMOftxv2PwlezG+YxszDpzq2n+NkkCtm+M2Gu
YpFtv/bQQ05RRzoh+ZgrZEPsb/JzzZSm/EbBW1GJidBaof7pE0wrLCbr24z5sgxo
7KIEWwpAAeknw/CJRi/Q8Dbtxc9ONM7yVr1ieB3izpotfTLr+LJJh3WZspn5exFh
wGyzJb9Tlgw4VluwZefRoeIJ0/N2fX865TWHTXg3wWCN3aQSgiGHIq2KEZuRcOwN
atpStWFysTtM0ykMdZ5htExcXnaAww5gIzcB90Y2Ap3hYtLUd/DTzcem3+D6zRHu
nCn5SOqIZMlgBTOvqjyypbiRT/q1Tha2EL2B0VubqYG7Ctd/q8zxqL2QV3Rlkaio
8HCQrEsDTFolfstJO9BYS4KsAsgrGKjhCUqaRyLVGeYvaQ2id2upvooahavSlSVC
M3SouOhFzHi2XdpWAmpI9W3C6c3HAsnngzFkYsZWNfYKlpsDCQbQHRRARr1eEY4i
j90h2ITEL8XEng3R/i9bXmoDGjyNNa/9lY0lTlmJyhzruJskt0mDuJK6aZ2YQGnA
JELq9W1/ewy/HQLiPd3OMuli8keaeIJ75zCY7l47/D/SC983iBArc98QpVUDrY4K
ZATZeLYQHGKdXSbCl765CR/USYOrvgyyXGvH9TUDxLXv+qSgw8lMzh9Dg6Hdoj9l
ApZraVyvVctITfvJs/X4f9vmVUZ01VZT80xNY+xyKcJFTY86Bd55ylkZPzI5Z3lz
2SJoJLlA1cQr4aH3D+z5kcbZE1iVufNgpM+hIo0UbVy/f4g0+zzKR6bFZnNfYmMU
tvmZysq7pvSe0rGeS+rzHSm3hEYF/kVzaxNwMUPqiQvCoEF9XDdplcmx9O7lf9g0
oOR57s8C6vgqQ90QnrcxKWHhX8qQoMKWBVbPkdZtzHniXTIgqQCHTzCM7MvK/1RU
A9oH8IGbQ3VAlNeZxB6XNd1Fl9uXFASB4gEH5X8Mx6XBIYyVskjGOPMhYQEIywkq
VlrQKqgYqBkoQnurzJH5v8XLaYmHDDwmQDyh5T65TC1Vfc3+oSumOnVqLvSW1wUZ
QfHZbMQ+XrlLxyTOYO3s0d5fNh/0MM2k1OBMf4/ZCPehh4d8Pd00kzPu+tIFI3lp
yl2t/T1SVDJ7UUfJ3rJoRs+mGKMvq3qUXWt3ydq7O2OlpdWwCcERrhNIRMqheVrA
GS4H+xIW/GYg6VStgkV5armbuK37UjnxHJ4U/AMNFa2K7OvYkS8iCZatTRB681d0
aFucaKzG7bP9cGeM+uwkLWcCFw4c3xgsCaqAzmXGDnBfsiVTGE7k222LmxOKQc45
476y/E+XZB6VAgr/Z01AjyR4Q6DJLZQMAZCSAHsgknmmTJaTMXNdQBh9K52IpELk
w17Jhw+S90hl1d6rs7d3ZkHN8Cxsne9HBCDL2fUDhgRCkunPWPyxp/WdmA8FHED0
ctY+ysgF+HScH/5dmS5Lwt2GzGVPyxXsubaGDYftRnRW1tmEVdESZBOeaRE9p0ff
eaVBDz5Gh70Qvdto9KLPGA3xbJNU97aSlnIJ89Q/nluOqU/gvCRwfcfFrbzZK0SM
ki76K1X6Nhj7Cl3g3iejJw1WCp/8DSzMtf2DIZ+eNMw8VSz7gfe/vouiS93t7UKy
u2+hAXlNE4vOtsS1BF/uzMPyHlW0fGMklRC1PFc+0xwLuRvyekiFjiqYONh73hch
4VpKYw2+uOSh9HXk1vqPZM/OwFava75ZH54Lg3AJYSVWsc+FCXvPp5QVgsotouEZ
I70wWJPgLgkFmRAUpaADGlSkKO9dWdtZeSPvOAYylrlluSbWthHBvSItzZ5htoZn
G4VPgJdZkkAO5hDmdOZdV8zPANdDQR3V5M2T7GmkTRONd8t8mk3rxNsh/xHxkoX7
Np7v+FHmSKnxBHBzS6hMYu0V4ELQ2DTrjYvHRcYUWzehqqYNJasPW9PeIjbAGU8I
IE1XNklsQ5luyYKEOUgE91IUcip1E1suXBRrz/xdl8W4F/CznaX9oMn/YJw0I8GC
J+wQqXgzkiVGLfgW1XlB3kDjJ1JnkFennc6gyZpQ3P+RjcksdhP6BgXIO83OiWB2
OaGdDmtRGzpEv3FMKC9WAyALNJJe1KqANT8qhMBLpkN6MJTHju3AOPf5bSvN4ggd
Ynx3jl3DzrsUW2yOiVuPrCRYCFnTuA3r1Wi08B+2UpQ7CPUfmIE0rFaxC+Y450v+
mWxGR7dEWisyW5kuNjiWakt7HKixLAoUBSwOL5WQtF+HheDOKitgY0Kixc74SLDy
sMjszCQx73hBkPAl/O8WoxHLi6KAywnVsnwNAsxoDr7ghKNIwYsNhEAmSRvqmNph
QW2MV5GHbun4VnREs/jGqdhtHHmbIQYGN23aqSFEUaoQ04CHrMKVCbnv9S48/ndU
BgcWaKJzmZPZya6DZwSFIpgrs4xhw7G/VWIVUNEkmUGWZrmoJXr0lKAp1hk0SU8f
myOSE4LMdZJdc9Gx5GZuTfFNJNU7e+k01F/AeDiVwXvFNbeoH4aOvTpv0BChMcIE
ODcc0L/NEfilihiXFXf66ilxepefALpSNN92iIRC7vCV4CIohSlo4ndeHnWxbvpi
c3pHNrztQ420k62LukDBfEvXU5njlj0DjQlkKI1p5l1ijrtsG+j3s9Y6ejGbwqql
XpHow5SgBKKg8uSLG8wP/otissVNgB8lKAvL24CW7/nfGD3Ytv6vChZtt4+jli34
dHHmGmOSym6QyJRw2Xwww205eC0silcPF5+x2um+sa7WytCLgcmdCu0hqb54L6sk
IeQP+miZMjHPrPFpCaf1GaJAnrrfaJZ14OU7fVsV/mC9isG/2gDkjP6sOsxZZc+8
4YDrW9KTXXz2gkpkFO8eDjrHRlkiSFbf6x50C0LdfoB3ei0ZsN8adpiaYjHpPx55
TW95R5PJjG53GB19FoGZ0zaHnZ4GEm7LsyyVVKR4l07V511Yr1MM1hK6ugAsJvo6
V8f3oBr8VFlhCwSOR9ohkCNLHW2G1m4y5GXG2+cd2rGkDmUmG9QEoJLcJJs00Jos
049XZxkqCr/YMIVhdxsvYX505eD/FawYOO1eqFkK0Q61IOYOnc4spr3e39gr5951
U9LFLP3GelIvLD3u6MbKIbSYfnUyeSdFln+ofpL/MAMjm+ygoZPkv9r4KnjaqzRf
My5ZrYvaNg9tMA0uraUdpNRUm1vdF2/cjlXvF5t/ogvZUbFNNKxFB+RAL8AdRYfX
CNVS715tuA/JORFszJIeKbYrAdvvhdOiFptKpUZM0eTeo2ZKqBe/FArFBHI2lg8i
i1fGCKFDmzvTaHaN7scWhYXpzi+/4nq4A1vsX60KexfKObpe2g41Awf3/gduTeSQ
yeR0Jf5gXYAU+58+5y3fH0wvaUdhClGTLwvIch+ZjpYVu7zIZNaSoOvB9RF2MO5K
7w34mred8bmc4kpekLNTol+nUuNHCNwuJBEzYWQEWNz8+4K/J+JBsfxYRCuaHIB7
gytgl1VX1/fi523xDiSaU+2Sp2ArJJgzLVf5heBPvNz0eKvkr48z4prycKqJht3H
C5f0307Imey+DagP+9fAFe2SWmqmFkvE1noeneKTacSUQg0A7cZIU014/O2gnZHD
4EIDxSbIqRjNfp4WdyNBTclTab1x/QVCEg86wrXWVW9twZEmLsKnnUJP5rRbXwtM
uMLTF2sI8nols/f8gLiain3QFNQPReQ6A6b5EAquQ1tBWci0uxtSxec6XKcUQmKk
pKvVNtI4qcgUB8AojoSV++91nklqYc80a3QQ8qCES00VQxCUv8YFewG4D4rOQRVo
w//Z+HqGd7qaGQypMaKczv4pV57FsuW3QVNATBYuBW9hqaodcUEbxzXT5WQZdgG6
AgP4wUNBNdpUp3AE+kAPu5n8GUjkA9G52A4PIuK5NHGRVh2XWa7lg2RdbhYQi2Ix
DyNz2tRVC9igFGMZ0gChriQsc/HtmbcH4imqCXubXKSfPj6OrkZHWCZ4AT7npmGh
dL+q7xpI/Dx0k77YZ/TQlsub1dLgTtKvIQycJpQRT/b0vEANm2irhAfC/0X56Oar
tkAieItlXTUoMv1jok/60DX5P5MVyieUbRYUGFAQ2RorvxzgKsMnbjZr+AJqCgy1
cSKrUyBaGUimLUmbcmeNL9dcCawpTxX0+rjL7c3R8ZEfBtkVVZVMSaT+HD8t+3Ao
NNcqi0s34334ibYnT/s7yQLSyn3JUHBDoV0CBM6eX6xXAekZ9IoDMvHJhlML4/l2
eyxBb+sPhXX/CZbnImToeOFZIFMFUbzuzkaUIjuAFwqnrP0HDFpDXjJdltRsdjsM
5s/UuqJtzV751yjZQ4AvyCI1+Sa35hK/95eD221meJQ/T2+s3t1qIpV90MOuW+rr
F5B5UFwflHEDNfRIyLbv+18yyn/zBq5fxF91nCpAr0vluSY1JQ+TAv4Ie0+qqQHF
HvbtPEepyp7WD0bAK1UhFqlK9VzAZFghtC9k4XliafoXGOj2An0r6Qx95vJZQYu2
0o1MHhp5E6/IQ8B5UiQ7bWcl/6kBotEgQ7sJyP3IUR1t9Pt9UrM1qzil+/TLMFS8
0jGjeI6qvrbKpM1dvULKKPw61EYe7ExypUEIkEVzmliDBT1M3aW/alx6qFQMmoXN
V2plYiVEwRpYZsEyMctQBiA1FiJL9jirNv5DhqRUpEIR+SrwVZ6kuBmR2u3sLX5j
AZklS0VJEZkfFWt1vWXseyDag23CT+JBwobDmQI/plq6o84ehpqWLBMio90Ozs7A
uCTCyCQ9rzCFsWrfMZHMULiAmVODy3QX9M9MKlzh8eW8UvSwC1EP2KhKbH4uCOKJ
h6jbBNRp1MjXP24/KYBzHzvp7Eecc2Ze1G35B//hvnS3obZZl/FiH1DtSb/v3Wd8
KRzkD0ma7nPjy16qPOVXohe8OD0OTzlwsi5M5t6LMi6ERh83JbDerSPkfWFaDx/y
O1N+z6yEHYD8rmgM7rNsMG6t3ik7VnuXPEYDaesgXVFn57qx8W9lez1r4YjF/WkI
avXqbB818UBIkY0hiXsKbvAw7xQufwlDTKn9lp8cF9Bnik8NoPwImREJUjrDsk2m
DgcWjwo6S2sK4x/bFoxciYfgLSXLr27SRBvYCUHHdm79B9MQE4KlAcmMICZfFS9g
T967VwQb/DxAAsLwlYLH2Y895jGqT0jSdofauGdIzMzWsyvaUnL5FT+XuF7+83RP
fG9/mCBLftA3sXfSsqOL19ZJGSscB3VAJ4FhhsJUs8qw8PUShCMavP05lJsJzWHH
e20t0C61C7Dcrhgx0yYz1dsYfZjbakL0wlGfaTbEXa0k4WOK3NvCCHUDrC5/g+Zp
dUg2kfaLyY3YWYkUfIQ0A7NMuPQx7eB9QGDiA8ojt12GAGBPCD5g8l7/w1Ovid7H
15p7o6Ir/6VNEnFhTBu61h8CV/FQ3T0jvgx0gXD1dp0v9HG7neJI63jyKeEUJ7IH
4uiT0t+zvr5rc0nviOkrR47wWyG+XLRodJAEX/o4vdsT2bnqorZIAaFqgH24U/D5
8tFhkmGNbsG5XFfs0IdbAjhvaKwuETNJET4ZZgmnYmuJTNOOhMfTpVJcCPaHLwjl
27VBinidIFzCoc6XGskGrCIK0rrTzI8f2K1ai8wRc9D3cphfh1eas8ZriLWhrbR+
RNnvGwtFNRMUXTq8PXuDS3n2TtO+yjEt0F4f4dY5zgKex983wNucxBLmFgOE4S6l
kOKK+CcjfToXsCAYDzJrChY0fuOmylhClo7V2Xb25TsT89rzUKSUltLuu7N9s1p3
Lth2j+UEvVDTmtV8sL7yYRbVvU+AVuwmhWUJsv6gXPSX+L6xr/F005x8QPkJWU82
esQ9JsCv2ibpICMBHXPIEHw0ReE+TVubkIP2yZSBsBFBWxmSs0ltSiUj8H3mhEIW
TT941d0LK1b4RtwnXzpLRMXiSBhm+RTQ6/8PHE9QpzL10ISxJxWgya91wj4BxK3D
itZw5+zUtZARNDpQG7T4u2uTd7uebklYKS0zh47P0isnOhcVGemyMzEyLlyQHMeC
jhYt+nc1sY2/VmmW6PfLKSDof12tH3fdUgXzxLmW9evmLbmsWIwHZpH38hYsT36M
UhVeyK8R0tflgXaVzOaToPeZ21nDj6kqBNDCxeYKHg3c+J/ZzPxN8cwcqbD5mXym
79evaHvOPDfDG6O7V4Gk9hqqr0qUaT6wRCl717o8WLXkiEQvzejeN3izzy5BeVzN
vp5ZyVJw/SYTkNN5h8L53CZZe/m+5hrxtjOP7+jRgtqoOWCsV/4QCsveLcQkRHG7
ZZzPGIP4jmlLtDZGearoh4hIagHuOJvA6zsPhH4kixsVvScIJ1YVUhBwpR4QrimG
g+g7ELzCj7WYqIdpfH+LIRoTDwljkX5f6wIWAvuM5wMLFVE0LsL2cKhXbFLWFPNx
j3GF8k7NohZ8gPePoU31AvMFrS+ZYGQlHfx7XS7TAz5e1vc122ksXarJx9opMhaE
CvbdNg1AoOWMtYhjsPTB2kO2ctgCls7mWip6cIe6Jfrn8JZqaVJzSsxnVfge9fyf
/trS501qZHG7A8zpCKMuyfj2tnJK3y39DExx1MXo7y4+mx03iVTDg+YBgRTpYlTP
mA+8CqJk8MtdBc7DY50SfcpO1B8j1SChFZqfYpqPmTOBvKCOG4xEdXmnul5u6nQk
wMUfgBps8TbGIrqecpCNz6O6OOsnOYi9effnb8I5uJG/mn1jQSr3kC7OWPxaQZfX
KgeoeedlxJbBSNo/ngHvsDYTFfxbN+H9sStRoS5iDa+7BaS2G12sXMkVB0we+46i
LrmKo6JEItoJSS/sAsH8/oRaPqEk94lhMY2rW9qKiU8PwTDalzLcjMWY7N2C2HTo
xd9QiIXWALOJ8TDmJePNqfCgftPxKcl1CIVpd3bUnJs0aSy+spqYRdOWHw7wWCmQ
qip/GThKYzBNbvtmbqE65vSSb+sQ72igAV8OW+SYndNhlwh/aAh7cSvASVTnQXM0
eqBK1ZalfyKA3OHcD4PTTrrIr4uunDOeXl2s02MddwzCz3d+JyInZ4ExaS/sZUnF
qqfQBgNteTaS+EsaT142aURvIx2e8BaAHiQ4T/4uzB/yb21jKwYvT41F90iwxddx
sZ5BwtvfHmUL5RfKLVPGbhNCklE2QH91yhTGdIfVEPfKMq1DUuDm0Oa5wQHHvOen
ek3QT4GmMMiTHfgzxWnBUpVTFLiz/4LCk5lINv6ibBUJU4x3MA4IjP/cMFAjA0/a
TnSMr+C2p5uZJmQWYdU1GHrqxfR68r840Y5tBaG0S5+APiPG+1y/oIN9MLaMXjku
nR2MghhMBnG8XBrEK1ad0+nFso1k0m+AFVMBzIMIjTP56i3AZhoxIojPXRo9Ys/P
lUyIsurwg0s/DWhIhK/amUsJCljsl/uxYqWZgmP9yrmKIXbJrfX7haWZ8isA9YVs
5WOSdpkmnThIPNPYjLEuUckotusEJ2XkmlW0p2w4SdcJWBnaRcMqt6PxbxOnrK3V
xLjVu112+vtGvdccZWW9KMcL+CLNUih9fZVTDjGt6E7439GsmfaMdUZWAvMU4CL4
UeQ+DrQtLYQBj8z1/06FptEMwz74LFJspYP72ja87UGgWqjiWWY77WsGNSiEokIf
CORHXgsoe/KiZ8wiZbt4DxTrijg8wFvD8rEySBvv9uVDJweLAIEDf32gpD8F4Wck
pI+cMNxKtN93Z0mWvX8wJQJ00Ldg8M0iRpUTWEI+NrnlBZLxdWo1Bcf/ZPg/VEiS
mA5LbJYfH242ioRhYGdW73D7aouYd+R54gD0JdtwgQGca2lGXGZ29zfsFqS4M3hJ
dIJoLrsCthoSUgMV2Jk0tFbeZjck/d30snmxOKzB8embz0EYIX0+SM/c4Isq1CVm
0a7vlFrnu6OuqAMHxWKbhFHc9EMQiBOWKpxUp6/pmn6yS8PEQcx/ENjqEm7HSWSb
mewPNm/15ceDxcRsIVDprkeFbBeTPCdqWDr04bylBiUpiU8S3vIxxqcxdmzCe1vH
t64W/LPl3PtJSS5CNKe3IE42jvUnsDPnVjYF5PjQOHQyyL8HkOHf4RoG5zI73eqY
EqsuwWmv9rFlCbqqQap9Sa1+uZZ/Y81DFeWLuy1Iek/2+26GoITvpI51jI2l8tsy
0StcBanamAa4MBGFaq6trAMg1JO2WQahIvsfRvIoXJR4CKByYgQI+SiIiE0ulMvk
zM6lDUoJ0Xa4GQ1kayDId2KEdhqoLw7wDdKoJJ3fnqBy1g9tWTHKhYs2/n34tZSc
5Rkaoag4t1PzYjbIYrZLeaqxFLsS7qkIzeVncc7QFrkfebdDTYbsydbbkKLZO2pT
caF1z3IJg0VbyZYb/FffsgBPhmb0KBRMpam1NSqs6ekI122CoD5SoUpiYtThjKOT
KEsaQgjvTs0iszYXNt1d6JkF5t8xKRtLNjGseXqX3m8CmDDwCH82KdEvnDU4gziK
+dv0Y++lHByPnUkQneHJ+SGXLZ1i+NqpaJhYfkZ6j0MvMjMLfktoyRZ+dm/j6STM
xpCJp0NjCG0Zgbp+FSE4f1I8kYNL6WGEzgvb8lXauW3g/K/evMoeSp4HjSAuViEp
734uxqDn6rzF3AwG+frMQjz9qmCGLjUfC9Vm6EzvmxcX8L9wIgGjNklZSF0emViU
ihqnxAbMrBV8ZXiiLhCx3ZF2d04trxjazvwiwMpZ5o8f8Py8z55WNk8b1YGQ31jU
ZONUuhFP6T0h4AewbsfNnRzrY6HUr8DPxncF7+RWlC1XS0FOmuTAXsVsYaMa+7zv
J86a42UBVeAAdj4qEvtKDIJIuEDJfcjxoYGN5jpx32NKVcLsgbZkcK6EK2fsGXtI
WGIck70At281U62fwNt7bqsIibyCkZy5skFVJznRVH+aCjF0nGTiMLs0M5Pcm+qT
HnS0hRZNRhQYpaHgOYCjDf9HHWBHaY9a6NvhI+mqVEvXG72U2k+SjxbNpX67BIR2
rrO84ENzvD9261lBxT1KuHbH7rTq9g5AsBHPcMLwNzjTl4qzeEY0ajSFOHS3ocRL
MPrKNb82kdifaq6TgWFAIybg0ZHJijA8U8e4O7IHQCePxQEgxrLs/ymX8utrKg7C
h0BvhlJx/MFDxOcRDH8ExQ92sAcD7lrmgkDHTvgrB+aGxM1nPZwntw9qFYMOtWyC
1k/scfWctrqgdHeqCVpymQPMvtbyCofMLl7jfP45KWBSicB2oO7i1HnIZITBFuIH
Ge1MY1OaQ8egUHzEC0KIOVUdTD1kFY3YOCFRPawKL/khSyMczHuczfjHPLqsmZDZ
bmlEl35aKHsj6J2rP7Wjl/8HH97Uag/9dKhzhJZrSXQs6oEeVrCdgHPd67gFmd9N
k+3cbCbEJNigIAabi7VgpkaZYoc0L0OK9bQnERg5KJLdXAOkHSKTafv0clsdWg8n
rjUn81R8+M7lFcpV16M2Kzw7iId16J5b12I8SGR4veN6JuYUO/58+jYs+RQzSllF
uYxIFYf8BZNzG6KpFSLkqQfgj+qMno9/Bqi7uARCQx9rUQUK8aANW1yQsNMaRUYd
CjPEgoDOHKwwYSnA3+br/ZLniibIH7V8oiXncMbrXHkgk0uCSLUCRhzV0LSvzra5
RKCinoeEQXNXqi4OF7Y2qKlqTwy0NyycZKoSWvR0xFGjeKWPF9sdV/zWp/kiDQC9
wzq6C715yzGVRS8wOyXpaab0SlE9+Al2wT70bFZAB9haudbyq7fBzFy8MnSawrnt
rMujS6NbAE21AG1MWHMLghOIu1KLI90+ot2H1yOvEaVu8XMwLHB3YTT7yL7NtQra
uAMMiNFocZ2IIuPcRzkCqzw4B4AhRCtU0pZwTNUDiTYt3fSXsP2g3ycaGAZQ5OZs
gFIkyX6cmEl/hpAMjxtQrVKbl55IdxppSjyi/oPIdlOwrcQZC2UPoNCxekK1xY+2
G6mPz7H9uvdJv0RW+JzAbj/DZfp4GwprQuQdJhRtD/eOjFqy1JafH6kXHGJgXo/z
VAe6BMgkc9GdKb3uVklxHGN7XqGWbheY0N1CFbExTEDP7P7rV1+SxgYrsnsEZHaj
66BND/hyq/0hF0+CMldzqOw5FWQUx4OlA+0Wfmy8f9TU2OwpjOcHf7MjMjUqX5a9
YZPdBlmojmdZCGuFNxS+NzZkLeGpE+Vj7r19/arpIt8RpiMZKIi1DFCOK5ezLorK
Kxfg6V9/uGZ9988LcmXvacck26w9DfcLkVtzDKhSOMvYHijFbKw7uOHZDde+NPsy
27DdURdcPzChRn2NznsOMkSaZ39be+S6jsdeoXLFkxqX2emkuzYeKJZPAM+CiD8H
JbREdRKaM3K1OFIOnHQ+LHJpvVRo2cuk8EvVJ1e/X8TJ0uEgrFvk1R9qyA8Sd69G
2m7nOnj5Pj+mTobLtZmCqrILBI2p8jsS0J22DXZw26TLhCJE0abNy6qZH4HKWWjc
2V/tfsMa9SxEheB2wKveHi0No2V3Tlu8SedsFnKHaFlaFtBDj94QHUdTGpToLDyJ
jF5MGJln2NjD+HwPOX4HhBoAsUovlXRtNv+4KjHpBx3G8MC7blipw9hNCakC4kBC
HUG6stIKwmyh81nOHo2AKc/t6KiBlE870B0hPwsSEC9CnpQAp3kqb7VvJIgmlSp1
lGhVYRvc6zbQIHp6rKqghTIi4QtFTPgDivUuvTo8i7TMwDPBdNR0hvMhQRPVq4QP
N5tNgpU57nJzuSUbFc7ibjcwRnJ+PHiCiN3MbseFoWBlbxY0xAoeuSv/xEgry9Ca
GI1/l6aGmhXUPEooSm0L3nieWgip/61WcyyjDrumkwm/DqZuHt+g37Bf547AzbCA
hTvnJ0mPtIYKNOT/V2uwUmKi80ShZ51MYAhmMRjAYITdP/e1dMb1PGulrxV8NR2V
BeZEJ+qA2S9uMyCePXdJF+quNuxTGYNSn6q01uNHU0UzO5j0kUE7wa5WHnQa06iy
FsdQggsGGI/rQfoPjTAM4lp0xCB6akNiaaMeu43BDuNW/byLSTSNLTpCszVRpEmF
Hdncn72YoZgPxJ315HTenrUioFTWbEZ21cBqHf0ZrhtPj1Exs22fd+7tLQvXnPMP
0+bZocN5n/0kegjkYqSyHSC/iXF+WBvY0tvwY9Xg/SpMbFTqz9DqtpE5VggDm79E
WMyG5tWDnxTcMsR3L0ai1BTNTBLMAFmW+JSq0YpvTzA2J4afy1xbRBOM3zuKCpnt
RCuVidzXBkmVdII/HJ1RmKJtSoEO/z7PiBSK9qozPgWyXwAhzbbB44CWma9m45Kk
m2BMCEKeHQFx9IHxOgHGiajFuX7EaEnjT6vyxbIEoMjU44IH39IMX/oY/vSKLZgg
bhk6As0jEglCXX1iwaB2RP/AVNoDyXuxj2Ds7nJzoUHZMY/V6LSsmhWn+f/iN9kh
5Xw9YmdfbrZPqRfTs9+oQh+3Nhgu9eNBTqqLXtp4DH+cn4tnQ+wVBixwBaSc3Et6
++ImPmofVoNxwVrkd1llE5CMUnKm6WFpFAvf+Po/J2vu82pA3ogdpWQQvtQmt6UM
9F3lZgfbM1uF+jbyf04aynwGPJBCSalKU5zQiCpedHNKvmbpVxY7rdU+cPohpcDU
hHNcieQM7HN8Af5kOXccCqzrAxG0pW7SVfJJgUI81LATaqYG+FSF3fp7Bw2yXQip
ww444G/1cKUy+J0mnQWrBsQtmA9tHO3w9K2iH3I8TtTFoCMx2vPcUTroYlZ0M8p7
lGI8BNuE5CPCOnLKrxZX9GDbidlkS0O25FUFOSga+GCMoUM9gFzHQxYd7s7j4Eqg
VTxQpGqWOwOQ2PFYuQINbYrCirxj2tNEcbe5OLntwEnStz3uzKXUF/G0jm9w2dvX
Qdf4q93hVO8IVVhb+KXbDZ7Z+D1J9nnIV07ga89jEBuO6fWsJorsFe9VSJ6TfKZ0
fD1qvXxyIW7Mb/5ioxVtW7uP5Am20fcWaerEbIHpxjI6nCe/nLYfq/2aq30mfGgP
7orp3uQ7Q0ZdYmKhSj1+37GRJ2/jU0G4w0CbstcHtHnJdUOXg7ne+c55AJRB8Icm
Qz7W6iRo9cGvzmsuaa2oSCgn+jA79AidfTlRGYy8Eox6/TAj6uThZrJMr1ZtEx78
KOD7ISij6BlwS0Zqc8QIAzcY/lhzOimACt7sY5cATHcpRRyWlaCn2zrXJCBzFoD0
lMWQ0RcR47imw6yXhPKY/YGWMEXhzNocLn3cKZKsDUK5NBQTDT3Bu82kg5y+jIra
0kXZlyP0iq2T1FCt2pIXP9VLiKsdgyJwB3jXPpdmFXcVcM3oci3pqRTVvaHPoOxr
69nTUcmXecXwwEnyKWg0Mo3tKq5Phv5nfVouT3JCBQND/m5Y3XaFGiufXT38rBfy
RtlI0ORt/JirybZesDU9rkYVn6jYZGBNS/bLLZf5bUsU5ypzOLTtOoqkLUK2SXoc
1LvgVbOb8ff+rlwaXJQ9TQ8EXjs6kwPJdzwKzZTLpOCcxjI+lG8E5L5G/EwwsUE5
VmWrjRdHfc3R95CyoMdRauDKjMcvona/Ec5QNvaZ+ScYTYXUZM5XV4P/lxdFXqXV
CoGCSSPozPycm4y6bSN7eydBmh0cAKDxR5YEGK2rvfnVAxe+hkKMOmI5M6LlbhUJ
xUCpko09dLQpfPHKVUcgfypjNV19iimmqFples809DlzsGXRqltOdN1qvrmZHwJP
bWhcSjKAabsTs8Jke0cMTg==
--pragma protect end_data_block
--pragma protect digest_block
SCrWLJpPuRkeZ68qZvykRCU+8Rw=
--pragma protect end_digest_block
--pragma protect end_protected
