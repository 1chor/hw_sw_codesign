-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
H6iGSWMrxseTw5eUu7dKPTqNcNOBkdr1ubrKrZqmsiVke/Mv0Szq0mCR6N4OSMLV
R9Lh/HWP/IGkKwiyGtYpYIfWvcR/mB5IV0AY83shryYGt6+cBBm/ieQ2usqEnxPu
KW2Dl8bEOEOdfbY4V6lRRUOO6djzzmvZrpHyrv9iGKIftStquBW0qA==
--pragma protect end_key_block
--pragma protect digest_block
Y+Aa3MYj7eavpIyZjUCtyRGNm20=
--pragma protect end_digest_block
--pragma protect data_block
1ieTiyOWfMgAlZwE87RN3ireBhL58vFc59Q8uZFWr4dPKnnYFoQ1uouFGWwid+0+
vB7ZpcPRLjNzCzghzwNPEwfzLCPwNcZNCpeH6yYlBtvbIsVGuosKv7yC135Yh5vB
6/snJct+agJYyQnMFCsgKSMfKRwbDWp+U2MLYueYZ69cJkmSo8+uI0d44vwwvPVE
+w1SnWYElqi/jBIZUGYcWFp0VPVcgn8+QZ3tVub52Dy8M0eUGXOYbdOhA8YTLeYT
lDRmrL/IAeRxL1+lYHoIgH2TDxW5XIOk8Tk11RG+GdnZlo3Ha+nD+HCGVPX4o2Op
naDXSlJyQtOBgoNRSmqLQA0v+jGMBZKR57up01GNTpIKMRC8HjZ4J4tpHIO8cylY
zBbykQHKxibkAQO8+93sL3xsn1LuCvjymruH3cq+YT8fRc3FCUnCyg/Xt5ZOTcB+
R+/DGb0p3GdlMrDMSFBZNUk7s5zPYHavpCiwfX+O8SAIwZ1Tv+v/8+9PDKl3qnOc
yZUPxo1pehjbNSpkF3MXEt0LiXVjruwHsyA1xPa5ptHyN+O0Mecor/smHhltEgo6
Jhbg1egj3EkfTR85Fygcp3Rhu7x3aDLzTSGtA8CSOyuiXDZ3YixLamUDHcyEb/Pm
gjvMkkaS4Nvb8m0TUYBXojkIfJOKhL8HObCxSc+oC5+NS3AfeiHtPzzXVPS67A3b
X8nOFj+q+aaAprSvoJq45AYvKu8jcbdZmzO1eyvQwXiDJFSahbDQnK/OhGpxATpq
XoxPBeNla4Axt0V7ZuMhCZKzbBQJaclxv011G6yP9WbQMqKa2dHH4ClSblbnpRB6
2Fq5IVCuqRtX6Xym+J3VY8tq5tilqut3TArNjlt9teOgeZbqYkVN2t90z2c1ZAJH
IaQGKtU4/a0haacCaJqn0TYThZyIqiMZi9C1kMy6eCYBgoDJI54cwCSxDcnD8kLd
32eCys8fIDe8VRuc8of2GeAfcNizreR64bl/BLla/3+3sXfzK3Zm9oruw4ahdx9S
7xs6ut/IVNT09ylHk6yeO2Jk/i/oIa4vldfEPglwuCgcrNf3+PrBYt6rSjuj5C+X
j5k4AFGpwU4S7rTcdrYftcFfEMsir0akK20II4kUURqvU1IgdTLiOP63/GyRk+Ho
H66zP+b9k4rRNipauQ+EAXACMGY4cO0FCBhStznhBMhG9AQmJ5YZz1TYoj4OPpAX
WBLM8G0DiXl9tPjnhS2DWMFwfzCE3dA5ypeJjpcFuG/3gtTBUE3I+07Piw9wFK0r
R1YafizkHamhvCTBI54d0Y6CeAtFMw9ta0w971Qou2kgIbfHVmYQMJONEhOycF2p
gp/6k0z8Avm0E2E/0kGkTggRl6iJp88ivyWCk1IoW0Isi0G+gX7Why7yN1VFR0SJ
92amBmkQu4ue1YR2uetxih+FqtgoiKzFl21bKoMHEzOSTJp01Pn9WDKFZC27cxmo
ZvDZKvWtbY2+q4hJvHwmLTjjoABuuW9YSKHFQa7+MnDEyzGMH43X9Yoz5NkNHDfh
Uc93Lnm/uMC3hc/iazMMK68F3G+fiOLrzg2Q/Ko8N0fn7PpKZKp0QKJRljVGluwY
jc30QSl8PUiFw0m5LFcwsunrhSYUvQa9cKgyjLDAkYWespeMGQ1qkP6ciM95WqlL
XBe3ESJyEu2ASomKSGeQUTK5ax+tJ/pCXk7C10cp1zSB+ZbG84eJVKpaCXBIociI
ja3RHjuEJKs7SLcbAn0nQWH42W6s57yMMGdXtwT6JR9jlxoK7O6cm78vIqqfUYsw
RpuAtE9ji11WDMIe+TPT8XGiUX9iSCn2vMsPogiMikgtaUxAzU+xem/GPCFsQ4p7
uuP0bqPdo/TMz0HY6DjfKsSDTKg5ph5Q2UykcELBpSSGrmKRsc9tgxtCZcqfKyr3
+H51+XvE+JiWb9aqS5hVGmckZH8TTFPlDSPWRN/5PxgZl3CYmw6NUPiV7FIAIgzj
yIzhJHN33I7xtC/jmcKKvjeZH8vhxJ68M8UmEMTz1/qAZcP0fQAIRLFxqCMm3Vx2
0x1PKHnci74iKJxbP6jC6WoMS5ycceSeO3vmaNtlmLpKMRnsMeb8xpOSycxUvYXE
OfItM5hVrJvAksPEzIocoKGH+tOwc7c4S0u5lWtUSoCCMURN9DYDaHLDiNOSRk0e
5IwWGnTbW0PkVjgjK2Wiuv/Jj6IiqzyiCyhLcytaAD0LCbulnplYX9vFU/wCpYsu
FLxmQtflwRjDmOE7KzA4Xrj9W4Jd2SB6YaYK+bCarkqCIU+XcbsxLmNpMY/HGEST
Darf09MsH+xkYIwRMaf0LvBG+sgn572U7SCw49AWmwZKU8p/+e6atLKnYt5Ome2A
u8Knxwzf0Z1v6CSmN5IUS+7mC2DYe+JkpDAitMNgnF3kCw22d3ObVUF/Dx7bwhFl
4bd0seTRx+moPD4Qg0CmIEhsdzyffVH10uVGr+ymT/0qnnt64Iz1rX9bDAwGacdm
DvJbgCtBZVBqJIjsqGh6lTOJOv7kD4cGGvvJSbU8bgtDrh7smgaMunPMk/R5sBuP
Keu0x6Pn1pALFEhrsTiufYCnrfskhu09zJl/rE7+oxwnwh7q2kfRXztb92/OTJEE
6iTGNjLKMS4vPWOd7BkKMIZMevVWO2ppz4F4tpcwIoZyjQfBRSYJp8RRIsF/3Los
TnyyfG7Tcuoa+ekD6lD5J1cUBfAemhz0kfySqcIz365sXUFJxjcgiBEGCcFJg7VT
AjV+pUbRvLjRTBPiXHvBG2Bwl+3zXcm5YKILqqStpycT++Xc3HIyhJ1ZiB3mvU/p
qTLA/5yoHEniIfFnFiw5qrTnnCML2qLYycQ4miMBaSr4DmLj5+Ikw/Nqw1y1RQWv
Kt/zGawZkJBYYZPhGyAWWamhmxO7tIBDm9BWwEyA7WjFHaH53LnIJnoHR4GzlPWr
GkEUdEoltttJ9+0RqD+fyeRMmSKGAjtKJQrVAeV/K+lA0EDRPrBdrBJ1eLiKDsFD
iH9pJwYETiW0WlsxoEVZRqSMp9pcih5RqF7Ar9TUUU2P7neNDUSE9DJ66wpbRiLX
GQT7o9JRxjfS2dkNrGmCUI3H0i0rvTkRgf0Dbm6Y6oOYXUVspMtWkR/Pq66DkhN2
6yQ1aN/sxn5FwR1i/qvGEbpWlmKbjLPzGGFLh8XeuhsiTTe8bDMlzEHJkACuNdL6
4ubrOoH82Ji1qt1Tz2h0Ui3PaxdgspVp2VdjtqaG6ccEoSRJnSCzwgGScxXLRUa1
N5WZaPGG5PB7tMvxdUNYCjQc3lI0hM+l0DaOttzZ3rygl5FqIZWAKuKMz4us/WvA
WpvAUMM9MBSPd4+LlZA2cSEMR1sKnTA7EI8P+b7lbbryeYXmXilpwIrSSyCD8cUl
yq+gflA9zXJxZiEwdtXIBglpaNTwlXUGDIcveAqMM0mDofjAvhg3wiGml2oc4BsT
8hyOSlUpuc4eBepLAMj0Nq7DXj5CBMcYz1Kjd7n0CHFcNb53ybpWLKfuc8HH83vc
6DR71PNIBlcrvTcsnNJ/lVtnuxvmUysxVtqWWosqu/e1Fa+d9x0ZPA1HI2jqdtX1
2TKTRulF0Z7daT8URqbfZ12K54EzXAx7Aq0cKPuNkDKK8RiLdvTWIdzX6Ku90G5u
A7aML+3+WenStlatzs+012jGr6ChQKw7PDsyin+ESnKYjbGQO7DvfjfIcup+2frD
Dxo92ONzjTs+llW1YzIRB0mecfZLlOviXw/Wqu6TiQQQwVl4pFnGYqQpfPp/Snqf
2v8i1otOAG7/CcyeePpsWs++UBIBap6bd5MJOvWHEaQ9ELK+GmVm2NzZtYub6T9F
tW1K/j+WVSgCVXhrIE7OVvxFakAQtwyuHEHj0gG70V0P+c0+FU10rXN7zFmKxvqP
8UCVels0XZY/zm+438ZtXFSBnMw1INd6dk9FMKFij288sYictEfT59zaRf6Wr3bA
aeW88/X26KM26LJr7zAXE5mmhkkwjosfig1KKgXtEyjqjXVTCK+vOgiAJ6E9W0N0
/7zlgMsueKsAwhW0XucXaJXYa4NV9tj6a9Mw7d3vKHgoivEwnLK3oJ2Qs3mIpGPc
P5jnxBp07zl84rQ4svqCvuLTSFKAwdWySlIExqZkyqbGM3zNQW73OQq2AMgHCPWT
QKpmKmGRK8ESLu6ZjF+Q7fOSqczA4H4QByMjpNw/fJSKygxcd0BykoXWUN93xGxY
zNvfm1icsFwNW8br6evAvT3Z+zWHfE/1aZ4wvgrwpjH1fnjpwYBsxJmNViPpB8io
QuWGDgTZYqFjwb4EkN4PEiFiznWlEGuefBOyuEXDnxSyRoaiNHPgBHZuR0U1aQIC
/GdSTBeVXUXeWs55VCQs+y0MOLuHKbTt5zjEf8ExAxMMwe3aImjSgiLcp7wTTwDz
hTsQ10MzwCoNKMRKFhDyTVdqLdiI0HOHKEhHrZBm6gKbeSEt/882uUYSTa72Pdnz
dFYdeWcayFHSV/RYn3AQuKWkHG0VcSIHoqqWMbgJoNsIRlMDW6MTjaOW40HhCh9j
iAu+REHP45De9uePvFm6azCLpQChrm3ewWCiXmYIT+dAUbPGKoH1UJ+er+24AZcY
yYdwAb1OP4eE3KLagmddSf9KDNYE0Harf74iRp9+iJDYnt90i2PBKFTHJRmuk9Kr
//fIPaCtXG2055FNEKt6eez32JNFRjjZres0wzOl46EvwUNKKVo5E36HRD0ea2lu
Hu4Y7A/8V2K6VPkpfGFiUeHXih2NMLPsNIJ2Eb6TtAGmbAPOgy/swX8zl+0rMhF8
d9AH4huKytHlUA4Od4FV0x6V29qu+8ruFKDMQ10pSaf7qU/hIas0ZyxMkFbgTo6+
a23x2/difyizswE2vB0RCig0vGAM68aEcEJma0Yg7TSva1W8zBnkn1mFWtkWMaPZ
0hJFU2cbOQyiXhZUi6+kN+Td+Hs3BOMpsaXVA8Wzo6sF5uYQQAXWVlxLGGWZBbsh
YFoo334kREs7GLnl0cp+YKkRlw5ABksMDIbFuARWAwRNJ/B7eLuMwz2PbGmqRHZp
Ed2VpWUU0j4TyofdumhW6t8dc/+nK5c09raeU6fhDFhrt7lua2hNmzBWRoKLu0lw
7ujVMZyOnuv811vkZngcgEYOjJaZdZWrMeq74I5938UBnMC3+EB7mwyWsYHpn3Xq
OF5go518fh3IBlgw0oW7y7oheGLdGSrXrp/nUXTnGmfEdHH46vMEpxyNrM9MmYR+
Moe4TsxtqwO6T3evpN+WRtbp5/3OgUBtvnw7gbngpaHkQGyrzvuku0jxHZqURJJ3
/qHGTA//i4lJvGPdCILnbEUQQ2mbg5Z2zW4CGICNeScjHwJD/rm+4wfS2RKhI352
NR9lONhKbnvhcdvyi9YEsN2yHXj43vjGPVptyhQkFDJ+HCWlTdKImREeVCWWxdLt
s8q/g8KGlG/o28zowdEh9wVpcjA6fdUnnkC+xiJBdvfQdXmYp+dsSTiK5JZEp0pk
k9Ye7NC1KRks8cet1rgdqhP2su+0vn/87PoyXEsGfkbvHr+O4SvYlJLz9H3Bl5Xp
Fa9xtcbCWZdIigxXt+YX7pj8H8FDwrhJz1OfUrYMiHJP6hJUIa+tTE0Zjbh26TBq
ar0T2407I5cn6YiWffQVukOLVlKyAx6bAS/qrbv0CDp0deFh9Zz+DtYvB9VOAOcB
rt+4GGWr4Sqv452ZDbwnHSu2UoFr4D4oEcAjp4C255iTJhdJlU08gXhtQ1+6+Ya8
fbasJz3e1hcd2fPLJudY8XJpiMjgoStUP/4/7Wnl63A4iJ+2qBnWxTBDN7pHclXn
A5Fcu80dvoyDhPhvMLSsOpg9yG2oDdzNgzB48dLkeA8cG4R9d0SkMWycm7D9xW7S
2oMyQZoTLbFjpiT3LmvOK4WUkPr18p0GA8qHwq4DmUo48jJ73N0Perrl+sSmz46E
jiiMYp2NQUmNcng78xHN91coFn1AAMwwsPfWXC4qdJ4b71W06DuR1Q/vcmXmjmvm
xz5utKJlL0e39ZdWSOIYMEPgknq7FyUGgVmTtzFW3MjuV0Yvrth7uaORhYACIPxG
JcG9DtGKpLlwf2YTxQ6myB5eFRFQR9deaXAwb8thWAlWjl3+U7zE3Jwk3WTTKN8h
cDs+mCUzo8EELWNmicoa9yjwpuMzzVs5L9nJxBKIwif0FHJmsziI88PNUVedIaMX
e8tipdJEgJek+yaXh96U6g+hWWlT4Nn7vtqiH+ySYLiNQlW/terjVv5jbZx8xiUu
5RvpCJMuO7Eg+nb77rZknvThJK/h2ya1IHCwPop0bZI69d3I8VynEEDl7AdCJ9sJ
sX/TDEiiuV0/leF1n7td95nlWxRVG7JxBPPmkoRyiUkEg7UGu6vAJL95as8GUmv5
0l5l8UpZUQuyHCKKjhoGJNqsMtHcAUZ38bckDT74cvQ8yoiZ4KEeimaFjd9fVUy2
LGfAnpJhck+Fa/08xVJ/x3mi0JzxWAqHeifrIXhSE7MUc+rkROU/R4H7xqAm4sbV
BKo71fxlx+UMc3RYXOv4YflVhD8nqKlxw9GIac/LCiW+EfPaJ/NI+VyS7KtFqEnG
aonU+dB8hqDrhiU+EMVXtGRBgnNi9D5B/hHaVRF1+n9rSAWqVglWvKADCKGMBzZ8
VgyL+vVLRIdE2AFEBqJZXYJsUskBfw5BP/TcJ1da2lwk05xCc/lq6leT2m0pzRoa
Ll+rZi1UQmTozRUm35GIv4O+6uv96H0uXHVt43PXpmHPSnURqad8TtfRJyV4qhNo
/vrctg7Z21Cnm3wKTgoOhkd1MkChga5rMnei1p/UO2YGKdPW69lsEel61GkYjOX0
DFLo4n2N0WJw8icU0EsR9qdLbWhjN6r5siiF8+k8Lr6VKtIcjYekCouZd9oV5pwL
ygUlqil80ZK/cm+j8Hrb9U8TbRJ7YvkKMo/PiNbKt+x0usuPrfuoU+Ykl+gXhdtg
F+2Alxhmr9GJHnWRH81cPAWPiRmBnhqgibS7tTcWTJXpFH9GFvrqp95+ntSsGYBa
lE2pdXgv6C35ek44TJRdWNkBjrA41H7wi5e/95Ug3C4rNxMMJ2r09lPqQz5948cV
X+6WnecszVbe/d3WDQ+PFAG+3eMx4LILmC5sDwcOOOoCM3mPZkh8G/lQ7TtSUijg
crabwcvxwYTVkDCOT/TOP86b/Ok+XQR1WyaJ0Onq1Vz4QN9aR9QXw/oe3Tzfex0B
oM43oLMR8OCZekGOh85KNrjxjEpgGAvztlrNK5v2RR+xLc4Z7jNZagAo9h10qAgR
j0DpvgGg9toGgw9G68HL43NTNwaoQ4kyb5PrxdKOUerSOU8tWYUnEqWLn5L6JM5A
W1DNRuv/x/ucXXHG4tEJL9ly9LJdRB1YOCHaY4CwRDgoNojPOZSBH1y2jY7Nyg9I
5Lf5PVnkAjFWWuQv9bfrvtPtsMujpt2ybHNnkY3rtWBgU2PO3Amf0Opw0Tu7Ira0
Ev6I9DCKF6R1/pX2/rwszVdbwZI6/Y/y/bBBSabWezlJ5MffjMvuIfwI3imcWzXz
M/10QgCJ016GvdIrdDpmFFpG//SqD2FiKFQc22ufC3QOxRaeqjTijfEdS4K568AT
661gQzqcKRpKO2FSmivoZaF6JoVB5FQ1GgT4df4wy08CyExZ1/pwp/KM9bzNxEqN
XtQb5SQ6/6th1OFJJ36AyYf9+3+HOX/RX37W1I5sjTCUD/3Y+zsJPmErsG7gViS7
bZQkne1T8dgcGiNgVFFSwKby5xlfMUlTPiGtitnQsAavFseUEljgDSRqikR+4HwC
yrSIrizmFtkd81SwUvVGwJdfZaZ2SDH9mHoxVzZi3vpMLFyocGOdvU9B+mSfTPsw
I12ss4R9CYhqPm5MZw3lTqlH3Of9933JLh7fR4JJbuPSqlH+OkaRXVaLsgi4hA0x
WGCsYkZzM7OkWErrGQTgxt4NnCvnO1DYnvy6frL/SnoVS94o2QSGkIi2MsE2IOFa
SI0a5K1SOB9pXV0Wwb3CNuVOL0AfHc55CmM+9rZ+I9/riuYmAPevN+voSUQkc/MS
CUpUS1z9dHfiQelpuv+nJdzY6xTdZBy6TF8Hf5mcwAvtNNMHgpKgb+wZUJhJbqqr
nd+018uF4uT0RNRwsPqtRLLDV1+K1UqxKms/8qu9B9tuuasACJ8f1huBfrgIsT12
W62e4ZOwm6M/aagoojuNAdoy0uTbLmkyzzZXaUTjChf9UqLIWuA9h5U8zpVuFyhF
evK0X/QVJo3YS9kRewxBaICrl4e+08c63ZO9jn1KGfClB+NLlYMSLehpq5r6YRdj
CHoyzW2UZr/OBxBLAkt8fF9ivVOmomMkk/xs1/k0vOo+fdRfhZiCO6cuzpc3SkfF
WB414bSznPH88lzcLRRCS6yDNsOpcfPEih6TYlotrsWua1GK4/lphtJd0p3PsmMX
XBgF8188I4j4XPoUgQ622TW8PkAf8vVT1tCYA168qL5LcYUXSPpDti87X7P0PH5B
m1EBFlJJsD3w2Zfzvhz8Poy9ilHMZ7PqBlfob4ZDvX1ECF6N9UuVEsnjeGAUBpAZ
irvnCzHKJsVBNIFdslrJ1yI/N9YvMP0voJHX/jemu8Jq9zf83Z2J0OecBxt2EN0n
G8NlZahv4A+Dvpkr6K9uLYWL6XQuP0yg5qGQCIoHmyUc3NTctTBFqAXXsfXnSJz/
SHzKB4aPpwwfKDhl1Qrj08jlwvV87EaQuKgy7dwmt1ZUQLaJebFE1YcrXCPVmWUw
nKAmQEz7z55Ac9tfgmHEEs8yF0iUMW86dqziYXuygCw6W31qDahD0natyYb1pW5p
fB9N+aBrIAAFC/dJBYyqkrV3HFZrGg43OrhsSiW5YnAd3peQ/UJaHEX9CTLODqAl
O4z3LZEkekDivTzfp3+Q1W4W4+/d8olYmdDAcjKTbnoK0kMQgaG73/tUvPdhqwuA
skRkhUxGbGh5H9/PzzopBuiRF6PtI862PiltX1sdcLPsczy9lRhn25sHZULtdFmH
0pv370oZoWE8N8On4rzFGNCdxZ9sWqn4RYLPHe2wHKqgUOravdeeywZhBrvqdBdN
9wUtD4wkFnRlPucrKu+B668DQAXzusebQFRJI3TtVScGKXsdgciAIYIaglrlUCsO
n90eyvoCiBT/Vc7P2jEOsoWm6HVvcQs4NPjoneAaB4mdz9UA5NX/sUO1AV3ahx2N
5rbbYfmpX7G7Qri6cKhK1xJGgrVkerK1NQyVsd1UFORlHomH3T1oTjtOdp4RYr5X
cst7YZifR5LuBZxBQ2IGgVxsnISSt/dIdg42NEByMVg/sWl/cv/2vyhIr7SOT52y
VXSkn+toTCIxybvldJQs1PVN4LOYUWerwSqhaP8IvigIg4ZKkYcu7SexAwkI2Sua
XlPOPNzfEEciI86W5HG1hhXIFLbg1/d0VxWuWGyLAq49+457Kg/RIVlZkLSn8AVq
OZYAZ1y+/n15O1GEVuF3Sbcj42G5Hg1NO+jJe5oSFr9Y2Hs1zLNlBVpiwzH+B65V
D5F5nhgIASXJ844SnKm6NN/0tWpiO02ojt1DJd97P9J1BOd3uKdnRWsM0alUwTYp
M85VVuh4W5MvwgGwYhQduw1tb7xr5/M54DIonWtsIZUdkGa+IgN9YnCkeYJlQLDL
T5oeWqqSfH2yBriw/4dj6wV80x69Rcuph8rNrjjjwkcuJKo1AuR70TpsjFApZegq
QpXAFvmDv92vr+LWTqWxMyOoL4zS43eyAuJM+CateiWb/576OnKDHocHKdqn8A6a
RXzo2DGz5F8NHM6FYZkvvQYGV76jcPS15qMcVOUV9zFwFLMeuDjRD41+MaEChzTk
GyElTaJDYU77nUI1tG7jvL8g8m8o3dB8iRNaH7PGd5paBbxZ5SlbDsyfarNJrOvd
l/IOO2L6wv0X5K8egwgvmOysmN72voXZQ2MRXgc5vCZKvhfvPX8Qvf88/H6GTNF1
+LCY44YXW3ENfjlaeI1MdjQBqBc3OJdZYa6+HP4aGYLotIvA/xujJ9RgLSvhaLx5
3jncubvlYrSgwF/yGiNmuBR2PyO4mfwSaHRLzEv7On/r7UQDXbJmcLKPyUr9J3TS
b630Fb1Rna+4sXMEhvT0DytF2ktv3wZN2jOwF6kgxn/Ba0hQX+azUxGBTok9suYy
2Z7kyPmOuJgV3BbqpbO05nFp2w6SMFOhSQLZjj3la45paYNhofGED447eisxfdoB
Pb2jp472M4qAh5mr+6RgFb1yHe6Z5o0GOj4DyPwU/Llw7u8aXc/SJLcrlJg+HK6b
1tx0xgC78bNuyKpzmSDHQfr7tXWEcUtDUaSDrJS+56kmtUoZEv4r3B4vNuEQ0Yh4
5broL2zwL/3Ld6S+c5ujCtg/7HTF1AOc8WQEDLIRvxkx9YW6VhRkE5iOhpuYm+3x
Q/IZUOpAvRH9y6qKm7EbqaLKrLutjS+Pnhop7/dh72hK3yImW0NnP1I4voI94Lob
2gl+wEmZ4tU2EhPzMb7TBfocRXcPFQxnfp86dJVZwreT+01o8znMgWK67nRm0Djw
6GF7nqOCNmqSK8yHr6W5kd1JVivUUVYHP5JOW2RM/sb8IRgwhomHNTgTXnpmqE29
y5CZPxt42XSyVmQkPcfRmi5+wn8T1+C6+z0jgHeUJ1M77fjF73gyoDcCQ3wZ8ZZV
X5SnmrT4K4uOpRNffEX0XJ2Cm2lpBCd5F3Yof7Xzc3lKuP/3o4KDhDo6oKhJBKDk
Q4t3IhmfT0y2tFdJr5WMNKHyXLtmca2bo/p+wW7MDg8xBbuNV0bfK3sK7yg37e5B
48wvjYmLEWprFGeCNIMgvDS56mv9KsPiKseTgonQxO+G8uWZqTdTfyZmgPSpKYAw
v9I9QWTuzdCLwQKIsFVqXhWUE8z4B5KeYu1GPFeQ61u+KqE1fpcTfX66ugiXGvEn
PxsI3DxpKhtBFhdon8MkVaOQufzNWboKs8f5TU6i+RIx9LIwqMh+/XYgqORgg/tc
uOuHVkX2IChICM5nJYZKcWo3qu4JvvE2PmUjqHS0OMT3Pa1y0ARjkz2U63+BmCGZ
pPpZJy2+JLRKm7HhBIX82liEDNJEbceSltIYkbXGJRhp87LLecuIUw9+X/YlwkmR
Y1pXkONyGOtpJ8BJVFlDEXVglT0Yf56aW0/2GnNpNMP3fIsusPATEslt0pe4UyAo
A98eG33yWD6YztFdWwWLcYXp8Nx/x5OvhY066rGLqBdc8bHR7KO5tX4bjBt4fMyy
F/yzQkTD98OXjN/qdzYgzNiMUoE8fTicn1hFMss1MCY+bFQCDv5D6/AHyhtaVX9C
7R5WwGszt9dYiKj9jchGue79RsyL0hT7eLERaYx/yiOHn+qCcIa4dpGRHae0o0LU
4gCJldLK8EyUiS7maoiHrbYgXBG6NZS5MzcbkdnWwJ3TCwuGXde8h5hJjdJ84X9w
T/fbDXnd69Nfizo0Pfb2uh5V45QyOtvJF5+/3EPUn1OY/pRpCMPdmrASsF7xn2Dv
WAENsyv93r0KjAMiylHLdo19co10/9W4CE30MdY1nKNUn1N64rZzXWrJXplLLQPE
VvlmMhY+uSVsiFq8JVA0AMSadgPEyEm51CM2eZ925xudvrnE8Cw79/kC43xyvEGS
TAzp3omxn/mmh8g4iqYrut4/eEbsAr+aJzyb/Y/yxHIOmxiWuDmdoBjYuTrusY1v
BzbZud7FU/P6jB57vFBro1QE83Xxl9a02JSmZPO82EHHiFYUSJsvv1bZ5LZeiDpv
uG+X719Y+xUaWdtFju2UqiN5XIkauUEsl4vY2ODut/oH2zpC7C89aAk9rymteoxm
54mY1wHHgyC4Hk9cpNVgwNrHr0MmMHVb+CuUxeeQF+68UhU8tXwfSKYtJlbdI/d+
FL9+Bj6n3ud/SQc1TlHSIu5q17JQOF/wOhClCf5cN1ael7VcN00nUhEtmiptVKaN
K68ciNiopavilI+6RQrJRYw3WcQ3mrvhGFzAuu+DZSAMx0BgTyVDlV7OPRwqwcSW
66OC9FgVzt49W75YFq5ry0mjtFLKEqWvebz8G/4z5ZL1BoyFjRd+tt8vihU7Fiii
lesUZztL/6KtX1d+yXjHHv3F+7wgoH5LHOKiGCmWoApOZLYrN778nWm+4WErsqf7
GgQ+GD8O4mvmi1fPbpEjtXK9EsPk6T+yWDBvZypR9Oj7tC9+eo2+WU3zez5fMhGp
iRO2WmEJOfRmsqGrzNapl5zTQSypJdB/23f4ww4BfescN8zyNaBsJxl0IQ/GvGwv
lVEOJQcKBROqZFpWDxJCsKgx83BQcNxSWDX8p6z+WADu1aGGO5yVsx1JAWqFQBBs
QilOMEMxg2OD43gceRx0oRpWerwCRNQDGsicV0Ed85GtieWvhqWRX1jpLhxjMrFE
zMwrmx79TnKbZA4YutD4vIQ98+Ht6t99MrtEcTrXb8CvERAoS7E7YKQTLPwttqVD
t0syHz4Fq90+gM79wSahaqmhH2MQn/KDL07WLrjXmJb7+7tWHqHuQ6kJYLxaXeqf
VNlV52c3n9St6kslbZ9QgtIt83FwbBjvH0d3v2oMoJxmo4C/iYe/rdjJjl6mV0gy
pZbpbJOk43en6SGKw8TdznraHi2S9BqCkOcXpmBpDNx76dmrUAY14jr8cbk8okiP
Mm3bC1ENeUl2dacrjElALORSmUDhfCv09h6NQ5UqM/mNl0vw8ZPC0yRoLBMFJxy+
D8E5NdMKrzLaVsIGMp52VI2x/b6Qf4xx07p1mfd1kMrfqdkPoXoewjMCMWi883jR
6gefVYYruxx0PFilQCgwiyor7Pvdfg4IBgTWNAUeCckMPmozqBWzgHq7r0XKhc42
yTFJbv+B63CSPKTHb/n9pNFckdhUaz6rlwrbea6shOzqtURxrXtgJMpfdopkuHc7
Q4DgCySGeadl0po8/MOwOtNDOKWYMBemwHUatxq0rV4Q1ksHy7RlbTX9nY3Lzrcn
bBS8ui2qSa4ia7PfexvhaMjK8Q49Elw/c/rGr1rIg37DS6OCaJ3s2XLECeUTbnfS
PM0SzbET7PXn/ZGn17zObMiAzR7/Mbh3cTzwMHoBxlyvK9NpjCZeyAdt+WSE64uS
u3CrRAskMjAqTfBJDklO9LFDYqNR0eQszXH03LAIOPOfaxuOYdETED9vJJrUmv4D
iyG08xH6epCqczQ5RPB5PVS7jziFdt2VbsJozX9tJE0o3o4BOeOVPaMaP+dJSR8n
OJXsnbupK2RZV3baE/vkaLl8JhVA9af5Fo0LixbsJoIKe+DhddyiCLY8xjb6ADAT
H1AECeKQ4Kvl4tMDjQT/DNSq+aiokqXyfbsHKLWe7P3/3arVv3qLNhIEW5SB2k5l
QblNKxNPq8MTi3efd0MVtdwoAOuQd6pW94KMPyoeMxeGwAKMb4Ascqz6V5HpL4EC
2RkxV9aLgbRpJp9CzIuBxS+rKFXrnzetfE2w+rtpkgpHY8h1YaMcAtebekw17AFo
lKZc9TcyLruLbt1LcufIyc9IIpnzDt5XG1ofdjxs0y8+SfSSN6e8en4ppSUj0Us0
WOfhCJUFbyh1wL3qQ1KqtpGM6FBYJxAvGFhi0ZBJrYjHJwIyTPAAs6tsLUi4klqJ
u0Gh6aqwf/uby0qhhBhubr1Vv35fW6C4SoLUTey1FWoTzL8uP2+jguXOZHhrt3Ic
Y8Lj4Z/hT8hniCoi9rEsAado1blNJn8WtwSLz9m4BXfDXcn1S8Hk4aN47QIY4APQ
w0tkWXSDhel0nBfoWFdVWViHwH4HXMB1NKoodSjyD49Y4e8sWGvFsafFTVbSaQWj
E9CgAeHnoYNvjMya1yt74JLvdg3QYtbf76dgpPpUVjPKpvU0X+OSy8tHLTxbyrto
nIsI186YqD4Zu0iB8OZ1qLsmj1VqUB/WcNwqlEefJJX8W79T6LTgyG6h40MfTYv6
/5/l13kYuY1r0UvTpasvS6xLuiKF5l4UXHeRxkgzb8txHU50nHwa+Eiq6kTHC9Hi
uQH+4P/PCU7hfXjYdZPR05czTKAp2bJZ3cyi9lzKuyc93vvKpRTWAYy0v7BCSVTC
ZJws9PVaOn6VlNnHR96EbkHPS3O9DA2iCuxCmuv1lHY+rel34nD4ICnxVXSTr9WE
/zJ8CumOQwqy3UWwp23bFmxPQvYTssQ+DsPtTkeWepMKOr0aKsJyiHnwxrSN1n6N
7YkwQS3frwXC8z4b/bdMhuzQnWo2ymSbARF/Z2cAm80jWvky/+mKfBceHw63Q5rl
S8rOC9+JB7fc/pfNPrspTYLxWxDCKd2hEnefwKLWoTPkJ/2k4oTf7lhn+6dQGylc
mSkMcpgyZXm3iBPoG6y82AgxKQiqA9u/cNY458JlT6K309ISf+1NMmTFZor3idA5
ct6Hn6LTfV6YCdRGB/r+YKxaqca5tJlYgBZLcBgdumIMr6/5VS94WPdjS1MWIVn+
KQzjeR5HAhZnwL3s7EXBTD1EhyA3n4lEiCbZTDGy98CN9aU+H1CXVkEHJcbOYKwe
lgZC5Zs8U8kagN0Sb3Z+pRaHUny0wy2oKap8cncxLx9sVX23pqGFnd2EbX0WEIcf
UHliOhL0JoQwy+Nt0x8RiNoHQBlgFoCcMtZH1jW64Ai51LdJCiO6wOFGbhZkBWVe
xyBPC4RrKpB9+6IZKBx4rUPZmNMm/9s47y1BTFtwjiKSZduabzxj9w7GgiABYYo7
dWwJOMhOCtezonjWYne4kllsuFDhGOxhdbi5ToeNBWNz3yv6cn9YE7uuEYpFv7GJ
PDwVGageX+yXRYQLMR+KeYKdOYBQq/N6on80ptT60g0CRr1arC5T7NOWrvh6Utgd
KPUT4ppOVQ73k3/EKjo0/PltHj7XLWj4QYwAGuQgq12n+MRpQ7sYEXkF/byjo3Qt
i//eClHdnDhTkdMWT/A9sYuMjjrf3wOQAv2PbCD6ZSwDyKKFwQgGXH7bAwvRqwJA
d/NE+4qzpmXNzzeqATHSCYPb5BFyf8j0QnT24FvKcMSyNcUtQpVEcRLGYorti+y+
HWM1JpiTgVMHjIhlf2RQxbPGGxZfXSQ9twyKR3w9n3D1qwCdFQ/wUNGeXISq+fKp
bc1hIBJDzl2+G6J7HRbeW8SIh+HwWA7MO0tLhkUv0xXA1kDrGLpNGkFaYIVS5CgG
Zsxe6stv/jPR4wTGI9/RcRvD5J51Fk/4CW37URDxhknqyE6ppTL4vQY0B9iR0Qwe
D4eOsO8LUNGZOMbOVdZ7rYbi6rqKmS0EN9XsvpLFr9YAVzTC63AqAnE7klqgyBvQ
r4xWfwGfyog95/w9mRm+VtjNX7UfebUjfZxHFZPv69We9ku4zHK/kh8xBRLTo9Qa
/2q4/kZ+6EITJkVJH4zKMZyD5GNH3rH+ZQAMXlNJqZ6QEoq+x4FLoZdEBta9/A30
CJBmf0vsoC381Ft4AwhtmF2riMFXcB3xQq7oLfaeRA7gM+4w1B6loAPlYWW0p2NI
Yqqfzy5L1GuNq66THRMmlWCb5pl9fFIH+HOSfVx3YV3Bbs652fRYeVaJKq2op4sm
GEmYLrcNesj+dFna/GtJ7WH4qpu20Cn8dM+1H1nLOvw8QQf1yX17sbjYNFI73HFP
YjLtGUkwl12LpxN2OOk2WCtuyNs4c5fNJI+oAvO4dbVlkZmeHGnNRlu3S2CDjwU4
7B2deZPQGzsqwwPP3040yQh0giN43HLq5QmaheOWim1RRmsuBZ4Szxd8ES9fEJMg
6rikC3YWSMk3/lyolWkDDMKPY33mShOfD4PO3Dn5P7CIMCefcVnh4NypKo4DbJaE
B1GpKQYyzzhYHQ4pURvjUghBX6i0pyq/d6EOZHpUSrg79lKknKdBI4FvMSPdobt4
jeZ+dSRqoF3VyECA+CagJJ/9K4NjBOpoktySxt3WSmOJxeU0NIUqwrJOvdnlQAQE
VLVCNOhzT/p6Ulk38ogdxvIyVsqGHtC6fN5v7F23oInOrMjUTyrdObWWrA3mT0if
iCjT+/QdosHQT5ynSysbs04xWY3TkF1u+J8ZYKmN1fiQbzVZNZ81SANOgxNayX0Z
r1T2e4wXfEK2/kXCxDeAK2Gev/5Vry/iQcRK5p7gJVFST0oTfLeToFpqnVXFMrq8
uYEVAD0Pu3e1gk865I1Jyqq5ViVUh19Tt3tBPypaxbXl5Zyfp5MH+oX9HqPMjmn/
XFm6t7RpBZMWwj6ToGVS783g/ymteX3puJU+fWOPDDQ/wxzef2xLnpf2NC94Hn4c
YuapvOv2ofJz638YQ3FLFp/R5uhZ5WWy7/8wCYM2nDkC0WsFIEaDOXV/OJ3rBnDx
KJDIzSdCh03dJvTvFIs13F/TanxsIg5Llq/JKNfcGTCHiutsR3aOYviK+6sW4hWp
mzmJ23lo0mpPnLLrOd0JIawEN63Y1TPGmxX5ocwzQay9hNTHIJBwk/45WDDCGDSV
O1DuximQGxQ3cs/pMzz6dvwdL60Hu0icy6wFBjyPA28qz0ZC+wRNHBCFXYH8YCLS
uV6t0o2lvXJxIHEWOjaoDTx7SiXTz+vmpBo3UhCxVi6zwNIBOyykwyg67X/E8KEx
MDBbbER3LRI0ww7Do4o7ePcSN/UR8+NTXpmAvRjwBbHDBSGe2PCV6brBPSOPCRCg
zgsB9COC1gqKHLsR4rpNkbzVCHD01U8DAQeYQPf/Esh0tuHJg64WNnHQnsACXshh
lQuzKG1M0oj/vGmFpO3XZ2ftBDaRE3kiqKePRIS2UdwT6qxvDzCsjwLrU50RoGbu
vV/mRluAMeqabfgPbgnHWuBQmDkVMVeJq9O3yT2zwOcsogUWsCOP9NHdxFvCw3h1
YsfIGrduEkRkesyxKqvnQvHJvO9LcyatUk6DneTC/i2GcC9meCOgtjeJuhULAKd1
JfDh+kzo9OUETGTcYpJZJR8YFMCo8M6wIC3Rc1D6n3ASe3nLtXzjp/jm/2HllWfp
W7gyFQ6yPnSRww3N3YqW1wJN2TpK4E3WMFgZd32xCMwNRaOINN8VpGcUFAP4DSCJ
Iul/1hvPtCfdoaLUZw1uzTYrDQu03H7xftxGrDmqbWJwFPxMuhPbujgyI7Af/4Wi
BPdwE3ClNohe7hzIxgXBl5xcgjvCfVtSoX0lSjpX2QaKKIpU6W1naPLVgXCvgtOq
1VWUf5mF+rLoraeqcujMVlaCUUetjTxQA+kdcNSir7t9Iw3K9vobApzrhmyQzdh6
ZXFKlPqukTSu0I0/QggqXrtL9v8as9Malwm74HTcCQL8ofRkJpxI3S0RMXAMZrL8
ld1PCMVZ6hWCBeIyQffNk6xRQ3FshR1uhAv5uXv8lcD/NdlEHacAnmlc0wsm6wQv
x3beq7de7iA329CEvKujy+RbWEOSi3Vpfg+D4oS4ii/hKp68g5UG1YvpE7VwyIqC
Z4qYXaBxjIdCDDJP4wFvgL1OIrENNdOoXScKqrIruvCDRr3pOBNxx6EER350IQ+c
MMfLNc+uxTJclD1B950FI9b+oSGWrgUsMfqV+yb8mGGZQzXRhvQKmSl87OuOz8m0
GsI1vSP5Af8ymcbZ+nXMMkme5vvUxNqLspp39wmcwrcedd6cFAJMgGrRwqiYTrAV
CMA0TTdJ6y9DzOlrOd+8WZFqggyMqldWJdUxlQQjqXHY+N+19aQem3/uCDbeS5j6
tKY85HFXsSZozXq1dlHaZPLbiLkYZBJW+8TgUOA32Ri7bsuovOgPOp4vOVGdWBDr
2TlBxMt1vfT9+ice4Wogh35g+BYiqXnDgMnfZ05DXqs8gucLV+9/brWgHgHwiU+G
sftXWO1A6RfHiIjPmP/4qq0w7x1OyWA4gNWhs23vVsLSwH6zZxAhOUkW7D5+4vKb
9QeFTgOpmUNwMBDVTzLmx+CzoCl/hjxLl6crwatuLAKFHfEcm5E6IoRhaxSERxUC
dmiPD63hfEp1sqNeX6bpi4DY7cikRvTBqT7ixaSh3DbiBg4ot3DCnIdmFR3iqduc
ZHJTbUcEVBypSjpjrIf3yodz/zbHHuSymW0tJ+qA7z53Xjpo/Er/PpMmdZtWPaIx
G3cFlfWN6CajbrKUhyHC8nP611kfGB0HjRYhWH5b8K/Dem6aVMY2Bnd50obvTCl2
xKj01HJcQDDjUNgNYG19Al23iNu5y/mllCQvH6KFG7embMxDJvTbXmsLeH6vuCdp
09nUTJ6uOSenQRBLmZ7h81ugqpQKbOdHo5lwlKJZDfkqfcGJtGgClalx/g5RvMRz
gm9ulJovUl36tmLIMySzjj/5zF/e9SklhqRILmNGccu0hg7AhXH5yNrqh2HJa7E9
JOcRxn5P0a8i1LoHxo5Hf3z8TCtqvmTdkERJVRSG3jDqjS0c2nRKGywZeu5yuvkg
hQuw5CtSs1f4InAqJaG1CMnN1M/AZ3ulK2cr9CDZwsvD015CNZZ0Ze9S2UhArXOk
IiGX+ka4yFgXwbjmofeItRzwRaaLnkDUXnxE6d2Yxsx+jJu0HS1eoqT9vIAeDlun
JhecDFXoNsQJRoB4aKTYMiCbHGNUgWB5zBZGVU++SvdoABPqZCi3Rx7VHFdKG6Ng
J6rdYoVQUOHbPAckmLklIuCmNueFSScYqBFg5jqkbSbt23NYW1OBg39xpaXPcRJH
3ao3U8o/z8T93d04nj0D0YrsgDGIGRuTwAadkoKFI7linvhR9T6LLWaL6Q6zugyF
R7UkxBFPzsDdobvTtoXuTcTomwr3iyUU5ntKCSxZSkzzevunniN9F29yiE9YLzLL
0UkvmcmEbDfE13BJ9Qblzs32iG3DurCuO5eKuIZjbAmzakMDnt9PRhz7XnJJ7N4C
ijendP7LLFICuzA6tKKf1Uge3Z5oKiljk/RN0UjN1MnZE8fu06t5mhXvcbdd366A
Ix3T4zmIoAyYF/gO54x2oYeS6OJyTKQFsLgfZ2/z02+KJHNhd4DeGtZm3ueAc9xA
4NAlOalBq6qt7jYJjm9s40IMbX8utZfK/p0QLngS7wJ4j/9T5lsJqQrRBf1qdPnF
CqsSKdNi/gJ4cK3MDSu0hSkdg5fG0vRsPm/4GdlXz4MMZ4hUPjq31hItzX4rlvyn
Y12MxAUC4NrHUVAndZpkVgV8L9GlX7NOxp7NvgUHMsNIiAYe7IHRJ99VKkMVbJYU
S0xBAT+D78k9Iw0xTA1NXY+5RrB79RGoyq7Oe6PNDyrnlplHE6OLklwpFcLJ9nzL
m3nEDdOAlIxTTWkogpvI2iKD69XVE/T8azeMZ06Kb8vjZaITWVXb+6AHHeNycTc3
e6cQIjX3JEeV4u0OKfC4l08oWaW8phoSZ4l3sAMDTGRSMF3lKdZTlYA0QkAkrvy2
9emc2AJ9ArJNhFsxGAtTNDEp6Hm1P7c/mRmbcMYDJJGtPR63k/Au0kGXlol/GTW0
oX4VbPjmKU1Fy2YCXfoZZltyU76XddwLtSj/M+yob16gre1QTK3/5S9KDfsJmB85
XzLrXgJ5+XMhgCZPxg193dnFzyCSndTH+EKpVXrXQ6tUF8YxerglBefvSxGkPNvm
RN7YP/LBDtS/DzCkYPptd+LXGpCpQ7FT47aATMWrPd7vZFsrJPoZk8iXRS1Nq8rp
GbEiuTqfY/4Gzf8gJ5rmzXESjknpkIlNvMsnVV3S7vd+vyku+AXiP49eIPsmLRyg
QU0hfuPDUQBqWvTJ+sqLdPIBQR0l95BCfFE7SfO2fX0fZrbBWoobiS/HVtq+0+Hv
gbLcnEMJaBEvA3rcEpOICw9wBqPjJ0sV+A6DA2wduOiQkUbrxP+yF0UnduXE8H+H
FTfr9BLVVMgDSDCI8V4mmnDQqS5w6kJbOb2Rpa6TH/IimfyWFjf5sK1Rfdt0ob5z
RigFuMqE/TjtuDyXVmkld9ZXSb99yjzype6ksCconNtwet4BxJU7jk7v8qkyJ+dS
9OJcky07GxS6erFGNTzBmsO4lYCOcDJzBgVuX+810NXLMLIjXhGW2ERaxbnyH5KB
jyPtq4JiN4rWVj7lMIQpsqQJwr8jMNgrKzTHDFBSjPqrs4wLWAl88KrTEBtESC2D
PntPLmZ67pGdgPhIKMIlabkGKS8QllcGS0fVt2EYWQpmweG9e0PTy15bKu+uVljb
TEHuPL0L2ziAul+Fp+oOX6q8IzG9u+YG0fDAtEPXKuygx38vAkwhk+82E6FfkObf
SZHJ7+bnYkklvjw1L01hy4Mh7ARgM/2h4le1+Ck9ez/lrHS2Yr+ErnwN3dZIF7cf
yatRm149CXlyWdstZxTZV0mrg/iDXnHkU9jza/VtsKpw61+bUrxe5MUOXNo1M9Ah
s/H6O66ZKI3hSktSO3rMPV+kwjyXFtXf/u4DzMCqrlD50pdJtObdvpNcuz7mU0aF
ReDW7XW01WbfIofTHLSJkgs5yHgp6fQisNQabrLvVNII4CC0j8pB/0GmAa2Zag4K
nNaVULt21jKD3OdyJamYiYhlbkJfsxTGM0MfC3Ira78dYTwDUclxaruq/XOe7ZnP
8Xtfls/OlqKA7QpErQ8/9TTZrxV/JsFYNcs+fIw+uPeR0z/RTXjMs/fPNyl9zWzP
EyBIFUpfX9iYtMI/1py2tpgdM5r4zofApfyXhsPPyxuc0V3M4uW0+o4YepjB6NqI
u2JdW33OxiShCYuxqru4A2bIrIrNmYBZwHvOeof5fasOVXy6l8JuOlQZc5sSUzxj
M05+poiA4zjwzL0qbift//xQqHk/34cA7GdVRqnkUuQ1shMp8Lx6PE0ecQz1tQjK
wzGc5sFcaq7/5v47d2ddVwB2WsJt/uHFkJ9S/t5ti4oqh1rr9dQbp+NhJ0IIp1PA
Dvbuf1SjsvzRdySeqvQE/65GTyFemQSdtmcqVuJaSFtgyxqNd31sAPiL6jRtf5Ca
8eAANr7c3H2+ktY3RYp6H6RAjn8MRWjZ8nDCPWb9dBzgxldvEbA7pFTubxwj0vd3
MW5rnSB2SeEPAjE/DpABA0yC/ov86moCE2+AE192DVnJdICMzp/bOPYH6S4YByRo
ccjLkmZbiK60lq73Q+3UaV69DJVlwC7Y21yGTnnrnqekXFb1JqjeyOo+Ldtsya+g
walCTLetheH+YLWjurBEdqIADxvlXVI6KKQP8lWG5IXKclubE7I6zw9gdNQnOuII
d/ZRrknxV4bD0zPRprVRYp5WzNCMb97CTvNwaJUcUw4EROAADQtBLSrcZtMDwYWD
0htjzUFtZL2AhZAKN3FF7vi3AlFDIRrJ1jvkwGedEHiL2maPRUHropc0xsOzjPyc
qhMZDToDq38BqqzLNXNpqRDMDQ1rOeeP8H4dggeZiUZdiRUhKufVWeaxz4f0RwpR
3lBGZ9MTdUHHeQ2Efhn5KOD27dSHrc5CJkuq9n1EazBrtqMSISFcRH4f3DXHi5qR
jD1PjwGUMGpqeZfVw+urtOTiCCrWR+8QWoW+iNxZEFGjgd7Z2WwbCrHTvtwqQWyC
D6H6CtDgDbsCao9j/mz6/2tvPctu3EFshrdw9t58H1RIWTl/fzTVC3oBUIrnka+z
gtVcItsvq6sF1PphSHSgdRPQMPGi+E2GNGe+FwcfsU4wILto9RFomh7XYAkNOhTv
Q1iVajTDf5MeFFqqYcQoVjDRAIkUuFJ2/yZtd5Q5xXDo16wCw0aRRjGcNYCRv7bL
UjmLGMpR+buwrYY7NUVcJvLnH50TOv6MvpOUy36HI0JdQX0ON6jnoBnTRDvbAA63
82sZS/zI8/Ez0HTDkT0N8PefuIfONzdkh02hRGehVySEXMUZUsGu8MD/gE3fQtlE
DbdJQl0q4j2nu9quigbjKR0pedDLK6+D6RzG1xkt8drhSB/4jHsRFs/mPJ8Nep86
8fZNLQqAVEcpf/YEShpzNfpOeRn+YRQgZhOIPM5OHgpH1hd7JXF8L1RzWsqyg4pL
If40bqWXfAHJTmJLvEeS1oAbVXg4wblrrMJ/WD6mApRcoaiCgYqWlFJuscBuFgiq
+mSy3tU90+di21D/Fe+StuQD6P0vvJ2Rv7nZzqtUCOhb1hKIeDDzIDt9NsO2cCCU
YZEXOhVLSo7ynkpe9MuZs8JpWPOee1LfHoR5FcJgB/ykARrVH/fCiKU7Aur38Wrh
9WvnXRPJc++EIDvUYFkwIJgRgaFb2Oeh3cMHDuIgkjrlCM5xOpXoxFmneFimGtQL
nwl6GkN4IOXUv0Bc5xaKJ5nz0t3juo08oNvx1RM+Kz+grThRkKldqSee6Skt/1ke
RkKmLG76/Q+xklZrZS9tyfKzF5b9D0MbO9YcogPXxojNOaFWnakWkVYMxLCaKqN8
8GOM+EP17y6C+Im3pO7aC8OVEwNdF3nSV2C+iRE5a254NB+nO97CWdQqzcqzP8V6
/KBYOMZ4SRaFSZgVQusJe60MoiWAIjxoIsWhJ7vA8ee5Dd4EI/htUFkpGpiDyvU3
Un/RS5hcPGd161DBLr3bwZeLX3X0+aKTXERswEKxX/ZyPsfKf4V+Rm/0IzAFlZ45
4hHjOAX+vqoQ8nSB0spaNFUXvkbG0z5mShgR4+EzSgxYnJjWyGpgkduuDBIJLplH
Eblzn1iCcm+YPgyuLQGGvdw7X0JLywGN6v9b/ttKWMtecslG5rxIjd2DHyKJJVQw
uktke3C4zntll1NRXVk0HqOMJOgW9jiXKMUh86SCkvgcuJcTXncFGvQQmNn0Wn+V
SH7F4nxUZE4LPclz8pQ9ktB6/+X8xh+BStPcpVBabHYt5LoEtjgy7qLWzj6jRVd3
JHCdh3wsE2Pjwej9c3lvKUPlWZducJXcqL56Rj71+QYqaWEZDxSBKsO0FPxwS1oG
7UP+Xq7b018rcM0d3/V2lYARm754TJPhJ574bzzq4xCPHvOTMqibMZWdAgIdat2N
i/FeZtTgl+k6n5+u4VNPnuCiQLkx4Y8TsY3jQ8y9Glgt8icky8LcWm7bflS+iNEi
LnZY1Bgc+6AICO1wmsVTNz3CU02YKpbDaAyy+mBJ5RF1T6XOwYLvKh/p09mDIz0E
+UJYO1ed23gWvra0bRR+s9FioRJQQRNkkK95+SWkyGjsguEIhqM5yoKpkoL8xIN0
pRj7oJeHEiMlPs9KF4xXUQWugU9P0j6WKDPMZe0QqpXUVpv6ltvqqhP5r4A890kY
ak/BAVn1/cPGqEAnW4CzVVok6Mx7L/SNC9AtxtE7K431m55jfgAv619yKhFZOssJ
Ws7P1Lz4YyPJtbWr1BVsbT24uOWgqffSm6nUStmtLF6m99ElAYWvhGPbg4Ga2H6n
idwgrZQvndKOCzcRylS9ls6ggDvMuZYWjxQIUhlUKUMrz1pA0xnC8SIcr0oAhjLB
HTU1V/qwNj44e/Cet0eFQN3OftfkHKj8vDiwpjYzp+t4AFdrUC/iBL9BNGTuoZZu
qFRAGNsKTult95c07VfOcZ02UKUoaSiYhzkdvhU9/NlwSeys9ydniPr0DbFzTdI8
ie8x89HraaP8XoEnOrduonTIO6MkLF5HgmyA5HPSVjotJH0qCljEsTxX6z7sq1mp
L+AeGxLMEqWclQ3YJ3hBD5ROWVY1Vqsm6kD+YnL/vOHtUydYaNBIF8cI5yDasrnO
7ckT2iitt1cfyj+k/fI7cEmB+F15i1ptdMcyDBc8EEKSxsn7z5dZ4tH193LXQ7is
u5SgDdqHMTdSb2tPPogPmX3ML2dPNzbAoDTkULAm+jtfVw15BM0C914ghwdpZb5r
CRAhjE9ug2B2Ps53AzXjrnBQFq1o+t0IB9d/eiepAhLVMZ/IqMRSzylwBPLrEWFh
WveyKZXYb+YGlxpAI1XjYGuxgP35acRNITOFYMvTb01Yx1E2rVyn9mDY1X2VIGdy
2XVYMuw+K5AExEQPLk2Q6IFkVwylf+vQTiQe0nl+VKVqxDO1qXUO2VBUS+ycdSsL
TmhbF0H7F6ZGAoSWaV3ydo/jNuu3so5B9zOytwXNsmBoznGb/IuNulRMOb8nYZn+
IZeXaYTqJq9yryBZH7ZJSCqSnH2SPlTD745elsBGw50yWoYftzh6pzS+ZqaMYbef
Wo7M3P9HDxO3G3laGQqfL/8kKzs59hWfDZBmWbYFELIWGUKdq/SpXRMaNimnRe52
mENQmuVUo0h6es0ta4gfxKV51DGgj/aTGIgkB2kf8l/Poj8tJM4Za/AFOSjPHkT7
f0ZD3d0C4MTTmRgrJANRWMOtULLfRXPprx43enC7YcwopE9YAqBkZwR1xJ50a/ZW
/nn0iUwnZCRwulUolacyQ43B4DWcbMs2u6HxD6D6VvaR2hpIux52rgdjt0z9n2Mx
eL6uckJSHXGkbAuYrTpulyL7pgar2BCpIZoorarGyxPH9mHL0VR2lDqZYziOwF8C
fdZwOKlOMBPg0S5puDg2/t3Tn6L4Q2xAc1Nj/rW9ty8ZTU1bv59FM78jWgM1KFax
AfWwjZxD6ZnfncFTTEX1BqZ73adawZJiiZ0D2o7XD3qJstClh9wJw0pWwp3Uzj1q
TO9RQ2KaukMBbJfnFFMFNfsqDA6xt85NKbzT56IESyLlVr1dNlChHGakWinzCv4b
IYG6nK/F5fUC7LmVOCiEqu3Zd3J7g63MF1kUSEk7JjjaZ0qkg/76S7zHdxwfCI6s
fDNDjxCbmIMR+MKc1dDcGYPyLtqg4ytYN+yQRL+IK3vqrR4kMdn8bQyudcpf3U4A
A52unWTU4ITmiwZYsxXxqDMcLBmP/Zll1EF5KMCyOwqKCpgdI8fzut9qMuo+YZ0c
bxJx5p5UJjRa3O2FVyVIrE71dGFpQh5HiDGVybXGLmHmLdK1aRfKgVO1JzgHKK0F
knPb3uSrNy8G4sjm7d9W4WIFBbeiB6Xv3xygyJJOl5izoVHJcz7KUZQ869ImJjy2
ZlzeINNnBr4PNpuVzbpwHV78TmMqNjfwCPhoY9hTyEGeYkycLbz8aWbqc89JKDiJ
AAHTYrGoNBuWuCKGiChX6NXMwrPQ6juNlsbetabNmOc4gMHpc59cJWhIBW8+zXDc
Kai5VySI/+QxXSpfq0riJapvFh79U5e4m2zh0LnaEdc2G531HX+wNA3bLnd+OhrJ
rSFFs13jK9QMfNGOJELqvHxJd0A0sRBSXEsf3u43OH8QkK2U34bluQWcG2Wc9RqM
WoClFJIlOngIScoATY3x9yLkmLJq3wjg5GC1yY5ogmWHv2Oxm34NLzKuuYe9jlmv
ARI8DLWyw7SnTx81vazZiwuepbAOM+JhVcc85ti7S+JoxCcDQvoh8bP8tDwhkLtC
pXzcbe9X+xCM5bTj4zDdlMmYTsCAvkeDTLfWspHvRHq3QY5yU903QEE7Z/kyad6P
cXvoNmx1g8zqAVrL23HDDeODxtHPhXM70ZH8Pmd8kVs9QG5Y0eBjbF0Jw2j7j25k
TeZbSQ9RzA/52/rv384Wi7P35fD6S+EL0iyb2bBx7F1zbygTLSeaagpzr87lNTmI
e7Dl56md0ow8yh9y0Ke+0QzXkTDOFtMbSH1b/WX2O4vHy8boQyRRGG5edAJbKacS
sr+4X8tZattZdab1t+9jk1k7EedXbwjZ7L4I38076EkzGI9K3wA0hg0ECZcKgWwW
W1BwjK0b9Oi6yXCJKZFs5/p4uuYSBoYMqyXaIzEGZ2idsnGnLWQFzyJttcelxk4p
eTzQrODDwoiNS6NU2pezNSau3g4sxpa0Iq5v5aD6hug4L1abXVftURjZ7/VG6Bgv
SZs5ct/G275kx0KfGztx1LqEpolHLD0ACUTm7svhWhHwSVbfeaCS2Q4Aipg36CxS
xxJKY69GBQ5qu6i1ty1IaFtcIIJfkuMc0PtGjmzhcX8gWXg8jcpUggAzd+/WEVi3
Q1OtquO038pOwCWFv1uaUgwKh8H84N3vkTzcDZAvD/TpMbI+4ABZ18twc5kD2SUY
SgKLLdYvrtFZs1nDwaTLPuxH7Buf1rpGrRFpq1Ja5+xLdUOd/HcHyYuoabaZ4sI7
hwGr7hy0mEDJSnHCKhoaC7iHGCuuIqJn7isXzHhQi5lGwJbRNnUMABUV4xRW5cl/
dmwofC9ru7Yo8t2uuADrgrrAdhXUeb5KGs0OxQq54FOvrB0iW5vOnHgnoJxzCchw
aPL3mgx2N5UP2i8ChuwjDLI3quLjEnGIba8n+41sivyo6By70Qr+0oiL9SQuxKGM
ixa9fhmEUvM6408rCbVQ2FJiXmmRK5fc5Tej3HoUQY/MjeFbtIH15Oqgvz3uLjMY
cNIgWwgMLVX/wyKT+2q84WGfySw5WqcAVFNs7V23NvYsxrBBF4TH8DY3OQp02B7G
G8364X28TLJKBgErXygtxp5QNhtt+0MdMcwAUkz/WH6chup+/WBh+gX+MiLLNMa4
NyJZsrarTTkBPf2EN7SRMA0OrhRhNvvseWRWxqTKHJXE4mIYgXJLvf5jM0zJ+/vv
R+mKCk13nQ4fLdM9k911Hrn5z07NSlBbcbsRXKeBRmyvyYstCMNcNHTYmj4KCMop
pW/R7baPPIR2uV4voMwyVpc8pnmLqemlGttp6W8FG5BkgULabZZ2NxprtT2dXYdb
j/8Z/bVC7MCZwaQvdr74SQmRCssyeQ0whC0FU15WR1thw9iHWYjbJX4fdnpNp4Q3
YGIX5ASs2xz9JmaTRyt6qJb32njwACw4+oUo6hFBTtMznPzLGkqHOFQtr7eG0VVZ
8IQg2e3KUG5P1hEfLUnWzKx7g3nhkA+kj+OONbEA8aXto84I9EmksJl0YARhHrLB
aVKytYThN/uz+vHaUG8uQMFTHlQ/WrmysX+5bmlfgOiHYUxPA1Qv2FQhy3JdjrbY
qbJ7422mnFp+Ut6r+Epb3t8eqbYWAVB3NIQ2SCMu31DACgW0zhJWB+qmcU7VIh9b
xhKfhfHtgf+VgMxQ83WgNgHENF3jbJ3Vu6WAkOCIm1GYBGKNqtT+ulo+ZkL+BPNX
8MLT4P4gp2EVYmBRpT0kEYtqrwonEHPDoRSbw06c2QqMQkDZRwKYIwYjR/MwwGXl
V08YT3a8UHXsZl7fmr12j9JRZ/WUhDdIg+PN4L65kfx3uGucqrggUZaStrpEGCPr
FWS3M01z/ajofWZzGN5zotXI5Ff3XVRivaH5P39SfCHyzx2bFl1zfG4hDzwTGT7D
v4e1pU7XkRfWxPGvYwi/9EKXiNlvRY0Ygs+Nfp3Z0ECYzyMtkFqW99gs9yZ/N8rY
KF9XKPLrk6va3lWflThpToJ6/985goHxV11nrmqeCLdH1StgqixTzKPv5ab0Xq25
QiE/4l1EfNR7tm//h3oOx+WElbxhcUn+QgNaUeGjPOGQlK7nurc2V6yrDdYAtFj2
KTTNw/JuCNEFhFU28eSSWUweylfPqm1GjJcHDjwd0A7ztGNYBRIFWyiSY06fyPJg
8vlsIEr+ehs0uHgrX9gmefP9aHHZ3cIrIg1nZPDOEjHZ9kKCihG87Ss33px5Zrc7
2JuwZIoq3sHts99TZsFfw43e6cqAWPYoeNASFsUA5nbmeAFfnM2cOw3/X8rno1T3
OIwMNnwP3wef01HFT+88isjPyceXhQ67cnVs1YBVyg7HiqRamaymdpXorzKKYvHM
zhdxm/XqQrobnrHy4r83Qzcv83WGBhTtHLfith7CDjm/cUOtTc4bnzJzzjpJ8v7W
GSw2YLorTWhRsaC7iuf9HZz+wJ88uOhmLMOG3N4qIiS8EgLm5rYOiyQAdENul32j
he+7TnayuFP+xMf8wOQiNvmg8dGIrz9nxcdZ4X1iaZtPbn/y7Cnj0SVy8L0isOar
PfXLoIIQlGkMtZnzUyXn/mvn1n0TXHnQeNfSdf4m0i+Vn+EeVcqV+UHYNNQPXx2x
d+UTkRfK6QWpGSfXVMl6H4Wm/0Eg8eP4eVq1BJPiYfRcZeMGI9Oh1O9Xd5u7NtQr
L0QJX96kDHnjbglC2LhhMYMo/8Jx/JK5ZASTZZT83gSW27cWB/ZoB/cc94UOZsVE
4BcbHgh138lRWJDgNnlkPcR+QNvJJUecnc6zbwZ+mJr8fdxJdlL+m6HfZrjgQvqD
mxBuIwLcMao2tnSsGqKP4Snur75nBPjfanmB2JZLsT9kShQotizwRF6eYXtEhh+r
tTSzVqHAN1RDJOPTPyEugfWbDRyhyph3/ysdhF6BPdLy20agVG3IJkLQhQ4a1jxH
UHh8URC1bXXRJwQfZMGljKwSvP3DIHamSCHIXZsItwKfhK/Gj21mkUAnxziwscyr
cYqSJw+Ewell0+b+npPB98pj0DAJJlv4Rr1HoFjNPoF4uh5XgW2gWnB+1mO/kaP3
l5SVL0ifdaNb7C75WT1DC5TfMZF6HMac8q+hN8bnTO8hydO8wfRsakPkbTGC6WrN
eX7+WVg/InbNgglJTjkiBZDjOCUe5fYe/6t7vCu5VXAE6kBBbhBUnI7Cur2LHu5l
1nI8ljKZyLQMLCLg9MhP8P+OGsmtq6PhDiplVex1ZiTWpHgtua6dI/bWFDt9ksVR
kj9QeylvVkkuBfdrEcSGXpyfuybr3rtZU6rfp2WM7QIDv3ftFVH4ys3J/0ClGshC
qsaJPHE492X6xBV3jBTA2C0W2sfgR79j5w1DOKKHNf2ZeIUslDOu7xZgX7HhXv0+
Z0zkQZXkrYAH9Ak6swwBFrPEgD9WRVkZABT+ZkvZif0Up0R5QK4KVBReC2wwI5v7
EaIeLMbPjn7nq8Njs3A+YgGSFOK3ae5WMnGwko7IfKjWwPTuAxG0VgvPc1TLuixL
GudNsR4XIc1KYGOHqtG9ORlcM1uoB848DbJZ7H8AhF+cgD+8rvFw8XIxRxFRLx03
0M18EZSujGlGVYeKKEjtGNby+LbJqr1IiQYIs/bhcPZ3kZHz5SAhCPeIVkYTskpU
+JxGLznUBDm0Ay2WtbjWkuMCxA7iauXOAdvA8HcP4KUmQ+tz3rglg2BkPW9gKxi1
e8h3ow4ekOJ2WJ/m3Asfg5OaMgeVdYbApb+i6+hDCDGy1+IxpYEQtmz1waxQVYn0
0Clj51BqlHHgUujrGVXeP1j1Gc/f+Q8p65HC1o2E/JJAMwSv9sziUiGsY2ZDptza
o33ky5cRX0722mG5DAfAbKLG6gx3RAc4TA0l40pq01o+EZ+G3u/LpD0rwxQ0gNQ9
M1qHzTtlbJ8UvKuZGLRvRUE5JW9P1h0weZDVW8PmY0G9S3u3iu6lf2+xnUnL+wxu
E81jjCG4dIMT/4FqrEntxkrrWyEtixjVECzR+kimKmQvb/ClZVRhxCRURnj+X3Vs
syaUn1BgWY6lsJJWzVWDZ1ST4cADT8mv/xok2H+cCXlipmq5OTdCC00GDe9WxqxM
6wGlSedukvePiuFLd23V1Qd4WW7hnQFU2dB+vQyhz3RMijICwZycTVs7601FiHCJ
ogDMJ60CkmyJRZoSOiTQruaVfKX+U3lJrkaCjBBMUJXNTWFpCaKnixrYdi91EQqh
ZNhpfaiT4POW3aiRgcCws1nllIey2Ame5Y63MLPV4skB6dEVZ3byi1qFvPQudQxb
IAbFYu8A8MYpPskqf1wKAzLHhYj2E41Lzc1h5cwve61mryxzNx6GvUs71YksDjSH
IUoICQ3QH2wzwAbFh+QvprmMtB+uegB+q7035E7TP2MWhQwu7/qBZ+aZ/sEniIwx
egth3BfTaHAu95rhm2oBf1jfqjHCmuxrltKiB3CoIDWWY6/ZWgitBhg+W6r+HIIR
dOaM81m8PGCcfedDYsQyU+mE3wpWEq1XE06x2kFY3kA/SRfzUiJN0vS8ZURbfxbg
hSMymAS9xSDgSSpb88Y0PHMdvPdN2OSt5PlfBeGBk5CYOZsgHwnK9c4cPmwwd5TT
qZP7xCSRSGzLCxC4PS9/UDX81llTzDM6l4MPb6cQm/iXPGHetHR+aqcwz5z0teW1
rl1xJ2SUiirMD0wWkbSqZjQYPGUGU96RFK+CXX2titW5KPiOdUWeBDoSh2ljsjBF
3ucWNqg8b6X4UZBPw98vGyb98rypT1oE3XdCYTdkjN83vK/srtedKMJZ8SfhZaBH
0wMaXbmkTlqxb8xjz4gAa9fm3dUSehDG5vh2kQbagg19ZCkkK4QDeqZSoPQPCQwn
V1kuYwKcksv9V1Y4DHMyQY6tk48ausa+b4QD3wRFdE1ExAEoAdbnHB+WGoVFLZ1S
hfVPFCpdccS+ZB6e/je+rxYodoN4XkXJW6ac/izJFSSkiPWhXzy7f6aVgfy0nYiP
u1i9+I4B+xK1kYb+mGnmNG8MpaVSjuJn5Gd8TLoPW3pcNLr+7LOwgFhAImjXWdIt
xkpfDaL/jxNf2G/wbwn4nc4ah94CU4CwQRQ3ivGLXqy6kzXBnEElvBB/L+/eImcA
C/lbAGUK/lC6+uPghyCZBrbDk2VJcVutlVQmEaypcKBQfWG7R599mS8cqpP7ajZR
9oB/Zelcv63znA+iqXTl0cJeaQxD8BF7ZDNPlxCdPZTs9MaCacOKSlAp7dbPa/MT
CKnPMZa5eH4V7tOOK7N34FNfWdz2BYlpcaCYeL5WVxDCEyq0oPK+KNZiHT/ZCSc6
9KeKJtegR+TdiZzxQSFaYmPRUefgAENCa/edoQxCMw2lc4eM0m9xe/wFWH2k4xoc
AKCFNBc8f7mC0akoc/kP8DUID3bohHbxHch4lJtK2kNJ8dZemquaxEgnRsyANSWT
/qcL7qpNRyr9jpG52y85p9r8IwrBLnVcU8sBH+JGc+GDA1hHrCNq/N8k3Dnz0vj4
pDNPFVxMGUTWD/mRLVO+5cIX2qtxmlP/oqOcaDrJUjC1RmQC5Cvjgoequ6U2HBSL
W5Sm+v3K99fDD5MAZ3UskpeYDRahIo5bL73GifzAubpF9f8dQ9sysCOvUJbmYCyf
P4JwaEvJ0ZRJPeFp+P63yvCQVtg4vzLsi77/aM5xj2gWuMHQQxqNlTxCulg4NWnB
vRClj6pcFESNkXC+X8mxsGRYqBfYhVN6225BQ+3/d+VaoFcoy+5AShPpG8JOHjbG
55rau63lBMS3ys0JGIkDR1nUWnGi1iCHFWDiez65xYL2iZcKIBrPLHgVJ2aAPGqx
J09B7WDB7uPUFqPlhT8vDCh1vGMNEE1qBdFoTJIpYxns3WKhbu8WAFKjKTNGjgbW
H0Z6VPrzmpHy9Vr8fbrTSDjxCQe/VSBKQbu8acR7jtx/n9qZoTl4GlRcHFvRj3CD
wjhz9HcXggkynXOkuMgippfc1KdJkEkTd/E10jHlVVXe6yHJFi9RzUvU4pgqhVWx
p/efFMlj3aC5vtkm1jNLsAc9ScvKrKm3PIjSrx0t/VA+ns2suylM3PCUZZLjJYnX
zbC2pEmfKYMuzjILmwSwFTU3IPoRgXiRMFSGm7cV1AkkRZF4P0aOcH62cHYwXNcP
RWSGDHbDvZKNRBQPoDJTRF0Btnfb5vLbA6lR6gklrv1fgmA1JYmvQa5zAmERL+TW
/vz0dZDqSBLsnshuEosO1OApvwAYEmY18jt8xIeD/MZO3+cEJwMJcWWm09JoJq1p
N7NIeHYPTBTaPGV0pcfYvTEKrKt0ymZ5ImU7eL4HF1SKCfXJDIq5XZHnUrIgqCeS
zz3zeO2JPKWhmJtKN8sRHebQwe3CfPgyWNnInqma3prlhj6hUZ6HxrdZhuSyTgKl
9rMK/Lr5hvpD9HJAMKCKZY/xMcodm8/iRuoIey50/oURZQc4FV+um4wa3surm+mG
3cNyz51WTQjeiqgnbhXAzjlA/108uy/uyUVABtUSXbuvXC2yBRoAzx2pvSCuV+t8
akfVzcSqpWFsjJk1IbPKKsvcHug4agfHFq8PODZF5Dl/8DH2oxHOnWweFzu+oZpd
UyytqLje0RSsaOh9JtNE+q1vrxbaBrtNAh2vBFryXpsIXjhVQtzwP+m3rYuFpOiE
tsYlnRSGtdKFrejlBywD0IXv0hzG0Ls1EVOpmcFZN9ObVWULZpPdwiTUZDaU39x2
wd5/+lYXDn5bKFHLqIZ+uosBq2/066Xrq8QSM4+gyMHaLeLumS3LydkRU0wS1emq
qJ/i/SKBcw66k7KmPtnbM5geqKg0HGT3R+zANJCMiry6K9ygreESzX8J4iEZqGsn
+NuBV3YLP3Qi4Hr+t1huW1qc2Mw9NhwRuyu1jKcMGqH8xJxPsfhtfOEOqwuYJC6a
4PoLwgmrwhoQef9DwkNBdzzP3XT1VYAPf/5UmKJtCLSFlff3XCzcW+NdemeeTF5O
HClqlp9lkz015XYq6tp6DQ8QfEFfyQx89dGRF44d2rEM1FjNHWz3JK9tqfgNNLGH
YTKQTFagY4ByqwzOHXB0ssp+hSBYFG5yEC4VU+caRfQ4uQUpfImYXjit+b8TnFGR
4/AP2o7FkFipdaI7p7IS/eqVzZJBvfxLbqLj2cC+pWubBt6DS58aE8wTnjHI9xhU
DezkZaozqmyxdzjivY+ThPzxTZOA9WYPC12kFnZaP68+96iGgT0yc6xQaWGP5CL9
LqdxtaZrNajINxvsQ5GnExl3RgezaNSpZNpdRD74sw8NLNbztf3W/4e5cW4sNkoU
cegOjMgDT1pX7VTk9+F2djQi/8aXii27PGfw3h785K3GKcn9usQ4Yq1Ukt4jQStC
LB6eUZ+gShdmAW7CbD7gjXZ+XAOcyaEDIllL9Ud4dTkq/zB5+/PyTQds6mKY8Mu7
TdQJD6Nhvjj50SobZY/yfRUCLUZRtNzMbM3suA/nWcrQzlVucVe8vSGLGp7A6iAo
f+V3YVh53cPL5n9Mi6S+DMVMYjfDm3Ckrj9crhevPo4PvFkIALe3RwyfbfOqouz9
9CQJEPJ1Xs/IfeJ5wFiCjenvh+M6Ykd2VZHoFdergJKz++VIhJGVnop4Bc5+Cavt
5Dlco1epfiUxlOjTCrysyjhzC1TePL33aT8lOumcOqvkTayw/lvg57OJfzY6py0K
h0NzNA4q2dyN3autONFw/dbRj0MO9njdw52ftCcJvOavpEuxyHhzBLvC5u86YzZk
N3BeHdpQUIh6+aW3PSnGypOscljJ1cfqKCWjrlyR50dfpDtRq0zLEsd/+qrguZ6i
yNRJ+ZAvUz9tBm4WhFlmA092c4IwQBMC7Ba7yrH1sEiR6AvYwa0KrtebJFEeKMbB
hIjtFEQa+irmAK3hVq31qVU0Qm8c8Nk3Mbf0Fedh5InP44qO9Qgh/8lcEFADHLRe
Oliwt+XaZ4aB+r0e4N88DSQRBhFjWzcMUTOd0+s0OgYZW8GI3BO2candVNG5U8Hy
FNHc5EmQY8h/EYlYR2XrOShvbvrXgXGjKYFx7JQNQCXBIobGGEOxepdCqNXtOvv1
434p/hB7wCPq02ZVOQWAqz53R3SaQhbGlavZ+V56ajZvmCdve/CWdn4NVRVzNSvJ
4Hajy7rZpQbB0huaCwiI4snjg1wDRXe2lv66U7oEhbPI2EU3NKvvd/suR5vJR8Br
+dABOo8z9RnfRLj07Hd2qruyMSvbhus4pIHFqSI59DtN/GqTiLVd2Cy3hirFLQPH
Ag4QNhPKwxl5brXfp1lT4jIbpN5W73l7BbqwP/5c3HegfQwWNmF2qialhEWOc9hE
jvtAn5d0/vmcNsLZdBxt4ITmBknZedNaSj1sycPCi3XBwbr+qNDCC0l8GA1P+r9p
m1+teN8Wtb+WE0VzPgHnDEuM+qsjEzaVG5sNS5159aR5rd/gkIvADZHkK6h5nzlR
Vg1XjdtZTr+K7StItZ7fZObPQUQcriTKS4iQUYdJqWoPy49ESyLg7Z/DrR5jjJtc
XeeEE4peGX172xB+NhrVzbpjQJoY42WtqkQTZZ156Y9G5+2bEcv7PD1R/8qg/enb
t8yHAVdNraQM7uCrO8i1eMEEbl22pRkcAHYST+zgaEZf/Qe2ADX/kakABEvGh3Iu
BZ6wp25IkoK08SeeRW3VX18XdvgdmM5lNXkhrBbNBscbssXkpe4ulxJx0EuVjg4Q
mMFrDVscOhFb7tslzqoHYKBkW6ibohlbKEYltQJG+0jy3sCb/vSusFcZKePkRM43
qnigc/4kYid64sPvIcdJZ/XwP7VDilBBX5GU61q12Hk27sR6WhhK8w4fi1huOVj6
0WnxdUHyZdO7AIPr6ShV/SSoc740zdvMPAVfb5uVcF6h3Ow5ChpdFROCWA9lQnOX
VseTPLAlgxZqFjxSicPTY0q3QddIl7pt8LZxf48FTCMTSMBPYc9KznzqqhvOj3RR
OJG9zrYsuxqZ8Kz3gWwj/885DIpbIOZGINljyuMa//dIMz2YsWIsbQiE0doPdVZw
ksOtGGH1wW6BIFXSg4keMwaIavMq9vcsL8gZlk5DbUI3mAd5KSrI/Z0BDa9ss9XD
ejYbe60vnSaxs3OR0qpfmhaFBylLeyuZ3h6Q+OoC0kQX2Ue9MzvOKm+8LV6fCwOH
hyrcqF/DgejuABE/xCZYOgLfM85X0Gz66bavt/TYdAkBEN1cwv7ZAUb2gXADsYBg
5Uv0fFUyktJ6oelck3zRPXSCLY8qbSL1OYZCz3xNqwvEk2gSy3EyZDkqeA7UTbkF
D69pxLcjVSg6EM3o5LPbvy7jqEuJZCtJ0goriI8JPX7V0PY3v6qL6tkAPs22QOb4
/ps7NNUs/B20buCJOskxE/daMEqPBPMlrQ4MHRraEOrVu3OKMSjB43mNrcAH8+75
h0AMYb89tAutKwJoqUaW/3dE3GdjaVmoN4krWhjIz5jwV9yKsCSUZ5K2poMOYV3u
qRJ9CPkFcXjrjsSrh+h/bjRQGq8sa15G53UlfWBEt04nrAMrcq9DyygJV9joEoD9
oqau3icvtYsx2Ty4hFc6inqTSnQdeN6ZejQaZDdgnjwjTlWDzZNg2XFP5zxqru3A
Hk5Qmp7y3ViA4Ue3TFhI3nXeXOFBi83CIHPFmewN9mUfRv3hDljqtcjsGxdTEMYU
fnoe1v5XfyZI5A4F70R7YH+3zSeEYE0H0IkrUrs4m5MpirIyF5RGOphtJttSYZyW
4Q+7oS5twCI6o4LypNRE4gyVR88BrqdmDnGarEqZgmyHJEFMI8UJyjayfeQ0q0+q
D5hdjYJttf8DjeMWsGyW4NE92CQCUknvS/JqtIrlEwF3eocM54wOIu2WTNogubOp
A20y/ZQV2mquupic4fWvECATM4fPT0kJ/OI8KgbLSGKA9g1wY6BrEo2Sm3nC0Nr5
yj/PuzUVW+gYgx4nB/YcapejXJnOH9JNu7Ia1MZxrBrNpuQZ9HkzIVhNSZOnQebg
0yqCEnYD8q739HRv/7+99j6/Tw/XOTuMjkpccu4ZIvBL00Y/G8WOMKpRy1Zn08EI
Tw+MUotPkIMwZEIn+gHFXeg6/FPfwywXgQav6eQDrNcZNyVdgoJNmYyQIqSQM1WT
Y5R2uScgFiKxGnqHmjSw6hivkrvv6issphlsBWU0vArDALj0VgarhG77qRItpEzt
9h0vPcSpqxi0WJ23pk2WKLCvUoQhogW2MtZuTwr01BvjTM5pRuR6G4AURs7QhRHy
lhxvf6BmOx8XPKZo10AC3wrXYL5tUz6BQkaHwk5PznXO7JanDqGWvf1E59a8x9VC
ifFxp1qgOSu+ehbSOOtceWMxuE2U3VHFDJ+4IwGEF337JKQdQ4JyZ2kyVzpFjc+x
6EQmqGE8VVLbaX47yq7ji+eO4s4oJ9rMin780JGNEWiO8me1Kik/igarawR+bG5H
K/GnYB3S+E/xmSD8PCkIx1YjBVxMBQhyJMOwh7tIugXUhjhmfItzp1bDHPmCgH0p
/yvTWISf8ZKVvgZuTbb7s6AHo9QDaPAl4ayD2I0tIQNQFSjrplWOsyr92AOUW8d9
my+0HTWAoTG+aTftTXhNCKtVzBJMZVUke1SMLsgsI0ERwPBWBZw/Ki1a+dYdJqfT
Mp+H1+1xZ9xQOPaN9ALOrzvvijMWTW8Fryg9tBWUmALLlalc1Wj7Kg35ie/zHU5t
L9m++YKGdoxvUyTrvyzLru6g02KVCtvOomQy9VW3VZlR8NXeHXNRAgugnCENieUK
iVyEyJXTG+U4Z0AMYv18scMuQNfohbmIsIAEgdKdqdAQ8x38YEKgK1553X4MMuqN
wvF8f3T5l+EMhS8vQ08Ewx9OaTsWssFI9KIZgu0IzqLCfjr18sjZENlgG/RqYlts
TGCIBn5WNq+tQgurhATwptqy3eSL0Nyx4hfB481CdZ/Qb8eWJGCdW7Y0+LcvOQkQ
OhLb+iBwlMF0lJr9rA/AsQsFNXrATn0aMx3J6jjKXXisifRfR9h5G9GseJwtyb2G
y5Lj63apDJJC58nyMMC7IDShkTegD3fhqfwoeItQfwrua3uDptJ6efVNjonhPyrX
KnMD1Rguds22YcVwikl7XRIfvUDeHVL6uG9m8gHDq7lzdQEn2fsb2r6gUNaUnbys
gVzjmE+0yeMBvmSmvTjfdMqDl+rUB+MKHJgJTvv8us0X1z3KzUpyn4IQly2FBv1s
1Dr9IjJqAF2hozfmEoDN8AqZPjuewr0qL6Wi9QQfxEiFtGMuNFXfvyvVBijwGDZu
fOao2BaZuK5uFDa+pyQUEKI2aSNYocRP6huEfoJ11ZDUefYRsLZSIa1JJi6ImVNK
dcKejwiMXdk01bpCf0KhX88Azc26zl+nXE+E3WV6hNpxUU/ptWw7blYd2+ZTvUwJ
zOc41SVtlGBF22aB0V2N65ZtHb1ovcaAKV5/kqjK2Vzfn0NS484Y2z0H9TZ5ttaQ
8GOfk44T71U6RPSI3M8U3KrCv1Vkt1sQDnqqh/RqCx00Fpk0QGBxPQXq/a3FQ7pb
5G9n0v8abMOdmPzi2No5/QJJS5YDPwhz9YHoXGUe8pyiicGoUsavLoALflm0JdUc
KTwEhQjkj4b21Z2wvQ7M00dV0evYjoOnOmPxV3ugKXYnAJJkBSnCzDdEgHqj03Cg
c1tMimPCVyS7f2PQ+G5yJH+ow+5t/lJwb0AS0ug6DXPQVsZBjr6T77iLsJ+7oNet
dNT8PqhGgtiM30gmxp/R7zuqlSfCisU1lgRLUAqpc5qQnoSwKiKlQn9jKE/PyWrr
YZQrLnoTqj8e0eQv2iEs96UyhdC/5I2M81g2IW2r+BovRyXERUOCJVTLtEY4S+lw
bB1C5rbaYgyKwviutAKzmPwEyeFqdCr9kQKdgQpleGG2ytMZ2qKxTK3kTKfgYKSe
aKRhoOH+bMvgdSAe3er5tfdYoZ4Xsbzs6ZbD+lesqBTv8Og1Hx5qwk4scKf2szOU
vuUPYddtpYRpYWKowzTH/W0nd+mQacoOzP9uLWfLpJicyQ2vRnnAa9AvOPCY3gGD
JGqBDhoDSBoAEI2PkH2P9s0v61BNvsZrqFKzlewvHFdWTLWVExFQy7ZAxI4bPAh1
krCSTaB12l6GcAzW15vNBgORj1F2xVsv5DxpJUY98dccdwVb1wpffhewaj/4tPYj
NFZ3P7l5tFVQ++63NS6U+0D52UUCWoERV1xkCASS2B/79xTe7pxAs1CZe6q1oMEX
ISPigKyVsAtlsUmy7bC11I3xhvFqVWVxTJJLMHXiBZKPt2gtlLhivxi8raLt8+VP
tr9fSms0Tjmqj1KZnwP46Hx9mGmnLQrjM/bw20FQYqw43l7mvBsXN6gWwwBseyr0
35z4aeFFv2NU0Hnz1x2v5BNA5jGTcGeKhte0imkiHyqEyN8Hf+LPXSaDppNDBqSo
k24c3kv2WDeDxIaPBCLiNCOtWy3kctXb10c1fy7e/PHXhTyOc2VTPryLQ3zqKgTP
za+J0roRKX5K9D63B2GIL3Zu6FfIHx8I8BP2H9yxxgzixvYnCKi/fp+voW57clBX
HjrNTyYWxykMfQEkAe4RyD3PoTYJtqvfWqVfDtwd4n1v+vrAQRuChbK0ufknFKaA
reanM7peMReoUi7/l+fLMVKOepk+14V6wDa83aU79qrRpIFsC+6Q6pQs0fxHvU9Z
UNJf1Lr/CWZfKbmAtXQiSQNW32Fsnc66IDJ1oCo2zI+cKkfE9qwD0UEGdH+08Au8
AToL9rDMBWm0+3phGdsf2XvAW2hJGhpQO3fWrbTtOQn4unSsnymGt6zV3FMXnczA
ciIPOyrH+sQFSUpKBrXd/hG/Dy69+lyg6Z/dG/jaJlHIWU6eVtoSpisR/ANeY51K
omG3wdwQBDhfMFOgpcreSseENSKS8EJ0SGkiwuKkr8KlSwperJq2zEMBpz+h647G
VMZ8atypvXIuxZELGlzx1nTCrBeEwY2Mvma4rOBIVy5BP8AYw8xIriEn8ys4xhso
t/i1kPLR/Oth9VRdelUPViZixTgc1BKIaATqa4oaV+VMszu7Icd74a/IcQ9iNaK/
ftOtv22141qlYgY9FQoI4AsmmZ1MtdPzzCH7hH3QjZsnwgO+9RGRkH4nv2l1JRFQ
RcCnmg/U9aMRF7MILngf4yZyW5loWs2WwqQN3QpxHCWi/z5lTIxjs4OL1YfPYazC
U9pLzgUl8+iBSxY26i/CUsUrG/X3dndearaOZAbm18w0jg+q4WI6lUzkmSFx5TqX
lYtNDp3UvxhgcM3mdaHa2GeJgXPF9dkdgYtliTebDx/ttyJQlXGcbTD00G2TkXxl
A74chUJUW7YOsjPSaLmHx4XI2WVNnKefVixBNjFt7B0zzwWHUOPS6Izyr0yw2AIB
SU7bVN8+Czk1pE9rNFYPj6UR5GkVgKxN1bPc9K9j2qXgOcVAjjuQWl0HCksfN4pP
praWZHQHVWitBfzs/3RXdClU0s8/01qDojXOQO9IFsXTzvJbgQkdus1mMoUL4ba4
AMmja6w22Zpm8G0QOiNw2j3ULoNvUBSmirsH6DxBN1KZhf/v4DaQsXESfeT/e1Cb
492HJ2MycO6GsakdintTQHt5eB/f/tD/UvMaOk/0WpWYaxVivUo3jx92kkDbJhbG
3rwZ8a/W0PUEBDDG39F3o7MT+UcwW0LeG+HPl4S/QXKrua/WN/zKZOWkWhzaSahQ
Mlv43cZywCA88dbO4HuvSzaaGaRGXtPWtMN9ZfvOv3xGg+tAR+KHmh7zcWX+9OkT
gwO4BY00tx+4POxbDM7e7VpBPZ+hPuJTcdKtKQyE1l+qTna6VfvyeBUeJO8JhD9x
KSKagGlDE1i8pu9AD9NjRcVgWle0iVvZ5hJEM36Bx11LGtFPqRKtoXoEPqp7MF7w
9yGuBH7yVmo8Q6PdrjE78wBRHbxeBijt5QCGJj/ti1q1A8OFR/UXXuRw3CCQwR19
/CY2RywwGOtyBs1kTSRpd83kxGuVdiENzyvLJxuxmpCfnoZvx0h8/KXthXTeJFzg
GiVkDUqKKfW4U2Fsexq3lrsek1rCODyNMZYKFjavCdJDJOamDTTSxUsFZTsAW6hE
sGzwjeQ+wh7lEQeS2OQB4S8SOvzZYQYqwYgeegL72Ohw7ep8or+gK7PnOo1MlILC
cncdHRVsAOqAD2tFkJaRdxJKLqZzcOjDIG99Uk4P5Tdm2HVkD/fa51XfIt4o3BVw
2twrvEXPCWIRcXbS5ZmPE73hC7tI0saT4dIb5O6As0Tse5r8z8RrTo5qQi5HXO+v
7+1+wO96g5ac5PYu98/QrkyHstNsafV7bCJoFDhO1jNeW/E/SYhaUaigBwRIiMv2
hF1XyHmAVQFm8J+4epFaWBMYiq4flUmX1QU74XbwnyqSkH+6DkfFAVZp6+aLsVMT
IuPhuUFl8bcXSaeKkbEKSH9LYuwYrJLf9gFQ9+/v3zUlOVo9PzzCqw5Z93VQyTY3
M6qQGoAD1ZdIeQ/iAcRRqFRGPYldRzflgyFAGTMw5z++GUARI5kONmzLA7xjyb7q
7d/juOMvuCaEL9s6wdNrB80sGsVAKlZw3Vg77KjvS70oCfHtYelIa2mVW5K3xxiz
9/nehU+FlthKcmRhYRkzcRDGkS/KGiIydv57Xn4Jvvf8sp0kj+o1teHkBzY6tO6r
Eu/Wa613WPJT9w+/iGXZ28YbEyFCU/SCWuVouzW3CBAtutNIxFMTEZ/35QjVdDBl
IjlX4QAAOjyYRV+Q/999E9hdscbmd6trfRrFRsbdgBZCCBLOUfeTkW30slpz48HF
HUAZLo9flCalKudOYoHEeuC8P4e8Za8iunAeWTavmwVq9NV0VgTbvMstf1JtGDK8
kMxe9x1bDSeqz3D1W2xXUCtZ96gWy2A2CeuwjD1bt9Dg/Ah+PFI/druhCgpAS07S
JD/h2fhuk2xD6z54YttHOkGOu2eqgPMhu9frYoZl2kRcYIozFpxR7PgotYvADO+T
cNXsDAPtGAJcRRmLfH4+x6mDFn9iTg9uX9gWgk0P7MAX8AbwZIAmyTzrKen+qXAc
hSMujONWBXSnkCR1e/gJ7OmqvXNFLROjceciYnHgwgt+llnqmQOgU+zKZAHPAqJl
OpJve5QSA6n1HD8XNUep+/BcXsLax48pwIJSeFheXFiRRddfyvKNxwrj/dGSaDKL
XQH/JmXCcS7AigmNBJ6lc4qjUR0wSAHZiZOzwffY/fqb2LAFurlTMBy0cOJ98lku
GmBXrdiiSc+yv2qL8Z6xWpMoKNbRhA7SN77S3k7iMseOwQGyPEL6N0iV9Qm2+M95
oe2Cw6DqmRs3DwQkZRAhE58O2mVEO3WOTll/R7bGtSB0+i1wMJB9w4qGr5HhuCXY
NwJCsXl3ugv3pgTXVEBClOe4P5slBnWmm4MP8b3/Gk27Vhrdcs14dHE5xIBuGAmZ
68Eoxu/Bto9k9xNul0ztbVf8IL4NqSpZWiLpGR/f6deI+X4qm7QPLQ99QoGsyAkE
fjUJDfWolMBZk54uF+0X9nxTXsNBIhUOCosyOYOnxa43g+X0QQ6wqG7C2K8b3Hn/
QsBLe4TupXN0X5BI8HETlknovBAR9+IJMgPPGKBxIX5LGlO1Xcs2hK33waZYpBlc
jLtZsS1JUk9GP3dl4bOlFfRtvi4SCvwiB3tnzbhD25srWFQtVVttXbaK6ZAFrMO5
ik9DtNdF3CjtWmj3HmmT9Sok9Zt5uTL73lf6kApW07LRSxi1SkzykUIPSXMQXlik
+eYgIIcbNMMqqQ0PpMuQAIsxXsgktMzkZtZUjBvW1+5qBX1r53P4USE7XDar/b3B
Rl6FRqPKuSqcmO8ZuV4tX/H9Re/bz1Kmgx2WVXlCmdUgT9nJgnRgORBTTk0Rs147
dtNvyO/0ji5QnIhBeO5Rd54KENcfqDh60v9wSUvEGUhfoWV+25vPlAVH6xssCBqZ
x1l/G/77TSvKP7JteUlLpYbg2upCm6/MbgI0i/rVYvwlAjemtdtPPwnwwOXPPe40
Y+gt8bYogh7ZbaEstZj2LewcKCL+tPa2+3pz662zE3qQlPy8lQHJeBOiy/miZet9
//jy1CVq0Fj/GXSb1AyM/8zxki7rOgNIVzJsJW3fAqt6uTbM8XwD3UzqRH62zX4b
HX6Z4lYFttFoDpxZLCIi1/ADTA7ykt0YluZVCd9rPMPgKqPyKJlZ8tHGpObgVQWT
rK4xCTV5Fr1NOMLOvH/XxRIB9Z6isp5/o8Ysylg9Sr6JMLUsYtoNIBXzoPXC9RBx
xwZl+c2DA1TcEYsqvWwq992fP/k8XyBvB3VEvBtcX6d4YKheNv8J1ifpro67s3fU
Rj/7HMsxeHVE2ysOKp6pwE4QS27cEONhcKXbgQ71ERFmvJ3TgiV2zQMSV47eEEVq
qjTcgLgZcCLWn2ujT1RYhbfwXAZwfyUxMkC4EHgqfwJhkOygHzq1lO2/MwH4FAB4
/c7zUFon7CsPuh7V+EsJQ+kL4dIGTvzNwZ3KWM4GXLSvj8RDsy7gJhbnbiUxp6lR
J5CRZFJan0FTSpXn8OGYGnknnUE08OZ/6t++vxnnu/k934NVFbwwPCwe3oreUZxO
8dFqXQwVhY22eZNvwF7ohuA7DmRlR60lJRn/mgaGNFpgAcbU2+no0mjsAgPW7gGp
s/Ok3QVHUiK29kYAMg/MLxe6FdQei9TEnl2wswn+Leq5QEfEf5AoqD/Xm2FdDifX
elra5CnijaJieuaDA/ioKyLIa3XNtBwqKBqXfSF/Xlprs/X658T1pJrYIRe1QmX6
CGg59LOmfFyK/5MGYcGSO1XvYTY1sUd424xA1iwStGlGYgyyo3hqL1jZCe0hwpIc
d5t3ljRJNTZsmUbr1v2qpRXrh+oCC9wUJG/l7lHSN+R2WeetlnjIrsipOBoF0Ep3
i24lWA+CBe3EqBuRsTCL8B6fPE1g8FyA6ViTvHzoJWqmm5CGPrnbqG3lLgZq9fnx
meP4KPaG82Ulm4F1W7T8ZP4Rxz3wb1OfSb4ZetozqKED+DOyh5roeIiY9UAz17+t
sLBtBbhwioS0c2VrxAfWx8XC9trVry6TLkmOOa9yXAROR27cKbg8VhdRZ+UkO5cR
VzsT03kL3KH6gmZYFLkfx4zwQC7wFEnJDhGRydKhfhPwNtSKH8mAHMhRP3OSw3UQ
O54p74HYFzVYdFNrn0hvoPW1WTYzne1RFZjvMAXBE9//PWajLtA1pfd2bVwvwQte
M1KScfOAv1Z6f0VLpDzyKeMNKm1sOGGV1gxJX1DiW34oKQPDtda1P+lP9A8EWDeY
tJcEitqs1aNEHmiV09tZVnvTKSjn+xazrmhu6XpFq1VxByQybICaT1KI62zpHQpK
FCXKXxaENiOZ/GqjPT5JcyRr9Gwt8isfAwl6QpBy21O28vUv4K0828iL+hSX1669
VyqtHWn3Au5bfP2zag/CGvGTqijlIYg/ltgvnXxe5GXc1kFElnzKiuRpLShWb2zL
HJR/q7FlEah+5ZNNqRHqQz+S2NNW0g9Ug7sPP89NItxAfF123vLAkOBUE6KdC6z6
gYdhghaBjs3EmhhA0uDrvSxjYWpl5RU2HcisV7DmccBz/+HEvY7tH9vrBStIslkd
bYdUfq6YrsLWXYYLHpAulkqQB8VAx0b+wEAWgSFh2uyDdMGTp9jjlsWBJIxkKi5u
qrXYaRW1P12+ctZEC7aMe6a4b6O4MUI/mO4kR6jGD0ilv+oN+WqCATf1rb+nCKAL
hdBbs25i5m/xmHJwzp8KyUEVTsBWGSNNswtURoVv6Z63o0EhG+p4TZgCnZb3SKnv
x2VHa+aVHFdIZErGXSgn0cFZv/HdscsmdkmbLxzG13Z9w2wmvHld7av01gwGcNFA
rV1q49x6sARSfXKqBb0KfC8Gm5QIf2EcEzgS2g4iMG0LUbgMHj/5ebOj71iREWdQ
SIPQMn756SEuhNkn4sHtS8WlGCpurrZLHNi8j6Q31ZjTJA/u6EdjqrjP1yFo5xLf
8FH/h1Zp+irPQYNRbeWUJNc6ALgBY21Shhaky0EMAbzWhYS9XrBL0PDrHwSQcoON
m65WbSsOp8aP5TQr7WqSq2qcJVeIDNO8BBHB5/0nrDMZOWitruYm9Zb2jVwGTBV9
wl+J4Rj4JXL2SdZyz1SXZ3e07aIqpbkgKY33q85qLG+WP+PSqwf8cMiZLA3qiPbt
9SbYiczLZufZ1vSOLqJvD6CaHZ9Ht28JZF5gp/ggt1tgLIVaPaes8fzTMFwmtQmY
VB3dvkF49s6N5nq+cBntEuteSP9tZ4lpD3oAGcVtxyv303684VLP31k+jB4+IBZs
AaohuMDkXGKOq8Yuk0WScN9Av/mca5hwcdnaM/3kgtGdA3Ju0SSzWpaoR3TFfuH5
d9KUCCnEyFNKnZUxRS3eFymWXXDxIbJmg2Kih5VmScilLdql4Ql8iLQfpq82ETcc
+f2/ydvRVN7g4gPfWR9FK/1AGIztvlZZxlRJksr3Mazp2/n0Jn9dZZ51uqWzHHnM
e5Ral+ZgCcIj4PVIV21M7makM/+eRbVlD8MrnwX1Jn/EQ9j2UJKcUImN5tny+Y2K
NW9ddZzg0XPv6Ohm2WSDy23oUQgD3QvVuN6KEjKDgVooZzGxkVTR9/tJ13fGsEQc
leRPo7sarA70SyX9eTKcVFEvpzEXcgp35gfkWabY8D1IIh38E1V4422MHE5mFu+2
kxqAbHynx+ZgktV3tSi3YpgtpEmI56TMI2xgluARIlkGjFj2ksVWtZS0nA9ZBvda
ISL5LzSJ0hE7soPZ5WyffP7th5dLTiPKy5k42wT6g5c0TVgfyz5A/Anfg4BbMiuf
oJTLREuQO/VGBKZaVfnJnGqaDTxps3ypjjMXPd9zi7AAA9jUIv7CbW3HYDPyJ8dH
vYmY54cnZ9mWTy0963OxUSPCa1F+3tstx8uAQqwTHlnFsLy2JWVrtjxDca62VsAu
RipfX1Dv0zReVxOYAdw2RcK/U+kzCFoZjObsggOVCkoCFFq2J8nrDK+IVGL1xQoH
k+LhVnjRGbfMGsL3MyMXb5rwRxgT2g+jXcxmi5XVK3w88uJV+qDSrQncTLeZ76fM
RKXOvXjSJAEsvINauLh1YQ/wxfIrYY3HBkXqPWCL2btBvAI7U2HBjtGRqwSBgktz
mKdx6SY8b0XdQHYLL//XO1AByVriFWysoeMYLV9n1T4U+aebSydQtf2OMRzxpipe
T9zdYz8kZAisp/mvGu3U+aZ5UBMhNK+n0nT3xSX5WjaZJqOiiqZu//JG80Rsh761
NI5iWeYWZJNrdwNUBGF9ciZ1z39n+BJUnyLPO16Awdfwd7d6pjAft/Umu05Mobpf
7s/VXD8zak9toJU8IKR+zX1ZwTDKuTwPZ4vnP+iB2sfJ0N7U906MECK2ysbwxDRd
L9tHEOraEkBDBG+XKb/s/1biMO2lZrLLaWhgNy2EdgxwqwpHm8VEFCqx4FRIPxQh
AvOMmd3W2yw4/VHXhWD668oEKqPfdwUOuFZbIDvmNm7K54CxCwFQ3YGpW3J7AEZ+
RDsKk3Yd0RZlxYK9jZfXv+uLixXFxnVBvkX5P3M+Y7OmaC3IeDljCiHeptnQLs5+
3i5/WYINz3UrRtelmTqslQOpUKB7zfieeKJotZ9aQ3ZYYHP2kewsL2MfCjePGACY
HOEYiVMo895XYak4J9MpsYBFdZ49x3laNfRyKELNpMP7d+9P5g/cbxTo3ltSz/do
XS0yzPqWfYfpFD79Y1/FEY/ODwlR/c89QegaOUOjp6ZQtQHvhHSeqdxIUAH3hDIa
Fqgi0ZKPNei3mFiMdzdmXf+0WTUB8aV8Xk9dLvuQlSf00maZIoeg7bnzuCuOYYy4
XubsJzQxCfmtsc3IVpdNbMFR2s20r2d8u+MR8WmGR0JqyrtQP/HIZdMIoZ7auvYV
0W3DwRG/Eu4Fdq4lOLqKwRLf2i/wA2LD2I2dHAvtMk96jjiDbAcCc7KbquCiFEuh
9CYMNq4RRdW1iwIaV5ZAUNkciTkcjjzHqsb+T4/1J83zyjpdJP131iMcWy2gi72z
FeEgFrdvnLiYGy+FxeOgt/jpIimNmW6+HGTDtoIZXGQ0qC2CdZxWI+dNMypMib6x
Of5NN95yyRadZ/EoZannXnYzfAF8tgC8YSQAn/2nqCvt85UIuy1O0Xtqxp5Q3cDp
D6IlmFZypRnwHVvFOd9RE0h45c3qFNAy6/n4nUcbnzYAreuDSAL6lsb/8SrQn8YY
wkHJCBciXM16eaD0StoIpXiLEKiAhqvL9ScKs5LwgPi1mJ/Hp/eTo799klBtGFZZ
d2O2LN2uyDyuv+kC5Q9Xd5EfqYUR+tOzPMTPY4fZJo/xg38CNu4XstY8C33Qu4MD
S2DEG37Fa0LMlg+sV+Z5hbUDUIbRtEMduFKEc/qDHhBqaDYKyNOTecungSuM/STG
lh23Ids49J6175GzVpOYVVWBDmTOHd+JZ5J3sx+O8qj3ljSxpSReUv+KdCQpvKbN
ocbboF4EPQ2oghsQYcUqLGKrO++0Q2agU2r3orq+gsKms8SdP77dHU4FvO8ienGn
A/OnXulR/I5XUJyQ/qTUKsLY0Ob0j4uDa7dNi9/4/pJa4S547gDb93Wbu7TjPawg
fs6pqCPOJXBbf1x/Z4zwcZ3DF0sHtefIsI3xDTmbX1kSAvd5oR77HvmI2mTVWxk8
EcxFq23HaeYHBXNsaaLSJ17o4RI1ZjzxFkwPafBJtq7K6JFHxt5E8Q5RYVHMYykN
n6MgIpGGyOw8sxu1tmnmqMlDRdMqf548TzJ8LV3Cx+GOddDYo5uYAv10EtG+Iphb
/4Sqc9bdOYPNMuJ09RHirT09As7lJwb60Min2TqTJav05R04GrKpBgDC+G0ugjlU
8WXxXbCAIqHMS2aYJOfVLm7f7EohlgEnQeyp2uqRwl/nRgryozdl49t9qUcaOtU0
7QM0PyrGEahUFNk851siTDHt8/lF+E+B4td91wwcj/VswxcFfF+jNXojEvNxtmnb
9mCBT08f/OOgi/MPbRctZnsAR+BlJfdZSvKwhyp0CkfceaTDVjflfQVHrUZKoc/n
u3LQYs1TlzvWJ+8mchO4tHaqZotu6JUKUaB4QviC39BBoO4LWipZwMGFVzZmu5Q4
WUPWK6AlhzDbaEJfcFKXPM7srctTYz4aHZ/wHWC9R8xmCYOLSJDZeszvNPUnoKVo
nRqyFWvd2z/4qwwBRd7HkgpP9r6gIt18g5QWE4DQsjqKGr1Uep9MSzGM3FVw9QEr
7WEti+BYH7QA9EGRslc4fBg0xf0TR2goaCM/wuIfbseJvfOBI0STLW/Akr6jpKgi
zFc2/A7Ti0yy9HtFHB7IcYhDivaSRqSe2KTLAhh53Bwj2owp+v56G/FNq8HRHfNo
1l/oJRTZGQE7mxyd5sEw+1LS/8l3kLBVtVoVVY8yYecNOSLB4IKl8IOUZUeJdwM/
nzf4K5VGXzxbfTi+2pRx7Edi5MVyzDkq8O3nRtz9sYDlfOtbu0j3KKvr6pq6M8EN
Dl1BLn59YY5iLBAiaRCbrx1vPH0YJvNHWNmGWGzJgowv6GyT12fGDwAaiILzsOco
oMFo7S2Gv5x20AzUaxaJXPTc3ScLZeP0NEr9Ztb4sD60d12+t8plziMylIUL4+/B
2ziCcBm7H6SjT+LQ9oLVnUugRuo9MVZ1huREN4Flg4CVR/xUB+IMJWnNlamyv4jZ
mHzoJ0H8Io8ECd7fviufVzPzRxson/R5DB0HhZqOLgGXLX/CMZ3V9S7lWgtso6g9
Pa/hIw+kekaZ10jjvcKwSafe01MCYncwXq+544qV/2bGbxn8rZOFygYqs43q+Lnn
D6DFzrW1khqvNF5/P5bxYsvDFYs9RrBlS2ZNZCwgyzbJAGmDMf7JHHuFnGz674fZ
/j8hGbjP0sv+1cfShASD5qXZwtP7gLmK98BMjoT0yGVAKUC8ktOLljNxHROxyXnx
LaRBXkypv6nek7e4yDzC3IXM8t8LTNUNH4rHKLRCVBs0waRkU9chaSHosDQpakfP
hcRB/Rx9tW/qRlHv8GMjgI9V3elL1D/VIu3AcGkeEjT+vzNXghSFnnoIqEFdApkh
Y8RuT0dudxvoG81sTkZYZC5p91iIbfyjkm5Mu6gllFMrkeq1T95Wgej2/BzaZTiJ
Saeoh9+LSJSW1Ld/G8nXjpPQmMAT8vB7BMdPYAHJYxPY3OGCYcCk4Bxxr1AhFwDo
vILN9yZ/5oP2BoaVXCARU+PJ14aumoU+Cb//X+kMV38efsXPSL8bha2wmrJvbGuV
PQdKcSva/nV1SHQCuyuNWCvDLyxwpBqiXo54DHGgRfLgi67sXxpgSGUBaumrYpo0
uELqo0eB35j7Jrwt/pXwf7qSo+MWFaFbiOeiokdBm2gV16pTF/n0aVtysbPWxIZm
QnGxnh0NfGoNLQIRBqVFRqIVrYEHqe/J7TGMGxnIh0JDhGZBWryl5zGw4XkR1Yx1
KcRN7LuJjsgJhWHqbXoWSd3XwVH4IvG2F9OWCjiAVuzxUzoIu8jj7XCXqns0czWq
GV9RHHOauj+XmTl04d+RVxXT7fYYp/M87lAmKphByw8RIDz7GLo9TLV1F/wJyyW6
nSoRFWKGGnLKKC7MOPoIxHXlw7jceacjAwYqvWi/78rHJFuqtGCPJ5TewQKJgVcP
fAmF0g8T4QlOtH/9ayQUNfqih0A8gqZLCTyK8Drw0YdtvKlUvsSGs/rUOkl6Zs4T
sjilTMfWktk0UJX2d643kgi2YVYOMoUKRtvq6C1Zrd21TtKW8uCV859+fMXCv53v
EN1M0E+fTw9Hj9jP99MfWggs/8/g0n+53llIgxJUliSwO3VK6SzI4rtJGljSYPwW
faQzUaZbmPlNLKpnpYCw4e0hFOJc8xvXgXFSd6nHKxCINc0fDkelUDHokR3bTKea
rSc314chwb+HbAXPGGSbUFnz5ry4CEpZwRtauWjITHARK2VGgZPuyj7H0vW49OK7
YwCdNMEK075e3dirL9E9ovLuk6J3xpp/dZxtIbzOQu0IiwCmvQyWDzfptpBfQFQ3
c4W6U9X/MRNDan4bx7pBrQu5jlPdwCj2BlQLXc6kni1qAB+AYyJx7s/pVyjm0fV9
YfZhoAU7qZCgMgm8qdoZoOud48JTF+iMlYGuUhIxndPEBy8/y5g5P1ck6slFMvrd
oRsRUzmpSplKyORxRaxVoHR/AunkJOfLRRcYE5Fymv3UNqeceesrDFDYg8OcIykr
c+gBcTyKRALwaCJYypoqmPI9rxwmbJeIIF3tBSXwCueHtpe8pMHtLXBPIo85NrC0
xqk9FjmZKYn8f2M7c5IYfJWzq5HH83kwFOgWnl0eu/Nw/y5YEmm0X77Cf/KtebQW
A5NfClbRpUZtE7St5HMiVBNoSKXZxIYUs6Intalm2NXIZpAju/ShbxxVMM6IHhke
+jikSlGqY0+xoHZAJik0gys0heQKpGxaV2D1XOfKzADJjEsPLbeqfEaHC9t/zW7U
nmjFAdVd8BbTTKsXyQ6u/nQjCovbs5hnf7TJ/Sdt2j/LCdnXPjeVXg8GubuvinxT
X+aIZbfUgzCpVS3TTkox0E0zMN+Ju8HeSq0hvNc92WMJI/+VKyCn7dbWfTo452Ol
W4/CD54h62j4P8M2Jmyro4VHsaIzPTL7mnPY7czs4xSq7q5EvxVSNBmV9BusRfRy
HKiftfRuwHcYGo8mH6j+w1jdfv22UO3uMdfkKt6EFsiNvegVvCg6IfcPm8Fq8gU4
gCxhTZk1MP7kLrBy/nXgtuhcJYIGPG211XgtPEnHLbpkOKkYF6+2kkMbdPH1DBsK
UCWQ+RBFF28GLXu1kpnVA8WrQ9MaNkm0m2DrvJFP55hH11C7U+fAtfygPo0WC/TX
HSmKWX8phwlGezvEA9JYFK25FB+O02kUJepmLr/7pXJODtWn1LFbYyid6jFQ1pq7
vsNiy6q2zh1fZjfdi0uyEq/lYUauAeru+jd1mUxgexPwfeJQf1Itv9owWO/wSzEg
LqgDv8pAQJDb4NDx/orRU8780TSe33NHayhjaL3jL7CbQcQDCRf2PucEc7yPn2cL
/4/CKZqMBDjhyPY+PxC0rlCBiydKQ5eyDens4h+e+ZlgJFgynPVqYgfhTgRK8RSO
7uCkM8bFxJ7z6ovzVzNaB+PjhPSU4+0QVgqBfto9iNMLpiHa80WRlWgTwigpScHW
Jkb8Y5JWMM4hn/SjZ4rmyK2w5Yl4drIyBwNpntV0hWsPj/gvAYLACvsTrabVIp7h
259z2Y9v5+zraKgI3N1+/6jHZA2PkUgEP4ZIplma4ctYh9P3kOA4OlnBwoK2uKLG
FwhsoBpkMpJlm8uIlor6sdZIdY/cUHdrEkXBJybmOPaQO+NOJPAQz+Se/15AvLIV
Hp6ZOwUPGq4N3KsBUStRzyIGUn/xbG6Rjgm45FNItyeQWVgjyfmuJ6GYkJ06hLpq
GL1dR9YO/2PNf3d6tNCtTzXPpgwL2IZBrzkd7J/NeKSS0Iuay4qXHDXZtYgjc77w
MNetxWcOHh5CiGCikqtynYoOnDox0gIgu+dw6myFub6YEIOBLYETjDvFR0Srio2U
gny9k7u8vvTu7XV4W2c5XPtGoPGlDWzrpDIrLdioHj3WlG3qI79pk+w6/HVtHjXR
S8jIPtKyWt15woagJzgR28yY81xdtMzR2lkY/X77FpmLo4mwOHDwcL/IXGlBp8x6
pbkyUHEee1ek7jYHYlADU6IaMCp+3nQSRzVN2jEttD0Cw2Sg5aOK1puUm3inSy+h
FAl1mcb3WYNVcoC43+LcZiAHuCXHc4E1vb4UHjb2fmenokYb6s/2NFouky/kHit1
pZAa8We2h8mWZm2tym0w3Id3iMQLUvbALbYC6eYCAOoTA8rw5/JoyI80hMgP1Pl4
I8PVj+S0tz4AOfK4d1epR66tVsE5vvddEMKlQGecsJbWg10yuZlLNb5SSl4l684G
8t2vhmQKsjFdxzNonFARoGXFKowg/jhS6Em2SJDljm5XvLTCXC12FYKDs5I1zQQN
NRKqPcDHM6p9BzuM6nVZuOXES1Paa5YloREQL3U/uFvheHN3PDLM9Re5p/to2V4c
SBoe56kk9KwID1MJ41WyBUFH0RSapUZE1RXqzChiSgDk42hjPtyWRMgz4fSnzskg
hYhNkQqZc1CaVZzOpYqnuGM+2gDnmJNdLkVF6FCYZC/CIIw3Ew/HH3Zvo+777U7a
6zW7ocN27dr4gZpxoP4AJqRgmkyMXphpErY97sOXrZ7diRwPPmbhu5Oyo865bb+h
YKvrlAx1Z7KRfPcnnD8sbeO58cofb+K3NxskeIGwfvTIDKIBvy4GydnEu7hk3f13
TVwjNMthQb5H4d43X14dBy0O2jAAmAecW0RyxmU0fzske/uZhKexoNlRAXFFXcNL
48RQYR33OvTJqmEtC/ZmOC6rmWlVfF3bOni5LsPt8OO4m4ecFJkQ7Y1ailgIRWY0
pr+P//hlIEaQ51LeSCtF0ckFSI8TumszMVnoLBf6uSf5eye2U0sIFSmKs01b2tZV
iy2LpREorYGKLxTuQ1NhdsNY9UvhNW08LMxqRVVdnilxlgmNeDKsvmN5BmRfJPnZ
2w1nPuXEPg93XjtBIPljmlcFZcnv0zbRBi5EHRtYnQndGvxZL22S20yoe7C3wmWR
mVQmI4yEYWFWWcbGZAgHA630WsW0MzBEpCuvu4kmzIkYuP0VV63Umsp5OMtIBNzX
EA2YhKXBMUrGfrJ/7onznLUf5CjUuC3CPScxepwQkCUTjPO7Kv24W2hCje0sa48L
sq0cgdy099Z9NCxgIPY/LCPB0x74D1YCHJPHVKn1wHJXNm0gkMGHHPR+b9M0pkZw
espv3T4lYEY3N3GB3jw5ZreQpYrBloBQCNt4lRGalfk7YbqYX8x6paftRH3odncr
mcpHKy8MY085Jipdl9cmTz/x5QqMhTSWKYeCrVPNiogFazJYl0LE7fL5OOhcI0qq
p6hIXjHzt4qt/1roju5NOZ0+Zf3EvUVOA8q+SI6M2V7JIsWR67VzZ3zQDfVXvkhY
IEk2YuRnJBgS7W6VUhxfzT84SPI9p2XPbUeTOSnN3w6MaQoGamLNs4rlPZKryqdG
mZ7bHbs6ji9heFYLEyLr1HvF2sdXtkYgW1jM3Px7nLI4vy/7I0LwNDXYuPZOEKwo
yxiFKbDMSVONtTa8s0BPHXGyjZtG+Y3ZDJiewL7bkioEmuRbwSl6oYIE6MVeLcbL
88rfrBinKnnWwWbIVjUlBnJ1m9jt8RNEHltyq4tJa1MfowCm2tMd5IwZlrdeLK6z
PAhKCDKqTHMZWzefywdXq1FsmeM4X52bVWfUQT5Y64MZoM6/YsM0stQYO7JNdrC6
RF/e6f4UmomOxhtaZRilUpIcnKyazY49Nro0OARd1nzI0bPFmhc40N6aw3er+zia
YgBWRV5GmxQ9E3ni3GiOtxenC/mhd+XzLMDfqIUR6iCldRv9mi5RSnbBAe+NMoVa
7h/Qvmokw3YGSdwA+8zLZoUAJFtJfiR3rqkR3JXXoFlSRUGbGGKStQKW3++DyEhk
ZF7RToaVq4w7ux7yKELK6dfs5mJlFJdgh+O4qcUb7dKeV/B8nAX5d8AMCK+FEXfY
XFdaefLqtn13NiBF1UQvc1AhCJ06e6LWiOAXi/gcfk0F+88ypBZ14FNv5EwlFr6R
CJenMYrQ+9BXZL9Q9eZ0ca8N+MygRQWYYV1l+ABLuo7+ON5dk8Aq6ifzLA73h7KT
H7G5jzOdL2uHgofhSA1uuPEgZrTtpwH1tccEKPVuzonOLUMQPvuj0joBcp+ElcbS
XLyy9XicW3K2KMMNE3Nm+UKTElrjy+mawPcwlEmdgDTIN8Z7r74PO9UuSGB4gOYa
fU/fOABcGh64UhIlU/qc/TtiOVatyrFJSSCgAdOPhOGTVrAh8BV9eNoqGQqPmzIO
3MkhtMQF06EBatiXUhD2OcDgl0oJD/+EhnDyft8y3reeCVIaPhT2UvID4cNk7y+I
uaX2eTLS8dGaWhJ8mNil1PNIkvaq7jgPyvDviFbsubFRWnuSg0u7kmC/uO7MzPPS
T2RgxyrNCWy1mxymqvDB+D75utLNBU96ji+rm6z9E87yT/IBEiObKsV61uh+HiUO
cayWzc0tGGoSiQyco1BdkxXqAVJXU98JhDLtBj+D396EBfcKW8ERmLuAA8B++pRp
pInGMPVGgFKJJtph949UC7O7cONaGq0/UCvCqbnNxQHQ8f7ZXKV4T9WwIJnyN9u9
YuuU+BWkDGX+CGMyzeJFY8ZRZ1Hb/CFOnPr+GriXsrOL104Kv5RY/QlsK+9UraRL
iCxwdAiQnFIM0XM2HYbjql5Mf49KueQI3QSWVSQmhdLWQd+5m5+Qts3mMVe39XBQ
BYJqQYkfxCIrZxZCkkMvcba5dGh97bk91QsOkJLkLAs3nu1tM23CkKmA8h3QEYAr
rMHYNLGhZ3m6pnvMfSFIj6XI3Pjonhlq4tGmM1Q+f9uvV3+dCBOfwOQeoQkss/wP
V1hYgJuxQ0BsqebHJTcS5g7eTrWTosASSOAviiFGCKOJyj6RoegkzkQXLhJmeALK
MgyTF0tadE29BUcldhAo/iVRBVc6/gauX5/LdG3ewhS+wxS7odWUoK18HA+v/5Jx
7mHsMgRfTrSckmdlkLnsH0k893nqrJuFgm888MrCodiP8mT5qthCBQVs2wzBJjM1
cDLQBcWuUJTjv9Hd20Lk5yASub1Hh3nzUchSIGAsvzV+s4u2BSY6cir24JVqHVb7
10RSDBE64U31U9PoFIJZF5yw5ofYHlIt9XpWrM+jaod6Cba5aIdB47OeHSt6Z7il
ijyxJfa8u9Qqd6zHqy61zKrqicyc7a9cqfqLbyMzrfywj3egmQshufAJaBIM9xjr
64AlDIu4xyfEKcxNjozfwwN0ScN+2os2NiKEjP/jxeAKKNOT5QHyDJXASKtFRscv
LAlcxG9yWe5FbbLvF7IEDJBpe+p30X4NSgUJdm4RgHvg1Yy9v5/ykkCPThL0Lj0b
7yM/0mRf3yU43K/nfhhQRIDBG9kaX5mNBkdEpHAx/jskX7aLkLdzLNEZaRddaG5Y
YTlrDXMjQDGWY44kLb/6PMy5/VguttyilN9H+XK45Aw2BRbrpop2G1iiMuImW/X3
2YBAGtO4TLmc532gbPGX5Yykj725h6vLh1yO9sfMq7pTefaRKwKyfe2NQkMbJBVx
SMZicJldm0Q+fq8b95RNMrsQzpr6TihyNlPTAzGZGh8/nM/rgU+t7zEOgFQHdAE6
oNBIKe99weV8tQrtOig13IURzmTZcqjWQAgNUe9D/vEy+uVLJjD1mRRa1MJF+ApX
9dInk0urMqnHK3l80PUp5Jo9cduN+RjkmKrKlZ1DPJPYNjYWqMb+NOc6EBuwBVLE
3RivsdMEq/bl2IILzuf4OYS1FVZ/ENaJwt5f82GLGT28X8r42EbWFyB1OdshWT9H
U/1Mw9KxRI/6Joih1YIZFPT7/qP38bBMGzL/7HitwJZ5k9Zh2c3JwLYgFbf+FB2k
ciBURR92t0KbjOGEi6vBK+oSQi+A2YK46hf9ebsdH4T42+1l1FmBlr3AQXUg+Q3C
oeiyxxXEhNyqS1UiJZnuUOHYByxnAB2Sz4k83bIib63vlbTxw8/d6YaxOVRUpUMu
Df4AcXlpbQu06b35MA5GbGpH46+Z8RY0d2G//a86A7tH4/zznAixkquBsGDqN5qQ
D4ISWwVAeUkZEvgV7CFNL64neMZvOyms4qsITDw6xlj5C1tD0UF9RtVPQqqXfINg
i0bTq4Jyoog0D+RYKwFOH3/7aR7+nJCNrb5ttuacNIzCEt9PcSK7gwchVY0KlF85
kYXOj6zGGKaDoWBDUWpxNXkYixRvcu19ImZeCWxO5KE6AxyeQVDVSU5IrMdYAPcF
J2P/VCv0qIu9UuPtsl/fCg85zM5JFGKciwYn1lTEvtjFma9otB8rapWvuqjSPl2Y
upZCbOGPg81dZqJdm9CC40+gaMaQIv/RF1n+O7mlzXJUgHmfZEu8T3akxm8G8eig
Hqr9c6JKIIin0zKKgWYAqrinKl2znqPd1Gl43l1AVu049eU6nKy80yhmm1qhgxqC
hyqtZgWuLYa+OURHmtAbzIrneupcqwbxg6X790NDa/mQ/szrgtpjk4iMlDeQdyIK
7jmJRWw3CZlKZENjKupj2ZdkS8NsAyga8dD0zo0qYsICByCp+5zOK3WKEPFtdtQS
6wSH8XdmaVQ8warsDQjcbvbKj0JebihXymcVr2rXFK0q4hv0/k1c+WP9M/DZQFE0
dDzu9gStjLAbTdPuY9AXF4q5sTzZWolWS7qRnP0ZzWHwtrMvchfg3OBqyNixKVjz
8GllKAtoshE7ZFqDgJuHJhUPBjJBt8stIGn9tbjXVTTKSFT9LXuY7lkxIrdMWsCk
f2OKDaZ8ygpUTveJNq+J1c5avKxvr+A7wxNvj7fMdAeWSxsuBBDQho0V09NnEHWd
nA2G9IdNjK4aua2WY98fnCKxg03jWVU0yFGzCIBWu9QQxCAM6pJamsSQdI3jVaYL
n3tgdCLugQ+9V1gW8hy+1eZzAsbDFz5DB1dAhM4gzcSbzHR1/z4P1VQ2R5B0V43u
K45/KWlJ3wZSXmSMqf7Nvg9cRdOJsMCSUVo09pjm0/ult7wsYHhnjanMDZ5rut/I
AUwqqYFo48bKX7TBEd3VXCgNz1fIz8hAbWNTzxVe33w8oTooYu7beADjT3w7oygi
GZijSiTlgjKSfNg2CAHvj50Xbnrz19z8004uTows/EYrKpZeNoZBdFpTuo1ueQ43
fufSC2WQBWShf1+DVuNQGXpgtLrbltLmlW8tvDxMi8FZjhfJT+RQzyTzKFeV5e18
kJoH/Q9T9dGnoF8CqXAgVYsuM97ctkpUyV0v2jwtVVktl1CpjdX/nbNGAx1Nw7zH
LSdWv4PW+j8zbJ78jNPKXycIVOxI1pRsdKhu57SM3MYu0xUVzEgLxQ3LT3rWtmok
zAYzzZgi7qyfdgKqNT6ys4QC6sA70W8CBSOM3TMH8ivPPUaXsGxfVaM1Xev9PJtS
6ucMjxgeW3S0tcq+LOAuarzUevCtHArkYuQlu1UGBkTOtz/cBvwxGvk+R51/bZi6
nw6/m57YXrMAGTlSvaYAG/r4FZfXWPSjhujaVtl5KCa3hjpnb0czXL/8ho9Vl0Xk
KEv6RkATGw+xsr9EiFf+/DFzXVJQ5LEfPx+WedQknThDCXj9Z6hwF29v0a+MYVin
Z4xD31ZTYSdYR+IX74nhfQu8g5s0IFH5fyuMYS0S20hdpsQaPVoTe/hjNaDW6g7B
WG5EUvpjyyD0mIwmQ2+UeuZRPoZ1CIL5VdIdU9b3gdtobKLkH3a+fyz1yG6Dh/7S
XEVjRqzx8JWHruT5gIzADoYe48zFw8YxFfJP89tx/eawXtctEIhno8GM0Nx+MMGp
4M+gd8B5QbXMi2zxYWDzsB1LxF/0r06wgPq0mDZODMAwgtJnCd8jzqcEheO6Vhas
Uwo8VDZ3NOZax0bS2YCLLnTUId+a6ZjpCqRhVrUnoOObd/Agl79qv4M+vvyfydY6
BSwEEuuttn6wZ4i9qOM5hz4PWQPCoLQSu2cwgW2ar9U/HEfeUOKt686jvvglqsck
lYAm1hY3CZ0iLAg0nc+jrNC72l72NgpFxfRJE/0FtSojyqS3XNA7xsHfyMcfXu3k
+QY79sb8B/I9ChdyWWf38RZjCh9pFUd5bx7k6sVYcpGe+S4M52BILL6d/0xc8d3T
w3j6H5ZFtNzP+eXxjYiIufuTKFkhCtQ3jTrY2E+5pUicGIA5g03wYa5J723Zzcua
X8Orwzckdhm/WC2nOk2pbWP90yEXNb+waiaL8d8Sd4V1UIl9t9G6ENhsL4pttEHu
WXBI7P+prrKCQnDzyex0JNrEmmqJqs4YXhRQsA7lzDHcFxyRXSFyjecH7BCZWTya
BUwCbiHixzarkkl4mSN2ZUM95uF5leY4Tc1Xdbkt1CN3zR8EXheeq2fgxPq6R3Kp
bjArbdrMxMDLv+4PZa6Q/QjVIy3jWwQkbHNm1ZW+Xx9WH63iqX6SKfH1YVH2tP8Y
cM5O3JDJsLez/YHT1YzlxdmswXLukGF2MgFmueP7RyhAjNC6MUTTbertiMs6l0fC
F/Mk+xHc8R2ybDlLa8VrCGLjtY/gJJnyvADe1syJl7XBtfS+cc1js1B17ClQX6JP
P3VL3PT/UbfUARUI5okJx474y1rDEPx3JGkvXeJcxjhbDYHtvQZVPew0vC2Miyv6
/bp1GXhmBmr7Ir7Ud8d0iKN00FqJ5WkNvq+xdIHn+QExAgaoHzj9gfhLTeRdS8vG
pBSlfeFezWakcLNI5IIIXll2nAmTwh/xx33IdB+2g1SqT2q7+OpxGhb4WORM36HJ
nnuMH1821Nz3izPDuHBYfq5n5fy2gO+h+zFIbGg2sZmdPVyUJgHp5PAP9IMWWb7Q
h5kAQQjL+uf1JlVdxZOBNe6fb2lI6rMmxJgsnxMKc65cfP6ijHyR8SDXcc5Vnl+w
wnndXGZx+2SaKZxEAT661K6SIVA+dRa9NKJh2BNP4G+4SW59iE5i9rxxuSzgUJHo
/O/o6NOKIM5hfZx18MIB0ghHheb0G6Opp1aqTLeINoIw7ZOFUFrE5j5JipDNrWTn
at2ifGomjils9tXJcU/3Z/eTQ2d4N1GNuUq9sd7XmEuWIi+rxSaavSHVGT8C69MZ
v+fSCKK+uaMXJFC3uKxCEJlPBzvzsb4UigoIFrkTWF9dNwzWWNMF+d8RSSr/NzG6
vjkOi1Ejt1cgfzVL5d9QHt7I4sbmvi5pWKwam/ZxMsgfx2Gqrsk8pT6EYF6Y3M8m
ETPhqbHqNc9sD8P/dqWuhQyAkLbM6uuirt5/Xc1F+pYGmB1SiqxsGnbCfLV/cVx5
6aSmeMKz1R9BIDqWSaFGXiN1n4GzNHelYv74KhS2ZULWSlC90mcFJEFthu/6BGzV
OTUnPRrjhd6Zmi0djIlIWmS6eJ5rkZo+PhLWW5fFfDeZkQ0uVyPB6/OtjKrBckR2
VCDHygEpM/oJL4WD2uoYNL3egpPbEUnqIwdZVYK0DOqJ4qFJxwkZr5YpNH350Mn1
tgLhbBlWUQz7ifu78AY1jakL4ucrJF+3bwzUkMHwNVx3jQ+42KxmdJbFExhHOq/g
zSN18pZO12Vgar0ONWK3Nt7ifOc4u5GJBObiK3oEZiYgyKEcT5RDsInsF9JVcDXI
tNpT5MboRrXi08VFFMbnFzJCIjMeAt6ZZzOyg31XR8Vv24XZH+oPffftkiMs3xu9
53zyNxxRDr/82x9wi4N4AhBwE+/yCTphUAmAwzm+4rLsKvieWbhp+lYo6XYbNnnq
ARz/pRzjfpxd92kL00S89Mg2pNAgvTHJzcmaAvax8VyODjLpDC5QMVgAr9o8J8NJ
BqcyYM/lbZ+sBu0d98j/s3nAYTGm54ZSR0iIJ/XdIFzbdg/CaSMhAjTI6QffFcSg
zfNFhPbjJdhrxPTpHO6W8ABSn1HzSgvwrJTEsVA888tfSscS1CwNre+VMXxKIB1z
AeZgXyZaRDIh4NzsiuTdhdStfm1NLspHEbzxOzOinWupeALpulkY6rvUsCsFwtV+
qtQD919bkv7mX1KXSnihlwrJRaC2+rlC0ZKsifFA7xN4qW/3tJtRZCHxkRY87KgT
lmCZW/8LEjmnO0lK5OmZrmNxD7Q2DiZ+a2WULPddgpRmDfxSVEr1hbWkhcbldEQn
9iBfikPXWRWe4oQGxXj8NjxR0nRIgYyi5UNEVfaFU5xM71U3k0n6yVyMS92g9kdc
StjBBthwqtpryxIBtHZMHmaoAobzrPrQvkd1l0YS8GgbwcbOPVuPoFKvAYVogNox
EWlcKVu7kadd5gt7sfwP0E+cagZCJ49SFunje3MhpejshJW+Fw1U3tENPI8e9uTL
L9pvRj9NG17D1ydH6lxZ+igDlEj/OywXgww0fo51zBoK+oA91OM4E0+8je1EHfsR
wzTAmOtTJG8A7c2Fr8T/BfqquBqX7vcauWV/+jIK3RaBfFQchMQhhJE9U0KEnsLY
LZnw8kYh3qZbfVprHfJa8phKDYQzcM6Xs/Ki+T8c+IYVJXB9hneSraolLApULt/4
j0KrqnirR9/fQy2I55P2C8FKONIKDDC9ph/CnM7lf/uqnWgf/qenD+R9+hwDV2fB
YJ+BpZCSZxHWRX/cG8scj45Svrgi3IiMP83WMxssLhtya/8LsdGTifiBC4lyBzLc
eVFPLa6VDWbS8nXu8EfqpA7apaZyaf3jTCGaThpXoV5FdBnGVGle5a6rdYl1B4yc
dKFzI9wpBPNANifF+gIWPIGvO/NqXYRDYn9b9ZfnsFN1fQGH/zucvy5Ta4q5Fu9E
LheCuOCVreS00uesHSoddvmYbbo69ze9ymOsuBToeuFeHhAkiLAgCw4EdcZbsuql
8bebPe1u9xpl07QWeuiVUFO+jNCJOvaNEeryAlk83WQ8vUyHmsB/8zZsgsPLZBga
VumLGmXhYhzbCLPMHc8J5aa9+vIwro1UbCzp1XJKlfU5P1oigyQU+WU87FQMvtfH
uVrXQb4vYPgEgULC93/J9Hub5X/OfuluwbdFjRcRqyyqOgWn4PTFQBrsKlYj7J9c
4yIneHObd8nyUtp9HUM/hV6enmSKuxjQ2W5rmKZ9TZKo/vNtUgQgoPILtsqyOpEb
+ZXeNy9F+nkw6OaSZjASpC/ngCYG5ydI3Qxfte0xlO52sMnbzGbIx2rZPxO0lflP
+hd7xWDNoLQ6CvyZlHuwD/Fy+3q4KWDQFyzNDbAsaGezlKLfH2+ngA+zh4YD8XUt
dhIbXv+I1gNBbb/IIeIAy+gMX4fSyIJJgkOZ6s2NfXb/8mRKaCUpkyniqIH+yTKd
4TOE4vl0SVdDmjfDo6S766hpcJYSgwW6k/Epyx6sGUMhLoDaLfwoIxRfYXL69qgL
+o0x/FlgpK8rgnnx0oVn78T5YJkDj6YykOTLNGWoRtgOdQzrQUK8e963l0uyvm89
MVeMLku8OqrESq1Rh9w8mJki7iZP5o8HXQxqN3CtTmq91vhfgodanmpuYr5TC2SR
vxSzxwTecLQbYLXdBOL500mXmsFlCq4HUbQS6veGQdfl1LUxzQmCWoGNyil0vSVH
2OGVkLig/jRCK+l7pepskbu5JG+VNXv9q4sTTkWt5Hqs8oEjpEzaJ8Q1xkZKFIwC
xfoEh7kF0yn2q2FYVzdktuScAn7Q5zb4/DVDAWPk0lkeKh28joF9fEWn2ST2DWcq
VlkAD2z7XOZh4RUN+p+cLSlOsJYFjwN+J7iuwm+zfgkufvxHlYOVmJWpzwpIkZ8r
tqpXKbdg6inWTpWSVoFQ/jrs2Dk6M4rJYstUa1Eb628MgYklSycWzzXa2hM7r73B
lCleuZ/frfYpMxJCjbtGhNqY26zHjVkqaKnU6sluJorFHDSD/zshXsO6J/TOEV0v
zhrAs1GC5YpMF4/EEx4wd+T3VyhOfxoSKfCwK7u3kOILdKlwVI9QvsUnNHKBn1Zs
gdg3MBfhAo/7JKkf1ePi5vRU0S8OkOBJhIK+5+fOcb63JB6kM394gu1/DlU+9czb
k9wpaKh2NYXVzEo9RhTJ/Z0ZgMU/Xi6wy/AzT1Oh0Yi7XNSGiuBA2C01VQxZKb1f
eZkoHXCuqhz2Xe2Y4oVzk9zMr4AlHvg9jS8G+QBr88n+HXGWR9Pcju5iALhb5ns4
K20gupeDg7iLuXYrOx8q+WP7tYDpu82oVwdG08/KyJh4gOtE5G8Us67DaDOH9CwF
8v06c4bFW891Kenxyhff4CeGmRu9lTsoi/kKIjjNM1VqJzbxtYF44XkrOgaCFqLO
Y1drxeVflLc94N9JPAu0f1QIbhB3DF+q2CJJMfM0L/BVSBrFk5dBtd2RdMrTj2z0
EQoLix8x/TC9COFeivPMezGcVgV6WvnUQu/3iAmKz54oaOjV8KzOyg3nnaRyawUk
SwjZHeeb5/OHNUSuefhv2cE27M1Yab08gGyyJaIPsVVSK9ffTvTEVkL53gtyxCp2
L5nuRv/K6uPY3xKEYUclPRNXfuHNYfSUnG/HEJKzKZ+6aeD1NkoxrRxNoV3Hv5VT
XODxmLcdy3QmiZ8KN2VxqQVKJdMsGKFbNPAZDuOjahimUSPZVEXcrZNDdQz6q5z/
QQ9XoPSNTY8KEskvd4i/J76FBSAyRnpA5Ju2Tb9UfzWQEeTMk/s1G665/CkttNxH
uvpaT3r0Fj6eSfpaKeOXAR+TpykeHm3iuz/FZuHtSjncZUBs2MLm3d0RmvCBLT2n
W3oT//3/twmDi4RNpwtj+oS1RpRpZWPn1kjMBrNptBGvniGNQnnHb/eAqddMMu8O
NBz1uvScBHbc23Jkijrm9UYAqc3k/N+Iheem69xAkSUAwH78sdPhp3vkbvcJta1x
PanjmV8pzfBEH8oQ0iAsVIMO2IDzK2lQfh93zkA2ms23rEfuAJuyfIUp2se5bThz
JShmrRWY3iDOsMxNUgPyURDq9RBuE1Nuosp5vCIH38RZXq0IX2Mf5qp+IqEqtUyN
4hVbuBvSBF+Y7vS4S6kITeHds3jyokzDkhaXJfFnJ4vt/UoqIN3eC9isU7AMWyfn
/zRLn2PNQNK9O41C3imJ0B30W4EahgIBaPYcA64CARV4pdBwElghXLUttbuZXJSE
V0PoSYNse3zWojnRCkjRuOgE6hwt9pLccBCwmFiNLIjiELwo9AHLhvfPyQVqoxul
CtQQI75Z1vcZBeKxB0fXJw9ngp8tLE5OTQ4j6PpNNpynuvIeKS+4/9mOFTfLXCBy
sE4XoyktuFJ918qF0tZkZpY+wRCfIo950xzAHVklC4EgKVhq/0Lpb5NBwNmGGPX6
zKkfWY+J1dWGvpy0y0OBIRUzGJb5LFepD3nMObef6xtCS9LmDaLnSBk//3hEXLJ1
C8LXDgGQ2IO9qlPGWAFifoe9gj97kdc2QXn2llnrtJqHMjgPOm7vXkZj0T4eyG0F
UKT/TwtMN+cO6yxeSQMAbSXVk6D9AKWPiyIZTU2UmLfkdDvWDuHlj/vOi07MU7ir
VviaugAyJ+PBICZsA4V4lRBQDQ5BAd+ESnCx4PwuELj64W17iIDlV++C1qcf+LVs
ZcJUQ2DuShSiRCMNPXENivI02cL0A3syN/foYg34VCYiNuSYNUsJiY7FjzSewXVx
3JuNVwkjGVtM4llfSNQaqXpE+P3zLsWKgAu3GHggpCrSNyenEESomtGVtXzSJphA
LnCoU9XMYIDZ21bsyNZvR8fdYjGwdI/Ftg4u5r2u/obqQ7pPrRMS00mhA0/7f6Ji
jc0vdl8Dv2/Bew9rhspkvX9JvcSfMFvHj/Gyg7Mcup+pWMcfB55JLXGxuJabejoy
vPaVzn8xhPcvtniJCxwgliZ4PBNQbvKVPmslDTXlE3rwYAp7UBlkoqf3nCGd8zND
An8CTYz76XQw2j2mHtHzzloIZ7q1sl+D1kYvtNxmMQVL0zrJxo+Z4OE709aqPwxB
XtQsjFj1+5C65beVrv1s3xb7Q+CjoFBg/dhfCnJs7pmRgBXdnevayRY0Rp7Htwma
hFlaIrC1BTin/Pztw6sRR25CI9mVEI/VHyD+HnR9EArH9WyRc0eIEO6N/hxiA/31
+1+2C9lEXs+VkcQsAetmoa0wsRvkKom8wiChFxCkhEK7BW6rNpSEhcqhsgQ6wBnN
paeJdUaja7inQ+clYxeqspaDWMixk36C3MmEWP4L/SHF1dXlGA+C7ziIXvFYD0fQ
uPsHiRzw/bjnOau39f3G/Klt3DA2C+3ql+1vjsFTU85/o7oUyW7IncCyomo7V4AL
6V3w/jku0q36aV6f5mRzH/l+5UYmltuTKQL+o1GujAszUeGtT7iOoMlzdVE6v2oj
KeNQnbRYvyX+gXlRMkEJZ3jBn0PWX1m9d2LpSQtfV8thinGb38OuXJkT63U8+M6s
VRDquAO+V1qa8Gw3/1qXeciilo80526WheAgBpGXpUw03ASTOQOQpaOQAMP+7IgF
PgWLiTJnMqwcAyRCRU0iZ7e/bTPEVbJYAuS/HXOtLFWBIrDHD+SBiemu2RBcYZwN
+1TnCts9jsTv+jKVarCoYdZcvWaap5Lea51NfuhZAqICZciHKxhx+Y3XeWijsIO5
z7HEdbd9/bzObIMywQTIPYptx9w1Ht3lekfsC2fz6zq/niNQsLd8HOpdr+rU7qoC
Db/S3/9wzA0mKiX4nD+ASk9UKHHZ5/XCeKrtSrlY+N+p4UiJluAWwJ/t7NQAXVoo
tE4eKJf+elfYNKnM7Adan9rLPhN1hdyQyQ2w9jZ8SIbG1V/9NPO3hH/7cG/lwDa+
e/Z1RpIbagJA4T0kWFuwUhh15qGlZ+W4DBsg0rFVK3YEA25GG2VOMn6timHUJD4r
I0GVtvSIBznyLHWdGf4adCdh+8bWpXIINFLGNu6q3+THDNKMMYLroRyQYcj72Sni
I6FnTw7Ko8rfyuq7KcfS7A2QchPtmDRPz6bQGuyPEtlqFsCIPRGP2WF+gQ8oYMCZ
eCRgKkpa1x/905JtiENUGNm7xBNviKyN7RwS5GLM4RWlYZU2Kg8UDZG871m9GL7v
uLG9Au5reAn9uzswR/9XWwF/ngktTR8gKpjc/Iy1VPMdd5JcK3YKVISK2yx/oTvw
imy+lNEaPrOEEEuxqrnYb3Q8uYALj6tox9RkQX1RKz8W3fgX8sbsxEnI6swRaztC
8kiV3jIsqGFBrarDB3LJ4V9NUUavajQixockO1JbQ8SnvUDbA/tqEcQi+qFGve0f
74+qHQ+3ImRt9h3HWq4Eb4cQQMHGN1YrlL+1/zFdTa1kaV132xYW/E+v59Fl13gt
YHv1L30j78nYKdHmfrW0NT6/meEYbzfHgL56BE8phMLXc3FN29ubrJbALVLo9Eaa
mhV+0RA67nWP6y+GBOMkRoN52PE4XWh94G5bk5GZ9oqTGgJu+Vp2hh8Sk5acZJ1T
WfTHBAr6FJq1R3AAKL1H/bBJVtF0IVbDCUBZxlDsbRCv9Mx+/N8bMn3ej2vKsr/p
WpWv8ACQX4U/FHdUitYzKf5aIDGrr7uinEnrBBECwzAFGV6TSVH5kwIbeAPa4ymT
BJrLqqY6y+EWLHEXcb02/1UBj8TQZZX0Xm9I9HJIsNmahAfMtikELyj5Gd3WcDv+
CYX9uvKlJVkut05p7DiyxBnkLo1dIJnbplquFSoxG5Q5pBJhYKTCg0IXhqQKPE7Z
tBrxhxBQ136rdHEn7CSburZ6vuhQeUh63uMs2NiKllFkuZ6gPuS/PiGrp3FJuH9+
T4GjeOXzh3bVw7X8VP4foxQTfVp0hoWLFAGtii5b+0HDFDC6mbFVnlIMFF1sxUHq
p0EXCNjQGE+GhuSjkkoiBw6xpkA0LWABCLXkMcC3nq0GQNO3jI8fFa4//NvJEu/C
ako+PdZP1MgvsUlB0NVG/eMKz4jtl6euRPCbixUFkX2U3ko6N6Np6PWDyU+0YQoW
aD2y8psJm63ELVic2KkOls0WU76p5He+r5CtUxsP+s6FduaLoEGCCiJW/8qtovU3
9BeosjrxLcAQFU/0OmI6k8DpwXBRSOKhZ2riC/4nRO1+EexQFk5WPU6XW4SrrOYE
PzHfJ8BxPrIRKlMsBos/Z+fWXOMfYIoE9QO0s046jpxesempBILksQOTCyQt09Mg
J8ZDjkfsl/ekBSTg8ZJRVA9tOAChx7repmOBqZqjykHg1fkftfpZpYJfusk5nypP
icQjmrczrJv8SXTA79ctSfW/kMTe04ljPyaxT3BQcbuOXrDa43ZcdV8X7g9pYCzm
cw0akXYc0gtgOzs/Lc0T5EMnkJ85sAP2AfPZ5QHrRrNqSl/d3obLmbLpFecfneC7
5lNgMFbpIPCMdYdmzcQ+iS2UnnOoQfosub99NyJg8u2oIiy8n4iN/OnbTtaXBtFA
KL+Ft3FFuuV08y6Nbu21t31xiWJt0SkQyTKLB5c8tIg8f5yZW07SvEbqluHWGHVU
w0AYnLQid1vHv1r+N/Yz77MM/UxzOatJyqaoubR9+Ij370Z4qTKOP+dQHUjkv5gG
7Pg6P3E/LUvaoMqfXxpuorxCCPvV6kA9mf6D53DuDm5iveORMEi8vbIRm0S59IYT
k2Lf2aj4TpQQMAMjpYvAu3eQwq3/LjTDF+itoLysV4WpMiVKkZVBZtL87QTsV4/H
Qjs9kxt018dNtpFq5rBj8vR9Ft1OXPiE3U2ccAFZbfaTfY0gKC1Ht7YOHOAHIh26
g29WFDFYiaIqbzxBm3oBDfeHps5PJ4ElC7uH/JHqLLypvoKlhJ8MeTgWCizs0sgo
rhS5/E0xTPcVx/MSGe5m6qlTyZ8KdyvuO7sTln25FnMIAwf9oPgR//G0EcdsEcWX
MrNAWzgVTvk91u3rmEoQVKM3db2WMuPLQA38wqP7IVj67/cmJBB9DkeQ1QcFB6jI
9QgZaDB+WJUahstBYMsjJBWNXf3Sl4eo0jiY1I/qK5bx2Vw811jMKcq/9XWKX4Op
2BEqMX/gKhR/oDq7CWZgij9h3X6C0n50T/+KOPFihYmh7P9ZfVtEwPNLqwc+Q+Qr
ovTXKzeq8e56ryghKnCFbUb62+f0JNI4YEraJbj/EgmKgFBFprMi0LCFO13HKDk4
8liW9MdHyfBsfow605RolpTJloH637p3HjRhGqOAuzu3od3J9LgaEoK7iQ1BZJws
rNL1KHUeMNjUGQ1hsId2LZSpoqX+1v59aRED/8cts7sXbmS0KyoJot6Zu/ZDE2Tw
YLNcKpbmYDgIAiTt7gFp75l+7STIohUvBEdfrv4VnhhxPeBZ6Susew0w1XhTZ9Tp
OURMXepCXmaJUlsbdElPPtB8i7/6uXf+TmBCf83c6xa3Lsomt4COLQ7f7wzFOsmh
vsERXjBYlDlC6e0CusGauQFNJMvZfp0vT5uFCOgl+rw2EXAyD6CxV/b4N71/skXp
IBPW66MbxNfDNrsYC4J+OKqXZGLzLFJQrx2LqMZrCikCR5LusxcVFg/B6bT4MhNX
n+fdFZOHW+BiwIRqq9O+CO80rZX9M9igJi1kDlJdE1vVzm+Q6DV52mw1XHN5LOEq
wyDiyGZ3HVyeFCY0DcQ4FIUx+X6irZTdW2BSoeyFsF/EGGYOAQ0iohSZajsoglNb
H+sJMPHsDRsWoCtWEH62tbMQMD0NWax9bcEDas42SLKOdHBqJgJPzGt7uEDzyIew
w/2CeJepTS2knOgSUiSpmkh+4PMyRdHDL8EixOPhFRsHiSJoIDkyDsbrQu2SXw0P
ArMLy4qOi3brl+DXbxLvV+BAcKOktnkqxa296YidJGT/oJAaEcUKYbKSGzLDrMPm
CJ07/4NTeQ92VfK2Y5bCUohdxWWRsGBVpD5emd20qgMNd96EALL11CcFn/tLP6kT
yFrXy/Zp4Bl8Z4ubtGBkHpVscOqx1Nvv6YqnSEZOyhaIKs3QH4qNjhGuYTOxAJQH
mDTPXpgg4iLPifuiwEHuYnKWtiSMbRx0uI+e8QiL1y/E9FdVBiQdnZm0DlcCCvnu
LwQQpdp3pQyJATW1NjrZYTZpcnNO746lWnl1lFlXEv6rGNoOyxaBX2kYFlVQVSo3
qFjmASrRlLHmLr745rpn2kfKeFbPnPae7EtSLRWIwROkcd5P5KuCZiRVagZUSwM8
C9Tyl15PVnWWjEp0RUWWhJ/XALPJzkbtkoMIYgVH4FtCknMNog4trYk21273cw/f
OQ1GoY+lq9WQ2AQ6s+c7eT3mTu03Af8Yf1aawWVCT2cXUY+a7zzHj7NEgsCXlVP1
3se5zP2Pl3+51sWpZfKtxg7UlPTkVwvdGBoYRlicZ8DdC+XrFEVd1o7ZnVc/6w7z
CB4ycRkfccWDqH/gZqfn8HTVnkdUT0X4hIAcTNkihMANn7/RhiYtxRjT/st0Bhh/
D6OgURGk0fOu+ReOcsVSN+tabWNKaKhupy1QVjsFebgm2nY2X5WE9YgsvGd5CNhu
z2IYPrfetDh5wxYXbGiUxkd/tXH69YiQjdwlvh7a/xEBk3L+iHGwYQoj/Uj6s/6T
gGW7Tq0zEmg7kGEIXeXfCBjAVqp0tWTsOXYRR/KTDm7oLlNtJurzeggE1/9PPHLt
Irhy9Q6lMhW2yJ+jnU6KfuuaQ4f+SmSPGI4LKma2G6WGLeOk8iqFuzykVVcvTikY
sovwdXnyn/UrA2U2M3tuZTMy0jw1DV9CoTRKW2MH/HHLku4QXo+4gFQPWQxvJcEg
gHnJTO+k+4d5Ie/tR4mN0eCOA2Mz5quShNSeMycGaIwNC9ZFwC3/T2t0T4QinORN
H95JEp49Ff0jyrmYYvZ/x28l3oXmX3k1azVlemn+LEQteeGwM1y8DMMm1qgmXGMp
/XqECEoe/AIeu530h7eZdXRoWbKOVr6sn2N06mJXK+xbzmLfjfiuNUYZ15wDXY/l
+4WV7iY5xePvDHucTp4pUKAL317cLZwvGdaEMk97zW2b+JVUOUNnaYPa7SOwBhdY
MqYemwEl9A+jgMRXDz6V31AE7GMFpXftJLDJyv2KVoT9xbgRpTNiUwSDFXrtPgpo
g3RY3yNASD7PGcWwYSXhd0MA+Hj/OsAlC4GyGuVMtJprysE/78ecYQVHXIIg9DUf
OGrbe6l98NERxcF1/5LfPhX8juvt6imMOAEUyaBTB6oWQWEh6rOs+Z5UJNfqIHt3
UT1i9AW2OGm+epH4A2gYvU/s9F6u+iXPMZUGBSSpfIRhHp7534Co31g4vayp+q0K
23LP64vSThLERH+ACyjE1bIzUl1+/TDuO1BWGuvYnW20eMdmZ3i4oulIMHG2tbXv
N+BOgLzSv5TC4GhVXiHhPuBMMDr8QAm+5hgKS4hMlltzWONtVWPxq7JIYN4y3EsD
xNea+FzQg/9k9xkIZTevEe9imSWHUwH/ee6+tzew6MaiJSw1DPc9V22P2Q4RJKan
0FyV5FQrbqCqpM3lsbaMVc3J6D5nMZQ2bgWWu6wml0UMVBb762c+zjEUYFvJEOVl
BAFfMiR0yNSNqr/yC2BkMIV3Z36ZMKwtAIXjtHrKSLWCTd1dQKz65lJVJHTPOFqc
F+azrDAqltc7OkJe/3nP4mSecczQjSEaFiulZTPjUwcSQK2kZwGjwgyLfAu58C/V
rND8cLJ9cfwghsbSp2hJQSDbwJlPOD8iSsVmraaLywuZiqcnRwWbS0XlK+miibIL
T9tzUUWQ0uaQ1oCimklASR4x2Mb6LGNFrRI+6QFXdxJ3A5yPAa2uvvC2VFsrw2OX
RZgW00Z6SeLKVETxFd0koz+gVr+YuFpenGuPPq6RyqET2XSmn3Ia6fL9NFziuZYk
lgs7Wd80wYWzET7ffo+35Sko/o0P0TT+LdOzz6u9ILJbHejT4VicGHYa5Nx6+9Bs
5k3APp5auRC71PM5B5Shcn5M8iJZ/dnFIvHEcrJhO9NxUpQTYlo9tofPr/FMYrTh
SndY8rfanqUVNE40vFHls7tELc0UF3CO57/oXiJkuyei6PzGyta1TZ3mhoM2dv1C
Y+8Pj8hGQb3BKAoDIMX+cYv9u4+uDFtpAVrv/9opslMJcNjx/f7wBUaasMpHU0DN
lgS5gcLJSoqUlqS1j4TTMh16EyPe2UcCOmxLCrcN1kO3h2lv9YXaZp4rshPeGQkE
wwaz+gDzIdWSplquUtLAJBhLRFBLCnoRnuuQEW7oN3fq+mURnyOj1n2UCORuWPoq
d70+hB5o+XzC2DriltXx/KcO274S0KJKSKqMhjiQFudh/QVqZgJOeg70GWdhBYL6
mRo7PRBnIfv3w2RPFL4jyAh0GTqdLEaPVZJhUbiuXHwb1oH7mEO5ASLZIkkHk1qu
tKr+y9BVdNsjT5+z6sdwd6o59JYDPOw0jDZvY1IDFPUSAnIBwTYJDSYYnpDmvN3v
1wrJQF0ndIn7Cx+EjExvi0wS/yjBR/6DFBUjXrMudACIfMchYEqwObZt5lCXn8ot
DJUaOTUfxDD7Y1g7al8qjgn2hQD6/x/S09anILw7tnRKsvRAJzYNaEFTWUBdX2aQ
X4vBFZF7Pm+c6Vm01q/BQ2HpAPd8+q52GmOE81u1yGKAb3EAw/8kz+5bpVqZ+R+1
/H46xcWUtr0D1sMfYAmsj6kx/Gj6az53/dS3ds4pyPUZkLICvmhbqg6A6VpkFJNA
MZ0gJJYytTueqQuK5QxZFcRmU+ymXae4P2bkRvouu2V79m3tPCBdOoq3xvw4QrBI
9EF5zOEG63qq00HH08kS7vzFF7ptUgf/QLMIAiggc5TEd+tX8sKJQ5DTQzmMxhvI
uZHPmt61n/qT6NyjyetCbTkKnWtHBVxYD7RCSIyZkvgE3rXDhD4u91tCGO+d0xTJ
r3JaHjnRk2XnA18lPrPARHibzrB1Vh4MWN0oBE0i6eh9caH8wYDTLM3MfQOqzCiq
/4Iv00m2Y3wCw1LYHmcY0/6l0cK+k+6a1Od0A7edcvJ/MynCWmaXJHcAlPHlVWHx
A97ThMVzbCWXEzX8OlTyTz3Z4MLB3zCCesUlGB7OLQGbVRYU5p7O5H4I72qn/hrl
V4T3UTCPOYGE8qZZKVyZAketorZ0wqhrQtetChRqyFfJThKvMvVuCyxZnqE7AByh
4Xzdhh2MeA2OPZN/TRBMeKyy+XR+ZrlCbpzfL4XDhNpymd9tZ+jkd7hIIdEmM9vL
rER4yqSU0IPZF36WPoyT4XkQk5fHPdGJTYLbtTAHmK9dQUoRbj64vz7XBaKPX/tA
d985MASrUWe1LIJJuC4aAzkXkPWea4KkVJwLEc3zWS1PmPqlWso9SpIRDA59zOVc
FxnceFQcScGFRsU26UvByP5Fty+467Yu/ASQLyXSsK8otYrVevt9hb1489qeMN9o
Wmh5FY+8DBfDS+cuE9Jee22JGRd1K4PboO+/sKW0QDcWxQjBKLJ+ORPUfpEvlU3k
CTVGi3HvjGa52UzApRokGW84p2X5wZlGXZJ3cIrdVH4j52LZzTbqzrx7KaexTMyj
YejUP6Dli9LOMh/IlT68P4b6l3mHMTCBAd8v2lBgOMZhgw1wRzEEYoC0sIR8OdB+
kpSJf15XqEscrl1Pfcwva/OuXm1tqFllHw3cS0aVYwTo3jf1fd2MeHOFcF04xKqB
Owoeh15VpP22l1PdnUXTzwk/xvlSnQNiiG1LNk9tYLngtcOdImmbPVH4txGqTV8v
kC50UUs1hcR622tW0AQxV+A8DKPFdVofQ1iNv9mcG3RsTFLahvZRJNKV0uPOoQVH
Z+zS1T/IsChIDuKvbnP0TKodmrEVImwehk/bsmDtsKXKmzTMIaykcsn2AipIP76u
aeZsdD/uL9D8iqUD8EDSdfqwaUeB3C2LCCvZyGc7Rvx9wWK+GKtA2EC1TXt9PBEy
RYgnt18CxNwOJUERSpLgVJjgl6VebMWTBSp9hoOrkEG8pZhXDe8S7nHbgXJwCQqB
QTWKivl2lfCylaaHf3ICPa7T/y5JTRIBhDsCNKlbanvwapqR/Gcicdl7Vjke1cOZ
FDFmTmn33p+yuHS4So54prMewhg8LJpomlrd+bt/c1tHTsB8zOZcpUTwUwdawu/s
6p7Kob2jnQv9mY4EF3d50RQsrt6px0gaeUvHPU8DXUVy6OXY4Vm3G7MTuyQiQUqs
r5vytwDEN70nOYbJkZ3fFpv3ONivxsyt+qkzAFgyFS3KmX5kMUs8MsLkN3gZRpv/
h1fJoIaccuyvdDzOZUTGnTxPtp/SUue1Ftqp5CI+UcOO/rYU/B/noVIWZV53VuVs
HbTL4Yzxrnn5rWQ/p10kf9x2nTsqDbr41Ms35Wgc/z4fRVz7kh6kJ15vq6ebYXuc
da4slg3++bUYqs0te6qByFxbofFHtPNz2Tu31235WI/b93AZEZEXOlcUlPC5FZfz
fzbKEu8HiHOnKpZJ8cVsgMeJn92rgIrJFnlAGORwDK0w0iCx7cHaE1zOJfgb6i3p
CMH3Wfz5sHixZHxN49Zi7KqVc6tvcPvkaVrfA3ZDS64NLAiA5EqvrL8OExUGVz3g
DJum80CcDMzK/uLjqmxgbNKBR88FgILiZdrLRiX39ajqTakvvnUlb/HFfMKfFwpt
Ekn9VHdzwohsqADu4xbg90dA7x7UyW4RIw4kejnjk9PXUorhBYdPeJBDCMrOdKf/
mMLI6xCGCNeZwNjb6qaYn7vnJPgJiO4iA7Ub10lN67UYNHR6pkWzMLL3SfKrhGkf
MBrSw8mALsp9n4VOy9KnAD+dxOS5dRVYVvYFxeSR+sGgL57Fdxdu/p8Hs/Kwk5+B
m0GI5TiT0Gm91np5GzHUZ2bZPTNjiSCMxNMicYEBXvy6cbwD9G9tE4DqbEH1Komg
N8kwRO+xbS+MTEpi19EkLV4jrPTxCwGMBq3DKj+SQVWDxZ12A0W6Ew2E3pv8l2Co
ZooPlNJvTexFokXPYCjrbykfodtuMo9h/rRE6drCqchGe52CVQFvZzaxen5yEfcs
ziiov63gb20Xb4py5pchSgtNVejSk4jex8k+MpynSDCjoeTAzGY3bMwGJgaAzDkQ
+WjrTTafNmlcN4kyhwB6uLUt5SGj3thKXXl6pDRFdeaod7ZONSDvQGVHaZvRIcTO
oc+5MyyT4TRvYAyR6MvA65pWwR+RQCooH3Xx3btrPBGFziuQ+bguE2Xetd8Iuc3N
RBMqiZ3hG2bjmdFVQlT9C/i1TIkLvRfn9P2v/QIjVHHr1JUuXLW/TUeWtS4sH7q+
ztWGr9cw9fKjry9NiNuHaGdAK2vvq4UvFZzonn5gBj2jHu45lWIZkQ05IprOaCoW
FnS+mIboxNUE2x+BXufRrzrgpP4ueFq0Vuvy4qsIjmygACSDk+quegejFWuzBDGA
GoCl35w/yyEMrXJsKBB4rDwxvGNvBXydW6bxHKiiLD02G9DgLFyAWkl7Z+8wDXEh
4Z3Yr6xi42ouZ7Tsq9zM789YLuwSOfW7ra5LaOpjmGNi0L06bPxgdf9OzzM9ZQz0
GTrreRfh5X7lrYTcfXrJkziekEPuVQZZiQz/xxH6MUHneLO3e5g6dYow64K3kJrf
5KAifenQlk+mLealZ03oWmilYQXsCfcnrhQzuWT/A9XYa64jBbxIq0CGQ6RApQUS
8iWOq/Fcx5itCLoKNBqfy5bn/Cm1xbNs+1nHkylfnXX4XCYgl/c8yrjBcyu08AhT
xZLBEeGcEd9Miy3pFNOs1z0AeJM2X3G07Mur1F9tCXH/b8/poAoLT8qZAHmzKJ4A
fIGLzR8JkDk23caVTEYK/V6/B0LEfcghXsZ9REjiirY9T+wUvtl/kIKn1Q3AO+xQ
4RocfKhs50T1PFH+bNJ+Jqun5sVEFkdKdV4tt4P7s7jWmuBXO4FmIA6T/09qQQWA
3fN5hr/UgGqUG2A/aPAs5MtIGL051akqjXIQiJ4QpRNHk4mgDy2V4IA5M19nHqzt
Rtp7dR+wco3OVMtSh947FLtfdpi3e5BKKDYV9ho1DvwgwlQE2L6rNLkg32BBm74w
n+hpFlDQhCyQ7n9og81ZFSc++Ny7EOAVPsQPwPB/UaseknkSx5LaahbKJfM3S4GG
XU1cTjXgwi2I9AUNoKPS4dg3k0smBxBOwjM5Y+5Nt/0d6MeG6JlsVYzONbgN9ltH
Q+FGTjUorcpcPeGG2qVKAoFmXgYrv/h8ERuAA9Qg7NE5W50sxIoWTqaQFD0s9K6l
CXwP/o689WC6unmwajHXHLqwiFHEWrKy2mmgCnf/zHl9PsIc3ugOv/R3X1zd+Flg
V2M+CvCuiWGVoUDmaTGLfNlNc8hXFvNX0YrQDNVAnmBeAUoNXgxuHLOVC2D5t+pj
iilMO6qBP5J0jlJRUDsp+fRc6nqmnpJn3ETy7hcqbAvdBHQv+Ey3zFIOpu+uoVv5
HAbxdTMIkER/xoOn/KoXMRHyCL0IoFqktZEBpu6SW04B+D6bHDOcxOlNnwA0HNFf
bRyJWFm8AYDSfA1OSO+FzDio0QcJqSJjHf+HYj09fUj6pN7ljMY8ATAtLXyXjfDf
fYbEuTySfZuWJtDvVgsLxLQOvO4BrpA/HbHMNcSmzvjhvYUJomWMvhe+Gyl25m9r
T/qiv+857t0ED2deYgNYdy8L+4fhdB0ASs43EuwMxanOmtyojSGSA09Ugdqzn11s
0Fjs92MMBV5EAgpfk/idEhPBsfLbf7CQb7iVxMeU4IMyHTBVJE9j2suWG2lVXdsR
Vh0e7vqAIsI0wMwNnEHAgE4Yaf8z8qjFdxOKYdhW0jZ84vC9jMTDW3vafWmSlkDc
LvEzXICE6fyQ3I+xXfQc1XU0mejKRXHBH1056RfJJFdj/OZ1QQ/E0Y/g4mV5DSZs
Qg8PLBmBzcKsuq/mrhJs7lrh0T5hVqGLPN1Swy3BYc95UCE4zjCL0t8kJsUC/T98
EFZCU8BgnvYG4DnEiH6sVHul08xkPqqYadg9UiFcXYF8iaGkeryF+NsMIyh3TxlB
gssHtRVIuZBnnBwzCdbJxbDY16wduA9iWxlEImE9HhNhUkRwG5CllqtKsg60KQuZ
sPT6QR9oSVg8IWHkeJ1gq6G4o4SPjAgyacJ9pyCrhtXknL7YyvsyRwtv8tUb5RJh
QUPewwc+HRJyQ74jVxC1MIK+I8CgLz4ZW7/6r2pnEfy78M/MiDcITusc6o15IXLP
9KgacoN70jakJ02WO6jSj0FK5n74yfuhl+Epb3a8f1eJGEwj5/ysjuJLj8dCEFCZ
EzVCtlKdlb5aI2omsx8d3M1tR6fO8WIXobeeB+PIY29RL01rsmlVgy2NhNOKWpqR
8OSI+4VTBUfC/Y1yinpcRdVsDpn0S/MZZ7TAu8AL9HnA4ghEjBDKFT5fYksoML/v
TBG66YJ+kdD6yfUnyYBGpseGVmF6nTwRcMAbyW11lHTtjbGiZsVuQdDILSCN8h7v
e1IzAj2asWQYuG/yqDEZXd23cLsxFMQcN7zVrWxdxGJMoOmQQfp2amWI0UdQInmt
latslP5e7s0+fWjg0D5Mif5pAPdXmwfKeYGPRpehGQGHb7k1tZxS1twTd15QHwNU
asQF+7AghHpP11EWaNv63BGyuKV2Ec274lwDjG2O+VOn34H74RUQ8X5yb4F2cpBG
GS6ixa+N0NDXWaUzEkjHz++4U0VhTF341C2ngW49LuNsoby5WM8y0ZB8jOEpfHHN
8Y8OJQ0G49uHgguuwDPvC4QKpnxL1FXZy2IGTfOuvAnNOZhjBtL0atdY5AQK/7oV
CGCoC3D20P7HijKuMULqMoFn4cbk9P/b/ULziKVWbTPaxcWIIZEN67yGQPigxb8r
Wu5PfDxTgjzjkuNs5zjluubANjkujP28YEGQInBIELeFKlMBtY6DjMN7NnxNMdAZ
rmnMH3G/IZyUs6VYnk5tOHr/bp+et4xsmrDUYT1SV76bbQS/0jbfIKC93KsSve1d
NOlgfPlBhSkXM+n1QRLevfrTfpNCXB/B0YsQzrCdT8CRCCMMyOTUID9dcFl6sjXx
eyvVWQQb5uzN3KmRPn5bvMeplF37v7haHNmMWA1wqopst1vNqOP/EcMAWT2C7LWr
al8dHYb6b0iFlorfsptBYRbUyeCzPhbCFpC2YqcDcvvIbSPooOizaK0DRTYmQkGJ
1+F1GRj+Buz69MY81dWyzUB8rdHx4iMdtStiqAwAYe5CTOAO6s/Bs1ZVRp6FycW+
xFxtBK+dHJIzhf77eCb8PQzlrvElqXHF5vunFeCuNxU17I7d863XV22vNtaC0bdC
CXHXTG+QxkPG7arlP1K+SgIXB1mdrahYretoGsJ6iFa8a0wiN8d5mAJkBFzEoIYy
b7lJOl/fQ+nCOiyX6GWSDjnuD+3opAHAMYRA5o8r+Ux9vjo6tBxl7iyckssZHtc3
eBB08BfEgEUK0h5Mv7p7QsEHmQatB0hzK/TKF7Wb6Qi+BqsBiunracw6ue7JLAiR
VfhZdaI5jY8FCv4CfxDnmU0iF0wvVdBWYmJMNr8FJK8RPKwzKY8VxQFGn2igDK0J
QsH11UUXBUqtSNZYbLjqHBnaYxtkUw6zDQj5ev9WIZNELnQIVeTDTZgjChKXgaN9
trxJ8W69HVpThFFovb5lp6Yc9TvYnrnTpy3cfONlofhokSE5t5diLlrqv1LxNQIB
Gpkccg8Kwq1Dw6aiuZjt57YgoEbySEIT1wf10+AAT+yaW92ZhxlDVq6wqOatlSUS
P1e6hT/UXGWZXORNM44KtJBcuutc+n6bpE4BavR5FAuXXVm8uUHLjv3ppfj63Xyu
4GqoCliU1xyRdLsZG3w3gMQ86EVIMcmb2PcT+03+5owSh+yVIAeXdlvLvPhjBMUf
SrcKFMqm1k5WS/JZCkSpU6wvS7YJ05uYmEHVTiYOCGBjyqIz8mcIvr87rP/nnH+p
Pg8hkr8kAG4XKnZ1ZgTeu/LOMocVv7oUneRyASO+4k0FDnFnJJJE7evMklnvqRS1
M5RbDLLNG29Gv9VUJP2Q0FbRMMgsLtJNE66W1G+yMg+xunXTwpGxoQYnMYsYON2V
wj0vbAvsU2cKe+LgVA+du5fLvC/hcdIh83u9DSqfRzXR/OjS4wlx/zdYvIKO8/87
KfvdBk4Vymv+4A04dN6tI3QLxlDRX06+70fPzilIkPcILfkdztm/VnMEpJgGpVhC
XeS7S9OrSALjkddXdggbattE216axajxF95bBMNEC3FcGxm3+Mt2lslO/5o/zka0
W9t/7+2HaAJzy9tFA4JJED8CTsr9qL9ZAq6WiFq6QtNj6pwguvGmO7WzYSD+xqzZ
oBqoQ5rc5zRtzcZ6MCVudOQZCSyQlHbOb/zb3pan0CWsKG+ujAYmDmPdmjAQTv3v
th9R9Amvv+hFEQATCWQFbG+gE8zumapKQmrDydvOpD1mXtj+iDPxBWI/6Y2hTPDX
vBw5Cyu0Mt6fGa9rEFRtr7yU451pT1jv3rt4QFP1PfxW0o4/r/eYjlFkvST4SEmM
6aNwJxGd8w46yxWS2Ll3NfkqjCImDK+VMsLjVnKeb3GJLre5vTnbx9pnlAnYWA2b
ujrgfdr+i4VRgNh+The6tP0dDn/TilCwyl93X+q7Iar3yKRvorZMWoQWAOcA0l4l
YpVLkjyI6qDef09nVKxDUMoZ4NzzAzgwpbKrlYZSSRjAqt19ddqaFEeLb2DBvW3P
dbiMJfqoT7eeoDL95/XzZu1nBXbOxHuB0Yyn2rz7x1PsZ68ivdMA6Pzb+8Y/LKIQ
UY9bVv74xr2weP920TTcWrY/6NibYlq9vscboJ97M5GGA4wLXwgxjZeJe+mTXESk
lNYPFHFxP+fIJjKuFrwizFOOv2Hkek6DFzSAYOyehLaIxJAG1aL9ZT7+K/NC2VQI
UrKEQQRFoFGm23wMJIOozEP9OmselA5jv9MxEwoEyIdmkcgvdXQIAQ+Uw7UQrhBz
/G+ZZ31Ff/UtSmwR3guj6bDHULeOvX4I7LZLz6CMsL8friSjwQXyvBncMZLIIJkN
kXj0txHzqqIg/aBFIR4ymDNI9xYY7WeYkvkMVdyKrahINZIitPayzgJcj4PkzP6O
E5Y1poX4CJ0Dm4NcoYp8LDHFI3s+nW80AQb8OWy1gCjJHlb5aJcRdIf/eKHv7b2h
e6rp/Imr6hRuYBd4i7msJe1h29P6mAPWMXoOV+zSPOrz3wbEjWyp6oIvCFRSzjO9
OKxfml30gWemhAMU/NiWaiSNUB0wYK1noitUAVlgV/WKaCPDZWv4pYyHLoL5Vnt6
DW5HmlwUc4KYgeRa3mnBb92iHaF9f5aI7BgEl5nB1q0PjV9N3sM9A7nkye/+/uEc
ru4LpYdx+HYM7odzpFYVLo8AAsS82YFN5z5kwwrL8Z+3Le2IrJyVGTnZMq68gbDA
1rd4f2C20u00gtebIkWnctktjytrKc2z4TaV0qjw0iIL2cwS1yR9DlzHMNTgMbnN
Gk86UHKEoKPbJ6CoL7mdy1iW/Lx0K29LFTpD8du+nVwAdu8oV8YLdpa79FfuONCC
fgOgvgpoDGwKNw2nUwIrFoir7uaYKmn0zekH4yKNfUjW6FQ6kXgaNsVa5X1HWqmF
p3efdqb6g7FFoyd2U1rBRnkSc9LlBtESB12Voy0bf1tcfUynjOQ0HiRYVCWZo1vW
GSr1JxDwBxJOKVv8h6shtBF8EhSep9xL0ZizaOt2r22SQhqk5UO0n+dpDCcFdCT1
v2d62e9lh5YzT3USP1xrutl6K4/3lgkjLmfJ5DWIyShpqyRl8qWnIu2eZrkAMuWH
VkduLjWFNlQB6+Pv0GwERn/iAHYs+6IMCztOxBbWse7GuLvjSo+udFwojY1kxokE
b8d+1VRvmKthCDwLxqZqSSOSG/dJQaTFxmokkMqj1Cle3arubTIgo41uvzPzMjee
+80t0gYm2+9I1VeFrcSrsRdMViFaGNwY+vS5ZqsHBm6MGfeaJMwQCRjwuUiS8t0b
QbygONta7bG1eIqcd1RCqGHm09y/B+QjiTcoTRDW7X2afEJOBkJA2VKQALsuQKMm
EyMWKHDNNcCjSA483ijwJKk6zmS4wA2h4eue7J5wXSfyREMapVk1jmkA2Zrb1mA4
dgKHAkilOkonflWbrKR2yYCbngmk0dmE4r362BPovdsXRzmqC1UcwJgvqW/N6c8A
Z5zj4Vqk92OzbcMg3YRRzTkaZ6f+aer2KGuH9WNxWLkf+th+jJssaE/SbIWab/Mg
+q1LAC09dWFmtquizH+pz8vf4iXr6A1D4/tWo4IvZn6gdj71CBFhMCTy1S4RD/dy
oCKOlV+b0HLl8a+X6QaKAQSavxxcqlmkU99wco/irUrMm/G9jsOa/f9zFVroybwJ
LXvFMLRN06amEemeSBI/iWowomKlIvNuGbtB0miWaQA+Ub6zGYuaz0HNyQ0EuJya
HACqYNMUqFd9Lf9CYIDAzJgQEg7v2pr8mrkgg7qewExa07U6WCm4bJj5WOymBLhs
kIDYyfLkJ5eJJTTfiU4ghBrxDE7Xn80JnMakNBZ+4nKajgqXkl+825TZ49MfJ4l7
QORNlK9lWRiwHV7lzbj1t56zQierbEjBDL5ZSnj8PwbvToMBYwqSF5IHrsSatcIP
a8QcclSl8akmfkDuB/gqFb3pXIaX+3UdfxJqU/AhsYRTXmAKfUhNM6Y9P+Dt4Plt
Q0qQeyQFi4lDBqKwsG2lILFwFigoH/84HJ2MqPWWx26RXcD+Yrr15MXVfRXVuyEk
Un27T14mJh6KWEI4LyhKF1gDt3agvnwDpH7quKxilV0Dkq4GZuHDmdtXBrFCUTUs
H57WzOCsz8RMgEgz2G/JNk7tBkN3bKt5Ze9PaVNdISKZWaX3vCcOerlYrL+tfQ8d
jBXjOQF0DCU1hxas6dJvSYmRNdQGN/w83Gs/f25pNZuT58WFj1SN7RbA+l1B9bZu
W2OAqyMqHZYHvwTLJMQaUSt6dV6dlU+jCzc6ldcwVI9NhrT93rq1AEM9A5ykrwCh
TAsIbHD51Zy/aRbfMmfmJFQcfO95mtzRE9EEZCbsdoogyI5F26GJPw3DjzcJsukC
gVreZYacTsapgG9mIL37TCZHngM/osN4aKUr7ZJcGArDPp5Y5+NaatRssfyuvDiq
sHKhViF0NJHpjJp2e91ILj4zgy0O/SekvwqIlGJT5svuU9Tf8Co1Iut4Sipvi5fK
okf1JqWDr1p9FfkqKpdSNi8xgJ2thpsrlcq3eg86kt0xM1oXVMf5eV0yabDhKzjf
u0A92HeE3xpj7C9EP2wTw6TeeDyNnmur5Ndc6lXf7CiFL9z1edQiHEmpE9doAHKj
8PuhBE+zPQ6x38KM5/bjt5vX2wmUzH/k2xU6qjEitH+zjV/XQn6OpeFzG4VwAkbt
SgWJIJo9ZClHql1LVmVXdffaGPH6EPX171WyVkrhm139jhu+FGVDw1Jij5vCqH7a
e71PeDIzrzY8cjFfwi0ZXiV0wTQFzrWbCml9+603CJJC569G97FKpFLYUQUggHRy
GW6hZ3d1NwGDKEjp5STYxvrv8IUmNSWY6FN/5Fj1hxyOu5ccLx77eEu7ddFWnemS
HyXydtKirTBt+1mEia0upvEnpojZSy73z9J2Vg8NVXjm3xB8r11bRgkg4lIR6s1v
bTNFUiP+UcOOb8bYvEF2l7rSDVI1Q0TnbyGuQZe7O5OGMZAXpzC89cEubd6YKn+2
xkxl6n2iHSRgPMSr3voUa3Xbb4aD/pTnJRLlBuc3/f/w3bqXRfYuveNZCr373zV8
cg7IGXBW/qz8bOWv3H7TtgxV21W+MX8oXm0T5aN8A3+HVssWcU5eluZfUMohyLIC
6GFHKgnE1nfHuNeRXRubIp1S+XTe+cPfWZByfG91/blksePAfgjfenlELIKAS8qI
sj9NmSLiJhoNvC5SvJyaMJqO97pvRfVKyZc+wfMSwEcnaFt6lCIEDkMkp0grWonu
/A+gAo9tFUFYnLyK/YNSbhuXq5Ff9+DFWZJsT8n8smnFP9kVdHY2r6dyaE4V6pd9
/k4BRFw6L2kfzcBLw6UbMhaI+dMvAgfer4zuGJd8GPSYGAymc5BlFQElO6YhGFEr
X76yGZpd99m01nY8bgqyFDjGkAI9RdqqdNRDcDWlWp3l95hDmzSCCDOaqEGA0hPH
ELKYEPK1t1M0H2pE5KFzi4yacYvP7e0K6IlE8mPzEjM20J6hf+BrRaDAtpWPUaNu
4Ctu/q+t8uvOqjbGgYT5lizfKa2WAHDJ/Z38pMI+jOjLLlk4kFYi2RRXKS0M7APg
1uQ0Ag295nV0zuNHJO4/PPcY+GKAa5ANT2PVoL+t1NlX/CpYO4NXYAtXrZy6IVVz
bGffj2AZRPA7V0C2yE6P8Et/E1EgC1NZb8p8mqMam/26C1mvK5vmY01SAaQqb3bB
32N4dvSwyy12JtTUXvc/cKq/yswyuN0zmzh3/gTU4U/B8Hih2TwP00ZJ6wLa7ZF7
PrH2xdiVV7nKV0VSFwUEfR3EhpwslmSDBwLFpapRGY1JM1vvixNlXEALrdF0nwfe
w+nCXpJwOK/BJxg5zm0bwySpYpEWYNg8TLiwgVk6wgSEC0BIEKw+ftk3PI1yoJn5
UlFvvcAsfdKzjZlhGeKkj5N0s2U6k+AzAo9t52r45Z0K9CUmkuAbm9BHeho9i7Ql
J1qQ3/gaDoO1v3H3vHXzhPXqoT2mrRskMShwjNv3czDAK9sst7FO0f59W8FmwNoK
oJe6GHW/Lukug4jqCsZXHY6fg1HLuSmaOtYwJN4CeG3TTB8bq/aq7dVXiTZY46kM
UqOP8RyKTN7Tg91wYopSeRSUQ3SHlmEGJXN75lmD+cDvMuF8Otn+z6HBjilmibDK
Fyqb2fDnxN7wDXujzRseot0lZX6AjGV9OxmATRGElZSugeDtxTV1rJJT8jwtFRhY
6+cdyNsKFXElEMIfSVIgxcmwkYCFYgv00QhkAYcP6B3+XKYUWdaNxTNgo6IjYrY/
c40oBFLNmWMocAU0fT2uYKSPy53ZLyz7ckfPruUzFkFVFckAeXasmnErZ42YsJAi
uBlcwxMXli67NDWwD6ijT1juRtCaMENpQQy4VUkLVH7KFu0Udud6VmwvbqnmW/eJ
M09eRKxsIl0p9smWTxEJqiKE0MWaGNHM4nz5XteC3GgEPKeKYuZiCnhL4Klp0Sgr
+9f8xWWcYsIhVzs2j25I8t6EQy55NF+8qTp4se9Wxr21Bd7cRRV0OA1gvhIh/vCi
TuNA0UdXn+uHSCOcZHrnXaocZbVftEqoShlSdeUe+dGgxoLubD58xZP8/0rfawp+
3zX5xanykEMyYCvuaWEYj6Bv/qV6WWaGHbLEfz+3Xkoh9hbSbpVdGBb/sCQa+2mH
suwO+tidyee8NwnJCWj9VP6jU4Ir8xh+j8cLUW3x3gQTUCVGNmWV83ZslenEdp50
NQc5+FjcnpmXSDIPR57OxSPEnW19JNrGETBoRUwnn7P/aGq6TvkKGnVMoXL/t7qE
X2KcdikgEHNf7u1Are6YLWve77kkO0YNIg9AJxyJQwlYelvPlfifaI9pkFEbUaMn
YU9CkZbpdQ9XPFAWsDhkBfPxI9lnFQFJv+w5I/TaZj1u7/DcH3+em0bk2iU4FHON
WKelLHM4aBQcONzjjUvIGiH58Z96qeJ6fqJNWRoA6kBP0eDrz+8DmXLoNcOoyzk6
8MwWox3gHGmGD6Ki2AOcmpweFADg/qzLP4T8bXrzKaL2hqw2RGUNfNLF1h/3xF+f
btDR6luBT0zodCQEi6ULEarFifFk6YOwYHdgdOo0mXKtoeZF85nSvBYQaNSdLLI5
c/418aoi2iwncnwgmtF88CutAYXuAtdEXnJmlMCbk9kPxtqslQP3RvdF8KiRtLAb
zRTI9WCDSamAsgTrWQA/2ixvmqV1dl7t82hsaDTQubz2YGLmNYOi5myZCZLQRtYS
1UcGF9Pgq1Ompv9jEaJmCDbJ8L2XKej9mJ1Fasdm5fU38gsKrr726HxsCHMTeFrs
d72CvbIE8ZFhLgIB+dm8VbZj05ZLdzqkggl0pN7N+YUs1vf1u1pk6q/jSDTPzqmj
YW6HBp2yjbWGOkIdNwqp8U9Y4Yc3c4a3f7HIVluKC5bMKvX/z3AhJQiFoBDcaRV5
iJUzGQgN1Y1c8ScQZ8QULF+ACfaz67PMIB65OeWLsjyqUCfWoqgP8njVhEKH0sPs
o2Jh0oJEg/EqyTf3pXD9QoBnBcoDKlha+XT3HTrPxSukI+9oCGW3gHB6GUwbDijA
ewqpBFKKbcNgn+s5y00JQXqLMDCqlQXTOdCzTv2dxLwZhKgGmSFqth46lreRSFe5
iIQO00aFOnxv05fCFfM4JZPce2obnjyEaAEELFJ8X4Yc8WC6F87sQJNCtyCwbeg2
KzadgjZ5ASm6DBshLSyUrHt4AJJBre2hb9JcYwNYIV79w1JMd3RL78zbE9zZC3CT
TUCc8xFNv28noCBCW+/Ls8eKFKagob6qUpmSB6qynpheB7xSFCYk8u6P7RiyzcwN
3yMyTQS8EeHXumUxcpiiU/QXIVAw2P0jEURBhKFgOFptYOPE92m2HIOG1IIqgU9H
dQDEMw5IME14oXOe1w/M1n5Lhm+Dsx2BkvcPY3VncZbGU5EG2Z+4cTEI/evUDnkH
srTvTXe7ykWUYvRCRgdtrzElOwvBDGHsqBMOc+QaFBEzxXavMgEFB8gntDHkdxB/
wuViuC39h0LhQDRE6jsZ6e4bpzbBvvoifQ04EbjHE7KjoK/VNxxk7zQ5mBm6xFFY
c8gXVExGr9IZrs0xsu/eArNDuN+ZCIFEErs1PjN6i1kHKgiNV739Ed1eUhRnIUsW
hCP6peJlXN6JuM3XPsZdp9xLTK5JyDoKILS/Gpskj6mEjAMpnWGamhdbfYRgHFVw
n9oEP/tLrirXXwSM3VIELxcQrkanPEe4Tf90duG2vOXooocbGr7I1ahuP92eSukx
I703fYUfcQgRmd0QT/eZ4LsDhkzWovwO99AyockEI5mHFmOqC1N0CVfPEHrhSmRK
uA4+Vh7WMi6pYTSpyYMktLEU/cCSPMPWckWCfJfctG3BmFROvDMfr4EG4PRu9ca5
M4u1VALs4hQtPuRg09ZON7SjaXLIES6H367dv+WEOnlIoI0qNj0U7j5If9/OQ6kf
i8wCihYFjuLBik9BGBynss2SsHCv9Kkkz1+X10VbLy9yqS5uM6n8t5wXNA56aj8u
HtLOn+89XRz/dExxhyG405QZmK4yQs6IAmu/5K3/QQ0BHxsJl2LmjBjgwx66J36S
Dp8kpiioG1HFhZOuFuwFibEuWPZBXf9JL9zSKwhJQ/N8VX7eTqhY1wimxrkq6Wik
JvXYvZWp7HZFjyaEgaIBV3gRFkP55qXiUpPc8nJgQ90s+FOkA3ir8MGaEoWgwPgx
fQm5kmvELhfyFjnmrzc1jkXpjQMKMXFzl7XVbTfyAlzV0VdnkYUy786K7UwbIswO
zBOMIE3We/WSt4P4mR1BZLnjlAMkHkbHv9/+qNe5wjU3QlDNmI3hFcaFBhbtyULU
bvHZWJt3p5yTc0fTXtDGlkbv/UU00qsq30S0XHncQQA4ecKWQPBuIu6v9xN3GQ6J
KNKIbUogtp52pCoBmmuA2XV/3GiGORNP5lIOiTB3p2jnycRPrUWFQtBDcT31XhJw
iHg+Tm1TXRcCzXT2ZOedf4TvsWBHsUL9iFYP77ZaWvkllUrc/d9Y8ILuUY7T03Iv
2j6DgcE6zGFv5Vy+iH9H5H98Q6YLJOVXlv+algphTXLFFuPbJo9aPhFGm29KtciO
oBApmvg2W6AICK6AYkVktMG3WxfSVB4gOu31XO6tTXNJ7GMJ9uOBmDadvi50tO3p
JPFi7Bz5kchA+Qbd+1DZsIreY5LAgGiGdV3QdYzVZRq3nQNCUnZYdF1M0AkRfmvi
mjUXB1JXLNWbgmgyrB1F3u7ohmJJdww02pef6WpgUWIFGUwr7mcYXyk70Yvj/wjV
bTRrLbdDHJiY9Ip/9jW34blbr30QGX+u98tJIzuzCT68r98yJxcSpOyfAwzLMqbr
9KoMv+mtZwZo2ikxODX/ah9w8nthvZe4Nt/2trkZY442OS1/WfFP7Qy6xYGTQ+yy
k+oHWEc0qzivq/hvBZCcl7EBJyTBm18A1Gekifk6fO8ofYvmPBlmsmF4KqLbeb1C
Zkai2jV/bWLrDnySMRABHxTOgxk/YOBSrv96Hyk+u27l5mU3kuSOCAO/0ddcfzvO
7e+hCp9LVoL3fZQ19V3BrDTqjOYvdbTBC4qiLP1DDpRU8dWgArLv5kx8qQZNWgSO
atZDqbApIJJ0Lh9l/rIalGjiNZQ9mF/oVU//IH+EApZDEQbGTTJjVzXCWRWBa0zr
vwyYBc62x4y5hpe+5El3BDw+dfDj2LCPklgTo2VrWzaojrHqwaaf5RDQ6lBzoxIP
Bk68lpM4BafLbWwUzw1emykBJTEd13OVCuhepBIIXlK8RqZDJkj4IgIgjBm8bsIP
CjL9XsrSf/nLXyH5F0joB+FefrXgvEkdcUepQA969pzSGTmpMFKZktOebJKOGGbv
FA9hOT2O6blhIApXd+FvVEFob1Ya/vl24DsG4qDmPlXqyKf3gryLftW7eS3P7N79
oa/omjwYY/A2uLotVmRaCZCFLoil2H24Qc5aHg3kDh5KzkJbMIZahDEvuJk7du1B
B3AzLkJVt/Ydbj11aNwHjW5pkNtWRPJjnSgG15U2cd1lkrzu3SWOTLOeJpIVXpbo
hEp6qiwyRisphq0fOZDegyb3b4hdXILffzhVUphvKawbagzZe9fBnvZJcsCu43We
BvD7LoDGoXFA7+3TzTIdB/wYCXNgzTQ9xEQfcmZFz6dEcW8XcmcK5tkzgli3jymu
4rBgF8kRYkQDgjEh7/OVpy8AiqA6frRrwUM1HlPcL8VLedCirVb9hUDYivOGCybF
R4kkxJC0RoeqF65iW6jLsi7xPyGnQcw4EzJOSM/7QF82wd+RY97rxMM0iGDfOvEe
O9rcvUdMbmwlpQrQbSySMZU7Nqz9qQ5PHr5LcI1XFG6myc7bnvLVaaEBPx9naGY0
UEOCtZxtsVCpINCUOvDN74fAE884OmvrNbx9bPg+Z4FCR/pItD+Hw4MIcld2Z+pq
bh28ydr9/7uuv0AEyMCOCN2Mj8bNH85/jY39akaheA6gMsZbv7iU0ANSbnfYhVEX
G+/T2bqJJwCpU0D5k+Z6+QSB8n0uUXvkW8vsJ94v4F/qbFl1C5zBPZZJJdtAjHIW
Odjzadr5uWkU+mIONPLnqeOZfyT+Cmpvbb4ihVgAtqbxZ9s2JamOD4PY+8WaJ03V
AfhtL4NlFCFopGt5M7VtAzK7m67ghsP0zs8i0ByhfQsPfzOXyPH217t7JHOHsgN0
OnI3+MTG9J+zZYsimKQO7uuemHEvuTltZTt1OjBCP94LPvh9xSbozylWRR+iZCAm
G14Rf/aQ4KQs+s1qATYbPjh+CYIb9czujEObnlJkPGkGrIUNpj+4jt3Qw/Vfo6+X
K5EFzHprlq6GnRAiupcLKgG33udJHFYKvK6B3eax/3v1ekzVOj+0sAlBVAHkvXPK
pth7GZRcX69T5UfFNTtomezumsle50v5lg8L6pcQlDj8Z/wVgVFJxyuBR594DLEF
v1Zb1B68QTuFPcH/n8vspVlIXNFnsyfvCfrXMiLfwagRgXVSo2dndNxzFm3RFPU7
14um9iBtOBrGi3kLCOFa7lwESWH8rSejx2mphGZ3RwTIZt1M8o2ooclr8vdcwi3W
+5M4YIrMIidBvlcOzp+m+MCllHjCY8UKcUXOsGq9WkRgHY6CFWREkGDqGjcw41qF
kuGCl2RPamauXfy3Xrv3KzUW3GAGZJtdutVwqPcAL9Gpnd2WJJ3mqVOGPcVYqmYh
H3jA/wnL5dACj9XF/G/9MpMriBP/H5jagL+NOAmgnEfKDXh5yBQYwOiY3hkpiTub
avDPlxsoUfU4QaIAE2Sz+Ah4nLPC8ETy4mKYHIcpG4kjlque1xZBcXU39pg302D1
svW9sutfO9I8OAiWW2tZ22oec4gO7/ZECS1EqkJiMbLSpF6F7xPMHms7jzwEaTsk
rakFlg4Va1hOObwikXVhlWjfeE+CJBiWP7xWribDJ9DeQMkU44RXQ5ajwck7XQ4X
csP/ow1zd8Iv9Q5Myq+2V2m5Ybl8MuBwqR6tS+GjymXexRMjV9c5p0c6K+9S3m9V
XF8zlog9xeEhS/MhActi36Zvxggx+os5URjfExuim2pa956ibPVt4rpu1CTvbLv6
I5OMifwtF9hL9EadxgtjxkKUmDiBJF/boTrc/97AqdZE74hp5+QiHPzf0tjlHhfl
rb2LWTO5uZeP5v32M4Qh6tZwlgVJIj/rwOqU1WMvF8kdMfjbxDba7msFlSEj7Xei
hW+DKap1H/6jjNb+GPKgxtVyu9QG4PQBk58nNTOJkwwdj6VEfwXVePRGOS2sFK0P
onx95jyy8eHh6eT6R9Y8XpT//rltoPaPhCoCc/2Jon0rBnubaSFc9joX4hVAwWY7
MCbGDQK9xKxA/6hUxXegSwmEME0rtZwXD+OO3J0nG/ndsP7D74ymZlgTRXBqG68i
MnzfkcAFFbQakq9TTzqogO3vVWc8lPGoT1CvjFVNJRXXtel7B4mlNdQ5hBhtW33a
XG6dUXcm4nWhHxdrxXvWgsjbSlupLjiz0yL7xQtUtlT5NTxnfDwk5jagTPMcKq3P
lUEySXG2grI8m9CPD6R5CKTKPUgWFwlfQ1u5sPr5iXC6Yf0uLH6MagUPiivbjg5y
Sxt/+5It5pA1IBl64hCU7+0USZS+iGHsWi+fbHS5i89dVwl7BqnYHNb5P2NwJg15
2gvaAWRg+vUdnrZhNnGbLmGvTCNATij0Ae6ohn542Boy3sGF1WVRjilRZqOmOZ5Q
FS/MOagU0eIfOcbaErCGhWsnqV1Ud5dEX+tJDn8yXwBjD+ZMkjIo5TfMDW1BJZ8V
YK2IANqQe0bBji+HyAd95Z5pz0lB+4/OsVwxnohnibXcSxwjpn+vFUq91QlDkefs
FrrswXtlv6Ty9n2ceoziVuZ5AV191N1YGlzumf9OTP6jUusKomzbzS+px7VPTQ14
/jBiiIQWpy3i/VKBpL7kYtZX2I6/bzllLd9xmQJwZDSQICVJXQkmE8uHgnn8EY+n
9dJe01Iih+TscTn+rXTrNJ+BRaeSnUZXl9pe/y4pGY6k4+7w/fBI7dJ1kHlGLUbb
qBCFv5Jx5vqmsPSg19C55f7uVNU1kTFDmesBxKQXZHsQRBf/N4CZC6pQa6IdfHkU
Lg6Ph2UAAb6kx2c8acqbiuebeoDlVz0mIvBsZL3ImOv6wQcuSs+zcuyewvRbPH6b
6dYZ3rxg0OXQqtVLaW754z7MvA4khOAvxPM+0FNDMejGwRR+WbWQT5w85g2hVJM7
PQYGFRN2HBBXmMqmXhhP24nc+HT/unu9VT28BBoVUfwmxfwfWd77vkKRkX77hRW4
BLWGlgRo3jZ1d2KrEz/7iwzBLQOtbqJv1EFzRzzfVJOUtm/wGbg7JK1ZMSA3b4aB
GS7nvtOe7xmtIGCeD6q17g2mE3YcvtAKF+saWKC6ua12noxYITknbfxCyyDV9K9v
NudQvPXxJncUs2goz7kD5gRLj4AHv0QTtcMAeKkE4WM+U0pdTONnKaiEkoZ9hTTz
9Af01in3k18k8opf18zmkjQTR0tBJHf9llV4CNTt5tOBK69nZGcV7DarwtFmguYZ
Q33qm4XgTNekxJMyIbLIbFItKxJytVZRXtAvv7ERkjMCKp2PtTqvZvmThgxG2+UE
5fO93n60GZ0uoCP1JYYoeDdUMM99yZO7t5B2q6S/OTUbDJRQVH34srV/XWosmkYD
FvVdBsvXvG3pQ6kwXpT5FHWqHlQ8dorivAzzzmgZsUKj7VCcLJvmaIbZFZBw80Vo
jrcqWEp8+A7IancZ2JPnyhkuM1wTMDHBQj3V1RSC023g2XnBBgVl1ckCiw1Z+wA7
n/LAg3DyhIYr5Xzlf4fkGi4ARVm4L+/Wd/7kPpg9/BPypDpLGifn689sFp0yvg/D
aB+qijk6c/RxUgXG+XPaBfrLHWM0PnLTtcEKy1qPWuwn1L9X5LhYbm1C8Irt3X7z
tL/abyb/u2UWkDS56gqRWpw610RnN8uE0LbANP6brg65Uj6s0T4e2jOSKa96Yi+h
WUvoHOceQhWFI2wGI5QzgM93sr+fVdxw6fntPbvClV/IN8kfQuB9C5Ejsx9KHLAy
C2VADVFgi8e4kvZBf9GVzUlFKRZrfr2hxJSL/cTQJHQDY6eAqcu8XIFlo9ZbSLvt
YPdsaKmf/52tad7PppdEriSYYrHcs9js9pnVGWE2vBbzx0Gz4QRoFRAr5Q7UU+iS
E8Jaw8rN3tyu26aAnvNrn1xVboMBkM6kao7wgGSLV6qRnL2rqD7FT0fl6bXjFXC4
WTKVx4G3aEtVbK8bvlDk2xScf4tXjOMIDptdzo5meCfTDShTYtwUKtvJYCVO5sa/
gw9rU5Ia06hB06Oeg2AWS9QXeMOKcXCxaZJatxbmMaOYcQ9kkTLxH7NRCRS9oxhx
1SMkck8q/Xypi3vYnuNVWqSjEmguAZkmyU7AOLaBtBVJ2ELc98Ix394P4CXNxnoz
KtNjw4rczxQBhzG8eV0NP5NeisW5lnIdvgD6b4Y6QxBzPUSRCa1SprFBnldDoUBL
My3QBPAlnyau9CKbET3pKrywGO3Vg5ExqzqHPh4/t1VwZDArYl9G2sndkLenvq/N
uf7tPMfkG6aCDJNnpnaL6rmpiXnfiZnUwk/SAfjwRoyh5ekIoNDwWx7uu0puxvw+
pg2Z1H5HF9a4b0nA3++gsFQVupsLcuiR+V8bZdtKP+GMcdKaBv3/e7WUiAZI7EFF
xhfSfvrLg7G5CB4V1RNY2PS09nNJ7JQkffzDDLFGudduzu19yqv4gjlfAmgGy0QO
f/wri/ZVmB9cMZprh8iwxuTlxQc+70FQWz03vrO9ngotro8jnY21U/0wG/e2h4kU
SaL4E3PvEmdp1oWDYHXTUMmKuxuOuBIf1NMR+MgsJeRKnoWyXIVR3vSqLjHXURMH
brMYKeac9NQR8rGQMa7u57OpR9F5fJBhIn51FM1cgXFPCeKS1S5uoUaO6rV+oLMm
QO41EnxAiCvtL1umopZw3DQNaNy++jfRwWsyEfY72ZQKuQTzvC2cVMVr3T5GueOl
2VteYV/Eg8jTDKTFRR1JKywh9C95P9O4jfDzSxDest+A96IlERAQL526VXLxAxx0
DHYj6UM/Jn9JdZAqAfq0gpJboSYCMZj+ruXGvM6dNlg/lCfzgc0m5cIsuc0PMm83
5Qn2A++HofYqINOvqTdp9Y/oyI+Y/syo+M7StX7SOFHtjU/fnyDCc4IGbTAge/3R
0H+Ml6PmhWt4zaH2LeXKq4HBKgy8MvoUGMwnQbIDQsHbAf64Axx2xLX6QKwbkIeL
rymXVrVzCnp0k5OwPOd/eTM60vbDXetsxsqzKiYPtW2TFTyZtlqzC7REPWr8XoEp
NqWnFnyqayhGHgV8B/SPYC8B+deSGPOXPdnXVDv919wKI26lrovzsueuEv3tXlm1
A2pGSQul7i8vq3L0VRKG7Xj+yrn41g2gDmniqOjDDGX8/D1EyRgy6RZsnAU85kta
Ra8W1DTSBGduARDazJXNpYhCS39gbmUJcL2ZPlKWNIsWb9pjNHJ+BgGc4/0+8Fh/
58PJS0KsttQ54JDjwL2cDo1TAEGp9aSK0rBFKZUWnHTYA6uoWKvxBm8Bqc3kRyxs
TGx2TgNbKEUSa6kGpkKOeSFuUGKT/1JxLHIE2rGTcFY5Y2eBM6dzey8Ps16kXauL
252uHkLLQ/KNfi8rrXuj51e72xPzDNHNT3P8S7ZdN8CV9rsY+OBXvj7pg/olBuMA
FGSGdXJvCB9iM2fH354pgGSyUOywBElQTuHgdLNM9Q4Lx7gWWcESf3NXTwTRX+LT
RZc3Gp0bmnMIw/VzuV6Ur8OOpqRddbjyqnCmtOTRnn727BESYyqfQOfHuukaoyae
EpYX6DF5m+ZL2kkEcdRXCMteLylQ0xU37mwoERKYh6ukpGk2/j33nPM41qTvnOj+
kqnTMdODvSMxYaokTBm5+L1DrOYl9B9DS1Lu3DS5VLOYe9wX7SOBNsOHcChecwSi
m9gQ0OOeXUA0TdRNSrw6hxAbVBtKnhZS5TozzbJhApdvokuHmcNVQaPZhlaubjcX
y8Q1mlx6AKMUEyPYvRycutrC77V8OslngLAOmAPVhDwdkeSrPvd9rrtrw0fklRRA
oAvqfhXjLIsP8J53MNWZ6ABsKF/UFzZszdHnnitlzXnInSwvyrKHX6uMab/22cKm
ZzR/ja6WMxEp53YmJnDzkTq0udc7n5f+BCdgJ3pn4M7sLFmnsgUqlMW17OXxNkLc
7sYzjLDsbDJ2SO/FcJxMXSiPVQZ06JatS/JL0bf9CpNPGxJ4tD3T1YvrdSONfujT
VOQ7blqppimwY1z1E7enqaVPDH/9Ah1jUurt6zSUAwr5XCcrH3bMx+nDU2xS3aS4
xPajgsb4rmKtD8p6wJ5V0XR2B3JSOkM4qEgE9ljFoZb8GSpVUxu3wKXG0UrzZrYv
JpvlSeSIZjEIRgPRgPmqCuXwpNJtaRzKLN2sWyqj47rNYxH/HPXUXBXjRJzgL/Sy
KjJVlA2uARsjSwW9b63/F95R2/ot7PnjpY60Cz72QxFiwgR8kS9Eq7g1iM/w/eoL
oGih6KKLUuqZX03IM5qWZ0f1ZKWvNv2vaowoPiqQbLk2/CHmh2qSrhucZIPbQgGx
89/zl3j3P+/mmZyF2L9Gyr4Vt4AxqZSv+nI/pk4vVBdR/EkAsUgiB1Isp5p6+487
0LLtZYuCBYlEcmgeKZsP2L31juwAnyfwz0BRUWmpEEAwOyho13zo6jM/heAHrnbL
uN4c0MaRgGHq22W/kN0XKL6MVWK+ESV1RDpjGxw/9ISsTnC2UacUPRdeuB80Y4Xz
p0z90Y96Iu9D2Ut9Fa6QJ4DI/tf3E/tJGZLfZXzD59cAgF3LAPEfyeOmMiIkSxiS
xGh8ZLZiYtRqrADw1H136XujYHo4dyC76D/JsNB2pIfcgooFNreIfWG+GufGSEwB
6bG0upYvR8IrnwNn/yvS91iDG8lzjctnqk8NBNABGvgOAZrXj1zLoDJBLpiL/8qh
8K5IitajfVUr90CdphX88tzqA/3xOX3hX3PfZ6qb+90QRg0CTL8c0kgsr1LlKoO3
CtLt7Yd2xaUt/+Dk5FXrNCE6dDY4H4NrJFe2brwRiZaBIVLvVbVjz+4UrjBZyTTU
GoHxo3vE4nb0OCOTw/F30VQ5RPBHVsOiroFU9MjAOBNNJPLPkmkslpnMehZZk3vK
c6IZ7719igNE2EI0HgrU4+2ZHlCwpojC3I80pW96z5Gc4nJ3Kjc5NL/WywAomXIT
jWrrdgL0/t/3zSA+4SUGyTlHWhHOQmRRAPVNrVBfHTPsumL8ssmPGiYi+2gbn4Qh
FRW8Xz+IPJdZ/TiLGRB2eKIOEy0UTwVZiIr+xNRDPabcTCx7lNkr7xVfMKco+BXn
a4di82twEFuy2wyHS6FVlRZJFKwLG5+Yff5kEdvC6qaxGa4NdlDUQqAV+xLrP5eo
rkgwGTpElHsN30aPK76hKMDeot5sXFhcvHh7p+XYA+7AhiiCAEhPRS+Fx3ksOz4W
HBB4UVR4XLayiKVRpnhuSV5zw88Gq+VJtUuGTPI3ggc0yppOXiPkwdn2YYm3VYBi
GzIlDTZYEuTtM/Hvc//2c338FZ+3Xy+m27A5WCLVpaNSpQGIl28ge4NT42t+x67k
56CwFKOTXcV9NGqk6m9KB2HzGvJ7FGvApVxM2I693hGEetuamyGiAvSIq/76x0w3
9C7nDfc4AbsL65ky0rnPScQ+DTMh/AyszbNMHPAuFuqYJrAUFvvB+TYBZHrZG4ns
jjrklViT6DVp55NslKDqEmw4lP604FHPtoo89Fpb8ghY71/Q3ge5JEpgS2D+K3vq
7Hxk+mNLBkVrrT7OATgYtCA0Rp8P3HBcR8jUuKKNlVRYfr4ux5Zh+ma59o6v6IPo
QIRt8xOzyqU50C983LUt63LfxJ96US2avFXpNhwcQFWsZ4LdubNNMz7gTYQT9Bd4
u55aZ5yUn/GRh4CpFuhLJEWprTduhvk6S6Ag+4GQRJipjb/gxJrJSlKmBbuhU9H+
zj7HYibPK/zpqJVCk1cSEFP6fe+g8yoUX5a9J+6IpXpryFrkpdk8j9dfMlmzmCI3
ZOVsA1bFUwltTa2Hqkbt9pRQOW4afO2Gh5h7BLUKjzzY2PdR4/BUsfYv88JdR/CR
GPMHQLkTo/1BGCpzNukh+/GQI6Z3titVDpAvt/B3BvmrG3bMkUmfHOIxr6Re0lZ8
s7Xso92EQ809+aU1QD+E6roUnpQ2bWQ00/35tcE3hv/Vy0NxHI3Q1Yc/50q/pIbH
pzAYQJJ6HJ90Szdsl1Ic+3FYbhmNEXwIVMT7+XaF4bFzpyzhK/T9JX5G0dwPcECR
GaFEHyMN9VmxekdjGTyxSX+jQ3svyJ6qrBCpD7CL9TUqJmxt/IhH9zxTWnrO9hFr
gcm4RYK5Ia2KBrktzpaQhsh9bzalJJuh/oIEOxTUu5+/K3capi2usG9vQ4FC+71P
tMT7hFk0nash9aWUilMMfY5KV9bq3IzZ5akerijVEEwj1NqrjIQaMlmVVY0XsyG5
k6Az4z6EdKVpR0qpe+r4iMG4CsgYqjgfSijWFUZRNwgAuMwfvIxRRAJmV/dV/DgE
iQD6oXctgt9tBJj3EWvrnK80t5jzwPxzZqz3K9/TihqAN9EKq52XHMgGXN+en1s/
SW8P5Nqd1oHhi9SbG243nwZrfBwhEIoXxT0AT1QO6YuWW+YaQuJUFGsQnLIM5ZCd
BwU0j3TmozS0G3GBuwYIQt8Ef0ORxZoPhYQBfoi2lyz5VMLz4VPGl2B0/40/Jtb/
wIWfXD6ZFEveBrGh2GvdV1qNcQ7af/P0FsU0GBNOvo0bkmfmSq8dIQV6Hz2k3KMg
JmviZM6MULAOBp44ER4k7cVcU7vCucUIyUzLceJC2DUQpeixT4BKDcMgTmnh8Ahf
Ks7+Zcv5HAj4bGPyo97bO9a+Gg9OJWJZCmkB3tZbY03/Hxd14ZiVsnAp0xs30gpo
VF5IVoWt3HaXb3uJu6B1JDM7moEbUw2++1k14hpmoSrJUJV/2BCPRYfHc3vkyJBa
K+3LI3/gUohYIruKaZN/QIFWfof7r5qnkXer1aE9ainPEW3hut+PNlgP24ajgAvY
UK5RRkWc1UbsywaqYQfRCIkyZ+mZc/kzq1CACMGStr6ex5g6jDewsrE6FrL7RT5N
cxIyAFoFiv9IJeT/jxRirpp9Qaf5hNHFJRrnWu3xxBipB7Z4ppQR/0eR2iBxtiv2
iXY88v6cANicC3/K7ZaNF3fnm5zXipGXRyHVjzkVjqL/mPTn/rIH2V+V0oU/erwD
R4BFc70FDG75+eR4a5W4WulDxre/Kev51p0dbTEv6OT5ueFP6Oxle2Vtmz85Ofwr
3FrdkgA0HNQjYGYW6FF+xVmaFB4dHLGkEBsdFP2BMk0clxL0tvDNvROIIDY24+5X
6k9qMwEL69UTG40oUnEyDr9dlZel6usCDacCvZFOHeU8HIjsBAUsdzmAGIdZ09ZT
JAoS6S2gLGs5Xffz4g1A0t86WuvuJK1k9zOfcXZRi+TJFIjA2oJCL3mtmIurtQ7T
HcRPgaOjJy270pfCpD39thF+ivf7XEka+eY2N75Fjnzc9+m8YHztCV4LfGp0HM+V
34vgchmJ/mI0whuhCihiajXlI5f8wmoWnURL27lx6/dCL6GGWz2hiL+e66hsIV7u
VAW8rUbS/J8uR3a1nhU0UFRvN8uJXFpqLHuiwJr9yDEEh0HU5RoyT6fM5ULKODia
Khd+oR5iuA6NXjED8DyChXE2P+MJWy0NXCaDt5ga6EjCpU0YBjwXNkq+7QZEb0wW
NDim/Ga+Ex9xnMhItEwesp80Gfng7sU9LCFfg5SMc1PkS6L4pKXM+KYe3nsD43as
861VRTAdfsnUw3vOq1MYJuqfO+ixXEbBcqDfn+yMqkbRipi6avEL8Wt+zoFC3XkC
hDqSoPtwKzN+zWaQkmtQoXu+AZoV10ybUx0J2vux+oAFO2KxlhHSEaeFN59WMnF4
odq/nael1JCTPR6oz66sHlojRLC5PQxUx1gYhsCT8FQUcUessLgJ/HI7mA45SmUt
D4XrX5Xo+597av7S4PVRR6VmDvYIPoqje7sVfh7uY3G3R+UacwBtlFBaGra3PPwY
b2nFvKCYdSoffDeY7Kn1XEkI4IUhBJomcYDVN0RhpgnMVjGpFDYgutlF2ZSFalf6
EH+8ZL+c6v477ErKgD8qgyLqcvpo6T+W2wE4T1rNV6VWHRD0s6jiWXS+irdrQlBD
BF0R9VCmQobGz+RhiLmE1+MdGj+6rzqyq4YxQdlbAFwLL/Z8Ls2q3n97bIV3B4hk
BUVzLQ2TGb9Ggv9WNlWsvu6O+1vh5vX7AJLYv1lRIgtIPL4ej2lcDnXfLGHDtN2Z
VEqO1d3Ce+byL+fa1BIQ4NTXwSA2HAUa4XqVzeVW7DXhT/x4Pu83GLh3dbWe5TR6
zhcYZJCqRrTkSx6NvTvJBaZXKhkJD+wp1D1LL1CIDvKj3um48vAM3T/7buBrLXh6
k6aVttl+Cbk8oBua7RMs3GJZyo29HovxMqmkAQypVepE/6laL94J+b0QWk0cDAu1
ButGobJXEFtEApLkEKjx4ysmKOc5rRM0NU/adkbK/M17GAkMiuYDT56M1fEpfXdQ
1mNQNxl1TfpwwUolxQuqTqQ0I8KV9+7F1fLJXhuxk91nWbcGpiyez3WY2NrBOMMx
s4LlcqZDC6nTVIvPHAdS5HGhu8DrgJg6LBDMwDoB4odJ6fyCpl7FiRofKEPFDMyJ
IokkCpsJgLvqW16xpH7t9ZurYMXfofZh7g5sZphPEoFgE60n90tk339kZkGao2rB
7JEbkBkX7WcQBUaW7X+c3U08kLd/hQ8659bLm1xfNLOgdctbCg5crCDZgQg7K7mX
284VGsKZM+3Gtnk2stDtpXYcvmfvAR0eQW2qmIDZBGn7N5mDtxzF/vyhi5FeY2Vn
6iT0x/kCBZv1PswM1ZeIUT/K8yinScd3y+vt9J636qmZTFJD6bcsQf7y3q28sh3V
ocYYs3YDZCsDWcPykwM9gKmbxKNn+rSJdH8swA2zcwGZcLYkri3gOBB+ldcxBEtS
ZmMiOiP4jpk0VaNEIbti8KxllXWlAsk1yBdGtlHkdt85dPafm5gOo3geQ4JuiV0p
3OysRUIUwLQzg8A4eZ3uhc/sa5KlfNx/I5itrtBuMmJBjjbHY7kyzxvpyEN/XUGk
BMj1dOLJ5EEtyjIpNO6hICB1xXa4xpTsaQHEj90qUcocAlrLfqY0KkH5LLaCerPv
pk7KZb8l2lydYxDBCJdhI7J233IUC5StoJKAotN4fRetLqaPz0URDYmdP+grr2Vl
fb2xbKFF7BGbwHXzm1x3S3D0KHq7rb16ZitHxIcm3sSiIMjsiOJeqD71rzTfN0EM
w6okq6jmi5HvQiM41nBzZWk0wBosYMn4XPQ6w+5CuydmShSlbPaEyxc890Y03rDr
vY2ld2IIJtqi7D+5C4IqfIhMXVHIsqr46hwjt9EKYRSvTLjTprA+UD2RKAesXS4l
X/yILL8k7dLaatzXIsXlVvUgUz2mcUUVcu22ppTey3Bhr/WfE20WU/65yY17wywM
HrdRp6T/uXujUIn8xSGGGmNVKK8CxfgMlp3jqYeYDKhrz7D4DrRmyHKu7n6YObtr
TXlVPvxLEHLQK3jAEuVVAFStxPkRNTB1LWDsJ+9pwL/NXNbpPvRV56Y+XZGb9FLh
1rgZEDs20HdG52YSUnAQTRs9LmcGXpE0U/1LBXuUaPKLoiw/fQX2GXkmescISNMN
nsyI17rjAXHKIDrdgnTPKpGGsRpi6gsnAsRx3i9Tnq7pfkIRugHqzxQjIl3nDo0M
CWe7cOE3BwKoT3Nwd7qKGnMptJttlrI2JY7X7L+FI6GBeDV7HOnDQwnAEYbqzBzg
iJNos6hUW6eXvuQJcD3D/0SSM+w+nn406iMhZd5OcFg/DXKdaRrx7cyRj8gGo+6e
cU18PLHD6C3bW4tULhfBJhX0yF4Clqu5Ta70N/3hHoAZtFOOolhK4AtFmTFbfKau
TXShhpxKiiHIMBPFhukA61H8JG7Czm/tryRUPge88dUnnOZXqz8RSAq5DPmY5lII
zmBsiiqtkJURm95MVwez01+MyjBPyfQIpnI3R8OTcnCGYd83Mat6qu+pNj3ZduMM
tzL0gej9S0oT9Fzm2dDJdBeWhaVY4RLnd2J81QTr/b4tC3xt6IzkYSby6aiJtP99
rHBNcOOHkBNQ0X8rjxCZ/qB3eDzULMHKg7g30BZct6XCWhqPEttZk+QvKtXZLU/u
Bk4OiKQOS8/jX1db7WiuJ6BiDhVdzReFYVhANZ5gMuAl1kdul1gmkpD++DUIRqXI
IMYSOV4fUIuKkJ0KaKBTgrOUzMgyvL7fNb4lfXObr6b9rKqd14kwzSMNuQRIiA76
v6Rn3LLNCj1qjoLgK2JpcacujApxEMJjHf6723p0aWKHm7tTtSALmqZH0PnIc4vk
Q/JENjYpjBnEQs37eHnBkGsYVRxh5WMrYppZT/f+1F02Aw24o+dRX66lmZW6Z/r+
wh1/BjXU6KqN/iMGdTpx+a9Qt5u0iao8pjfuGmMKVfFCY994M7drwjNB1SFePGVq
A17n5wo0I6fa0LLqfOg1bXuS3fOJUA/LE2svaxkj3Opk03auqgW3KCedaanhJath
YS2wPJhdAtWmy1ixIDCXTOe9OAto2mYmmOsA/7kaTDRQSvjoYqqicr8ksuQLvSFt
C7H/vQugD2E08HwS3vMZ7hC9e/bOc1wn22vOQtA6YK4DUxO2oymEjpkpEGP5N8Kj
4wYNVz9CxNXM5V1A4azCuflzYLdSMEP88TSs9mU9NZMXVS3e3LXkA7h1cBgK4vge
lpp45OVwBoDq84KsW0KMzv2che7NPuho+bxrJ+LaqujLLMOz2Ox9ArKfowm7uvES
9yUICFikm0hH8XHSrPcC907dA9JJ1c2OaZHfmZRQP5TXd31GLhu5c18GWx75nIvI
d1aTA/VNgAObNmtWm+d19UdKVzACUIIolEphXAYUN815SOIeQMdtgmyXVfgC5usI
ybQyB5UzKszn8nOlB4zqfGXwt/AUJyAe5cMNAIG6S2MQLczZXXW/29YZZ9q2eyyN
4orkEAKH5u7m/X3l9vKnDND3u2DVgUGLs6CoGbxEPhIE43UUhobxa6fMQ+GhLWlZ
XU5LVcK1jYrxxtlpBMC8tBl4uMMcmaJq3HlQHffeCjKTfmpW0lrjB+6XTIVkfuqn
XewGp6EL+Hgft61c1Q5sHIkQCxVdMkKi9HkaYIBgPtWR0eYJX8tuRsF2tyFzOr6F
JKbl5QPziWM62/AYfb/oE1VjnZd/ThNhMCYMmyy395VSwQKLoSSNY0XpVT/Mi/We
AjwHEOW4Vnsg8FBAc6ElsSqTePTOF3Y/hKTjD0BQhIdBc73go4jJDwUpiaZXrQJ2
nOPSVcPDzrjcI049L7TyFaReP0w6U0V74ZthSsQ+woo67lcJtmr5SQKfU9k8fp6M
NBChBeHkxD/ZZZGco0T5d2O5HDk2O10hFYCbgo6ssIo6UCa8eu03r25+8GUdmyH7
xjzkpLRUxjXHCeToXJsoSX1/7Nkhou53ppUvtO+/sBxlXpZpngGPM9tu1GRL4M/x
PawURGRndshrDP6gNzyNeBdh4zO7zvkWTqMwnfOnzkyD9BfXk8vnxlGEfaLp3Di2
ESAUtcn4j+S0F2l1g3cNygkRkZawLR835qRQSeUE0QLitULjvRs0/IXnC88QJ3+P
qCXJqw3fDmKHEjmKsRDY1LQgNLmJctBgYCr5syFadk+7itfPVb2KJwwK8gyBs+bd
jGB25Q4ZYc/zdiQOX00NsWWscnPZl+FuJsAQWmXG4AsSVU8AcmLF7EdwmY4QyrlC
XHXUF/1/+UD54flkXL8EcA8DCUj8PQOpg/tCVT+C8CkWhUhusoe/kvKNTIlNZo/s
y48HRKuvYsM+xiNF9RoMmUChHFkEfgKGTe2W4sodCVRcEb5jcUEjDXfSC9atq6FH
OEDBwe3+HWi77A4tZbXSCGIwwzC975ZlL91YOCCBF01jpiBM/cDd37Z/iC26jPCQ
mb9KegrXEBACdBpWoR8x4qjPpDFgkYpg97MZJj/HGEe2zUCym8X1ywP7brMvVUv5
+I0TmWioj1yS/5d6NsoNnL1225t5jcP7l5MXjsRhHbeivXUo/u4uUpwTQ2QM8n2Q
lkrxyOr4X/rLXPTfV6cz8fQIzmyvaCfK5LgEWDHurbAZDxRd0eDAAiGddvMl4NKU
Jyglaqh95BTs8kCL45joNblhZYUpTwz2d28/PSRnOWG/ZRdlmJm66BwuDOfdPvbj
ukDEcCmzGAA6Fe3TtyTj63+ELINczN5DdLyR+d/SbralWe984Ea08X7Q3umRSVcf
jhXE7qfrFLTBWanXekhj8UOKLGvtKi39zabQid8OzkoU8mjeRf7/CA5lboner3oT
Ppo+C/gLIN3c4jRqml4IR+zqMKP8hiMOvYZQIPzKKKQlvjZg+NQics6LMshCG9ve
rSYLwh7a9PEk94eJ7tcYgix3qnOj8aHhgKO0RPpMs32DeQadFHC2KTye379ynR+U
7ntWkC5m3OQ/PrHJzWfYifGk1ggZohuhRsVdScLwFNu06fBYPrHiTMCgieHH1j2D
AaNBkoDALnrKtBw/LcSmEES3LUpoepUYh2uokIsjfpmJo1Rq6tOi3AgyX/aR5IWR
DJQVU3/tIvK/ftmWVc8aBp1S2tmiVk3gDYQCJKmD0QuOaoCyDgsPg/OnxRxXef56
3g1t+DvJMr9XDJF3Zsp13M5RNnK1DhB6Stl0yR2oyorFWrQv7RCI6AKIYZwYJVV8
ksUvWbdjSQYbbpyifOCdA+wP4AQXPjZic42+s1zWHLQjfF3CbqNG7YM52ab3DnLK
kvBbluC6junY97llhx+MX7c8UJe83+dm3HUp2swYTFHpC76zNOMmIpz8vLvWgoWJ
WocrRdnuunT2qD0uLXfsPrnUuPRAu27/7N1zMYnG4Q8B+BBgOAlq+lTQNEhk6fXG
PCm9i5bueUQA5t05Pgj/7q9tLmJrzCKZdwiEIqJ2TNAVgX+R8ke+F1xTAmXFQBfB
ymuH1n54MytwM9kQPP6iuQEbggsOrT328vQOIm80JOA8a1esSWRvgPsYbeEpZnzF
JW6VeUGaOKrDOutLL8ckbuWSAdhfXjI56X8atJ7udYkRuTmqqBn1evlcgt6dZRA1
JgPkKkcdoA/3zq3vJGynDYE6EV5hTgOX6qMjIAJJrOOjSZ9XZjGM8kmO2cJYJE1g
16fGSnX+ki5Rjg8mjfs12C3YJ2ioP+nqOUGkuGIw+6Z5C78Be8ta5qwVY9PwL+0D
KFjqqzdi7pxcQ06fbua5f9YmFhjkdrBx1aV+XHXVRz6E0DyQw5S+wXVJCd+IEST1
lKVjZGJJInKBiaMfGVq79yv64eKBKOhi2h8ixuTfJE7s7E3/Kk4TGxjZfKhrJQT8
e/oB30jJAnz5L2Y2XFD09yFLDZ6Id9U7wheHAYvHXpQ8t2oBJrplO3pBlyztg8m2
rIkqHAvFH2RYqc5HeI2HYVamoHh2aTQn4lEXR5LD208FyYdTYZK7CR8JnlfRAHFE
mjCKz83hVSC8db66Ph+6P7PDaSrietH00wMonNrxvuBkzz/LrpACg/+rHCWt2631
rsPCGbGqrVXmFyJtq1pz3w17vrTsjVGiuyJM2aANbAOisZQyNxRPaKXikwPOGcv+
JKmgjMivlJVEKCmHeUUtyXBOGujzYeLRmWojQQsm8Fvxl9ByoNP8P+BsSTuOqF5V
pDLtZzeex/0paow7SzCvbM5aXxrX5RkZmLCLGp2J8XkOrgJp7ch5UVZhcA/SskIc
hX4mMG8M0UdDlnTt3//ykPhjwziDBOUq+hTBDyf691/rw5EQp1NIimnXCS5Oo+rH
gMnxzPbB6MB/Jf7ILRhKNgY9JWPwhwXvXRI5ngcluP7UV5Elsnr0SuNLc3TL2ewA
RdEMR8c9kLN4iOG7eu6B3q/cIEmdqc6OtOJ/sDWhRDXKKdFwCMnFvuxTJSFsHQZX
VVuS8/DJDqqNB8JdriOntse/hJm8Fm5UxZul6KIJeUstDI13Xg57iFCb3kvm7DNw
XLcxn79jelLr9AIwOHN8wv+fWZLlhayn2BvqhRqi4RUuS7QPvyJhamGU6DMD0VQB
66C+CJ1vD0K5cTZDIR4BfvUNHpebuKXVbSI3kKltUprd2cqhr2V4Q9kA4/Pr+fKa
Bl4O1Wg/nxsYCj89wxd+1cvISavHVou06lPTjjaUPv5gA4HVVt5Zg069J0bRWvN3
f9BvmgYMfl2diuNUmgBxcxXMxsSJkbxo56GhpOUZFpEvvEFwPfvK6UhSapggjoY4
OsFcIGuSKGgEuBc0NCW1w8tdxFVqhkXxuI8wJsf7jdHxRaf4qfCklje14nMRU31j
YTbaBq2Soh36llRQXioJKCN/LU2kBx0aeJJ93d8alcWonlmHRaf1+DfI13gw1iXR
6x9hne/kxRwwumz6Y6jw2AHlTVszyKQUgCY2cu7uEmFde0InZMWgw+wP4nPxa2w1
R7UTF4aqrZ/aVGxTZdLAJnETFf7dE0u2G0cc67iZjkjlghaGT7+QjhE4E5RiS0Tb
X5u+S5mLYYbQbpp+PyHEFIKsLzTYITuLPfO6DHvCKKgl5EqUCwLbHZWGBQ328hn7
iGBzQ5NdCK2O1tWjGA0sPIitukdJKauh2CTeDWqSn0NEbzCp+Ay+A9AmYhmPNbCH
uFOONtRW4fkjC6mCB6F1yp2W9Q8HrVrB8q52WkNxr5ZG/DYoLQnBM2FqMy0D1JB2
mJWm7Y3cMpma9g+ItJoCZV++Rc4ylXHemGiK/pxqIadRzRFo7xobboXRs83NlZ2w
/HfGztKMpShlr82KTOZMqVLrlkaQ22r0ybsV+ce7wM+BgZyQkEHfMuV0pVJ6cKLW
0l7BzN09GnTbbdlCinj4KVwT0WEQ323MhnMhU9RV4qPJHYgVGxIIly6Xqko1B7Rt
2jdVEE2CPOYjwhR6e0+fVtnuOUYs7ZLqdHQpPi+GxN9UrVBBJOz9X32byLf3MJ9k
7j++PXJnlDLitgjVK8Z8TJnwicsS5FscUi/UGL1rSW33MJFc3t75J+7TpO4RuKCj
gIDKSeLritBuzOkJm8KyXh5AmIaDzW5wlfigEpe0M9qTELVQh6ipetC26VV2IQrr
ycZfi+58hXPGVdkeObruHLj/XrXfCk/YWdeY4jNQdSOK4KBc1ruyKGxcIEBdq/eo
EYlB/o3gauYbP359sgnsjaYL9HeAx2epPlkHSqagQtnyZj8WzySXyVSnmd1HdiR1
aMTF1PKkUUIyclEbn6GvhEGNHs0Ow7zZUdFlTJRtuK7Q2NKu7QiTXbmfjpHGgshC
PQRSe2g7ogJHJrVTzozqLlneSurGy3XFLgnl9rs1zBTaNBIYSw99VToamdl4GbBS
gdgQZrjvA31LwlbkhT7C7blqXRDZcy+3awnJhmVtA/fwP2reK3SOnK1ze8jj3Kdk
dmBsNGoErDsqk1WpNbliNSWTBPv9dEXG03QSL5x+lgqj6wdGOA+m3Nn/ouTtkQq4
TQUKIGEcefjJAh6VprBkxjOFurRTCO5XR5qmLK2nQ6qqQh41nW8UWJmAC8KdrAFo
vk2xcBN4gw1vebG+DZ0OOoARy0Kx7d4ny8UPjJuFC7YtB9AIDcrpkNW2jwSEfhNn
t9hYEVG7rP/W593AYFJjTKAhmNu2ewnSIg5MMgZ/vcuob6clE7y+eU2lOVon1gCT
wtxN+nW2wvW5Vow4W5uYMLBCL7+CORjOiobhkE+LMEFXQIZqDUKshaaZQxeujaHN
NdYQlF+9C+IF95wV5rnqlsBWafTstm9zk1bJMHQ/i+nTCBBN7Etx9eUoJtJykVIn
LYJKJMoOXzsj6WQHNOIc6DsH15N64S9qbQemjkr1XefbOCEd4fDbM9HKuX+JqQUO
GCbL4EQQRbX4s6dqnA3UtaxEGFLWPyVyRwiMFrz9b2fhqm2Y19lJZDiTFmu50oZF
PWNyq3CeJXtj4Sx8e1y34ZZSHNGrEPPwdQsyriYh5zwF0JtUkfhJFgGRpvDPI6Pj
ot+0lBXA3HgeZ9ImheN3pRhsrb0TtE51P86KHTxanhmb2Quc37EggLkGouklOAh+
YkjdvoAMOhzEvNhVTGqMtdkHCQLNman2UKo/hfeRpCSLzXFqsNoHOfKCl32Mg7aN
BughIXC/aJ3Z5+0u2kbm9DoimQKwhZGmrmE0EMRfJ/99UErc1NWuzi+sGu24W79S
qunKUsrOmW9EiseRSY5vMcg71UWUJVgQ9skfsdgCgEjgHW9jONZfGg+uQFstIPfJ
t2AZTX+T6rsseJap5FuM6jyBg8R3/rkn+iptwjB8PSgLKxgD/jbHr6foLiTK5EeT
U1wWdSP2fe+ClZ1K79GnBIOFS8NepnSbOveiVXER2ovFr4z2uaSVz1GtW97DTFaR
e04QJD90xBfEM14xGThNX0DZSIkkyF4aASsxeacwm0BBHyk6iulc2mVmVg+edQye
NQ9Hg4ze+toqtzjmkyMB0Bqbloz70E+ARCmQKISAyV4va3ttp+0jbxtuVLMsoLia
8iuYl1j2/8Ts5DbP61U1xI+n7GieWquBg7f60O69IIkzC75yBh8wFWD9gYoy+M7c
w3wTDdagDDPRmBrWfqDzoeqPtZmKdEM2pQW2CU4siiwrQg9Wn1zlulJYMHbm3x/7
wyivn32ulWajHTbAJFAFUJ8Kizp4xl5FfsEwI0khVslnmt/foXgz1b3Yv4S0FbOc
7htzrNRoN2jquOQW/hKWq1IGMxIgWgZjwtaZ/NbNAm7mbzAIoYbuaGkisaD2vdoc
FC5WjTHTGroj5nm19GZW+A0q60CXEB0oqwNjywMb3qGPCWpO8F9Dz1CrWRh37zDM
w7BvKTD1zHIos21xxs1PDQ98t7vOY5SuP/IlQLm7ALoWaZSu98Sd79U/hROss5pn
uIcaZ9vc9o3vPkngRXq9tD91trIVfrnLtKkLxo3cJEuRlZ7E1uNowanYEqffJCdi
Dn4ONVVKsMFZPNMVYz3/dScd0SsH+Q0hNENK/HBJF/h/8Q2X+yZteIy/7oNyamMG
BVE+zzDuAFbrW76O0K9euyChIlDjCpBmcMsd8jCrVX+19Oe9ky7/dCEdsjDjeDrg
jr/g0QfGrW91a7FcAy9o/s7AGNm8SDZ2FftisDwCJORlfmUEPJWrdljryfrevpG3
ao8ke2qNqTWD8qTpo11NC2G7mUJUVqKFwbI1z4kB7YSrmlp1ZeRPBynqzqdpJHlu
hqSj6gpKnrOnBkmF5vpsRX1tWjRdmrrEZm3Bsfhu+pVPN9UFWcrbf2z/64+1g/Bm
OsYx+2GALyDjtyLFSn9gKs4/0AQk6Gf2kKW8NZB9zcTj+AiLdg58Y5J+1Sh9KWZu
YdjLFPCKv7l3ovGDITfmDLXPPJa7sj8zaGlozj6r3uhj3qjnfwAR01MmjDXC9H7g
qaGcTzSsfVPoZHHxySHXfPu80GcKSnN3/NHG2+NRTzUy2cFUYO+m+5omVXFcAfyf
wdlE4832wMh4s68L0wWy1l9dL0TlwqulQehdfsTAbwAns+d/Be8T5t9b6cadxGAe
6QXcuqChQFDS3HSGrE7j9de7+eVlYbnSzX+xmMuJBWxGVwzxQpw9dcFCFqzckBFh
dod59O1cMOlFUh7tFMiuaJgXRD6MXtogkKV9csYErDJL47zAdFVsRcXzRbIEO6t4
QiNB5GO9S4kZw5pwAUL/DVhKdkjpMnocLYQTmfaFqfcNnh5C7IKLPiHB1BT5045R
cV0X/W5ZpN10er6BwRApageW/9GUnvey7HEZVHJbIVriGn1sCHzbcvRia24ZOd2r
ZLHE+NzrQrqDJNEpoXbSnUHT0KjrBZyAQVNLYzu+Vn9rbH1xBtvUclb6bjxb+rkM
e7/pUUSo4QiETFwItUDW+8Qn0fEGo/O4i6LbvqRvbB5mu00DW6yxzvur/GJbxWLS
sgs+mL+jI22idu3JTG2tZPGctr+mjWFDzZrqQm5xKoafd2rc3rfzXKASLWpCWxBD
l1m+wqb//e9tJq5wrkAgA7vwad6fKQC54p4JvmO1eDmohT/vjrzWFPjy6aikCgJt
RHIquOFUN30FWZQsFRmm0kPW7ShFBplwqskWuFcAXxtgv4eHoui7B8JIoqZ6WqRa
UthQyIpG2F088LBe3mGZjKwx8VtiGHDNG1kd8tIrlByUwqZ5j5tRaWhpw1rdECwW
5Q8+na2IzU8ja4P0H9RQGRdE+bJcak8E0OxBXYCMpYaKIHqg+9aFcuYTWHrp0Mhv
4cZg60HaIYXkCMjqBf2Ncoyaa4pRwUyayYQUcMdXJzRC7v23dKfuqddkpxvrroUi
uKhJp5GtXHBXOJ2Zefn67AwbkpYCuWOWY/G4XazjyS0oWr1TzHzI0hiU7QyOdW8u
QYfYi0OhNQCd9bikfaC6MV90we+/qNZVSjPSqGhYX93OBL4wh4hRQy+l+gtVR3UD
J7zMPcS+4Losl9TG2/YCylIrf8yDKow7poidoUSi2iKzkPZsQQszFfDD9QehVBrz
ZnU4SGy9/vUxtV97Aonc4/C7kf30tgKSLXkwm+dj8rcrMmDYEuEsAq6/Ep4jvw2Z
MKW5dLGYpMMyPkvlO10FjxAcKKTNeYg9fg/ldu7r57dqfIf8sisff6T6Nw1at98r
fnNqjul2I/L+fDVS2FeqjgLwc3nRgEvvcHK7YSn1gdHJXRHZfUHefECU1bHL7V+R
7Y0kwN33DZtFlNOt8ajB3n41lwijRRzJ1CDWMMF5bi7TF9Qq0qJLCfkl4LEfkIf+
rM76GDCoRhtf2VWACQErQ1L8OWC0Ulcx/Bt+XxCNeB6kKtww3cdT/rSw1d68HzFo
xhcKW9oIrrcJzHvr2K3mn5iiE4REZeH+Qgq/fHi8GnLbdYSBY2dkzyYoQeWlv8VE
bifpuduDSjDDovhecH2wAjEhpZu1jk60N8Sg010dP8ryo/wj3lCRgCbUEUkYaURI
suLPFfy6OwCoBJE3gWqekLgI9BJAq7A5gRkk394M9pw4f3ka+nymCOXrEfk2tmYf
zGWyz3U2yNaqv5hYM7PzdxO9b9BpUiw/hUqDTU8esQaFO4AXhbwrxjkdRt3hnRM9
GAemvNJhUnz/A/10wdVHiCHGY4+fE6+1ZxZIa7BRfBxn1ZqbxQzPrvQAb0Aqqxgn
2hu9srYPtCZYjwWY2mIQc2NfrgWmaL+P19o35d4KpDMp2g0WN2OhEyv0RLCvSmf4
b3lVH/IxFlMYkPdBodOqAvRyXqEFP0R8NaBWOcNDmor96BkUBxSbNwDTw4K6U9X/
Ab64erBhmsFEVZAriUEvSbp1K1kPtSZyT75z5eEahTTU6haMuYBEFrghzkG2gJM8
rESAxgaIIJL6Fi+3/oDMkieoXqlOM/kL3qjoCc1e121WuqfnOHW8Rd9p/EAX1t2n
b+1vTDtn5XbMpByC6K+WSaI2xn5k+R1YwKmlnYhqjhZ23y6agyKIOWXn9euqVf35
0GTevAnDaW6kdXZcr2iNTUbniulCtvJtz1YZ92ug/VIQGyRz0JzMGjYeLhXEyMeq
ovOJEcS4UYYARH+mB/KmFGM7rGvE3e+Z4GIOtie4ZMFecWIQ5vVQV65P5uAqj0KM
OnxwQv3kuZnnzRE9WW7i/VRvba2C9RAow5Y9yTirQihPPHdcnhjj8M4oSsROEfVG
GRELBBgLO6UoX3gFihWuREk8Y4aD2DTugiINpT4JdxIYDVnHE5MlgOUUbd4KTQVh
nVA54TAw2QCGFhw8yl8CJ5J0U0PhMbyKDftZNcVjARfr8isTYPE04eLoCgU3AMNW
oPq+4CdfbeT0xm7FVx1tDTaLYvJN1t/XaQb6KXX4zUXVJwrs4UI3PKmC+B8Uh6X2
wqSWVnSA+inqO5sztEVxtWlqrGNX3bHVGYe3FQ7kw4FjgonX/qAgBs7gTRqHhBAh
o1KXYNiB/rmrV9ihHY6bD7A+e1k3TwcD28GKcB566KwRUyvsryjG8hkLLX7VkHye
sCs58xrBEkYfVE1wt2oywoWQQlzVTsGvBydSIhr1KYH+FbmsRmoYtXaFmdYaEvFg
phrnD11xm5XUQyPhrU37J6nPLIEZdhIqdPTOdZu5icUyNOp1YLrFTyio/Wg6HRfr
8XbgDvClkiHCJsCNiWV37md7osKAhn++X6GlRs73ffzN/xarFLyNtFdp8RKw3OC9
pdFbHKhvNOylEGqJarEbzzANGAPcA6yl6D1yv8j1OPg2T3uzjc8GNCZsL/sPqlS9
pMkMbBAzE76NfTUIs2sXLW7vfs+JeP1kPO2jZ0faNvccSTB/AqpL2Z6TzOrWKVDn
QbgaUMleeb9TUMB9jZTzK4wRXyL+ctTeMvJZMcPhBGrUkUmQGGUWs+RsRKoF1quL
PE+AdOVoP7mOt7zY0XqQEF5I/VuE/CQtNIE5w77oRONBcALvED+LCGbColRXSFy0
ilX2j5sYdw/HzgxN9DmDrJNDVrzJIUVmCR+NfM39AEW1PUgh+7JWMmK+gSrOKm8N
U0RNSx0p+q58WrZ+XOQi/ByEXkuVLt1FyDtMgCqKHrLrEGC7x6ngSJM7RCZ5Ed2V
zWnZkcPSK+GpqMFGaVhl020FuMkubZTiSzUuo2Z5h+obiGDIRVPRxQnhs/U7YxIP
23tm1LUqEe1ZFwo4HdSnLztpvXRQz1Y2A3xhh009qvildzIuuzs4/1tNiK+5PO03
RXfMv7SkMN+uq6/CT0rvSGQ5WHmcqr6E6pgMQ5E4fvAnj/VKOqHLxK/cwBLOG49C
fQt8GSdNFWZCN3F4heRh5FvBzzQjey7QT3ObaZP9fMNEf/heh7D47XOlCAT2o2ZV
ReCv85OqPgpc3VDiGia1NQBqflAub7djPHmBqgc/6J/J10kngnzLOqw08rhcF5o+
SHy97CZwQjzsUe9J4BiwIvyXs19qKXK5XAFkooIeaG1MktwDW6VPlLrPjt07MvWm
YskmOeoXddgHcwhNNFUXxY4B4Zs2jftEomCOAGvEJnhUJa37o8t6FypjhMauFPkC
YDOhPn/n54mCekJQjRP8NIxnJGkBPqYv083tDfTwSI3WWaWlEr+mq+Bl2XXzoH6y
mFg+5mw3pQTKidHSQiAZ5kskDFIqgDdtE3E/jQQfIN4eulD34r9XwMgr8NkeHSB8
u3zsocZPvZVYIJDU0QQkBzZNHKdfZpY82YYpj6O9CfatsnjE/Xe3EzujVf/YpuLd
hLPMtXxsH0qp7bjwAoKRy+oSCWFfNNCbZI99koDCxGdG3boo7S9Q32B7J8f2NV9E
cBvGCEC+s9hY3aBMy462M8LtaikUn/OhssbO1PEtHiThEh/mJWqCiM6WVXL6rTlY
ZifX/S1Rsi42eHQjn7F2g4Wo7HHGfEPo1+lekSVzmCg78lbQE8Pbp2NFHt7cGN+T
QmrKUq7N5SG8nqW7sY3OBtMPDjbIxZd6RbwdQCLrYzXZRjwSeMOz1wf1h0sWaW5f
8op9f4GR4w/JjMeAxNHLCPI0r781upzKWwl55kzdtjATK0FjL+IDaTduS0As7uM4
rHK4dE+Uc7FUSnXwu7sqr2mu7ci2SQNiOij2gzZ4jLaZjXq9xcNSjYXM57vr3mUI
l7MRulm+7v6pG8Pt1Fe5ZU/HdbbduGgyb9jJ55mF8x45T3Oadl7/uwkPmjDrRTBo
xzWgHHDtc3J8Z/jWoTmRL/zIsL8kk1NYQ0BQcHmv6kawP8xmQpREsbUb9wz+WJ6F
SiUXlVEPM5pHts522Ki3QXTOV9t3fKfurNMHm0oDIXBiSAsC6BoxeWCTF+Sdef3P
8hKbspQElqJ0ifYcr0ynohlYjFBTXtAhVJMbUKdTtsPszkuGXQk1i5L8lG/umz2B
Tl0gODJu4q48yZnxUjZP+eIZRvJvdlTZxAmYBWvDoqfG0Qu3d42lk24YUzfJEJtS
nB3hqztZQqQyptwY1hEyDXeR42u53Lce3WKcC+O994FfE7ZQ57yEeeBIhQk0YaWO
o47Ue138g3sdM1efvlccEhQCv3Az9tQF9wm2pvDBiEP1Pz6Wzjh3F3o987Lo5nmM
Y4R21W2GyrsLmu1/X3Au4Ik49LUZ2ucdeXcXxSh/Bc7QT3/GxuOJ/qmp/hUSgTYf
RWwbbOUccxQEk1Q+vxsfaS9X88eZhj/2wEgG1+zSo0Cso5NuihiTgZCWBnfje0y4
oMZLtgaavgb1dOgHsGux9l4ngbM8vdUMWoL7nwa9BPVZXKcA0gb2I9e/43hss1EI
/OAIML0y6nN7wWGJ4HzonQOoJbLbbzywFFVi7mz1M1IkdlBTwVbvBJLXPLLK7gTp
hFsZPXSn2l4neMO3md8tEbJhdvuFg8kGvYCvSzU0pb62fhVAjx1meBkBAP92H5kX
6iU9u+zW4wqn4Hk8Gvcxi/OKwQVsoxJ1uf7Xcxmk2pDlUicTMNuUnp+UQUmvn4Qm
sRh6D7ItpKZ22DLFP7SXE8oD4srQEvn3AQLVRA7gWng2Xed5m/Vm+P7Z+0EyBT1D
N1a4aoGHPTmIGz/qLzX61SAwN+Pwa0/stRwP+U7+cImKtjKkUfBZHBucSAQ7qGU4
xTdXpY18jwxH9boVPMWX9shmzSO/onTkefctThE9XQDWbGFcBdYlqH0MXXef7beK
/kBrHK/3UZhEBMPDhERKdb2YzOGeCe9Mmp3q5/BYdBupuxrylD/nM1WiDonqKyVS
QG5S6BBXz+8mEeE6p8FPrN1JmLJwdDXuIzn2DaEEg9o3l3Xycgj3UGFsUqE0d5Ap
dTtNfetJp9hG8CEp+9carIOOOFNjSZ9lQ6HnnY4daBri2TXYLH2xpSgmA5zl1xNs
Qn/dO3oxWppKydyYL2mNqY1nukiZGEV2fseKjWQ//3WnxkmJXMnb/V03xPAlKb9g
F+Q+PwnN2J6LzsoVbLLoe1E9mwfg+How6MXF2hUNLYk/zC8P1CXbrRJOlFOxqlBO
gLU3OP5EGCAOr5o7XZ+zF35JVA/4N3Q8/JzeW3Kos1apb5FsujAdGNcWXis1FW2h
HRJT2RZ1Ak1Nes2/iYMYzV93HRiF+aooy0+T8At0+zxEG4u8DCW5a7WQHO1YKEFR
yjKUzP/pKrk5wBR4RJAtKyx8dusoeRZf29PtM3sb9d3fQoSw5M9coHbRksrv7C1/
MLCt1PgxREZVCNLn5TWamxbz8mIwH/A25/KiYC8U+638m5Ac+w0aOJeAW7aHm/vc
udxIySMxRCXUB0NZgEgH4MufaCRfki3Ke3V0Nr/fIo590oJfO1ZsxUrT7OGKa1Zr
5al6K2gImliD5kF7LBeGAl7PDbAzF6jEqleJEh0shmUiBD9L/vcO479/S+Dq79Rt
aTVT5KQ6smqdPFsX1F0pwW+233O+34vLVXtgwEEb1nCzqWaIgGyo4+cZuFcB9AJ3
iUzEagBy+haKXxUhgnyBveO9owU4XCzzIPFACFPXOIPiE+9TO+0uV4uLHxBRH/YC
ssbOmzNvka0Cgah9s8/mr5aOt3ITs+W6DV6DdD61LBAPp6IHFX6yeHCsEkG8mFVV
Aa5Wo0h6ni7q3gqfxj9RZFrcCm44JEvxjTuyj6Xu42hIEdoe3fUrciQ3TzVaKaz0
OwFXncEEqaVM26a1iHVI8naAt6oHqnnZHFXyC7YWj7Q4EiOUdnKGlsPhyHs9T/jV
OR/SKzAnttl5xEkIBEi35wIrZngq+IlsKNlOlBEQmt3bbJDafwGFLxQs9NAUBJw0
2/V0FmoZcQzq7cLiKrEomoxzj9XdGpUYL55rHRy7EjsQ04gaiusAFi83+bW3G29J
NKjNjbCj326XR2f12SnsQek9vsekZglsyfrE2gGutRh9GsZJsE1d8u6ltWWpsZ2U
o77t5rPXidGd5w4qnNIz3dOF+jz9RKTXdkLDCiIpU2dG23OuiigQI6iMG/faA48/
dDysXEMtZz25riPJjr7Vb/9nRz6iojfB16AiBJmZffNq2wuN7oanQkVhz40fcho1
I7MlRlx1I5usQkd2YtgEMqX39qNaZz5OrBN1th7ioKC96qUo/fSYA2E3caZjjAmZ
O9b+/k7sYTAHqksHq4WxHyvViNLk3sh47l+f2/dnPx0qDuTyUnPuu1si9Xbwn0Vy
7qMUcgHYoR2ISQKaCZhzRQ83nmj6X87jXMcD8QhV3jHLIuaa51LHDd/nwnnMzhWQ
cQeZ+pAZt+lRLMo5XB618dkR9djErlJF5mWH8aVjndT7PoYXlcdlaYBbPYvKR4sw
xYPatwFRUQT0hhDTONIB0YoJjSkb9+Fju8gkZYJYRYXMw8TGiLQ2WoV7I5vKLmOg
bMn3TmB/S/N6URbJTqe5Ox7zxR9vXryiUo15Yv9KmKf8V635gPV1noSasAytaSPN
fmtRp4pR87Bd8Y6hsTPN7QkUdHtf1dHNeVBXyrxAe+nGMOxcxjxKmZ2CuixH28I6
fHZWIY/UynG2lgyKwIamVoRtIhWFe34aIyirM8zOp7WbVmNlD28rpt9PFCipVyqk
bLxGzWvEUfje/Hv1+gQvRED3DExvc+nwPfq1WN1Xqq02zABO4uU4F4bfACo+b8wX
QcPGxOg8EOtRpVhFffSGwGUL74OCa0mCtqpXq2xW+0UFA+WKJ3FovzOJfIZxFvad
i0erXDDycc6fa2Yv/PSPPESvMFFSVNmKBGCBH1ZNwjaRbri3MAeethXs+nb3Okiv
4LPwUCO3EeD867Xoo/4EB+oPfMyONy+GMHnmFteEDclGKOq1Deeg4H0tz27UKyDT
fXazcg2y22I4fVBLjcNmAJ8lF9tMpSME6ppcYqM9zkIR7+atUNcXWJa51HkUDzNW
Dcry2I/079SAc57eBC3jeYNfHTozZf4PBv0ScGjZfPGJ5URo8DYqPHtefuNmg2Tr
FEg2LWByLd17+aHtaI7JACOWDPd6ETAcg/tRL3Pj6EHGNASHDP3bUxtW1OC6IxMz
n2+ZnCrpiXmhW9JoWBf5UvAg+82JPO/OCP8/vdBDPYHr3zpxwujgwSTAzHL14qei
JLolSFbcd0xNCfS4hAXV2ovuCx68rz3UW9ENRK17KbYyoWbvdsmu413vQI0rdMYA
RTpjgYZrx3P6m2pCNIWtsZtenk/lnvm840jySW3ecjaX82FD/tn7h6nTYRGMRwpz
3Dx0sYoKmhqRS/HlZWrFAc73mKwhnCTWMXqwZ7dI3aEFwY79iUZj6gnUUGcCP47D
PcxAHEMxlcSGFHSR5KKBrSSFfZDK32MZ/i7xATMl2INOtQvQSZFBug7R0gaw8ozc
kWrFH4wU1WLyvnsOd5W7Q0LO59CC6/Ci+glO6shCTnQgCuR/RMZW+xGG2WhI0nQ7
zvUrvyDNHdwBwRLaxw0IANcAhCDwmv79OMm7+i4MklBM0dOgZkpbNSLD6RY8axjg
urx9M0emkF6Xw9czgZm1yOBmeriW8aNIv/5zDgJha9V+Z02D6kTU/LcA4bt/uBlG
jIilfMj/1DrALn+xLM2JyK8KCH2EE5+2UBoq5w+Ym6ZEKA9OE71t5r2fd6NIhmk9
C/LMQQvkvfE97hEMnXrhnphYrpd++x5S2yE5IQCVc6nBy+TB1qBJhUYnWNmKv8mQ
icxHKodJ8rWh6WGXh9XJLvufXUFgGMELDFBaQBZixI8eqLydnJYbJUjUfx42MV9j
bx6UZRic5wcVisLqULioTC3BP+f+gQqEPvMXuQ30SRvg3Ljqjwyq4v51fnm20Yx/
4Ygp7ogbewZzHJ6AC6YkKDtwR4As6BG6pHcS7j+SMbuWMdUv5qPCI0q9sW1a1Qlr
kJpEA+P2ueBRMwxsxEYhdTVHsXLXX8PFB0W92eFEhRrhekd9ylRO/mQasncQAd+o
Xz/0D9nUbJPclf/TevnqQDbu3IRGbOO3/Ummr69ZUlWQX+t1rxDncoXzb33kUH4C
XAdbl7s4ltxjeKjHskxLh3a5joYnWGTnHpOnGMOJtvZZmUBF/DaqHabGEqY11fly
6tL868hPKXISZn2HXLF1TC6rtiNZa3M46lDK8N9ErFEplR7Z+dtFBh6ulq2W6WwF
hAcfeMFTYt7Kgc6cATyoQ/g3qqHRmda9FoMpchtPRheBeWw1nNiSHUvZJuZZJ90I
ZkXDmsOFc8KEfq0eGAzpuHrdqQQ+8e71tvs7aU5IH3KBV8H8uP+ttCFIBfIQ+miJ
X3b1syiUEVIY83T0Z/ZwTyvVEb4/qJ+N9DQCRjdjdwUeaCXA0x3yUSPcJQ/HHkqP
BZY+Bqn4o+yNW4qMmpO7jEsnGk1vzfhZPq31k/e695iswdKtEgNXa+N85mDCUKXe
2Za+/wZGTNrHP+sEdR7Dk73XWm5fHX1lrgNR4vSU8zwR7ntWbfQ1o9n9VR9TiQVA
6/anCk/8fP0Q2VxySeAW25y04GZB1vvLvaPSaOfy4PKmxoQNggB1XPM5jDM/e3wB
e+bRs5CZMSuGC8zOYGxw+lb+dyjO7eyas4jpjeufKnnLENS8NVE0ThEtv7kBpU46
Z6xE+BZXA8YP3RBjoR7uXIdcVmfVtV7h6a7iAm1IqWgzfD3WrLUDDTfRHuj1JVd2
2+SwDWDY9HcnHmmIiWLQZgP1nOz6+uzAdSsN3eDXMTMlcf0y5WbT+yUjIPnkt7n6
cB4I1MB0SjBVNlLxIXlvl4oz14GNiRMmNw80FC/fu0kZOQAq/pR4QB0PAlQQx5YQ
W1atrV3t34f0tfjg9Z+qLUG72CAny9amFvhLAQ0NeNQoRkO3O9AOuZkcv7p3qMQc
1XObGzqurV06ibqPLvmYSUob9RMzyRq11weoqqZDsn807z6bsT12puAj7FZytKlj
9rokx4QAeegvvXnKJBfNZWEWSoqP7SnjAy33EbA1D7V2s2m0NZU3ad8y/AsN1vX/
0NK6jHY+jgoFkw7BwDU56NzKG/gCRwAvbXRFhIr3Oj2siZuOCiYd2rsaH5khvpEw
VGINf7htz/pRT67/NGlkeJ14JPE5I6JOX9vsOfJxW7mWLYkKhtGLdxXF0HvitTf/
tMwg1uDPcK5xazK11Wz30rPI+EtRRhK1Cn/jjqiVj3gWRa/tw873cmV39NKzJ4t1
aybtCTdYUcfelJ58/jEregnlLjrga6kHtROWK9O6HD3n+NVy8IvbpxYV66fbAxfq
oHfqUELrLmUAnrJ2XwI4ldhCexAwB+0po5cFI49Um7DwRpQXUJQWi5VKpp9MZgLz
vuR5j8T47Yd9lYWrqDDVg38mkdv2721Tsv4FeTy+MQFPMc8GCjO9uQUwlddfxiHu
EZIaeHlWvrz4QFzeUcFdcqE7UCCPUKKAE9NbgX30GkogA4+v7SreofTlMAaRyeCr
tcBB38+BqhBIxfc9zQKjNEGYfsecn8ODhBqyK4/3cFESg176Eatm87VjBcQcrpnq
jfmM6npRse/6zL3DLGMkALM2/C1Ic/YP6RrZQCeQJbG//V9CXsWjsB1CKfshTCA9
re30/Ko5TG7e7HGn+cgm9Z4iTtSD8xzqVUlgCyvO6XRr2Ru44/P2rfCuGGvQmabx
t9EJU1PqKmdOE2xaM6ybkMKSbFUaqc2FAVet8GxW7zbM1PCozV1IE8Rx2Pi+hP/g
ZKhQyvu9PSeWdYDxopC4D2+MoVADmzuAZbD7tmyukZGgrUNyCbQ6EZIJo45+kWaV
nANtMYKs+u0Zdx5P4UJbEXo91sBlAZiqEhybpO4u/OCm3ZXy520rZ5yz88m8u6Cp
aVe2dnDohm+XbKgi4RiFS3DemSX3nOYvDNyAMYIzZyhOseG/ZE4cAE9q1dqWjIqq
PwDbc8c1KhAby8yKZD7Q7UWCPgI7pJTbLGdr3fjTPSitjpeJ19NHLhS+w+PNYjH3
KOWR9ITEeAeaQ7qtcFq49W3WnaY0qTBRY4YlqXCqIJ0PluWVnD3j2JJIUrY7205/
bQEVabV+x/Y5A0LxeKWEKDzZgw+pZqaNt9N33g5jhzrlTupT3dIpdxiGRn74Y2jj
LZY21wnnARRPXpD1bL17CxC0/4cmWjQAVLMWTnjKxc1139RtSJQT8VsABJPxrWTH
tVP+6nqGL/LqCMazwjmjM9YtAldRL7mHqZp8LrPavwXmfgOg/McI7xrI/zO+vZ9L
fjzJ+u2bfmD3v7Oxjod62DUkogx0NCD4Kjngwrqm2bXX2YvMPcbX2lDyWxVrD61F
qdMQv4167ZMdGuYixvQWbJKCWRjrkykYST5Z54snaf7AVNjVx9bVerDPPyHE6BEY
NsUDOi+9/6kSamcDcRwrwUMQ7iQcelB8dvK75kLzWiHF1kq6F3lokb1Lq9xrCBC2
93OuTp/9IlEkEn2JhnWJgAis3qE9HOnN3xz9IzYXCtxuKz6jvfe3eudxz73k1yzm
cHC7mlbE1UGcFxaM/xb1Rdm4/TpNql7YeG6RpKjB9M0QatUzNNCSI51uiNvYiraH
911YlE7a3JjgqGzN07Zt+NSeViqyKvd9amzaIcWqg+lx/7/QyxdMmOUmqM2CW2Aw
nqu8kWrnK20faKGZuksbcTjjcCF/p32iySKpvAXHaKA7FltrMn0eNGTTNZR+84VI
7TSI2MQuVe03SNHYds6xE+xdKUHWl5BUPKy6Cmv0FB0eIQv0Jwg68FS6VKI0Mp+M
RL89cggXtX8q5+ZooxvIo9BNJ0VtWsW6Gj96EgzbfNj57Eb6PNJpjgjnTIUPuEkj
BFbclJGE+ksjYI8Y06P5e9ps1il4CukcN9S217FwVezqxB18iF9e6UFPCisgpNVb
0oAepaBagEZAz8iphrQvG7HnBSrB4bNw6hhFXJyy+Ci9b/EdO5MT8b1WnRc+okUB
ruwV0N7kpRzXkeisi0lKeYGw8ggsKy61FfGsIEjiL5wjpPL16kdWTiMW5nWrPuyJ
huuAYdtAGR+eOAitQRX6SmRkYotEw4Pcc7TVuUJPXlx61Y899GRTIQW9bUtTls5r
QuI4E0uqyYcEQR6LL+LfYya+SCx2HHbZeuVXC92keETjsK8yqgUmIER8KjC/I2lY
v/kX1HO8VIerFfD3auCH4ManX5EnoJ1G+TddC9qjTha69KpM0M8CCOteh8fyna9Q
8OWllMKlZQdCckvV/cf/gYvQrRW+gFQHEXKS/2kUF/Tc7vwNX3xZfrMEdhEnbI2P
q6/83xylIVNT8l9z1T0+u7gzReR0a/udh0y54E5X1U5NrhAXVbe8sSD1IhfmyPpF
FP9P1IEK5kFnFfqUEnvbD5fxtzoqJVEKz5azjaI/n0WZoth7V2oPioLlBQE0P4lE
u4M07emcGjCGQ6YZHobA3tWbvkO7Pj/NVWmoa5XP0tToGx2bkqXQH3zhHLoMcUc0
w3VEsNRuA6YBNJSz32nIMeuY+YiM6eUHiQQ/QXVsQviwvqWudDODmD8KhHcBZgAe
Htb5hJPUfOKj2zlvitSyfT6GhsiTyjpTTmZB2uRcviANp0jkSaZI2EmKxOYgVFPx
cCpGQPQ0139LYkHev0dixDwMqGzxVaZ3S/RTj8pMbQKj5VnwgpgmHWwGN2YebanQ
LMzUL2MuxV9AxRvcCqc+We8otPQuLqSU+gk9Rc8aFa9ZMm1JdfH8z5FXi4z6AMbA
N83aQk/TocQnckg2sVuPlzY3ME04bU78YBIWc6R6UOPZLP14UYmFDbHJFapZbnG4
yCxu89ILZsZSNNbTUFlP4ZDkLRZq8MQ+puz+Pbal8SvziC6C0fzyWXnjp4gRqdaY
Xnu7CXS+t1fsdXHDgdO8l4YghfGNiC/kgt4r1PnkRY1A2mGHHKMS228ZsQsNhXgL
Wuvjs2vnTrjVhVJWKa1rFkspl3Dd6j5N7a3I1hncKD5fnXOD81BIXWJDdAaTJ+lS
jxIhWgJSiJjpkqzsc2AiO/Y+J0sqb79Go46VuhRT9YRNIJA/QJMMr89n0v6F/bh8
YgASX4m7zD8H6eR08wo2K+HTifllnywGxMV+EBrwVOAXLh5NcqoHPIclv5TmdvYE
5XCiuv5Th1ZeP4JbtXEd09ZNVvfHqI5DZmHx69YtGhgY21KYKiLJnddj1lfSZCRO
B2/No8KVpEI25hU65rWhWquxynzVkvm99dqMJqfVRDXTmruV+rwYmUHw+S7jAChD
wuoQgfiXqYBs0juovXTUZ0Hhq83TBCRh3ra9nZWt1oxjGl/ubmaXkyUpuMJzm+o5
/KFQsvquqzS54JcqqKjsYPHplwnjEm5PBayZWtJvah5iUZ9wd4GOrhUp7u25jjwe
bFgaOBrQKn231iGMCfTAOiGt5Vy4W4H5v7ndHe2lgGYSkQ+8/cKZBAiNyBxCOQh4
wwdvHBmhX4ru/Sd7FyQNU4Z42m0SofFbJq7UPLz5H9xr7GEjRW5yxkWFbbWqGi5d
7sd8zXJndH/7xf0YJ4eJopdlZGo933QPltdiZm/3hIWSvGWfFJrJNBcwoRZ1MS8K
5mEA3OacamhJSgQw+PSKHF+LlOD3Rn0oacgxYWLRyCKoP5Ehapk7spDw2KZN8Dwk
QvpGeBb+ehr30laAHdGpv/05KepENK94GBXW2HmWGzOd7Xw1Lmvb4ooVTkpatZaU
sESjBxp/XU4AYqfKBXASRxfvoRu9kQHW/n1uuBL8WFzLvoQ4s9IMczDzBhd3/A+c
ayfHfHqvhHfZtSCBAlxsCZ/0zeF5SmeavxSTEP800ahRZqHEUbDL/Gb6eDq7stOA
M1RAnhPJoez3G/wynSwT2Ft3Fr2gDGLegx/D5oCt9wXphpMTuqvFwRNWKbZ327Y6
3ivQ4q3bjZu67Uku4EK/iuICFBps03cIbnMemtGtZITRrnEtExfh+MRo10+1uCVv
+Q01QvYUlxg+x2TW8xw/435ds6NcaWxP7oYucFdGUUfk0nhPT6N9Hq6VPdzwQO0z
D8wNQI7HhvkQViN83q+nPB3JGcDiytTg583q5ioyXurP8OxHlIuNuB2+P7Q9YJQZ
sPuSNVAxWpEYLZwyrUHwDxk4xCyNuljBMXeDBG32arWpGbzYcuOY9idF97vdWNGh
6YZ8hLAppmWCiTiwaB4Y+JUxHxpqKhiEUGIHOZ50uyA3EpmktedG2vAMCn5dWJY9
bhRu8TocTolrroIOx09abzbBO+qxLaoFboX/DDKcmWofMbW249XCMvIuyBtaBMf8
KphE0EVA5GICzt2a/DtC2loncjuR1dDFV3M03omr2VV6yHKgJvEC0LcYrFls3n7K
PiR8LV1tsJ+FiWYU8J4PYb62u9FYG/etmaf6dXdSeXIvPUaf7E2Nw7R/bFF6p8/c
+DAvJrNv9dOx/2Ncy1ZvLk+xJH6awhOsv1qWwgfdhzLXF/QWshuSkqTyt7lIMVYN
EmOOv1bfB9ex2JUiXK6aPvzTaDqrXZ1L7p0Gj+RhgvIdtTU8gVBEkTGet7jAWWqj
W6zk8tlmf9FGxZgwhwLeEyEdf8kWWZ/JdZvM/kBmbkHwaUy0CovEAHPbNSLC21zC
BuKLLfwQ2VThrRL9kSLQZHDzNZjU/n7+1is7xrGCLtK34cLZME+x1SLeRvZ+TtbW
eh7hKHP1XADINbCfz09vaOvIuivn9jmYxeBC/morvJyMQtOhH+RsU6tAc8t6jy2P
UGvn3kt+eAsG7rJs9K1Z5963OMEEnTF+Yk8292JMrISE7sF00J94rXaZyM3EsSeX
/Jcv+JPlOCu7T9tTe7JbLC/sqksq6xrKojZxdcRY6UdheAY/ZKJtStSbOx2YTwku
NMmaf03tJSX/vIymyidQPZgKI+1CRZO2mx/GY77S/n476/GZkUxbN74m7BTQcUM8
TQdQbMjZGOxwDrGW3cGBm9EBVBWeaSa9vjG12bPXPAEpVWcxjc6ALt3b1BsPS2t/
uX7CiWWvcKaMRZchqrjRBdWXSAwqf87Y7EgVhS581QuJdEPmPMZvBCyEfdTFw50W
DVCnandEoUf3uwEZXvcH+DeOW54+k0OsztMy7EBBKAnogPLoGbnf2+Gc3F+rlBw8
+SuDroGW7R27puEu2kWiz+uUIB15P/q40tXkq/jNbPwtinpkvWv2BSnrMPqL0/4I
1LEr5sVwJBIJ+COsKimZfMFxMuA54rnHLaiCC757L0WbrUNodO3lBDaVbsZyncoX
5FVKSpWv9caNGuRD3UGi9W+1XYgX+h14a8Y6V6GH83NCdL7nKWpw/n73oM/Lrjf1
VjOnKLwVKeRcZ5yyM1XKnxj+kxmCklwJlQJFjyELpeWi/KHA1p6Wp0kxfnq/un/T
f/r5sw/96YW4yvV4rhBcK3MU8NhHebIQkv2Di2v3OR8tDSBXQdgzJTecYyM5vtZQ
soKWOuXf4XW+Rapn4qAyzxMR5EclBrqxeqoFWmoIJ+8BAuEJSSrs2DvkWPJMRRx5
Fzlt9b/graSUXYoGjqvlNS4Srw1EYMZRgmLo5Ue9DdLZ8dgR6aHpob/flI08EM78
C+09zFGsYtmmmJyemrPtKY6ZCjwrMDF2bZOuTCynyk/XdOhXDUgZujOezGYFfV5S
vZNb3/haefWNfaXCTRjDjq2P7ko8dhd+owzRZ7k2jtJRbZpNN0JczIgMTBvAOnjw
7PcMQWWNCsJV3WSihFFMvI9Bna1UZ740U7H0Y6aD0lvi9KlY7Bd2AelVSJGMxqyE
uO7iIojEA9c9dlDZ2WFTgG4/0jY3uOY9UXrJncBI9QFrKRMeKU6nRPttyGboXxi5
xBX+hFMtrl3rjcoKvCy+SKGFTxL+tUAUCPQ7QCxuo8h2vo/tGWhfmhXrckOqrC2h
0LTITf7IS0yqymVSTcv1wj4fkWl+Jle4WJGYJ7vKIDiJdvCYLDOkao9b6KaI5xJn
yDaorxH1mPY23gQxoduQv0iodhuGnVFve4qDTMQ5vgUBjY6yfzk5e8a2p1ShRJbs
FnWth0pzbFCv2vaMKjA+9Tqcs0yCNVCTznBc/KKWrL3HZwCwjZnV02JkrPCoRns6
WpL3aqHR7BPPLLaKfyBsTiAadE6DoU1GlcOWm+2Q71dPFCUABaFaSJvK6sGidscY
25C/sFXD7maqZCPh8Hx77pytIwoPff/veHsI2XbYYzSEl7Wb7CA7Bd/N4uEpYulj
xES3gVVabfEqoLnI0pL93pdGmdxjVZ4fkpe+q5akP4Qz5vBaSpo6n0koYky4l/mN
HsOpg0oG9xTb3pUQuY42jpqPtb6NaUNIb7qf4vc3H8f7sYZudF6wg3EWdn76xnYK
bT8IJw5Mm/DU1y16H7O49XMYNDyzRLTrCirSMzoxBtfxYPIbaSgPptGeGa2BwCRI
as0yY7xsDKlBhzDQlZOIAz17J9ioqCQr2zFWTTIY4SJmNPD/ivke9usvy17iTvmH

--pragma protect end_data_block
--pragma protect digest_block
rZTgeO2P2uUzETqoQmtZ5+Xuynk=
--pragma protect end_digest_block
--pragma protect end_protected
