-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mIF35AkV0MhMa2ibTmfBqKL+S/bf9Zpeh/dxOiUpFvwhpl43HfCEMFnrwADPnXz5yfkbHyp2gG4G
anmyxPQ+KOPiU5dE1vLDZOLSNWz4IhHIS3EPanL1yKAg2uxbBWuieg2MpUYA10/J8ehZAWJmcw0s
UC96W1MOkWJk2HeGzAp+sgQjO6/gTGNxYvIZNVDkGov9rONR2MFI0CxxZBJbfZwsPnGfS/QfGXip
yfU+DwzZHdz4ykVWH/D/3Ffef+ns7LhRCuFErBN8lCwbpqJDDE/0M7y32InbI3agN6C7nhRJRSa1
qxbUlaNWi8wgKvSaxofH0JHx6s2N4IloOXI8RQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8160)
`protect data_block
bNkkSPDg8X2yWXPZ0xsUqf+MCTtjm8QEd97YDJWNVoLSkYff0Q7tVv30U0/Wr4dOWHMih3dkPFYF
GlP4GfCYDm/ike0zaAffxKiEBcj6Y3NhftLyHdpxINys1TpCeXxLCjtphy2vi6U3wMf6PyFhE3wK
BgcPYEXfwcBGOBFxzHU7JYEaNuq+QVmLtmQPRacBJ4HMpX8GfV78uXNGBuN33TNTmRJEARLtP65X
ia5mfzOD++KmlsHYH30JCTEbZ0d+HyRmwux2W4hBkM4JJ+hClLm7ghQvyIOJsFHQRiH6Es992ULq
6LGKMZtlOArC1x64cXE1WN0/TM0R12P5LUShToe/SE3M7Olj9PU/Ivq2P2b+7qmPAes/qHS5ZJK8
mXhRyst6fd4T20JWxoWBuiphLmMXUMoej7RBfviZWdYnP4ZNyqFcbJQzgR6kVjI4xwCQdJyxcCHp
/0XKuIT7N8dtNxWpOKsRi3WVf+9voPCQFL9kqBFxIkZs67/s4uxqSwFDVYAPfP16oJe78ASYfJ9U
i3hKccumzKiikybWRf4qS4UyxxWPBkQ9tzt69RPNOpoqbjacOczg4r5EQcDPvOUfFr5DPRD3iHA/
ZNA600AFrsuMYnFbF+Emuy1wn/RMcinDqzXae7QQzWpif5Rg/HL25gwC4rDMgFIBbA2BQ3Vraz8S
p4JEnbjOUi+xwk5ZxM5GoB5g1V19dVo5BUy71g3wlnNDvyioJaIOlqQPXxUnvFrKSAZyoavW2LJf
YiK4fz0DNF5LUY8PLJlUas2IKFp/qieraW/gTe30vYJTQ2gTr7ZcuiH6FrFuXi0xiWtU6DRTDH1Z
inRF/B5wN7gtQI8c/VqjqkvnpCPolVSUf/bDtnOqRD0nvWK8sn2ODzNRoEoVOKJzrXFeFo/BzxIC
nHadrWpokAuR0FNiGsYqvR+JoRZRE3beCgJ4iBCCVPaCj1CIyJK11HN/Dw78V0SvorTJFo+/l/wH
xHGPrX+4vZelu9V0AMmhvrsCd9+3BkAoHc+YycQwIOcDs0DqT8tZqs0gDRe9ZGPHCcug90CN+N4P
PHqndkGJqkHkZNi0irZVMQUQURhchqfQ3nanlx1qA5ifpqCGRWoHAPCBB/3071RiZHsa271w8mY5
MfL5FnpcJBUVcoD5g9dC3vNbzcxnd7R2pDomoZ4I1O2Iavvh2pgUN0PJ5UITMP+mVH2DAhe75hEP
NsG7YvqMmj6ooQoOIehcBInrtQIS+2ga24sq2a34KitkB/hrWjsIYcnjeX0I+8HbvkyxZdpmV27d
wVUWCEDIpX/G8WvciLH6dOA3SHhSIoXb2jIZpfwDcgH4sOXxRnQu7t5g+TnxpOthK7kJxs1Pl0G7
BIMRV01n3lX+eidbucXTBOnDAIy7550uSVsHq6+7u2tKwxLwSe52CItJrrXEezB8rYNuBu/ulUQ0
HMnNndsIuOfe0/xGH5arziRwIMBafaWOT4922fUI49NdJ1LYY74Fz4aKCxIybywGYZhZk4WRj2Qc
LmNYlgH1gsB8QTNYZtR6jqXVXQrrlb/96nCmvAEIXPMK+zwU+vMRiLyDC5eWui9KiS0YYbmP/8F6
gUefVZiGmOgr8Yv++hBDgq+u8DE0sncFiEO9BtRdsnp+nDU+LidY/CItJZ3SHwD0dcmIsx9KBYLG
dXXOXxIxOHk70QNpwBho24zNoXio0V0yTTEmGB0mzHNGjRUesz1RZs39B5SwhN1Fmv1glwPQNIwl
J7HciKXFKZoQosOUHXr/lxss0VIVRDPFZJsYQemHzHeSWhXteIpmBJH669bsPdD+pAdnsjxi004O
zImpDd2fntWpFbJOtbWVon9y8IhiMikB7UI2P2y0GskoigrZX+G+tQyhy2bY2bKN30S0MqCF5e9i
6Ndiju/vejawv2zqVEhyrfnCqr0fIcgSzKvBmC3UAPAY9qkrfqJM9jXmVoPJVJ+zy+jjqDsKw5re
eNX0H32IQmGyfSDJXr3xEJvpG0WegNCSsCf7rusyFsLdgqp/hJC8A0rJfaCyzkU4Ovp6TDO1I3DU
XeBQIh+aBFB0TbLw9D1APInA9O/mUC3jkq5d60gs9zXnPTm0U3lSDLt8bJuyjF9vvhLsGkh66v9k
BgnpEjphoQQUs43JXsbOGfTbpIPMqfVJCEiobuWRJYcxhryfEa/0sTrpk2DG1eYnN8HWJQajtwBY
/PCfwDz82FDumwgJ1iQCqp1KWiFREdF1gJtxDahF6ZxOgrwsfltL2GB+1ItTvNH1bDh2HxsYgJ7y
lyVNp8QbKza6AwhoqjmxQZio6qDixKxBgcKn9aDeKxf7sRIhoAqJmwZAMT4M8NbnC+17AcG5b/jg
XCEhDKJ9yCzIsICvFmvvQkBKCzTww/ivIjLXRYIONu/Xbtjim2g6E8VNgG2bmJwy8ldqEi+BBe1m
wFfdldLfiIvLIG0MBYa9XMQaJcp87a3fRVvof1hfffiMZeh6LWNIPbfSgMKWW8HkdqiZFsu4vqmW
mf1/IGKM8/QSMDILfPA1nNF+KmKnmuQi/TukhdJQWAOILx6PqWW/mYpHcbjl7cnUvcT/l7Xck9pi
QVmIjh7VMIWx73zKrWT19ZkFPwB5ZOrwGFoU/cUyw987SNGF5sb0WOtIshPjzsZl4OwSwMJVy0XE
OwxKX0mkCZxv1GrMleBHNqdAwnLv0TpzlJyadDdvgxd90yCgQnc02WaXrF3vk9sEML+c0lj5RkrL
zYqzIXfi/qijfkj+WAmEQw7WPq0fcfum13T215RyJPrP0A3xdErsZur0bAiacFr7VwyGyQgKKZ9f
eN0Dzy0FyM1clbsV6y+skjZCnERABFldDnH8BrUwXQTi45DK5oOcUToJ6O+p3MPvxjS7gLp0JMgw
eMtiSkpcxM3jvQ6bOmmKKGEop85w7nxfzVlHNmt6R38jyvdb35p7oXzco0Vf/o2e9zpF2LZ+7OYd
ySGbEyLu+DQIay0h60HKS1ElrxDB4ukaTsclh3w7LLo/7IWnMdvMROCTtmSyzy9A4ECa0nC1hXK1
etyZD1NYdUegsMdS1qskwvJCDPUsnOok48X5FeeCF2Voxy7hKYOfxvYvk0acu9vRm5BiqWVimZie
uB/SfrGSdnR5lR4r3jw2QHmorvf3xamV6As6ESnGlHICrTA2OVQgtdniUR7BozCADlQ3aMCLQ6bV
JuTSobt5cQEjXckZtbSOhOA1u5aO7ZUTLoP58xW/2WbZKYjo5qB1KrzPATeRIjqs6GHyqptb7MnE
Cc+GX+cXoAGOqNGpRzFYQrEsCH117ZpcBnmq7SDoNSX3T4DonSFVjcDWHGX5re8umHP+MA6UBXS4
Nd4HHruE95KJDCNn5+yLdyHZB2cAANntz7YJqijC4lylxlsIZp6Caox+Sm9OnogEfOnps8cCfdec
YM6ybeE9PlETFlYbtu5hrw21VA/M3Ll75GyjTeW1HQq/pahWB/9MlXBb+GPLieYxO3Ia4ClSeF/P
UDgpQc9XM4FLfx4U2OPNQ9zUb+tovXpW/VD9AeTNxHQZzRZyVVo1UMGNCy7mgc3V8XrsIUusXPK4
4seS/JT9ydvcNmFaQVpSlzNG1nJCxRr1pfxvbsUgzXNhd4O1/RWr+gxGwFB28YQQoJp9HHuYFIT8
Q6NW16gTtLeB5SRlSuxGQxeqM4ONo74/Fih4rloYE1/0OTMFP8FnYshExwWHo0AaxNqAVqtNG0lw
xHeZUtQHj8ugndm4y5kaGU1/RbsWkecF+UFNWEihzDJjXMiYS1/Z9HECixqT201SI8RmE1TeHEp0
VN8KM9kVyIGCQGtuotuLtnNgGR89GMjaXx/W+gvaL4/M11Q+U/iGhBNyH8bDZfh7vSkIbnw8FbWN
xCK0Jqoa6vXQ6dgYFMj3//sS4AQ/zRWVzul43ZxGSOWFAuY103gbsfS9WazI8rKM4hHRW++AyYl2
MZessCcGqjk+PW6u0vyCC9pKJOkD/qnkETz6/6gzC5viG1pacUecW4pZrc8CS0UwDyJTEpm3nZg4
CzdB7T2nK1AugW2qVwIdqxe6B6vrN7SEV6vqfEJTktA9c1Ak/2H1qflWpnBH+T24EpEWZf1s5yG7
SaXM89QjEA3ek1J7NwKX3DQWTJnwhJzbbPZLYIhOXIereV90cIdWXGgjUJxS0VIoAYFTOOB3WbFB
vzSss9Dufi4wOPmqzhlhj2vq0TrHjhnEOllCvRWPYjNfXaTlm1V97Yug45AbOyR6lqpOxcupM2js
9Wmqi/xSx5XJedIp+u/v6z0HurfG/2WRvGbQhQwHoA0NY9djTDstfGtWin1fMWOz4MsMKvsER9gg
5mzF49rMP3n7q0NKBgxD4gTPIO7TE7qQJLP874GAsJuOUG5sAm8a2D5W1MK19J6dY8QK/iGOjG09
P+OkytWHEyhF8BqJdxx67lSnAR3ZkitXpXfHizKNNpIX91eyY0Aggt0JjLZpRCANp86VMW6s6f+B
lUUnvZouj6ygXXaKIj0KTJAADENXgpQXrBeVYQz68BcH8v/TQnxfMuAtPlrFXqo8gJyNkS+9DP/A
aVa0K8PI0FY0bc23i2tmFP5SKUpiYN9xcqTm0gXMdaTzwqa0DH24onEy4/Q8MqvpuWG0aRNakE1R
DosWY/TMBdhZJw2F1Lh1O185vHwWL9EpsxaIDUYEbOQAEoJpTYWKBUH96Iv6gzqMuSrQIEb0Ajkf
8eolra9fZl2opnn4N/8k8be6rJ83ecIWEGXs1tH5dm0arKwEkjDjaHxi7p3MPYN0TNitk/aWTgHd
LrZiLN6/UmHlAk6L74IgJ7ZxH4hiqHjtAL6qO21GX8zkuTPDp7LFNiqDKDPbELN0Up7+JIKBlYYD
Pwgr+BuKZIF80pdoUKvymzN9lpPpB262jt1TqOZ5F0g6wBHopbUJHKtl18FWCL3oeP+p0kiZqb3B
Vg9p8B2wbS1/DP8HHY6HspKq1TYESE2oZZ9zB5o/f2cQRl90aUiuNGg2nKUAuRTH+s77dTbaHJ7y
6JVoUwW59jeZqFwNl+axxGcX0gyL7BxYzkKJLXgN6fdOnFt4hjYWM3tKuhRGBxwGwSBFGsFSfFfE
LTqMniiQskiXkCmKo6I/BxVT3lFtR0R+r5I0Zwdb/HmB6NCAqvfOCs2vw03BDORwdxc/2gqWb80P
FDeJBBIlNWElOcWPhS8YVYpc9DdRD0mxDcN1YhTmrIEd4eVE4MmDDTC5O5o9VcGmBG+oPFlJp7mI
3roU2StAohN75B6mpGKNc2+vQRKhJPurr6hLOPcINzrKsM9/alKw6j43bN63EPZp0tBqPT8oFYQN
11e/d/77avqB7DQoGNG1Yt5pRu2eEzYLMMhMYQsfDKuCE5AMJYguw2NeLODz7J5lRlAZweJpuh0U
yEHa4smla28ZE+/C7/nBcRd2hbGrjWeBhXiqf1l9OYcNrN0hKNRGlLH4BsqCpFbKPugS2JdFE+zO
RmKH9KrGYv5CvlsZnh8afqWHoRTyyNHhsQQ/m2dCumbX1rksi/pMppwxpFkKi3GiA/NVvu1iI3bu
gwGCc/5IUM0XOQV50wcWk8ZRSROb+CUNlAxutXVZHPaNvFaORHRjUgj9I2f/rQuFxs6crrCGzfU2
w/X55Huv2ulk3/BFQ1+6aMAPEFG0NNZXBa2YdMVJMCkQv0f57aslENmxiRJ6YYRqg1wUpCfEbV/H
AlwD2+eoCJXmzSQj53onTFyY2/1LHo/r88cNHLeM/VmfNKNJn6EKLEEvLjV9lv13eWp/gudZ0VH0
04amCrHzNP3xJof/OTgf/YheAFGx0d67lR5tr7A1LETfGU3Kut0Jsexlcp/ouRl7GKiFxLcAYf8i
UDG5PECehcduXuUDC9gOSjbVPq70/C63tDeBIZ1wlyzqixwfxSAWJIJoYi5LpMVyBM9nLIQiTDVc
zvpNZ2vf7wcLclWqxR4dkMI7IvHaJYwA9U2CFrLEtCXP47imw0bhPx0rqZO7TYm9RxduP1e6Sl+/
T+lcahItBG0mIovMYhzZVxIkLMnD/mzSkBJtcJ5hhj7gIM909PPJjcn/sZyHYO0eEUc0sziz46TL
nIgX+8E+1gjf2uVm1iCy580z5cq+P8KQTIeMLlhAPF26C5bi4MPe2AKgLwb3xkSkPhVdq4ad9enq
I4pDtBZdwboAF9/6SM/uRRjFgb8Lw9gvB9dYGF28m1AhmDya8S3jLploygoW9l25Jswa8Kp3knrC
ZfnfSCRmlMrDsMJZagAv4P5vH6Ecqckbtq1AxjBE2Kckb0CC3ueU7PEonfz2PlSatQcccY4dos0t
mokDa4Yn3jRRw2s/1nk6B84BpReEwwDNTydqyY80KhIXmMH/+irw/tFAAhVYKq1XCOXNTswgQgqf
HwFQtowKwnwrpI30kARcEE2AdF+RkvYzB8wX5M8D62fqNU3YJwRRj6usY3D0Nd+uFRhYYLpEpuaB
/2RL7Caz6qvSzOuyfax1Q/snICYikywamXRVH0COKEuJCLafd3vFOs765d+T6NQxTLk6+YeqtNpW
yaV2PkUKRKnSfrOKGsNYQ/IhxTrL0v0tziTujZOuyhf/r4Isk6t3FF23j93z1xVpVxZk9l8ozwcb
lm62x0O/6jbqrzv/+UhHrEdIbpwCIaNbw3L2PEJpmhuTswz5GfhJy3TU1JqowOjFBQUpWcUk99iB
4Z+6DYImAYYl6glgERlYAybAWUNYEvlzDKFgAlrVCgCkEtgCkRGYO/1R0xC47zX7+HBiGHumP/7c
Of7aU1GIcj/rQwckHCczh68lQFaR3SH8rwSdAgXA8nSkVFH+3PNPg4ERqvyzbXX0pxX69j/Zj+S2
lFPgRYFPftIP4uoTWJCGBTa1SQAGj0IxoorHYW4R+d5c7II4z/9c1vWb055hlzcsISEKnla5pm9n
MMhGtHt0g4gztzLNJK4LhyOmj1Pig/tsYYgwM6BdSQ1U/V84DNV+HZIMLCO3TCUKsaih/eUjI1OO
s39wxnF95BvRiAE5n/cOIXAEl0N5TMjm48EDMpYHQyYZPuPPrYmGGziQ5zCrdvKCaADO+r+70qYK
lhOTZIFhn4rcT9pT3NQCJ1v/sB5svqngoV576000ZE7TrcGT6slYpICllgdOhIA2vtTOiv/Qf6po
JpJiAY6+rQL7SWmnJ01SsgvO/KIPR7uMT7HCy67jGNAE4M3Af5SaagYZguY0t4KFlOtlV3hiRJMI
xxSLzAxyQFPw33lWWHPmXZW3nsktHsP0BIeG2tZCo3KZLGk8yy6K8JsIRp+asUhs4nf5kb+Y6p/d
7xkgbLLT/fw2J/CAyJC5ISRaU4mXMDxuBAiT0UvDvVvMWXDoyQRtXdiSF2rYwxDo+6V/tyd/UBmi
FEzQywVJHsEjOrkZp7TFLY+FOS1IrwTdQqal1VYpIP80YaBI8ZOtrVdPC6SfWxYErr8z0A5Mk6tc
TuxxRXXqKN1UDQYyKMdRQzGoV+UJCqMrJyan2WDJ7lABF7llfSWfL8+mrUkHs3DtcgcqdwQoSkjC
wL4umskaXd8smR9uFgYao97D5uY1HbqEbMLU0Pf8yrDktAz1vOARgnR7QfKGkzVY2f6/E/FwHF49
5n6fXoLdpAM/2uk7to4kdLS/mT9qRgEx3l0afhQTlLjYA6/Jq6FzffgFUaTfcVaPagguEXXiG1bv
TgxU5n7wGB+b3JxK/nQejInXbQJgIRVLwZ6bbI+YlRJOOngta8MxPv/8p6CeinvD1j2GZFy6Rx4+
1cRT2WvpeOLRnw3dccTtwmBlFVqw+hgpN8J+7h+LoE7C3RjJep59ACUQRSw7jN2SbWy2bRXaLt/X
wYwFXcy9kVqbzjjKoe8IU3z2slX2kfG7eo79ljDnmi+IlIuSV7XXAKyfydsatYXgQAMw6Cfk9l1f
SKHmVutLhqrZEpxblR4tR/4oK8/lHnG09aGaJhsWXh+4pcRK8iapqB41hEfd6FL5Fuk0Vs2hYg0g
tlJjEVl+PBu3zRHlL+RUl0F/jeNpHR9HiXdgsKEdAnMt9sXimRDP7oZlWNQ7UWRLs58sZUklfyAN
xFsKLe4qUVvlO7sqSIsgnBMrOW8AGe9YHSxkgi8soBv9V1Yw1TOL8kXkWr/C9C3r9Q1bazxsCFDb
r1l6EAk2tX/M2Z3+yStvv8CfNxYsTsOYzfRqxp8beEj5fYf8psvTUTBITzBjy0VhIH3TpP0wI3JR
4flQr/Qcba9UiNl3wrFryVvP55iZt/cZIhN7j6DMpZ26YWD7qNv7AzK9LkaNbdj8Ewd7zwYVdFzy
I8i56dq0+SPfbZzkR/03R7b/gHYcPuGe1+NGQ8QmtZZZrZyUblaVkzMj+iQ1NyyMCOZQqSMiXutR
JCwF88BNaFUMLpglxsRm49Rs3WuQ9sz6m/V51c9159v2Du+t0YYH4Sfbh653okHoiJ3Rg4MbunVi
bbM12kKn8csE/Z8nEW8jnchvHxfXnnsC9sVtRWe7IGEP3Bi7VBd0y8xXy0pHpVFJLuwo+4p40ZF+
41UV4jDVKPkoy6MpaPZZSpEX/b1vrKQJG2ef72YLAtdFvopSKFyAy0MosHFswto8plJIryQfph9e
2m22lt1zuX1NotPUebZgPcmYn7bSRSlolnrL/UQ09L6ZKYTv89Kbw5bkG3mdBB8sZAMSebWAxtxg
BA0wMLt29knWJ/J9mSRffBl6oMFzT5Qt0krgOxNyGLMzaGts1KeVltPK4cdpNyiq7jyYduzP1jGP
V/qG0X5S7bRKhVetdd0RV2rjUsMmbXYVXxF1W+dqnKqPxferjusgSVgSUE//yhILr+MA1BM4xxVK
jZlo8Dh7/mqfIdpaQjIwdpKANsFrzM/fmPhBWnsaHHAjVASocOqxKynGJSduNUb6ySfrVkoXuEv2
zg93cRsDciJKkI6ZZ8RiSI9hzhaBM65zc4HqV9UMMm9NPbglR7kkZtvVI/oFgzL2m6uPEV3UBD+/
C85PrbnkgN6ArTIM5TY9bv4uZzwx8H30Ni7dlXikIu3c7W9bcNVAw0LlFFaEi8qqY/vsAAtogGQK
KEujG4pWdPK5LU6sJj3Lp4tGqSXnksi1HD79PPbrVoKHtZMD5RUAfxEU4X8RbdXNQ7LlZl0hBBQx
nbR4b0D6DYrOobgN0m2l32vvys9ATXMYOJX2FYHcy/PpIzj1TU0JpVjb380yPIYPQuvEkt6268I8
S1bh1yxUSBP9Z/dyZlx0orVmjbyn+7w+WYNK2KIi9G7zvdsc1kuEq57lVy5eQtjJs9/B5zqNC9/p
MX9X8X4Zt7xKyfv28gCUO3+hXaV9EcUQsMSc+PeHAIXAhdhhITXk07tEts4C+2UJO5MGVlZIQzAW
52pjWxGGt1aVJ3KuyF94aeN2tUFqFMXaWO5TZwwMHkBx5x6ZP5hyAUAmEiAoyJOdOQSygFriN/RE
T/xgZatbO6KBcwFWeTF87CtRxPYynIIEKKCGmDkT0JNuJhjvVIMJq7MzvCLezCk6cTN7GIqOSJDd
XFRyB+Pzzb8qCL9LRJCf0VtqeegC2rVs2HghnwsUiDFy78H+4LWUO4GLVwReQCh2aBC1PxM/KF1k
uWvLVfz1gmhXikli8kt2mJwnMr4+VsjnSi2UQIEtqxDa7D7MOnkgCL/Km376yj4PD08TqZJqBcOc
rZc8V7yTHvIBNzI9ffJcqG7sNvkMOcTg8h6uj8FT40V5Yh3f1KC0FkHVgkuga5p+hG0GcZ3B3iiT
SQEGwqy7rhETz0frGCIFfm0rsCuTx5xYlYT+BzOL4wfceA7sZyii6Sz3K5D+IlIZx4V3s4D+fieW
xLW3xZBup2C1O7dVdKuAzJ5T9jeY0IAGsVeeYKD9/aI4QUkD6cO55fG9lKx5c5fTfuJj+CFxBDeN
gTLSFxkg2CnjTnTd41Y6hpe4Q5zzBPbvcqDvy7p0QQpY1oQvMBQGrjg3n98YbvBUL9CXVO9+eSSW
nbLqHW3ZiXdg1d1/A2zbAIGnDPp0IEyx8fFsHEPeRvXjIKgu4d4xyCkv2soZkqHVVYTBp46pjEEW
YFrTOct03INDN22tYYUS85nl+zrbk8kDm9Z4u9nwV0JzH6Zb/xGXBn7Xv7dSGQqKcL+UpIPE6vVC
IQUg3XOtSVKP6N5PpoAu02SQvQLs9wGgz2e7ZeH6N2JOBhk8NIH6U6+Sv+CZPheYFT7aILQwBI4f
9BvVlaCnNNNj9bNddhToX16WRDTVGiRtcvyIis7FWvibkWHyqg463tEiLnPJQLB+xNqsyDXvQyLS
6IVtlm32dCoAPqYV8Cpp9KEFTz728SH1mFK+bvFfNvScvhoGut56cp1R8RVnNAag3HF497C8as3m
roNmKXRxVcz/NBOHqUMS4X2ObTeYTV3Gc8qCRey5LSPUAOfOefYbxKYS0DgwZ2qho70mSPK/qFwO
tWrjjRcODeuIKF/bWrXbEH6opxU2v2RBkzlTKjd7v1iYrlj4eGySWvgLb+lGP4kh/1cLSClZn8jS
E/c6QCMmlq5d6V4U94jjykGxAH0ts2H+BK6TL7JVsZ1Kz+zXNO7w+YHiFzrPNmfjFYUQXsValdR+
8oqCWrOTF2toOndBSrp7V/ttQc54u+0K155KLcmwdurb7gwSSEVCA/bn25jZ75hhg9eojJcs4BKk
AJ+Em/Jsbgupfz6Wtd/2soiJQEbEmbYUErM9IYtnGQTcsChQrW20CXJr+JD3jgolKE10woK7i09C
LMQxnVKRwTPlcCHZCqGZ9xR2A2VXoftTJEPWr6Ib+HLm3TrgN720jFksWxkcloKA2pEtC+nC9zYV
7tZ7vlLrFT1fbrYctjcHkO37U4yD6NP35RlYdWEqxyN59eKqxFbSUrUlpb2g8KTRuKBZVg9RjTQ3
AMn3AvwxyhDu
`protect end_protected
