-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
jJOg2Z0+TAJtGc7Hjl6JTctRUEWQwzLZ6ob0aGfdCgdm/ZgLUvICpcVrwHY66OiN
goyh/ktBqpKBcutiaQrCSohAQUOTZ5AFExLqCvOaOFumWbi+geXIIYkfqPQEMo14
vgHfb8mrcRoDZ16MFewWnXzQwAFyMa6+PLRlnBx9taY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 70960)
`protect data_block
aaNF8Pm1JCrsWn/PeuoPggp2RKm/3gPZxxsosLzkAC/RSrLRvt5sS/1CG51tULw9
OHcIRx5J2+yGMPyz2MeynI+L6grtgaEQODSOBGzwNbQxQ2hF5YyW4BV7t2ovoJq9
HxFBL/zUlDvxinBEbGq7laa6fFk770UC5PodpPsvpsaRmONF7NpYoqJwd3w8op2p
toBBVRh8weJeK3YFPvJUJG1SDJOz4e64cwObhytxihsHLAgPlZ8zmWrAhCpRpCbs
a2XzbPm7vdLG7wXq8AEtAh/B5WGQ7uYfpXo5zNHvyVe6OzQxju1mmT2+EInlKmZx
Xe+tFlVHQp5TduXsJ+/2HQo3gd8fCoIsSNs4w07F46O6z0HgC81ZBqv8a/C7EgnI
MNMHWFVYtWj2MEMhRqKQ8fEtJGvvAbOUec7jO0Jax3vdIAbMii35wYViXa1gnyLJ
JYaFRbTjNhmnaKB4Uzh+qF6lZzWCOVZkwfvZVIzv1F0yrSd6hH8CN9Xrr1OB9Zsq
TknwSuQXwE/0Kc4acTE+P9ZUHtBuE/abNI16FsDE4H7QkIYhGJq8MpPdVPcJ0Xu0
Fdo9vXEYxL8lXSVBNOdKFzBwhsW6q8T2qhgl/JS/0VJZhi44zQRQ9GpqI1O+cXvB
JcN+1N/cHUDfnW3wzPRsC+w70ztI7bg73blSBPruG2tYXIDcp9yKgHeXjTC4UQn/
wq9XDQIc/+flnJcVXhF2xeLWmFi0NpQY64PUE7yuE4LiFX4Kt9qYBA/BqqZB49c5
ilKQx8CDT1kN02i3k+k37KQN/wtQMtUSWuppwuXWhmFgE6tF7qvwQO4nY2ZRi3ry
EGiuF3mh5hzolL9XXg47C+bEwwOw/PT+J4vQSh6n8f6dmS3kNQb7BCluMtcpxpZj
B0LpFWD2ztvjg5R67dGp4IUPcMxaScw1bFOyycVaswwgVNdHROPRnZxjvdBhFhgA
sQi4kLdNN6b08P1Vrw7wjKrpJr/VGJwmh3biusNb5eG85UNNmJqVFuLjCAEw45zS
sGfyJ8O5Neud93LL8mEuuSa4pSX74jO+MLOD5Xx3GrTFRY9sKw7Ok3WYGcWlAEey
nt0KAH3Bd3zMB3lES1ckNJ7Mhi/l5o+GdPgK9YiKvNm34kvYpp8BFOvfP9zqmIa3
VqrcesiUHS2pdNMlhgumj8OFzfKFqMXGwmgWJK/zdhlxG/PxMuZJgusKx1cXxdwI
y+RQXluzAHEXPXH1Lxkpb7RVynJWY+DOCI1dkrx+xhbdYo5lJ4WMSJN/+7CNkHzO
1N/MpwNmVvlUhEf6humgkeZnRhaYv76r2BEmFClxznX9L8yimq7aatETkXZnK0KX
AkHi3dHn5CLjws3fFcrF5zlL+SCOZavafPHnxG+6nMnQ3ep4MjC56QUJloscgPiY
W+Kt/QczTMBmEHN3i+dq/8kjwIOEkwsrrDuq9LLs2rCFVJosVhiUHYRcC0W4oec+
ShGfNd1LDMTGfgqjqEbTTRaG3xwA7kYPrkM1w+XX9FddyPJw5/ELsSThxUIRYk7l
1a9Uh0j/hzryRMIKuJhwiv0Xkx29VDQYadskracGVQztkGwnbW05jFSWUXfq5JEP
oO3RdoG/e6W08FxR60vpRh/EWBFe8VdIcXRcfMGPdGQoAUTltavfoK+v+JwIS12p
GVKSK+3aJcRRDccafrhgI8FKAKFGuhkXVFQ3WHvRx2P1vXbW50nUW5uNlCU/JNcD
OfBHA3oeunzRWZYVUsf9mcqk6BddMTRXmeHNt3HBp3YAeU1E1qcfPXlRQjQh8RDr
IZonV8MzIz1aF9laJycydlgMiAfUiWzfFsyoiRaYX6XtvyY3EMHhoUS0gKlqgL8W
FmIGCmaiNEBt8ANNbm9qCTIQrVgDTCTF/EERHSnQ/s2OZVX4mI/LN6GJ6+q2l5IL
geJA3BUDz0bM1qMYo2C1U9KOby+HjyEDAMm8Ykr3U3g1dW1h/+l160d8pQ5V51/H
VTVOkalCPPL6v8hVBO+RGZ6KyS/dfz4X0P573znZjfMPd3KMdtme02YZGwcRzczl
WKYtSyKE3ZRu1I4Em3Bxi5AQZCied8B4IZfv/+kOCHg7+buVdPziveN5XCJ59ALn
IU2E1nROAVucvFxQMuOcjExzN1jD53o17ZAWWTrjXrmE1+H0M/hMp/B/nMF6+sGj
zNbDMot38F9wovO9nUOEjT+iZpfE7IDCfQyQF3EA5H3M0ANMocdKAMA3u7qltiOI
7aR29reTvEWOhFWmDPfFHqzgdt9ksajO7c7hYtaTCXUfNwNglxv+85DTEHQ5w7FQ
rfEVFsleHmB6LiFe2uIJgaDZHQkNppud9nGysM/c2NxAeDSIKFaq59mICrjiayuZ
gE0w9b4xKttP0UEcfY2Zs67X+xvsrCoKvrAGO6jEG6I47vIqtRiEiwGxJc0DA5kq
dxXhw0sX71OmP4gxDlZK0ULB2YZVlL5clFDzXlEeclxwY+bLLjCRU+xEPYmt8wnE
XS43BDlufhguL8Btp25/LzyZfrxS+iX2fvlh8ZxQIKDXIHuNdrQdEcxAKG1yZahd
9X3dQx0vnmNYbhsuOj7ZJ5tSaSgWAwMNW+jSEnqtzisWAchIv6drhSk2v8q00jAw
Pgzqn7s9IpN99ocnEn39mgn7GgVQg/Qr2IFbhhLYSqHc6iIHUKH6PwKqaxo1ehi3
w0A6BT5d/zGsGiaPTHVjHyNEEJBxSirs+DB9I9ot3uFF9Rv3QDTneDKKSTvxUYnm
tpzxUNIUaCk3hNIjhtzWPHsgodHRduQafGB+29cijlDhpZkN3Pdb9CpUbvbO6JH1
N7ah3dFAHBV/pySKVdgoelZOy1t4Xhr7YyZdOInD2AfzxSlOf4lIxTuu4tq0pzUJ
26vxzsLRs9v3WO61ACREe5eqWlbx25kncy9fImUwIncEl68JoMjjfEoY8P/lLFP6
sIatDnVxoxWP49TY8PtR4eIb9f+1xXzDfrGSkE487Qgka1ZZch4v/8ncbP2DMUSd
6JSHGrcf3ih769kEtfRzqgEvhZKaWBTkyUGlBCKACrZ1ZqO3gZC0ajySS6pvzSWM
+4mBXIraPH9nqOgJlJaDKgu/mW37Of8/QMARpnf6gAtrfzGzcG/jS9oxX6yxrNKM
bDiDMxYBMI33c6aCR2wI6XnOLDCrnvDfhHbPp0LjF02m2mzrjsg4pQ47WWCOQr37
L9w9uIk91HLcLU066weeDm/JdtKiJX7ZrS6Tw8CwlbFiA2PuDVCGI5XYT/rTm9Ay
U0skHegzzaOotQwWfoT5AlLfq6IjLnMM4GGpaZGNN1U/TMvaSpd2RxkrLuu5SIla
AgQXDguCpYuP0Ix5tIZK2rL4ijXmuqanMFyiWgYNjC6kQ9j6mO3fYT9GT8bdStlJ
7S3gOuheSz/GlA/lh/ip4wvUMZKpTw7qqiHlT8nlQJEFWWfGSb3BoPWUV09lAre9
gVWF9CpqRVn9/whog/N/CGjjWfdg/FQAY9bUBlY6JZzENuEIn5rnyA6zTHRIoHdW
R8+PSt2RgKomXPCfh9VVvi7fVsSmHsHGsaIW909DhgEGDlKtaJo/70uosSj7FaUv
df34GbjxEyVq6sUpjROvVyfdM1VtgbiYLMH/Kuu73/0ab5D4PzIf4hEFGTL5b9MA
q4E8rIIO2XtWFTf8ZRv5fwip2n2N/CExhXGgV7eLn3itVUOLOqQdFhaRDA+JDh0+
b56S0TfTrgRX5nhjJBqtIGgKdNP5BVB62AtS0iJ4L9BKiN0tyUmDlUeCftV/AVBO
AMzuua5iNY2YkHjHIG0msuAsOaPlxkzDeZUnDoLzLhLkNoK3VuOVvek3rhOhIu+y
ctV/qRxd4/o5UyzG3iB85A6zc5maIipueJHWzdQcOBXG4NroRHoHmyXjzK2TCYjV
cbqczsL6TBGc/FAzGNVKKz7dpGQIy0BrmbWQFf4yQutGTtmilzKM56pSgNBSItoc
7dfwIwADrd2hwVr4YjQcnKfQmfSgo4fbDJE9JtnTu03Q/CmroYLeqTV2mU4jGeeG
heJKkWGgm2fuO5QZK3GslNnThdcLH/3kFeYwuHXbFAMOkjw4A7ObpUkTF8yuo7XM
A8dOkrdIDTAwU4vEzjqK/Pr2hnQplxajZxaKcOFS2b6mI1/tUiYSFlaKscvVVcIZ
YcqPYsgtz6AZGadhIVst8e6AZPednn5EfwQ8PL0pEqrvFSndDhGZ0dknrGgnESCY
gIDqtV/q+w3scIE+B6dZhc8zrfZvytxV8zcneYDb+YaxToJY9J2zdmI5E4V6KY1p
7uWyHLsthNgUmGYiM6FNU/xd8ddNYuFY9eQ4AlKZwf7OnKoMxB3waZNeNxxaoGjJ
b8fzV6hIV+WK3VXafzTV8ckXGqBOH0Ke4vjnKg0RfVDvBd/V7NlQnScZ1Rreo8NB
C19aWUFVnDYu1Cv+HKVGGGje3WFzleoA324AH+eSA8/js7/jATkcqw93ZTBsknBh
NGEtIDcIHp8QZ0cwLt2IPklaUBmHN6cHrOITt8+lkP1QFvlRqO4DD6UUVZmoOOxc
e49KC/VoCoct7NN/1p42BDUTlljuQWjgM4xK0Mon+FgZ1xOqKNokvyHgdUBLbqBZ
6iKJ3T4/e7ksjCmlqGNX8gdA0184rah6qN6hAKdcQ0flDyqoeBpBkm/jrbvxzqp3
NdL1fc+4FsF2gopsu8degKBkVRsRh/8HmTWB/U1ggfPKb+TuuMyn5PqqHz4V3Ugv
xY8RPCSidfhccHsXRCwiE6JrrRmBlblKHV6dX+64Dz5fO2pJqoKY5n1YesgN7/m/
ahfAxTyrKy8aJJstjcy5QlP6uXJjejnMF139n2i+8inVuVdYuCWbEiVkotPwDmJj
XyP/CUwZdVwEVKwBdW2O4gVOJmqTSJupzpO39dKk+wmtE4VzaOQybjoGz6z1lXtJ
g2flKbqPh5rlodv9DmwRCWQKnAz9uO8JHYeLv3GuhRSWucx0DGMoS1zUosPtf5un
EamMca6OXGdFUGq0Uw++fPCNIUw4e4fy5Nxah9qyInvnb84Huh3yeHlL3nvPSH9e
swYeRtHFH6BhOirh5Axn+f7gWJotSschz8GpthUluWo25KV0MFTClM728X4lKWao
91CQiBj0Vz2LJhrHDUXCR0NoJDrMLyby2gMI1Nw0z8JS+6h/EPpG1uvRtwi6vyaD
5xdpqhiiXK+nK0HnbyIlPWRy0hf4pENh4xcXkoLcnei/7ah/+bIuUORBbuLPoIa6
7+PokGpkVir5ogrc6TNu3tUYH/vGzOHCKqUW7Sb3gMom0y2pJ4VYaQq+qrHTfHHi
d7dAGtbKW0oYIVLHT+FMgQeaBNnNU4VtGrZvjlWZBenffm90oY1lordFUkITs5Yx
egX+9Nq/xJVZWDvWHpplahX6kJAb7V/HQdJnA+5MXTZOlT+v0JXJntoaA5sHodDP
E/4DBmumNGym/5yZY5gOpTuF8gEE4WJu4FqXfb6m/o0h9RlUkUmGnLTvDtXQh7+W
oDI+IzsEL1Rk2i0yW+QCWE31R8kND3WC4bkBim3Aad5WCXHTs8SNgdeLi47jokCR
0pQqF3m6Xr3xVv9Dp/cnYMK3oybdOZBBEVBzgjwJDBeYEBbeu3tEeUOjAjb72NCv
WC0eFZ0DaHTdsDKCVJW1M6pP3Q+gCxberVbliIoyU4JpP6uxK05YGitAUQQ2rjOI
krfAN+so810CwMw0IzNnLpu9mOl455bm75yropPxAZw4Mc/EMh6pn8eqGI4HiPGi
mf3P6/EdH7FaR7x6gKyU75RloHjNmIFgYFytd3QPFTuk2qdqR1/WDKBtlDQ2dN1E
CrGz2+mnx2YIsOUrP/W0789JH5ZmL4GZ2f/hbAyEWY0G8foBrEmjdOQcIVsyr5WR
k5TLD8//qqIbgOWvrS/zv/uCcpo8fm2lPnDJcQqwF9aobceLPk9jk8OL3ueUZAdc
cfcBEio8xwijHaAKJ4KMUFAiLh+VHEqmbVEHsPMFjQaCRCg8wFSLrqqRwqyMPWBv
inYSwW5Nlq0u/0xVmOhKjCRjqo5jj+ktGsXMFKjaWw+CGD6bflY/m3Lx8XkLT4wp
42NQJOSc1cT4+bmNmsCevxcnaueVAeiLoqhC7/NXeXxE67oxpw46+Cn13MExtVCW
FXZoaDwo187UuU0rIyNHDNa1qIH/zPcOPEyP8j0UhQ9ZyHI6n/zvB3CORGKa4rtl
AZ8hjGk3UaW5QUkYMXY9j72CfSH+XnxOsI+OeCQs7moW8FYpQCVdrWRjRI4uqSKI
cD26W5pch6WYJbtSubI5AlkmMyGsRiN1WRuCcHzed/xk13SqF5P0SfUuSKHdpaRD
oIKvtDZqPp9FVh2v0NnAOjWhU7K1bNPZqUNMwl0laDK3D3PMkAVSxhAzYu1SV+Am
l2+uA5dbpz2pCKVsBG1lfFHG/pOMmEuxO7IjtchqS6tXjTUDQ1RGb48+fp2u7jr0
ZUyM9w0dP2wuKAqp8N5Yr+vtRDRDC/mZ8ZHnfFTVhJDmtSUGqg+QvEzGDrNOqa1H
040RB4S0iWThQGsEAW86TK6i1DdCrk4Z3Falio0p5vBzw3xoYHQXoucRjVAKMA5k
Nt9G4giMOQFdLVz8Ullro72V4GHrK4EbH3O5vDIGBaANpwiVDZcfuL4d1ohulovN
U8e9KcovzIl0hMT3FIdideCaLJBU/RQdzq/fQ2BYvXDMgWuhxhdgWXs41jckGier
0EFixgKku4hlTdSy8lp+4X7EyO/YgsgWX3Gk2NPPm/ICYyCsekk9MqMiIFbaoeL/
8/R/wbp4JUC3RHJQF6jIBc+Ta+J70Ax93LHzscXSru4LtVRJTukzzIKLm0wAjx3J
B8TbNT7UqJB0gmIk62/KmcPYR65VMkw1ICqNs3RP85iE2REOPRuPx+n4jJi/41FB
2uzM8gj0gfSsnkek+3PxrsfPf7Vbm8OZoodRB78oup7gkBYbazuKudW2BytDdG3E
aUFZ3Su5uvyYAoEJTPHwaSVTi04/stpFwP5J0Jl33MrfBl6iwcx98TVF4DjgQPJm
Kexlj8Wr9rrXkGpfU0vMhm3m3ZdNkrAGX56WTxM4dMvxWYB7+2ozBZD5vIVFaSdW
/rWTDet2r7tOewVNwl0rZ24ge2FGwlS/ueX2yaDHCpg8v/jHPE2jBMi1Nq0uDinj
1mck74yhWLwrZnEd0M8Df5nc1BBeS/aReOzEhfOA/i6wVgTE0gnpnlRXp2stCezn
8OQeJw73XitrY8JXSSGRtG6QfGwNO1IwuCBxi19LNaUHfpD40NgBKbt8cGgajVFW
S3rjb9gXF9tRIQINomNOq4mss/1I8vjKevRQ0Xdw4HdsXAlQasGYumn7Wz1Ely0/
naXu5Fk7Z30LWjB7MopkXkTCRurPGf5E7RTIQ8P19clRD1IDBikIzzEs7jQxoAPU
m8DbYaJP8jQkVznnSfJf2eCtZ2zTphhs8JgcjplX240YzxW9vveqfQKbgMPHmOc9
J3aOXDGoHyBrOx7F0Dqa3BDvIDpcHCYbyC8ROC5ynX0rBmJtOinF6hZlHEFhSmu5
MVPXrRvqoJjU/bQLLOlfyQvKaXZuJ9zOZJpBtIo+sEC3UlGjTaFQu7Gruh904rqA
YuY4pXelHqOSA/R59XwQFpg7tv6ttCBdGVHzq0H5K67bX62H6B0OL2ori60rHQgL
mE5klsS/MLCUo+eMEdL8zO/IQj36xW3vBcvH3QPt2uhmwbjV74V4+wrSmLNf9lcw
qsWG6eduUBxbbAReBjCmG0i0onyGZBHbMCFZokwEI/MWFuSBpOGNXDikBe8pDgbd
fQfHomqOVtQibKfdM0IL/PqYyTWQJt0lYqjw9MZtb43RfshD1Eyt9HjLZB1lHDj/
3IYsFs0TQZol6pdV36UkgzJW39hLEoc2EqQ7MsiwqsPvfw64eiMxTrH2Q32xiqvc
q8eKz9/9GND8Zqf0MLfdkPaw6YONeNmV/FTmZYBVmrv9JDvhj0Sh2G/i99tO6UtC
naXXqb8t3FurJIDNq9zDnkQZSFKTGPbwGIS5z35Yn9Zcb7819YPle4nLBcqu1SAB
97GspkQAM82I1Ex340SIse44llYNspD5CKdQOJREGvy2Yk7/c20EsDQ2iH3zu7e8
hDLQS6pjZLe9AArxwVbdnS9+ZxsYwh4+5+cpIeg+HGUDmaWOBcUHvLLs1nDcMLib
+4qyoba1SwgSEiN3DBiUiaKbo0fvby6+xkhdwp6lQXY1dfce0zZnrr03NjEPneUo
4bQFYY/izAb9FrSfcMkfP5L4tz4M7n7KRLUh3rpGOx7nYAgL9dUnRuy62JTfvrGw
fgxzQEwuwQyWfTknULuSrVD5zXYwgXTAWScCqEMDrCKigG+bl/CqSeoBffGGZSsE
cliQ76ifVQikY4q38xX4N0NWEYzvZX4D1eRBKxCJNtRmANFx0Uh9OFyBf+oyOI8G
4LRKRbYRT7h7HcoSUu9a/XeKE6JV/8VHCfo8eC7soCEFG/GgIilygbcJUTITvQPR
AbA1DJx3JKBp3fBBLUZ/l4LVRBDMlN42Vs5HETZruGMIVYsO2Pf5k9HaWsmQxnOx
7Mm655fZv73Wa6Ec4lY0Ib3RRRjWEcc1unhiQyzbfRohU1gVcNc67woEtnZnLPvN
baFEAH+CYn3Qr5TLLMDmtbjO9Gyv55Snr8nRyA50k7hjCokGXwDTxxPyy6qPKuwz
KtMPa97Ylg+xeDLya8BMi1I7HgTjzbGJcC6pxtFYKZxz6WNn0MTAJBYiQaBJQQsW
eAB8ohIV13R/Ja0TP/fgHKkqFzARgiE+o/KVsE/xYr/08/Zm0xpd4qQSCdNGiUhh
YToeMtlj9DHje2wrcPH4TXQcaGiTnIiKxYPUjbZPmuzR+2K63bkgiujKwruqU72S
dR0IDMauNtTE9J1e83rpEjCUV5yRPpsSnk908m5BjDdauz3/bpzpjEE3Q9b8Nsjw
SQ+azouexJMldY3KM8z7Nyrt7mI1atv17NkJHiNBVFG9lfs9cgMmos+83UIDSOFI
0T2eBgii0D4tasbulaM4zrCjEsPNy22VFOeA26VcnjnaBTsswXYorrRq+dNMEFpo
+GTvlnLGhOcerLKKhM3u1Do5gMKaekDNg3dlJOckkZLuo4zgu8id/MsCD4F84zea
uABdSqfQBjC57tWTICmSjKJYGCnxu6caKtJhW38bzduMkTMDRcfuEHwISkMW+rX2
TryoVwQdCfS1zeZQEa9NADyqmMhBjm+8XQLiMjTOg3jDyzvmHxIACWAQwbWkwepb
WLdByP7w4nyuUkTF+oQ8PrAfqDeRWI98/kEMShvL1pgHo0rce0fqyNSwPDHxsYX4
xOqQ5dIkm4l8vHfpuWbeeB3GDvmwCnLVyLhWbOQAC7y8nngmA+t03AvsRK50Zb45
rZi6UZZFS7HbRdnOyGwyb6KXB1ifNBQEg8mRPCWyFGSlNW9zcolxm2z9SKpXdebb
Bm/7YKjhWA1cUeIE/0OHRSIThgbjsGm3lD9WvuK3FzLEX9a8YGUGyc6JH9FUaiFO
xveIRWTsPfxNAJ1BOdiGa/vzQ8DRp9VsvXvDniqUhITq4BXrYlKtozvzwUgR3mB4
m3bwwbB/gRuN4zIiPOnHbNOHBq3uOVt5O7b3dhrflebPh8J27zHORpkMUkieVFj3
Gj+GIXkXdjYdjXki7SuN59mVUD/X3QHq7NsS0JVfXISomCeJX1TmkEldrazVpY5K
jYWX3FfRYBYudaPlnadcIoZf2z6z9uaiti5d06GSKRWsd+LMULrrYL4ECS+jSdVv
PqioZgTENGLjSCBkfkhINB34QZkjOGWCAJEVrMNKcBr2hRZLEjIWprTMfXE3u2Mo
vxRRwkYVCW9TzHELDaKaF8Caa9KsQItxMwWkxbjaqTiPpAlhO6pkXl9FnXyFkE9c
+mOAhB+WW/A+tf17a1D2EjoqNhFnlEXOzBkveqHCv8pZkXsl3ZZIFBR3d2IKObOP
0XPLYbyw7rNrgZiPdxdjTquL9D1jblcV03Ksq4tIV7jbFx5jcpPNwK+lzznCKCLD
5W4pT6nuvQChbu17gmpxz3zZk5cizhcON4coOwp085foIY4sn7gVlEZ2IesxqYrB
LRHzgZv5v4uyZCN2nstq84u1ndMXZZarqZHSmlGGfaJAXkDUVuNvX0R6iu1FmD1U
E1+av2l+6XgUtwqyE+bvA1BNlf+zOwHBigKUwSN8pfuCHyYrj+Ee5orPlhjmoAXS
rELm2PNo6jNhRZtMaTwhMm1YHidV72Dco7vwHGVz6RG0eq2xQco4bQkeoYaG+k0A
CU1FjfugQj9eo5hDTvQ5Kxux9Wj5iRIXZl21/IxN8OA5ZknAa51Z4DOfFm3wVzJ9
dHuezju56OuCjdzGmG4LLrhURwc6JmbDpFpSWdy7kF5HmYnrwsDuMxj/MW0/6rfD
wGpcRsej10c5SvqBX2PtPKv8o7g3ugAh3Ri6mjCzCrBt3xDRqsSemyZxw/CvwYq0
nzUbumZt1Cc4UKCZNWFgOjLuq7WGycaxa+1KAuwQGcb8oFsbjFnXG3R1luPhGfT5
vZqMcW+fzGUAaJqRd+1ImBE79tgfDVu1LruC5CVnkl8vZMbpPBUP2ASOVV+Ar/k1
mA68lR3SePRGg8HUw3CfNDjychyypja6JF8aSsr7xUWHLz7hP++A/hkV7eiWKBPR
26/UqoMUcHQR7Lr0tXi50dm+xf9eT83PTSAc9/4+SpPH6p7dw2PcohN6VEmH42bd
lPmAa184+INQXjbw28JTq4AfUO2ue+30QxndxTvvqZa96G+Yg4XI9o00OhwYQxcC
EzDtfAUSeubkPE/QWMhj60DeDDfwCFzOsFv+Tke6ixXAMsenxkEKo3XzZdSGKvuC
ELqMvit76b9S2gLvPA937GL52Dl+HmF95LA1ZdkBwelb+l+72zXrqnieV+DlQqmj
VjylwHKEYG0CJPQTISfLCttJ2vrBdoBSEn8uAX2/NTu3i4rE776+M2ZwgnOhl0am
NYl386Yd2qoU0j6iRR+UuwnCl2bHf2gv4kGWd0yZiRsT4Hp7Oxrp1TVyALscmLSj
d9w0Prc7KlIeGi38UFCwiYboEy6qo2+ckxvxR6d1kJ88GF47eZcMrjCQC2n+h66g
Wz/rWPazeThruLVv8sJTJ7wau0txwsBEpxHvvWF95cmkFu/1jGpLmK7qcSLpnODh
OjTNQ+iUkeeHEBOwQNiymac8QEWxqDq5p1Nt79CzPQGD/ZlDY0AyhMkHFci53TCm
PFRSYP24Eky3HhHCaiSdSjojaZSIY/tuKOf9dssQ5Tt02SL5iMzxb09NnGKbvG5N
dXtDyJibzg6fHPXTR4RGPbVfq9HCqUBE8nfUOcNFhsQBdPqboEh4ixPRtSqi3TIQ
LXxpRzkVOvtWQ65mGUJdwsuabrC4WLXsOb4yqa4F192qD2JyZuB5U1ThccY/wfB8
oT4QNHsCmd8XtL+wr+Q6XBkTP36WgZDEOcmNqUNvQfNLlXqsji0UrZZA6ll4HYK6
u/SCHikeW9n7Tp6Jhx/DZIim5bvIpJW7ufLuyaUkgUyD7vFLL0ha9IDRRXAUR1lS
h5V8ADEUrDXuvS+GdgVWwFyud3og74LyNA66WaYR2m5nfKojD+XULqTwAOjiD8MP
XMnUZG3ErFmeD35zetlPAj20NgcY9oTDaJKHpBVuVgQjcefXVjz3tne6CdIxGg1o
CReCZkqlmZi4mh19UK0Wi3FrFcBlMCV1kttcniWTj9ByH/nCT1euRlaRCJHB0KDr
yUtrx5bpVpSfLoTdYaR3Q5UrFYZARdhIJJ3DiWq3icDFXQaODHXDRn6H8IpsVYyA
flkX1qjfzh2aPHVJGNADkNU8VHuvZSbIxr3UvpfqZvoEvKBEEfVylN3EJArqL8KY
DAaPW+u/2VGM7DXPEuqfrTM4GDRTlleY2oJdyemO7LLN0X+Hnywnyl7/Av07KAI7
HpxnwUSR41DU4UNu+iwCTNqwRNDIkNJ9XP78brgHa+1fBiXP4TB2Tk+RpGR8Srxv
h4k5YMmS7rSvxTfBwdO/Ks2NnyLSkdi7qOfgzb8q+B87+6GZ7UTIMQRWIYVcNr0J
sD6CoSPpSconRlNDEjVvrBtIOqHFlK8ePKqx6mtd8bAjWF4FbV804aFnGas8XlrP
0xIyMUe3NUrb4E7raeI8292r0G12b67uM265cxMaEDp1CcjBNL99cZRAE4Wrt6T3
tJBkxYgdIBG2Y9mfPCW4PU0VSYMbIWHx1qXXbYirjVfB0zsy0rjCL9FIzr3mGLyW
OOvxoIA9gr7h982bjNlWv4/NZzrS246RKFhVoHGRxrn5+g9wkD19okcUZ6sNUIlT
YOUI7F0LRlwrHYIvoihFKZnFIYkx9XrPYMQXRNhUej9D7oUxBsOPKbYY/ap6oBlc
9IWKpUdwYNgXMVxpZ3CGZj5lxAsVvC2cACEDb3C2fc4z0bkXgTvSWu9r/Zvd8JBN
ad7a6yTqM1PIwPHTtDJHqRmqgR/mF3USB5ih2NTFgo3/O5Cb1HU/X8aenZUsLmKU
FL1A/quJ7nBfgs2yzLljZtft8kl+OAEHq8fN7Qu+QsuyA6OzeI8il/9wbgfd0lYU
vbQ+hYU7TnoSHOHAV5OHfVCIOHLsb46WdzZqihk1dtuoqvfIW/cJxRtBgmvNAelj
bb/zqFevBB7FEeq5nW4ZcJ+BXvgSm7g3CSZIz3v//FUNTkw+h5zBWqKuoskGNKtZ
O/q/xw7xWkpsV3oYkx4yEXc54veeI4VCHvAaYtL6bfbWF+/DU3k+z8Uv7FD79A+1
DpJqV6fcP+6G2/eVUk0YoFEDuZKRkgeASCYZ+36TSFZn6WEQ3YyZ2YXvjYVvWvs6
TpCUWzYjkTFuTOVHbLetoQ40/cA/wwZz+juDaj5nCnDyMTQsvLUGGRvVGDdZfPt1
OZaEPGkffmj6fCVTRIu7YfY5PZWSyPfILlpX9B5b9w/pVrclcJ/2yrtmBsbF+T6W
xvcxujR0P+ASBd+JDyvjcHkSP3X3h5xV17mwPRciSAGu+2xB+y/ixNeJhi1rIfUq
4ftKwtroc3KcN1yvdQ3HEM8b100QU/G6NSqajqziHa+Ed4xIXZjV3KCGnuGftxwR
uV1YswcsHlGbVGKVynEgEVk37e0jY5WnkoOsjWrpRveeybiS4sgGyY7d1ZSFWzqp
As9wDKaiUgHOKY/ZF9j/L4c0jsZNb+NARSlbyzyyMTHj78kyurjLWaDLuQzMbBVK
U482Cd4k++FHhC9LNu9mv3m4u0FhXNjNO4DNIpmpBaB6PB8WCcbC4q0zfFnoumT3
3ZPretlgY3NZ9NTrb86pgG6LFGhi9uhqdHge8FIJQY12vEcG/U/N+9ztGLdxiFr6
zwwx97cZwAzj7YS1zkc6phjq9+CsVwmDZnn2qENKh4n5KpRnhmR26w5sB+U2/CMc
ESKwmYfe1h1QitDFPqvEAFoYNqKCmRFh6+8T/EAAwGAWJ0MjSVBJWFS7L5QE1uYO
8s4HKFUVhxxXeCAPk6CchIiTmqhNMNSfEa0su+zMHPchWNea3NMdKkBTi7KU2NiA
zp1VEIr1878FJngr7Q3OvgLcSij7hPOxuJ3BW4BM9SJvpv+WgsHUf8h51oroV+nM
9Cd14955h9evsPLAiiWk/DNsYGku6RKZ49yPYkOJSn/S0xlhsSZdD/ijQb+M0oDD
jYIHEhI1tDZEPQchTbS2dJE5W7K61Gkl39R14wzNe1mAAoReFWJRdBPpxjpYO54Y
IORp7q25ue3UbLdseVMqBQRRgrsd8XmQRtqCnLo4w9T1xt226Q3HfSnyJZzmmJy+
dcM41kAsCgvNPpV0iMsnF7Bv6Z9Uy2u+Qa6ZNv8N5KpAkD6uZjEocL0u7yP4FA5G
XZ7L8eVbq90lHgO5BO4+cHdfRSeBNq1JHgEDR4ePWOdJ59xVReNh4UyKH5VCdzXQ
E+SAIePuXeWYaPEnjWhziKsI9aTvt3tbWpf0pNva+Duc8vB6tjZYqic1dCpYY22l
5S0xuIRj0EA94FWFOG/++qe+T5yoqTDrwbU5qqbvg9HzNxKY7fmI0bC1AlpMBp0P
SnufQlhbCDIT7Vzg4QJQNvAwYz7ESpHKmuQu29C3O9Y9qh4qbiDK1UpH5NV0q3OI
cw+AjUfSErHJLjdLS+r0NOLXFkkLsrba6ajWFannRa9FrRKg+ayTHEFzKqORd+TR
Q5TzYOX8xr1sS2bDj9z0FifqomAIrgSsF2fDpdDCJVUot+rgwB3tyBsrdU5x7BVq
rY4Qq6d/W4vq32FaHV3U7nfnLqcDZCmeCzxNiYugJGtJMF/rP9t8aYT7TA0wrvlQ
5NgGbT+d5gpkCsu70CeiLwJ0aw9DG9KUB4QO1JA/f8H74khZmz5h9AbRRBRQ8q+P
Kz9XV7esr1nZ69xxuzeD0Ysnd8vjsxZUOwq3BaKSguBdR3AnJNB2yO5d9tOJ8QIv
njSel0rLOlmdU3m0D5EaP6gTjPeYrfFkXmFFQAYC7u1HaZfA9iAXcLLXMp7jwXYW
S09IYeo2nxl37JNUT6lZ1NbOY3igw9XiyUsNrYfmD5M9l5s6z4c+f72DlShy/fJM
9we8da9PgNvKyVARwEIkLOUWLGmPJGjheXF20PWtt6hQ8cptBbFWB3fkenf3LJhx
XpXS065401gt7dM2H1WXMFcOPkn5/G7VXKt+iV2lSD4doNPihLDcYxJ0JPEmJrZ0
pUJHEHLFTrJLkx/E2p6uUEX6tgp5/vHSkeTCDDLvwMLn5LS/kD1W1d5r7uR2KkOi
0W144PNllKLjEJiznGjP2Iw0uyL6wrRH/5Ykzf2kOYY/g5KZz6t3Lc76zLAzeQ3Z
anrAOkbCydQt+QE8qzR+nGyLywKJxKffTeF3Kh0KC95NLQfnrS4/2gbJkbdbB9x8
K9cawRVMOShLpD6YGVucmJsD3flOuFvDbKlbgFiBgdqNOTjtGmYbNJIXLSmqxjlX
tMAz30Imir65m9XiQcuJfdumtoUTrEeSwJ7j7fBXqWHdBei/aeV2JVRzByRdIpZr
IUJESYQuHzZOSbmqbu0PaHVvYLgqokn7THljPNKDsG0YoWy6Ubbbre7AuELdmgGV
lHqAJaDUL/8RV6LETKVWAgsFHsy0kVq9hAuyvGpzor0rBLB5yMwItYLBmaXYNsk6
RuEYLFG8S8R8uSzcYqZL1F+d2McSkvw1qEeRuyOBZ9zl8I9nef5AlsHhBknEN6+K
QOrR/zsPmBbh524mrH7tSVI/oAzpzv5dkhSVCWj/yQuAN/m5nvgM8hCEUwznw3RC
7+pK43P8NPTzEJGVw5mQVALZ3Hqrhlk8MGkDyRtT5yhMdqwiMypGOIWgJqVTifCC
PHWEJwth9vOA6HT60Dr65O5UiCIdZXTQJSmTuJSMklc0Ud1nsrTpzGIiBDB0MWej
xyXPSnEFw6UYahYvGVkhSL5dPWqkCqRtNyA520IHE5oKx4jkUEcfE6TLBx8eCfhZ
G112GUQU1s8cJ7M04U9gCMJsN7zNIrhYWS8QulAbAHxyaQnnvXIRZbEwlTnMi2Qc
Go/4lgiajn+vTipFpXA/moM0/H9biAzzOXlPIaWxOv2lcqGz1Hm94Ij8Ks/g02zV
qXnZfmeBS/BG6uemUb3SN2TIMpsaBsAMXw2bOfwhI70bPmPVX01r8iqMgZQstDEv
qcvyj4V5zEk2+sMY27zlM2XqNEx83iaGxP7zfW/gQr3emF9v49On/jUh+dA2TwVX
D/9Fep86QtUqWwEtdgfNB5qMmeIBBQ89hxp+7MhN91feTuhEVd4TYDS9Tgi5ciU/
po2SrM4PpwI52ep6gb03MwkefspO4DNJmHw7rwWM614RPAcG9LJYcmyHxmg5e4G5
mCfQwzd41yfZdm2b3PaUK8X4f9gRYl3qYMWt+18rBiy/nmsYYhKCMUeKWKrKenlm
lBMiCb0kg1bb+ejS1rSM2H+0MozJ4rTxKSr4G/77LQ78qaHrX5taGBr1LCTAnD0s
74HgxNsRsf+G+kGbtycMkDXUb05g57ZND5MUIh0aS9aW/VEHUUieCTEhEjJ+9ZGN
p93lf1HfPCkeIet9AFOeAc0kAZ+Krk+pae2ZxHfXSOVPDCofK2zRU8w9ILm1nU43
WhDEphNGnMaKppnZFGxMDfkoRq3wGZav8PC0jFBKyXdOnx+Eh3aWWRn4/RqP4eF1
qT6WHgkJDbjusBryT3lNupIeXMHAunYcj0Yi2MQBF3NeokOGiSshYO2HpDdOGThv
Kh5FzXApEF7Gz3uEEkVheLa/qAPcl5kqM4zRmmY5GFhxrwvZSP+NhOXIAkKYrTWl
YRszhMPU3TXql7eC+EpYBngVmG14Su1nrbgCgobRQG/zw4MDUv8wEO7VDo/XXTel
/huTZTYIXbZLn+U92PZBCED/q45m8xxYV5XG8Vwl3h0ON8xEh/ZV6D4PcaS2Utnb
UuM5L7jEBec1E6NNEcHlBvFp1OaqhESzZIJ2RNX5SD/X5oWsQh1h+KsEDiRGdTgB
eW/PbNeHLA8rOJQI5EATdnNjJ/vJbZFXaUX9sCyFDSWUCXzcsZBPm81dutjAmvmi
Muo/VMGZf0iGwQRxbLxdC5MEuZ4cdhFHta9UMd186bEVc0LmtT0WR5yhsEDp2lbM
pTu4KWEta1pldlMSpIi+BrwDtOMcFTdNaEh7EO+CL1/jiZlWOAyZVabZhCecgPJI
+8uEa+1FgxIcjwDIOFSAQkBhFcYsyNiA8y818NUNPhiNim6Xyb/KQsN49e1sXeZb
ThcuUYRPpKj2IcaogfM8nltagu57FXa155ycJMlEM4Fc+PKd1viHPP6UcYtXuQZ7
k5o+ExSEECkv30rRo4mQ4aPucz6te8o1lnNt30ufTbTYsfIayGi8fPNZXNXTx0K6
weuegm7TTXhRWW3pla0N2GTuMKI69V1ROwQLcwNNobLamUc+FDbyFyHWlWyNzZz6
eFy74rwH+eRp7BO9B/C12qYE9I7awOi6tpgPvaW1gdg91LOhzLDy4LQLJpNMzps5
p+nufsq5Cjk5UAvrT4rh4phiZGEzLZzyhykoI6lhTfAyuImUhcj+wxm0sfMt8ag6
fTgwWp2qDN9VfvESeZGOvSyXD/Mj3PC94env2i2rKbwsuWVBQGrkdK6x+M2tXiZ1
TEBbTA+A+fX35Ybod3fnNM4shn/sbmJg2VatETUUF9O35ffOd2nd9rD3UDKQX95U
A/Ps3fkMCn/2AikOYX651121QNbo6DI7PR7JVDuGFC3mAwRKB3Wiwg12aRUPwAN0
KJLf5qUEmWXQMQ6yhUZTYy5yPpMpAlGO4tefYB32sQFFN0V+nyYLs7E7uBtb5she
ITPXZZSW0+ZWY1Ov6N3efjQdWA7EPP29A0YCaFSqPs28hhZAWTupxXI0aL9ezK4O
5QB5q+lQCzlzcmiLU6inZ9Zb+ihHw4+MLG/QD2Pr9/FKdTBeBrAwshz/qMSKQNiz
K7CEyXrpaD1GvJ8ct7P0UXK7OuUTj0h5GH6HprPSzpmkWB1xl36uY5NFvpWy33jF
08d58p56oi2XL1Fw54CUyvVHW1qJbv1sUdoUFXk86XZ7PaxWt2TVxBwcH9ix3+y7
ClZ3mkwc45f5qh3u71RVvMxR6oPwp5NtV+kYksbi82j1pu5X1cZl9NGLI5dWZbf4
vdUP7Hchp/etuq7hiNWE7K0MKz6357mvSgUy2XaPJFFMWiWL2wgxi2Epjp1puf8U
sLUy+vAMWLiNo2dp9d0b/aDD4rL2vnIqST48NrsXFUCVbSFaD8PJqikSrPkBly3C
6lgxR2UQBBpMC2IUYT/4FtL1SnTGvmKV0kJyG096FbZ8kq1j2Ui9+/4EVtIZZDLu
F2awpCuM9rJFJroMtDQcczKbHuMwikGJPSq4AEQn7DvmhJnDQl7RqKAR0iXkcD37
B86KHvL1mYysEuPy8tANIWVwaBVJmTQdFm5c/1mh1LwNbszwdHgPUsYLvGRQqMEj
0pQSj9m5FfW0mqpJEFTDIMYATGmNT2sJ+wxj5SnVM2xHks3C+Voay9V71cTd3wOH
MIElWZ4CNjJDm9aerfTINZUErpSeBiz3gc4mem+ftpbsbJ/FsxN7tb5/FH3huG8X
7xS4FSIOApl0gfnS3P8eVUOeHHG5/BQV9I+W2RQorS9j5Xn9fpfsIIMAgzMlqKoM
ced/k4dM9LXe8tPJJU9gGyOmKgFoAMy1Ar5ZjYICcQxwvUV5FppT2uPl7rp2rWO1
jaT/XYvc9PRdBCF0gGm0kr3j8oEKrM/oRd1EtOCvjf/f49mnSuZeXgyhOy+fAiRz
FJG3J9DOMzFcBwiyhnKtQZyi/vFC3GUDAf8O/yrmTtkG2RpzT67ullxvgLDESq9q
wpsdhFWSKZ4ga11P4E0tKjjkvPlCJ1zn1vL49EwXzF52iurb3wCh2I2vRKonLg+4
dhvEmm9FRTeVGtiNfjLjF0s/ykJdNTlCjL1M5LbfPY2rIGXdLYhCxdSNqhm/RzuN
UjE3v1ejFAgQ+cfFg/Dlvp8nTiV8tzugn5uDmeW+41VC+9GIXwKEcq1gcPDuTAH9
E2I/hEX1HL45qd9UXtOAzInU9D3rDycesWVYV2TzgaV/oDRDsdz30SU8tstaAnpU
oclkewd/Msg7hTK8aEuP2WE3X5HwcsU8oRzkl9g/H+N4M6KnXjgX37ZTmKuSnUnx
CUoeu19npkm7UiRZP2PKtx1TozsDgwy1IuwgUFsz7vDWl0ee6DH6eAMbpXUUBvNq
xQ/rkyUlRMwt/Muc2w6nh6Ica7KvQGu0GIXdRxRfk4olGd/PfxaFxomKj8PRhKZi
UC5deRjb052vCcVxWhhztMOeGduqOOe+GQO6JHLScW+7qt0OgsU5mPcE30JPhYW5
REdCilrXMeI8Wrlh9h/NT8STm84PypSKhNH9GMt1H8D0virl5slWLBXN7eNdjp3b
xEazgEeVUcMpFQATSzINhtG1YrqjAJKd/WMy8f6tVf/q2dysD0D/5TAsNHq3XHCo
TjGkygYUx/14XYETeu+QnPsC0aXk4BUJDhNKRnXwHtTbuowNDDiCQYg9VJL6RBju
YpleL4GxaTZYuB6h4uMNmSAieJELpBdkNJyt/fJhPSuOBRQD2dfJYC5evpAT4VD6
+SId94ZR0YWkRfi5DsQbZ3KNyp5H2mAFzf67tjnKyDucU5kNMP/V0pn+yHylhe3v
AFO2PPTKba/lJDOqWKZAbjfbKi9FzSE6k+wBx5dEEZmw3WRYjQgrRb/EQ7wl9hj7
N0FpBoAh/CGPIgJ14/adLu1Hc5qhh/XJ9yPgjujKT08H43+Bo5KTg7xv2FCwvpEO
evCm11FZDc41zJqnxcsApjHal2JERw9vL3obcm3LuCN3v+ETeWFuBWuxeZVx7Kc5
URk5wcyhLykmBbA8/0oS3RveO7z8/IQk80qqdn9nK2ZvWR/m1+a82IKnzzjM/vvs
dYPEQFd/JIkc9KK6TEUKXt0h+5y6G5+NhWVStheSZzjcmiKajQCcUKOwW1C7K8bk
6lrqO2qzpjtZTTrZRqIyPGOIbyl4oVkiQpeWWQo8FQVvI4hittEH+ulTYFowOVNx
vCB1mrQdWIBTrDMN0Ft1G2dyWsk0s6/FDVxZbeZgIk4ZKTbFb2ckbHgrXBzqhsul
c8VdHsVCo3XRpMzHIjQSY6iPYEef1Mq0CLGCLvFES7FKB+0t1Ba0kjzTxi8E0KEz
2i23LIgeQkmnUBTjCAjzvQi5f2ej0T7Ud86R/ObtLUc1LAKu9wFiZhl4rAMwsRNW
pCZFoxYbVGgQCTfbBzb/LUyxwm0LVZTKI9hpR5zayWNs1efKgA9t4+81xxpE3nq+
ZZKRM0pdc/heRK7T4xUikN1R6UE8s5id5RZVLYxUzZvquUOKaKkOc8/+zMpWxHLq
tIBMDMgq2ZzTe3h9mik0zcWc2TAEKxcgChQ/vuz2kwbIHmyBuwYnQon9yAO7nAOu
sFYb1lmAOcRqIywFglaCQ2KqeGy7umPVFZ16g2xndSiNC9IJuG5LpSC1+/m7JZZV
70+emb0ee1huKqJxjWHO+KSwPJph3qSMwkKr1s5k1TejpVkHy5KnOCZjZPIXk2U5
oJ+tF0C8Gm/Jr7VOYT8xPL47pV6zy5wVJQ9ESBbc06kEZLDZtqBFNwWNGSs0Ck/r
UCDEwqYx7FgrR5jNT+VTpK4xHRKIT/9/L9Icdek9Mg2n9ezRLetetf0/IbJ5S5R5
LuBePIfVCMk2EWD4/Wvbz3llyeNRfdTEc2ZqhUqPTyMJ6LQDE6WlR4mhOP9W5VDj
4Q8WJFEOyps5hVWcwj6XGfB5ittPDcBkSxHnXhq9rwyxNXIKNGhvdGMVMXSYGjCc
Y6wjUM7Zdk7v3SX36FE3ZF1R+ohYCmS9eH2keLY5whkUsStuQBMcakHEM3UD1FRQ
MfPvFgJhv4luNPs1txdNtmciyW8OQ/PmXZ7ErLeTpjHrp+QctVwi586ooQhOKDs8
TJpTfyQlhofzyF5EgR7rbXZ7vk7N+lGT7EbXJUhdxmShshCm1YUAy7h6nNi7Vtoh
VqNa7qq0bHUXatJf3XEb1bt7GS1b4dHYoFaH4eA1T4oTOcdg3h3yk1P5PD6lB8FG
oi8b+wFwfk1rf7ZhcOxZ5/wVG0+c7zsgg2hDptjFvs1M6FB8bEu2zer3+HdHirpY
t5bTl1gLTHduQKRHESQITOr61oUn3PzLcBBLol46QFcX79jIqEcxXRucsvHneJgX
m7uNlxGcREgx+HTX30LHHoB5Od8NbBNApj11sfG0LhM0KpkfYAiu5r30FUoR8wMs
4s+8rDIfEIRLn2Nx8iBIJT4gXUyk2aIziIqRpRhl4ml3JG2vN4pxAEd3vzYou2uB
csuMd1hZnBuQKN2zW+O8H9elkBKJzcjINntJ8B4LXTfr86ylwe0M5I1R8+l1mrzH
4Ag4Du2aKMhJEeW7NUlKuJmsoGxPThRrFZ0eJ1eKDs2EGaoh2e7LceObv4gp8c6o
Mulea4622z8dbJYU8h9vB7KODzJZypUb+ZqS5LkJ63sHbvlp+OMKOVWoBMD7TH+G
uiqvaBar/9kNvX1VO9KLM7XuIDgh0zoswI5X/7hVSHlPQtDR+H0MP5XeKxpJBagM
y54xO2LWFqUkVNmzdJhQB1fHB8uisEbBlAJJHsFypNqHR0eiVZs8P5113bnuz23h
Rznp8Sm/J+NUeSW8AWSMpC707ss+cQcPq3WktHHUH8ixNtjRkfQGSkwSX6yWuuF6
FlKFe/CFGqQfGod1CxTdj5sS+xSY5B3ofL8OwhOtmbxMFJtVYy04P4RpFQExxt09
QHYhYJffHBRVBuKL9HhkEwxTxECPnABIa94UJvYwYcmxPG8RYRfSQo9DsXhFaKQh
veejkO6DsnLdxEgeVQ4f8mJq2/eeSV77h79GbmyF7jYaqDTMfg/PFG9QIaTy5jwp
fO4N/czL1u7eIaosNjs+GR8vM7HiVfsIXkb0h2d91vto1iyAeYE7Uk/sX4zO0OFB
DsywhxIodgHGqx6KVHsRXlo51rxtWV2a9gEpLJ6diz9wK1QL864pcprwQFazjs77
T/YXT9rI5GatnDVJj7zn1b5UVwcIJONrSBDucrF1BuPUObyMi89PrTYSFcx4kfne
3sYw2XactkAETZJZ7nfKN1I6bRzuDK/w2pMnYJec63Q3L8mChGJTpMxCqrt5pL7m
2v6Kl6EaozPWLOpNUk8lj5vd8DmO7Rg2muId7sSMYOY230ugNhmlcNkL20Elet7e
uZ+gIk8DetTZu1lO3P9DWyweg8nnRSmiata/Ul3f0c8oYW2giIhkXKNBfCGqhjE0
gfMFlTOCX164BcyEwRZfgrms1OVjwgMH2pUEv3DiaIOPf+Is0NGBweCNYIi+vDsl
YP9nAamA3fhtDNF1434c041DAU48uNnjy/7a9kTNmvNQ2+3ZpBa6/G70ZmaI58AN
RrYI5hpDDVKmUxSHGq2a0jnycepRKZpdVRwaG1NnCjGd2uNJxjzy/G06tawnlhSN
jYPLWzELzQ4aaGEzO0ZhxHZcmRSKQfdgeuEQimoRs4dD9J/Uh2lzgSKLfsqEfQbG
IGQNr219GbcJ0TvuqUn/Vm8UnD9d/KUDKaMsuWmYLVecupP69oS9RR6gH5Iu3AiX
LvP1kFDzOnA846lTG7blw7eA11nsCqsb/9SOlfZ5qVfYreLxorAPB1Q7czIgtvZ2
QgR9Zs9EDrVYJd2PhUIan4LXkGrRgyR3cmItzOIMP+esvN9vYsW0WIIRJR6gkYXK
x0kUNirxWtHmHGJgmGfX/KKHd6NfnK3Eb5DkKwbIr/pAeYwOSCpK9joRbbBNYcpW
YhbTL/lOAM4l+u8psrbzG8BriDF0nze1ZUr19IfRao1nXbDELZLPyqbyHs6bWIGw
D2z1A+kr2GaIg7n2q/DUysPLapnGkh+UoR0kvYNqJ258u+qRVvCZMrkH1dnZW/5S
bwggxR43vHU/4ecVJd/3tMhsyMBGJTI7eS56J5TquQy8So1eF2rYqrAyUEHQBuAF
APCQ9xD0DyyRVDeE+3yEY7vpOPeYMhVPluT3DeuNQkbl1NHvvQzncxJSSy/nVcD1
XZMEwOho/3oE/wp3inE3dwTcCr0X2F5bpakMvNWbjjuOLrdKpob+X20liL8oQO30
05H5fXJG7Jxc6qUNqnYi9HfeVqpgASsDocxIPZVc5M9xoQq5Obo8qkT1W9ZzOC4u
MblFtWzLaqbx+GKWjrYgL3TUKgp+sHvfgZbDF72KJpY8ZQJY/LIUad0L/je5cUOo
cDZjlPdZLcoqbCBhYGixT2jvk03K0RlOWG149wFfEF96griimCQ3uvixLsEA5e/d
tlPMNpgKkMLMHyDOXoGKdoDfq+pAvqz7dRHjTMxvkX/YQQwFzRXTDEI+kC3ePtHu
HSJTM3pmmoYq5XTctWmCGTWuQJzKPG9Y8jixF9U0v1bKjavAQg66wYyfLikvVZVD
k6PHZsMVyMRQJWfUL4VVkbU1QO3AkKVuQwUwmijqkeMinvnoQvM+iLHW+BbGtUHG
63k2zRTg7iXZeJ5TAWFeIWUn/7PHPBuin0gzdEmOicj0CMsjaMR05QfjtFBtpDDY
kk9oU2RaynMZ9cIk0Cz6HQv1nXqK1th0xXy8OlvDgiwxxnIsuk1mht1vKNg31frg
Xfv07HAVmicglAmoO88Pril5ISYhqnRmz3TfTC1nL2Us29Kxp+UOhTGXdDtwjnDA
baWbD8iroX+rn9jbp9Z3qPriGkAMSOEVkV43+MnzMzdiSZw0rnGrNvoYtVJ6vHvJ
rpNkmvkaycUL5VK64To9wFS82SFk4FZSaOVZjFVGodRvzPOeRGeKVRoSRRGu6k3E
EhJfNKtJ5EQXJxTlm4H5Rhsk267hZC/1A5SlFbhNPSOK0gZJ88BGG1B2GxDLkfvH
MFt/yWkFe3KVQ6V834smBFqM9T4PVMeAQjMFX2sL9xsOm2a5TFFQ7+Eu0sFo3YK/
gqAmCkJFR0qWTJpqrKkAzknsLN+vWJPWneO6acQSsTtUv8GtkPZZ7/dwahQhhxdt
92E3BuxXk8/PsQ2K9bjd0LKoTujcv3lODlEWFtn/zrjxQD0lOqM+lzGiE5V9JXWH
VN1TSUpFd6oIuDjcmV0/3VJGZY5BcuAbZSwUfsdBmvuJ+36jXCxWo+hSAO0Vn+8B
Ch/5SxMEeDBH0Wged4DiSNexD31E/FMuopuwmEK8bnTnh6aM/+sYWwrdrPDHmiuc
4Kll3TUFDBvibPxQnWbFAfw8g0btggTKkNGG9lgFtoE5yktAyoLVpM5reNKAif67
W2Qo22cDjcsMt+UJ/aMcyxlU0WvtaXwR/HhlCx45XSOkGV7GaTLyAlOTtXPxcDEo
WZ9KrQk+SZ9jVvA91CJymWAP/naSTbVovHyppb5bRYjmHIgJgJl+Wcqvwxt2dqNC
ANh26/Q8fqZ+nuRQ7SKLxrDtZ+wfHRe/1RpkZ8pE6mJhyemZVYdARDREkNfOwRBc
1UvfahhKi2RHMWgVtOutDwv31xlTAZ1nM52ktd6FemMD0tytT7137dXDcTWGVsvU
IPHvyUzzBsY3lSc5DCq9KvcfG9Ld4I5XKwdECWHcifEWmTVAhwHBLV8GfltgzSu6
7ndjLOej9xKo+ZD52mBn+5PuEQ+WafrdaMqQ1+Ucq+J4Ea62D78uHSRPvV8SaHnr
fGvvFPCKTaK9Ba+gDemE0rCpvS4UgaJJPi2K5HHaI8/rkfGNgO+0X76fWPTNKDbE
ijFTZQ6K0PsY/abrZyRpSn7fGE0n02+x2dIV8afElxWNWa3u4QhAxChb95nWCPMo
CuBdR9Os+W2JIuWAVyotTq+tuRXjRC6OgjbZTrc6OEQvYTBKaL0UUP+xZwSDuLpx
Psn8e2cuE5nYk7yMeitykajrZBRbgAxPIpTMVO/k68WblN/n04KPfHYhukZXR0j3
UAlzl9l1NcUNuR53b2RETEB/QWfQpyZZZ4Iv3xVZkMzc88rf2bm+59VKaCFFXcB5
VFkYLbAgeUYWjhKP6vuk2jT6wTe6/NkANrdGhiHsHmeQ+PFmURhgv1xPgnVIPegC
B55Q0fcnOKS9g8sdkR1YrNgJDX+gW2KvoKziz62MACn/F3gave5WENI2wwfA4wf7
HnnAoLZdDIdkBSnnAHO/0Rf+5ipGYtf45dkGfW0d3VsQsX0s1aAUiVDOoe504NUb
eLwWKlER7coIzW5BpGeofPK6NRtaQiIMgVLGL5G5rzX+zUKNiRcCP54DL9NJ+Pks
u8zq814j26lnA+gPIx8BQAGDdH5wSQldGyQmBplVjrCGP3+5ZzXCd/mgoPAF0VP2
BaPjfMD0K4IVRg8I5uV81UJsm8+seO8tIcsp/fz0loQfN6mH3B6A0saxQM9UBI3A
RjY3JLqh4DI4HLUZADrpLnX707QQcaK1584NHbU76Vm3J3Dz8K9O1jFoqba9PBRg
J3D5S0UMOLsbz01eZDkOIhHTaTs44JmRkdAeUFn2YEKr/8NZdosPiQQ/R6qpzXCI
R9iFCw82PEzqseocyXlCoxvB+RxwdvvHtT825559wY8G6JvSrVgoFWQOszZ79XsJ
l429F8c0zIAk+hbyDYAboBQD3TRWgj5tVEsbHBPnZNdSVdPV9ZkFcKgm3e8HFpgX
BNOlJ9yT18N+Ea68jOAxoo5W18fZ13S2fC/UV8TEHlwTln5NOYxD04RIMY1Umnde
GDNLe4m1hKYJuOUteC1wrkBD9Ej+ZG2jap3A/e00J2fxZdYvDKwgbiv4jttaj9ik
XRaeisHIqSvS4EopL2gPtPglBk7R5SQOZUADTK6Bm720WRLeNNA65cD/qF0eYbjR
2uofVBaiHbaN3tm+OWds9yp/0PwP1t7SbALwGCwsZHdMifJuCLVGLrHQQRfA3Na9
MPQlLwkKGJpxMybwPxuaW0UHZKPfn4r1Zt/8IYgDaH6l39yhltx+y9D1BYhnXL8y
ZRwl3Mj/Q/sLs/qL8HktZ+2bmHWK/lT+NN2DtjR1XYKFN05rk1tTfO0K2RaCB6/z
HJA6dFQRXy5qSzWKheUzxKFgxg+4rHik4kvDvtQuzvtQsAfuNd4CYQDKaxFf/UA6
yZ3e53QGtELBRCeqfW7K1mx4B9Tr4hihXLE0HNh/w8uDAZ7rBg+prBFeyksNygct
vUYQHOte1p13mN7pqFw/K6tzo7B8lZ0m3bxIRnNQR1KF8ZFnF7txgm7ZeBISDcIe
a6LNE4afe8+IE9DRIyB9sEL9hm6pA6ZfnbHzpmS6itfxkQo+DqBZVy+aPj5L0mFr
AFXAAZSNYzYHBC6JdVrQbyvxtf8e7mpwS1cDV/uDg7p8l2qzila9euHrRwmXSCzk
VdxJhTzrpUwlbNUl9JtnfrTFgS7ZU84RnoHah91YeI67Bb3Di3vTwi368NJySqku
pu5FxQXem3oEHD+IXPVfskfLqQpzobROGELImz6UhHILo8mh7SPRVLRYIcyHN+fa
TmHp6C11u0Jf7S3KEd6tRO03zF59nDHc1QWYkHpg4xWdVJYYQMcHfPt2J1ptTXfE
SqaXLpPTOGqzwKegTb9dzesI/p7I8aZrWLMg8o5TomAxdEoUVnRwhlrPhqLnAjSO
d4DhBS3viRQyUMKYk8t2Z4NmU38wAeL5mmYVM1vLv9kpvyMyNmPNm5pp07bDYBEC
2uXv47FYIMWmQkQ2MDTovNzq5bxDn0A4m1DPM5JHBoDboCTU5Z1826wEWRG/Wxlo
Ym68+x0FBV5xgeMrY+plxADX4hLPaIcVDaGVlXkhWC2K+1n1qown+H1YZhjqAeXw
gKneX3pzogHnRIxgaGVrkhRBx2Bj0l+yfHn5fsW2QiJ9P7oUuQ1yGWdPBdKZOnq1
alzMjdSLyiCDfehjo8PhVKR6cQ6UBbYDnQXQSi8/VIDZVwrmkHJwxRA4B1vjpcXQ
SZLGRBCRZ1Cz9OogLkKOGtdU+LajGe+e36XCuZtaT+zqTG3TqpDevj3Oacm6QpER
k8CGF8rrTtPorcCHY93Y7JKCa9wjd9WiheIJ2PHZeibDJ3sLtcMozqzbfjFVf4m6
K2Uy3IonEI2PizET5AvTjCtMKF3AfJo3lOkTcCBLdGq0HTRNkWkjt+kIxt/NyIwf
/vlRQaua0c54v1eW6Okffkt7vSwBwpeGga/Cw/jSyu5OtFE2KXrvowa90HGp3q/Y
Ee1652nFWeMl8DPUj3q0f7SK51bdp38yYD2bHRv88mRx3GetRVeCAmm9wP6slIeL
82l6WaRhCyiL88dvj3XqsCgE83+VDCt7KQQcRbO5uExwB+Tt9ANz3fNvhrU7Kezs
K4tIQE4+0Y1upbl6dpNkSjoYXp4Ex4CKTGsnJW5UjlN+MjWq4HibkRs44xzmJhAr
aoI6YxlbF9WyddHZGvkiH28LrvJGiNpSyjv5rKUyeDkf7s5C2hWLQMkUvciDQIK8
jXhMyOaUb6hVwb8ycuAj/9APui3sVa8BB/ZsOnC6vexsQtotDzk9no2gCPxXV33R
ZItYGpHbbfJ9fueiDQNMFk9D6uDCGdvWBFfQ/cqEkIqRbWRaycVuY2452oNxDwmP
+Ed/pC/cR/U3gZQghx9pQI07mpKxlMiV7UBSgF5eeEjnJHsMufBtMcjR+4gLNTny
jkJuLSfe3lRBx0YfIH7H6F2LnxoArGSZcGimRcJx9daPZoZxFR/0XLrWRnoNooEt
S7Viss/tOMCj6mu/nRhi59VranmBLnB6JPbDl7zGpLdP94Zi6wuQgLqHdmeh8Fsm
oB+xDNofDqFTjOR5nbgSXTlnr/gYvOsmPm3E00ASa4BVCvaoQdhNzoqHBpw45PsH
+PYbBHNORdPKTM8gyMl1CMogwmDjlCgFT0oBNyxLPcJtpchh0a6BZeA7BbtplTa2
zILMpyqYqoRVIsqxWcJR4Z/XJzI1Tt3DJnKnagH9i9xPa95YrfMueDREjaryt51g
hUpN7DeAO1W/c3F5O9J11fLRW5b5bFjdtKRcDCwUw73SbT538K/hFZa3jCBw6L8x
ioq+maj/BwO8WIjnKD2cMrSzGy0S8NB8/0vLWMqFvG9Blzi8CBHjJvGAKnY988GN
NiIi0Ga5QRZXZU7KYiRKmRrDS6U64OrWTYg+4xiTpXcEM3UnVf99MNlqBRpmZTj8
nGfFUWmgJXjfs9iegScvC4/Ze3ZIkiMyMDPflzMxykiCbyfa8MOk9noSdH9mLutH
cDYY6C3llM9TnL23+fKBBiWf7WRAAPzbDWOrkA9hbi+fa9RhXKGUTidosFV/Etvi
SNOHB/JfQz7IXern1cheDeMjVtjzT7YgGUjRRm/qGfrcNddw0Q8Wu2e0rYZ/da4O
qR09TZVf+Fl6JrpF/CVP3pLMHXQ8+8qv5GKDdxd5boXQku0MbQPDb8IINMHo7Yjb
GAPRL6ldlpMNrz+FCutEkAdxQd32gKJe7gM6aFGhDwEBMHuJkFRS6YpFaymvQo3h
M73TIwz9Rl5L4oJQcKiKLmvS7IiTcHD/PU4/zv+buyeHQxayNJegpsLllabUemcR
LTo0arHOinm50sjW+1YEcTYaSiz8S0Qx2FgXnGPwGmbqr21gIwo/G/Z6JOCxkJb2
OvW2C3lhrz7zWyy9SAR/eR1JBAKqnAdI7mDlrFgf1Evb+jXXF9Kcy61n/4gKHpH6
XBCgCQdwGPm7FxkLETvpAh3eda7c9/82w3fwwmVSoEaF9WVrVhuzH/+oAMOQcAgT
q5twyL6c7dluNdkxF7u+mcXNIWhEZUmnOFufOfTwDaH1oSsNv9HQEEOf+zb8OuSz
VKY3SGhuzTmoqkULP4cbllqY8jqhTbZW5Lc7Nqb6eZrz7f3NRKlmwpKIxcUvChZ6
AAc+0tzzbkdHR8amuyM8XtQzBCLFPPv0jtW+rgGqiFZBt8eTDwMNZSFNhAXGQSCb
exsJGLRVIIVQmndm8XMIy2t5jw9/Z/+y9mX9cY9CsFPAR5lt+tc5GLF7/iu8Vdvs
P/+8F89Q6eL2HOrymRvXJX490ivDiwJUj69hYe4JpljEYLJh2vC5dWr3jjWPvG1Q
IFtwxRV88z3lXRf1242JX+Ijmc76DlxOrGgnO7hWhrFjBqR6Hye7OBNL2irjimiO
au9YTXa7RR3gSf1Mqei/E7nLRnhEtrLCNthGa1vZI7YCeQACyJCOAwfb4jeTMgVA
ggQ1KBjbwgo+OE5HZ6bgP0A5KopBMv7pOZaYfW1k1vkuw3Um9hkE4S3cxxWi/iRq
xqHVdiOHlG2jvaDHVVggUPQPSmQ/q/xch2VGKWeeZiRXbhAmxihQydl+ZEBEUsCG
cmPfbQ7pCOsIULlkLcfPEc+mr6W/Y526TTdou9mvsrC7wzsD8kDKQjjbH+Qp0DHC
0n8LRmhkCeH8l0NGbIoMNWlxt1wICIaOSN7jy8UoqLuLlvoOFPi1qQB91bF4VjdW
wh15oYyYyWUnL/1KWl8427Sc92D0EvzkGjDpnfQhSUp/q3FZLIS9jaIFQ5cipCgD
leVXUqngBmKUiypwr+UUszsSDvx8/43JWpieQCcd7vlkwZTfWsAmtnhP4q1lL2GE
jGN9vBThMKkIuN16M4MOfnBxRiOMaHp0mgZlWpBoF7qhjVITvFVVKEUU4bLGaU7S
V16uK6WEnnfHGr+xO3aZbk4mmhtjK7R0wAMl3JbaYyFWA5dMBTKruJrsGzoFNeO0
eEhl1cqZ9vmUH8BcgxweydoHkd82e1IbQrcr7Tpl9SChwTtV3mE8tOIcODNRUWCP
EAk6J8Sc+ZqQ3eqcF+wA5MLFoJfkci11G+pt1naQPyRhRfhVTkTHz0yL2wPup9D0
FzWFYffJm8OamUu0RKulnP0TTE6pM2VvesIcC6NDhkbNTZ/8sS+9cXFTI1ZFRldb
gsXm92Yk13kij+cnD0vdeELdokwprfpF71aq5EZuOubzeSDdziwd6/LuqeCIlWqT
r2F9DAmF4lUvrRENiFwqrfAMuJsTwfmgboSKMOCqRkkMK5mAvg0XAtr/vc/24Ggu
1oMmcnllUtHNBJAUpvHvIku7ijf4yH43xAT6jy7GCy+yCldbAhMXKDV7OIzOsu5/
Z9KFb4zvRNdSE0xFih5C6hbhJH1PD0RpmGLVSywBl21TDqZKG95/M1oXE2yc1VnY
8zhp1OXpg+e99sDWoEjRSgR5veeQPM1MJSJ7fFO3otydfrFl2IeeyKtRJESrflCj
wTz1Bfponli7+zuJvEOc5yxrbJn60Rz4ZFNP9n/E7NO+ARUEREW6KPbA4Pj2U+rV
tQ/4CI7urX5n6LJgmRz/xumq7+0IBsruwDCDJBpd82/fVBxrMwhwS17wmHaymO6/
mMmYXYq8w0gXApkRL+2PNpVPPDrbcxxRxKS7V6ltW1ZJb6BC5BYl3FjWVAXeQ4rN
hWdOPUIoOyZ8g9hGAHctLT1zmiEl4h4wIQmKY9jqzkKf53VRrUYbHTQm7rzXBEve
TBaGy6J1PikfhROur+i9Z/P0EOy4XM9Dq9jXGvM61RJyZdHs8KjOA1VhpmhE9JhD
KWgUTp6+znrsSj4bxPqjZGsBDKqnpTPZ0HbNHaEw1xTd1TKFhSJUysk26cmmhJtg
U7YdXk51FOQdVKpAUvinE0AUMOfDffgskfX8icoqOXXkmz/m4gOkJlgJjRobpP14
czvK7MxVI4kdboGONQujxJtKSNZ+C8vCAeGY4HQJgWugzm1rH9fhz6H04PFD9EWP
mAbRZgAEkr0PtV3OxTcL+2eMPuKk5i96CnilPxdGVjZTadNtQXHGQ997ruS/N9f1
46hr0Z8ZViVLgzOKd87DWX0AI1PN2BuIf/KHHYGi5e3n5DAnn2k+8qY0A4vupPQh
AY49CV/a0Ork5H8Mdm7dNRUEfXjX0rnJ4tvCzUSx+M5M+hjWKLcOQx0dASz6dQvc
TPcZr17LC/SaZgGoxRMvuXkZN9jop17jLhTPWm2im0Yf2jZd25pW351OKDrGXMVa
OW853GQuq3OQpXdvcrcwmO3PuXlCMCCSS+ecp99wfSIz4M99aIBxCyIvPYR0rFwc
SIphnXqMEhlxKbwLsxSkjkfBfzF1naAA3OxRPlViuCYM8EjRWVgdTCueV5adC/iC
6G31qEfGhuGLgtY/B0b4RqG4yEHiq2Q9XUctbQ882NNe8ZllnnrR97R0OY6SMXgj
87zEDIgFJubHdOOpsZsteZCpFWYTTiSw82DO3If7T1wg1Q316xXxREREHN4OsFEp
lp6l60HVNMabFoFwnH+Iehooy7orWktNzZHuP83strUdJmdtcpoNkFUp7MVHVYyx
settnBmb7zPUCsnK+IkxCwGCJlWoR/UPxnaJKBhfUBi2TJHYsV5gfQTn3zOVHINl
Oj0+TpA/9hgmCf/6RAf3zxNHJrUrxaAMnChXgo+9OLFgEWbZVi0vw2qlI8UUu1JN
Ppv1Nyhsnt51WMRv/HRfCHznn7671GpH3kQ2POJJSyRHPy6tIo70jCdVu0aQpBVG
eZfLQj3jIClR+8sdTTaMYOh1juwecsOdaFaDBR8pIaER5f6tVgpi+rzzkEh/4RGu
h1+d3ixesoyt+1BFhXGxrAvTVZds2AaDbRyNN67Z3Sblt3q2Jq1Zq+DE5XaTvMIA
MwP6rxoUj7rV2OUURgy2vhGzTfl3ONTlvTFm/U1l/AlBQM/Ir0s1K6dYN7FmHGX2
RZ4yI1JnhSh5fbinJBJCGu7f6XvilRncS97pFs60+nu3SOVSxTUkr0ETLJ8osp6O
Rb6Hs9yRtp5PFKp5fVLgSyEOMGBSv5bTTKFdQ/0R++FX9/w2X10m46FaqsDZihdR
DcuYfeN5BOyauZPU1tEv3pK7hT9GsagauAlasrZZOIwSXf8qRFdS0OeyhpwNRFkB
2lCgFaI6tP/ghpbSNKHK4rPE3StwaSgCscDJTrUwpRecoqBHck4FDSQ52eKGC+w9
ag6LMmn12U2M+VyfLtL9XYoalZlDjaEZudaA/gPSVuktt0YLPVqt/GVXEnd8m0cm
WhN7wtyhYcPtV8vwODk53tobR4r/Z6OCPo7kVSLRxW/92zYG/mVWLpCANCuVh6Rn
Nw1ygCRuwYjm9qubaONEcDPbWLLq4ZLUrFkvo2CcjZSqQsR7j8f1u7iV9s4Ao3/z
zl7IqxpPNNrjjvr8aBIPeNBpD40uKLwR02ONgyZj83Ka97LgeC3DZ6EPIkGowJf9
+im0c48aK+A8sDk3rBAlJYoLvxoUEdbY7rmTQclHaqTl2Aemg17qpdCQ/4DQw+1/
xlO245I0jmdFjoBzKJe7hJApiyKXQSEfZuQETABfex9FDx5raBwAohjtnVcOvdGc
biwRhl6pb88bq8m31jTXDUzNDL1g70tFTm9/XpCMBfis3nbNOOoeFkh7+yiz11hP
pPGMfnJ8cKNhTnsB2dU27OkRMBZaxRDSbuwnmQko+Wi+kuu+RmTiLzcgc2hDnthx
xTfiaoGcvhIPJTejqIvW2o0MHqp/yksW8Um4aGTwSIu5RZ01sZnvbevzFRfFsq0J
MPkEsbq5rXdzZicYifyHYJe8K3rTx1Vu9rMyU6qS5T0E2/yG72xg6BDuSlRnjI1p
eC57qJ9RML92K13KhpZk2Hvz2b+D2UA5VzV2iPEGqPyrCAab1md2nY91EnSfjK7O
A7CiOdikrGear+Q4Q6+UHlTybWxtgpIwiaSd61wwF1tcRUHIO1wQaP11+b73xwik
iZK1qfNA7VV9NTK5phGlgzXh/99lWguStFnE52esSdBT7btuW+siHhhZeE7xRnJO
5GSjFKG+y98ImdajSb1r5jtdpA6ffyLbva/cSVmBmjmTcNiogam2hn2jZb2MVgl4
r+RJdYHzQKvRbIoYyxMQXArQYDu8LLog4SCMumMrtYYOtCKagHIrvdJ2Z4ddtI1O
iWwPYnihSzJOSmi44HTmPpOcvJ1LKW7Cpx+xdY5Kc4tdiDn37M8qZI78xnXin7yO
+OBYhjpeherA8wq2bLIXisRu2s3Klz0zF43GowM6yaYR542HHSqzG70uyUoAS/si
ZFH+zSBTTF331+KIXjRPtZOGRxVxhDZoWMkMbAGrR517OfIjY4RlTxvgNqRXFeVJ
wsI+z/8ihctSmnwP4uWWcMRLQcSSmVJSqNvqEHzF8T7T+TfzNicgndAbf8kSdPcn
7eSN3i5yOHYe2PqpdyGTg9HqkGg45DF9rFRq90WdEUSPtK2lKQ0t/hKX5cWZ3mIX
ytaKuNvW9LQI0lrYSmLJp4FmeS/che3DVYlp9DfIWQcolMv6zeRBnPgsuBhnDSio
b85iC+QZ6LYX/RdMoz8mzsVtG5gO7BclNt+vEvDyj8BnvZhr43wbUYhOCMgWqaAQ
0XGMAsZy7RChZ2PXl9G6DEtm6eahxJVcW2clDNq8y0R4/QZcppjywmWNAZSH+6hX
tHI86hNohFcZRmfFin8vUsw24h+nY2YEu7ehqpiF0WjkAi2nxbvHEK/EbfVINoY9
svobUxVqC4aZtkjhmzgUCqpGE4WgzuiLLnzGIPshdKY4L3Pq0FXNHfvi9Cyb7yIs
oM289kG2YFDzGord5mWw2hXuSTvIGj/CWxiLhZbUp2X2qg+xack5mjyQrsx4tJJU
XsBBmbtOaJdsC9izw8BPtsjOomxKIjXk87oeGDYR9zZl2+SDlf1wJEvdWimsdCxc
1issg0HoHRYHVYeDrCmTUKsv0ibGdYLqcykS4Rz9yZdgkQwVESW2QNIJo8Y+Z56l
sOlsS1NNsALJvv9J1WoIQZCOWybjtJLpIsuRpED0MxoKlZDffdWuxgdJwJ1fswrC
w4N+z4AeHxOIt86XI/u7QU3IUXhkgFS6QwIfYAD6g6N8TAS/Rxt2VV2r6aEFeEyo
CuFcHuYD/FlH0BKJtZTFiT8+3rH9XMA+yKdV7pDKaGkoSVeze69c6kIdE13ZkuZ1
FYOVsu8kpVa1asw0grhhVeZ8JZp7WSQVFgc2wLK1uAOosB/DczRQWTCi8/QO6u2+
F47Lm907ojlnhpa1v2ZD38bmVthORuQpkqA3DGH7DbASOIZBu8zp1I15ofNrPd3b
WUE3gHnyy5PUzoxMDWYVau/diOs2HKyedccFlmG4/mbuGIF9Y2rhowt2i3wKKjGG
8coI7Zy+Oc8b/AJZIAmLE2A0ZBX2i6N6ylD2vJHFrpUnr97/v4K7jfcLvrV4NNiD
e08lchMm+LAo0Y4XOz3P9eRXAMvdL4VGEr2xv9UZiZ6jGvlmwdP5NhZNb3BMYqMb
4M8jEncPF6t510RcoPHMVH7vLWDXnQarWROn0wML0JtLOmPwsK1m7OpYA2z5s3w+
oL2z62mMyvWIAb79sndWK3QnAQqIJsPyYeelPhMfOAPvemusKP6C1y7v+ETC925Z
ytkVehXRzAf8i1xK6cmLNlo4z1L6bKujkhq/FbV+55gHPkR4HEsO80bo3+NWv3AI
MYa7FWsGUiS8P8l9dO8ViKUlQLZQ1WVhkYXrzcURET7sruIytzx9fU+bnyEEissy
SaTCSEVktq3v6CUtowkFMwZOVY2CAbtKb9ErWlQh1eSV8dXKdGfmD2bXb6g5hysG
RuClpBPDtx0hEJ7Wu8Q2M9QGOg/pDmFPzzeZ/xaDgtQnh79VxN45S/JpvUXY/JxK
4StclAzCFZ26vLSSxhPSqJKxoGICmeMUxoIT1M5tCCsUDMoMNX8j0BAW19wy3dI9
RfuZUALcs5jjNneflmMraTtHB2jom1Fg9n1fSX39lzKm+p6vtKsRsGpYyK2KaJHa
KPmz8PLcEAmPEipGAHhVO4aaMLdQJO7brRZzpns7ciusPLdIiQ2SirG0jfL1sOUS
ro20mtPYpv7ZcUXc7XlbL0McHD6+2aKtH8kKHgy+64kgNb7QvTkMyF1Fi9SLx5Ys
ZN/n17p+qTEIpGofSLp2ptGQiOJCJfRDmCME7m9K/EXtFnifo2LaMD2s3j7AaVXf
WAH9Uko1BXnPvHb4jLA7L5cl3RF+Sl1v4W+u/NYgxoXQ+vR3XkKfHt7XFSbAHK9q
BxSM9QJ2pNg1J783P8rPeh5m1KJuubX7SAmujgzBpR/z2PPI+fuNVxym3kTRsGei
3UcFhsLNfc9cw6v1/Mw1hk6FA0Po22kADK+YJOUYKr0FPUuqHw7uf3mNIh5T6u23
Hj5qUzEfCgktSH8iem4CpxsRM0vAGmyc4rBqARs3KbKgn8wmfy1AIB4LX7yeBlHE
z1wWI2I1c/fQgpJyhEfi8HIF9YuOf1bKRg4FOYjbFh/4pq4Kd3STARZxzRBRaBhJ
VEYD3ciJbTRTfZw3rs2G/3sisptBCWuMGHLNZrbPgpiEXyR6qcMxzu+pTdgdtyMT
anDxcufolXzZLOsybQ7SRbvg7csrnzVQLHRY/ZBeOUfLvJRwV568n5GxIeqIbJ4/
VLaTsVpNBKEzTfzLyk5umXq89drDIrUX+z3/LTk7f4XsAngk85PLP7PR/ySXTuhL
q7VNcZe+58BrU/feNtOzzkUDJsNsyWUNR4VMfqJk8PwhNpE+OCGCwj7LOvgQ/y6k
drkO6Iy60AvM8OrAq404sRGuQrpuZqBKme9EZd39HY7J4+EzKw3ZaHbiy/XRFT5b
5usizpX3Ucw2Rzex0n/qcEYH0YOFcB/CBbRwzxaWxfiF1lW5U8mzoTTTH7uyPSqr
B9BcT3m+7yoFAtas+qWTVxxCfff6+j/XppVzUKy1hTTBhJ0poVnh6GEBuhLewB1G
cuiCuWHEf4BkAxfem9PxIAhmChRqzjq9rWXxEmy7lT54obcMeH0+IxUJApGhKECB
67DAy76LCghio+JrE0RIFqsJhRKqrSmTtw97aYRtoib9JxN+pkHPUKT8Emgpf6b4
fywbJoPxpu9DUhRADQgYFrWr6Wml5M1q9+hblsg/qiVWjBhH2c93J7Gguos3M+Mx
Q8h3e2rVSRbgt1U0blzX/ore0LahIgHyC/VZbDqlUggI34vAF6JRg+4k+zH6Qih7
w/7bWepua0TP5eBcz4kih6qQ5RX744cJyhhXc4WGHXl44Qf+cCkYe5IFzUhEZRxs
XNabOf/nP7nGBUf15UPK0qsXMi2mJ1f/ArxThnOYWXS6fQ2fftXv7LHre3r5Qady
Zc1P/kHnV78lG1THEJBBXUEVmYIvJJGx7qu4ULRrgvU9to5kIJ3RSIfdMDT9VV6B
txX90fuGsGMGtbRmkr3HGElvmaLnjl1U9Vd2aWtS2AggpPiNrQBHC48Mz6mrFkV9
wCzMNmjNTMAoDpQFhGC2M3FvMe3usu1avjMlwNaCL5YXt5QYc5Bw9oruI5m9kzha
G/VknCr++XFWruPnM4v7cU1iuBdX3K9E+8q1Z43xqXwrhp0uEGjP/XLL573powEB
1ywfLXPwPagSnGM9ZeB8Qhypj0/NGD8FolWLkl/zUHEzKa8mGY2NtrWIXJKipfIg
4SiGzj3D5Sn4/aJOEyYRHIED9lKrWTn5ixFCNJURWzc6kyUrCIwgm4E4tm4W3Hy0
xBarLo5PYe8cAsnj0/o0pkF71DaU3/u6IItQ8zMfHKdM+00gOEW0QGA82+WF0CF1
kFruHBU22J18yFT81Nwh9fYmPFys2lAQ28ms4lfRdxW36Co7mElITF8Q2uW38JqT
QqCpwA3ddU7LI1+XCc4d1O0PUisjbdutiXlkG5oeJp0yc1fEZ12zlUGslDlQ8d9t
Bt9c4FjfreysMOw53a19XbEvCEAXM5p3MVkv1HuQV1XOTeGCVzqV8qG/ewlWvfNf
/yvgC7F9632O+xd0FgvOCHcEXUdZxVmJfqeAPDRLTAagMZSJvI5r17wFFDjv+nxh
ezlib4eO3o3pkLunM9JEa3DKXuHQjkmpxdp8nWmAUX6kJ+WVBqxecsZEUeNy7u5D
k9eUJD+AwM0NUcjXJfdSycGjZ4AS1/7xrmf4E+loSBsamF5TCMQmT3U7I/mXN92O
fHDUQ7/qpMZEBLNC+zUpMoqcIqZ5Iv0bja9MKjS7iiTDFOBhaSkBYERsYkkDGAAv
UFvQOzKO4Hp90RRhzjfWn40Fs9n/E5XtOlUei/CymUS4XEnme9SJcCWWjYeMWao6
/WMrVpB9XxqfVXbSM7sfnXi1lV986gKoIVivs5HHxgxkz2gtC1MlOiS4HwM1Bn7N
Kh791fCGl89XpDRMabOlyteKMcCl1H48plPmvBR/PimoxVTvZZBKpoMke4rnfzPk
IEPYmvBKxDDqlJXIqAMo2DD40TVyXYRVe8XdTP9FPuQ7aiCAMhygC/Am18hFTZoV
hgyhXsIJUtfnOJFpD9KKAMAEsdpuFaVFyZAIMpOsfj/FovuNF4HqOoqBVwviLKtA
DYe/nT/H82znqRPYZ2DfwLMpBLCiloI0WqhYVJinLlEsfQg1W8Wa+DppFLXw9UGf
4qQGTzNWAO72Yr1LUL8a2aYXXpWiM0sxWFaKe8D/8B27S88zCeC2a/MPDpiD3dmU
mbNhjmGUlmaJzw+OmVgivp7JO8L2P6eSxvDbmS+8Vt5LPdz6ve4Hzegl9EXbhh1Q
uWm6t8g0sIY4YKJert0h317NoMcuiz04fBj5cjyffcJFlSTJ8ALe9sh6tPM93kZm
hAD9lMjh71YzwuE3duHGqlV9SWZjoeb/wbblOHM700IrdHY9aLZgmimDz9e5ZHNN
YK4YApJ+QcjyPCLp9bszITzX3H2/2hrXwJnyJjpYcXq4P9wfF5sLFsDIRd0VXEk/
hS9vuazApu5X8KmqoXlBa+V4yppZ+pCJXNngH33WwKvswiEbxxgOZH01esSMFJIP
uNqdnGZWJr68t7oJIqlZPtehnnvoaAqJ3NgTQC0A12i6tsdzpp07ZIfhv2gCYKHu
8QTUcR4dN8MWWdmmYCF7cqwjsvz4BCqU99exm/Qhg0gshxNBs3OsZCNAJnZpO8XI
ie5HNZaQx5zkWjKQbOXBUggZX7xMS1dzMlLMKrgXzV+M8FqrhOtJjMtPYwNBVjfp
0dxo55hVgd4ydtK9eDOFB2e/mGLq/qjr64iwRsDph5IjY0VYG+wqZI1cAt8GDOLh
L2/yhXCQMereLSe2oYalvz8i1H8h13rLtnB/y+gIKQeoZpDfSb867x1QR8xfpW5P
jbkBotqvLxyEI7lBkjEkFKjpxDaGxXMCwwoD15JcEf9q0q8+E6BL4E+EJUc2ZLXK
5+EOsBaFrLaS4tJ2MHCwoQWTsEIHdP0QD8OPQA+QlrUmW515VbLYHBt2NoC87UQp
aY3vp/S1TtWR4HKCMOiNLQVP4JlQt76aklw/BoDZx83XEFlTgo/rSA9Hl0D0FJbW
jujx75T5NVuBMoxelSPPJIEB5Ri21zUQpv4LWisrF4OMXU37K8+KG3iHewqDnV5U
ZUao2pTOFmwayVUiXoaW2omc7kB2c5RBpJ2NBOpdNuSL2H6C2PEUWL+d+PX9AttJ
UtDtdNZgp7kfGGx6Jz5IiwtsL/+laGLTsaDBP4wBuzlqATDmP9brgTJoEE4qOGK3
NBKe9n+BSNSk5MIW26avmgb2oQw7sxBlu+vrmJRpsSk1Ex/9xQq+4AS82tq8mnvr
wCXuRDWlOQ0VBTJD+rw/O/j3Qg/3Y8ngYYcNGIP+hPQPeRLGrGg3ALNb8x40Zy36
eJoehNlPy6zF7agcn/OgLn20m7n0KACfSuRx7f4ayv91xado2u5hq3ClwWWcYYk5
rQNRwSp6LlqHpmu04WLpT4AyJNrZli4rBODZ4/bkYABW1V8cysOO++DHpdDXUCiW
7ps/8Z3JOGfi1sBOyHZeVLCx+P6qGVFOAE2a4wyWkZw+ewXRIneXWgkiNEc6vebS
yF4ueRWwpFNEzaskII/E2BbEb/bu4fMEQ+Ov8OqNmArN6pssrGAAGsU9kYtwr0uI
7dxOPfpgn1o8cwlv7k9wWmeSwOItUMfMzmcsSAauPPUvKC7RBw8TyOY2mRMer1Gy
GuOyW+0yhpIeOcYp7UXiJJRKIt5oSLoPK9yf5EWoPBTwp65GYri6hOkcH07DeOAe
u2vHdcwtJvXNeXo32Ww0o2szB29qMOPVHSyCr5j+DuH4KWFUxFA7RwyRad+R9o1s
V2twocbH36+/2YJh/Ovq1qVTP5TohUAbDA2FdxkXkAL8RSthBWRoVX6w9wPT8xca
HH3r0Y98QOE1oXmtYNeaATET6PrKoYZg9i2z9PfQS7e+qGEFjiSYreIuKCkhnuXU
Aoow2uCfHMR9VgLVoeyzYwCU2QCtj8ZLymXveqlGtUv8Fenf3FoT4cELvHE90PrX
8nmK4OOjUI4dIWVh3qlQKjh0R/iX3YiAKnX0gZGlfJz61bMBoKgAe14pIGJTiffO
jaiDMlU1VywrCbrHhYO6VqPgfI+tdNowgtuxLOIJc1ani3kg99pCIoZn/Z0Di4ZF
Lk9NrnliqYOsrgf7BumtdphPIAPTRvE6VMC76z6g8aZeJrsTa5J2WdQNgUdVqqZo
0wk1e96Ktu3sQSz4HcWHwXHy3Jfgd66eAFWWPfu25UAv6TFdchE7aWjmyUjK86Kg
nJgIQVb2ZTeKCeE4CnQxT9+GX/c9H4yXV9EaU1JpFcCaxLHUZfRgQBp34VDNT+3K
5eTWcVUxD1ASdRO8zbP1F0eg0blSFyI+d2N1hNA7RbXG6ee3Mgbjsywkl5UX2KK4
yGcAeZJkC67VOPZ3mJn/FxdVap2RQ0/inM9XS1dU9RzzIrJrCo2ezWRpPYbwex06
ENJcx7KkQmH8LBYnAYno+WBfH9al/NVESX4ryek9PZSt5vBQtEfvC9B6QVLH2RSe
InYxp2pkK6RipIzYgo/SgOIS1Xg2jro6S7wNHmTFU1IqLhHsXpLFNo0F7h2yYuwb
mAy17tk1cLEaFGK3JkO6Eec5VhiHGb/o0ClPGivJhwPaIcTgTCkUidF8YWtlh8/K
RGpKXOQQ2c20UGdLPcq7JsGCM470Hl6k+TSHvw5a5DJ6pbpynWz/hyUtUWBQlLu4
nrGldY0Af/DFNLG4lbn+q7ix+LaGrJRjdvn5l2edQO1b5R3e6xjrG+JnLY2F74im
dDStG0cSLWIrqobqE4Mw4lEmsaFHqV6DFZQYowKaTFumvZJ6t1bG/2tIDuKRniCw
qwWWbS4dvCkmwOdC9A2u93nZmRMXVQIUbadm8Z4aL/bBUJDoa3s2lOUNInjWDP6D
zHtKlMbpTNr2GZ6jIFkZ+dTb+4ACPNT8hQDfP+ji7ZCnHPvOtpTsLqR8kKK7OYch
7Sk7ouiG6HMODUesY09YMSsM9Wi5dZXQCz5logqgTQ3qPAp1QHiLSuH9zQAJvFXn
UV5+kaHrbZPHNLeSYmGFiaYRXfTxH/+UsQcCQ7H5P5olXl4s0mZL4QGv5YX1R/rY
WRLenLYGS6O9KpOaipRjVP4QqrLxNxC1h/JTJjKpydKzbb13cZE6/vL7yD4OS33m
E6IoC2P6TV+EI1CcWU02A3slg9FxqGRYQjsQyoUE3kY8R5WlAVHwhjgxHg9Y4rhM
AiR328LimJtnSPQY9zj9t9zBiPW+SwUImjwUL8yTJoT1SiJlKE4MltLGbGviS4jp
k1f8s9hqUfYk/KIMLpg4NBCBNZ15fb0tZp30t0aT8GsEWjVzyVjfFm6mX+JfTC8D
mxu2/8iaDkleN6BtblseWwmjKcoKC6izWjy/attLUAQAt4S97fLnH3W1Dkd/JoDq
OWztsiraxIHQPJkFUnJhHsBT/FIct6iEmXQnOCwS9VR2JAAIQn63i728hYZ2a636
fOeLx5x6xDwK2/6e2M0fxbsR/5EKPSFZgJHPIab3YvUvVX8NxdCcdKTNPK/ORW8N
Mk4JBRhYqbDoDdXzSH6GbvDJXr6Zaf71Q+k/TiGTghs6l3oBJt61Q4YDSk1m/dGX
vZNKUK0OhCkLO6EE1BJaYD8NIIf9MvSFwE8ex8J/R+SmKQbzuCTCkQ8lfJuzhUPi
wOmGixpJw6cjuY8QF8hg6otHMdxWClqJox8JjJNnWDaa876gmmTNBmCVInEnfeMe
TpTUumzXyFhgzosLyN9d3xndk1wIxoWMFnh+dIB9R3iHhUKXMeIt0dl3kCN93sc7
bLkloc6+3NDPsBXO/CJOOxyy6YcN4JE++qMqRrZmpISQx1LudWzfGWoCeNgKrL9l
V7llvKDWiTiEU+A7VwvAFe7aPwy7t0s2F2FULD35T6FrkCYKhkylopSxsEA3xsBd
tfEGEg7bClqUuYWXEXE6z3yFZid+kMt4rebQxBg8GpCDem+KeDw1ItMewv4MCSvp
HxnUsR4RyLBcjcIjRClil21FXkXYuvZEeogR0igFkRZnt2/6zo/Y4ZIt2lppz+x4
UqGbA1ITlv6/Q7DdAdRNgrsOxuZYm6xAaYPLruJqH2aN6whrAAh8pkewrursbj9D
pbG9vghOsJ/S8NLr/MEho+gm2lVN1KDyitSo759TaAlGwCpagQpIBiWDLRAI4V+L
FcjKxf6O91IFVGzsdGz+TwbCyLbkdXoSOh0eWSGMDzk99EOFSl6QJKPmpp6GQzFM
NMRYdIKhGtNKKl3CJzvRyzn7+N45ZuJo5J3yb5BA9olehA4Q+wweenwiUafMGASJ
rPV3cU6dg+UYRgUEf+jbqeI9+0VG7aJS2iLE5piFwdb06d/9ljXTWieWmNqO9Lgh
o5Gzr5TYapEM5bTeX1BVDBTq6kynbnsk2rXqKvliMoUTXZunYx3Mz4jX4E79Lb2R
C2G2yU+RDRDuugtFUYz2VhiSLz4nhKIuBnomperFo99CbdM3xBakOvxG9Qghx9cP
SGb04sAaS4A4wDImimkk65VOYC+2ZyWjTBhMNX9Hrl4QZUmJ1vfXX/rw5UOsJ6Xu
cbNHzwfWfGX7TTKZw69DF60CE1sJ5H1HrRFGjuZUJEEeGvNUjAQZ2/px863AWurP
AhF+lNG1dDZuQBslk0TmaCByw6Wpc6zKAHKBXCl9x3geS13gLogi85/jrFleZ8IZ
q6L+kAI0cxgmkdQbIfIkdZ1POvjFQfppT7rkrB92I8lm1SWzAFWgOwhRR9+j4OEj
ZP8H8g45uBqSIHb2MjkLnA4IywbDhekgdcfaTeziZPlxabcrqbNwi8j33+wJDq2S
sq/bX8kxJ/XrgFl5r99Sersv85dENlt7F0hL2IMnoAY1GCmXDUDgk/jtYE49+Q2U
DQ/ahXAPfXfZtZXbWA73nBMlEzF+YWWjCPbyemc+OZFRSEUYJMV7mIXLym/aLCi/
yShXC5hKiBEzH3jEPX+Igxv7K/nrXdv8dd24ZmVwSnmqi3LELkv90iGZuJ7jW8zy
MDJEhtMqEprtWoidoz9NOz0Io1UMkcBc1ghAGaKMgeeIlGXn+BSkT4rAO1+fkvNl
HLpEq422+peYCoNW0mFjbdrZyRDLiHXLl5qLNnS++8+MX0ieh5U3VWHVuqmZ61jC
BPyhaSRu7aGlSXhc09/0VuwVMzwBGH25VKtn4zNZtTe0ad1RdsV07Ey398ecVTL0
wu9ODwx9J9quOJOHvedk8qgLGyY2z63si57yamAElcf1QcCNHo4FBb38gwlgNjWb
yTwwMes5uVNwA/GQUbcOzZfxFc/RtjRYe1s5nUOS59c4/KsHOXVT8RljCIVt/0NF
LI9S1ls2VevW5dKNhd/warv/4RQ5wkq1YtdKksGoxCKKEX6JKXXKKzAjOhM8VxK6
Z+mVyFizRbEGR/zj/+pBDZXejcNTeYUXwMAzURMkWiYQB9ZfPTBsKQ7ZaBnYpOC1
F5vLWpGv8CA3BHEmmBeXdHPXvF/WtFHReP+GNgAfFvGoZ9j1oLrqfT1KBCRJArwJ
lvBhtqkpe/zyHS9Ir+lQxAcaNS2VLcpJWeiznK1azgIJ8BGYid0BBpHVeGWncyP4
VkwxIhfjHDxX/xH6Ceqg+XYUpvmp9W8sAIY5E9rnmRvVJ5TgQc5Av8Ciy22Mtx0N
Uo154eajqMlTYi4YFUigOez3g1zbbOFr+NgMGSkQP7HHSQFiJffCiG9y7CoOd/od
FbLGkI2WqKKNS0CGB76vRWM1Vh9pFcTXI6GeCGjP9Tx5mkfdNAInHtGLUu20YLC2
knpSyUpkPkAaQ1hdvRyVaflRaU60imDliVa4Yt1MJWBX8cN00r5TIM0CDR1yqk0L
8lrRyW6fTzrN/wRXbkhm7ONoeE3mSLqu4DlvOV2yeaVA32gLy3YSCqWaLWOst591
o7x+U26hVNxXfkjTD5oNwTqCH3J7LBsOk7bKMaGwi7LgaDq1lumBBRkHogwW01RL
C5OAWDNvpP6fBoxSF6KRvtfpETk1meMNHCKRuaK7WcTAc+HYvuVg7fkNLgGxFrgs
2ih0Mn+AXcYsOdV8bR16HeTIVfMHoUoYnloV1cdtTjXgBuxPU2ZhuKj+t3e9K7vJ
4HHWu9cYUSTMBpc+zLk3UFWxMgtfpDazaFS92ib8Wwli/Gkk3+VQvnAhQSl+7p+7
LNo9T0y3Gur7gds1HhN8ltwkQWGHZVn+fbMq5U3JiIVJpNcuw7vg1vPzMHBn4BLm
Pwwr38WiZXXmP3IJu0LKNEld9aL+89qzrj6bWJgYgzXZyZJc1dTqEfTk1r9vgIxN
e+fjC+4fERqeuGfvEUdhYRgO0CNvIo/SFGzezWUM4QmbgqUAmrK58+Rpr26FoU/A
lL/vfet0wmjG9LJ5qTIXUcqdv/8G4BkgU4rgbfgULjDaxj5gbQ9aa9n+XTkLq6W3
EuUVEcL928z027DeYYNJcr7v1wP9XCg7blhOcdcm73JomedvA1Wa0bdnI0EdNlRl
AIHUCCNvdIWYn1IHw6Lt/DfVe5jRVvvYZrnbZuzOefM2KKNkXiauADTXYyYpA1no
fuEsoQQYQsuChczK5ZXgMMiWdnStqtg3F4p2HlCyXTLgvWMOMSZYQzOmJeyrDTbh
k0XeVG2JgkNHZBPO8taB6KeJMCdSdhNUCIbDbDCp4bwLPJFrM94mN95FcQfVtoH2
p7Hm4zfDpafBZSSoCcvjE3CwbqDeK6cBlpk2F0K3kVPN0gDetPpj3wXC+NqGD2Tk
JKdO4HxRNHFpg7sYgZZfqguV5ZW+5rU/J0aU7/l4BAg+tl5O0cyJCCPiRNXyJtNw
5j8dU10F72faDQnTuPSTqChUvF3O3ZUdI5pSl31LO35l/3WA36tjzSWwP6KLV87T
yjIAAEAE+5P7QsDNSIhDh8yCTT/qrFumMiBjAA6daVy3CPw/fUTbvk442swfBR/5
XSF1tIEPd4y2McxSoFUf8X7rcHZhH/pjrICuIh4xocy1XhYL3U/2JueAAID2xSHS
YFavy3hm0DhBzrSz6YOJT4A0n7U4rx3yO6c1WGIaqHXEPxjSS/ej0QlljdJadiF+
zWXVAoGhG4vI9z+gMiGJhXVSoQ7H9986UAkF9IiYhicPMt/lBhdad2DUjhvNs5Fz
NnminhXuWWhING8itmBZhdPX8rzBmDInfWFh7B47DSA5F/4PkX+2Xej6yv2uk3U6
ylHXYGVYSRXfihoFi4rV/yZmgOoY0hBlPf0iujgfYo+juQAzz1PE/OuqmfBOJf/3
AEgR3ZHVAGg3i+OybTDhQbk7y5aJeLEv+HF9zv/h77Q8q609a6WNA1R6FhYzqTL3
opz3OkgbOHJEiB0UCdO7D9IXqTzjWTdKcNicPpat+QVINfktw+HGAXthEtZzvj4F
LzXeWcyktFjsabK2Pv+TrHLqsh7lIaL8AQ4FNb1R5lMPkfN1X1/lZBXx55KkbkHR
hqmRepoBawZsKb3U9VOVGuZGJ243442T7BuRwFHbgsO8ZvFo3OmBzbPwhCzbrWg8
U9eSQSCB3qpAoUGsZFNIdrFqUvGRhdvCfkWIeVRXTZbt1YBkh7S5if9rFAed6ncl
V9Q3CG4kFRBkYPfJLqjPEcOgmitekQY/fYRf0Kr10oCP7OW6mtnuvt1Z4kN2oDJL
yU7/q/AKVBPlz5n+N44PwO9wr0fjhsq5jKHwx6q/8Jjh/YXq7/wI2A0kw7bN6Ags
W1W/A/kx0DCd0Nacv9cAXDiQo3oKWhZIq+Y6mD+eXFTe38lOI8KEsSRmFt/G7aAb
JQJJ3yFeKr5yOqDDDTr3zvv08xo2QYMEcu1vXby+n1keLRG+elrdXBOINcm1ue+e
qAG9vbKLBwEVlsz9ej6xLOiyjXLwnfLt+oPxLyKAUm+T6bjJlTZya01h4CmPNNJQ
kemloF8FcOXs93O/kNJ3xABI6wFP9mfdH7AeP9+udx6/iJN6ww6i9gGcC4j/pXNq
hWlhQ2o4aOyb0YnuRMfBUxhqXxNNhv9fZnifK997T1Mnya8fMeous1xI69pwTUJA
I4RqSaAkSZngWJ7TRYXx7tcl0IvKX0afdtfb7cdkwnmPmMV5u1/oeRkoQKYiQfqx
12sXstDc384l+/Zmg3BDGmkBXOgtMTQhw1z1PiSZWhDTZ0FfsEO3HEBwFJ+in/l3
OV6TuAqUWNtf/J9/h/9A2pyRI4DXiFMuBlscLvyB/8gMTKEx/k1EqXSOnU6PKYuj
rWgKUFNxSzQ+yKE/RGfxlYTuOS0JFArv+e1Nq7QCEZ6AjyxQzUT9Q4+DhuwqCEjI
ol6o7wb5eYcoYfmxUUfIaokdTl500A2OklUWTBHJIMo00vrzxFEBeXKlKsjygebl
4ziYJ38JiTHmtbkn5vsOoB8/JznRDDsLqCWUkFHBcUTpYso73rhQUbVeOrG+/JI2
D7OGaWmd9esTgwpLOeB7C7JdM2E74329w936tmoX9SlNjf1OE9MdSbFtFG0AbAhR
lSq9T94ULktUTcdERXKJdryvwHV8FT55/OrklFk1/BU4D7v4+0ep+OOY2mNqMjst
+cZPJWLQ3KavEl3IU2Ppp8Qt3kHI6vvMt0Of09aW83TEmRNhlpu+DffDWeLrmouT
zGPSsW0ddW68aVRoKdIBII8Gs0tGPdCVxAOQSVmv4cX14G2KhlZd5gCUWyVsNuhR
0Yqp88XPjPtLruKFtFypP3uZSAey2VsyAnkMjFpBnGuEXY4tGtLziOH8mzpa8+2D
De8ndGx6iVUMuwAK5yU6ic3uYimyBDiMWaLBDGllGXTiLx2A5db++KoqAaXT05NF
wfw9ooLtfJUmDzutg5uRZ+N5gMzO1FLIchQFyfw1X6+q6fCDnaxyIb+N4XTZUmot
1XOam62b65Id20VQR+N/LnEAetCQ1L00RkG81+hTlFR7N9Z1Xhsjw36zj/vNM+wo
+Hj8ZuZeUSqVuMS0RlG9dbVSJ7qXDpZ8MU+jpHg2TNk3mf8ayJnGa7ETsamuNXIb
0KBiCGyHyD/RZN+2x58nfcNvSmHEb3z6fs0HgryPDPP3lsoPA96T9hMVArch0ZAw
IqouUfDul7HI/cLgppVCO0r7ggSBjCLgXXfmOAGb5K/GWcDqsiPbdjnOQvwqiXYd
94OGRb/awevs7qaI5J9jgGPmnD7UaqFYEJaCeoIcrZdPIj2z/E1NnttWNCljoz8a
cfZU4Frn7eB97u60gZCPl5kTdV9GMFD3WWnJVxdbgP33lknu2x0zLej+U335GszY
TRsbV6xNN3q1D/p+c/Wz09IVei+GbRRUYuN05OjjbADqPfzvbaSWEqeqOuF9utin
+dRYBWv2qyDMJpvduIGtOv2HpThYUAu3cq88/C7YRJpqg7DfTHLWrKedRxYlGzGR
FrzrRIdf2OwQsHfps/t+QL05UllSoleGR2ebq5dB2jNa7/mZ6um7yGN6HILGuUrQ
sir2sBpvfTaghbpLutVgn6WmNmJwQ27QZBtQHgkMX0ZJN5cw/fQen8zxnEejFpjr
RM0KIKvEORNQguKfRJEtOTff6P8fLbf56ok1sZhmduew+z71++anqjRbY91poyMk
+odPmV/UrmJU74GIAd/swcocPgX4r1yn3fgkaf1kUgIY048qp4CJwXfx4zVTjBb/
iIFcTxwTF542XeacW2HdJqcy5uku2W2l5YhxtDUd53dAhJKkfuufMw1/o0EG67Vf
R8GjJTMtvoBpG9hCXEDOvcoifVJhOZ/1UmJ9p9i/l1ckf0ZJW5DpJfj24A9W8sg4
RjzWB3f+re2YVMEIKJd457ojyvbSivw76MII5smLZvVSJx2bYzfgDS2hE68+pWhv
f7Bvq8lHjgFYJO8FSvx7+byQTUM826RibmKV+MRl7nGhdYTzDOGGvPLYzN9td1AA
qgjDhLPkmrpU/0FXHZx4ukgyCyJcWfVAhNNoKaDtVnHWupkUNRJo32sjIdOf4Yu/
ThAEPnbUh6+w0CGiQqBEPWBfrC6AWp4MQaYqKmHRZoUf7SmhjR4cWOgxgLjfJOmr
m7cIVOZbmhzITJfU+LgKe2XogQTHuiWjP0BMfBxhMWC9ywm3EZhc0RVjIQJHfmHq
TdoJW2yaYqEaryAsfW5diF/SwAnRqBVikAhFM1rJxVBiz3rGYXmpMvFJ9yDM5zmm
nWw6uKD7gF8ivYarX8tsnD2s8vCordc7TjTcToiC6CnSs4+/pdm2pwlBysfg9c90
A9XvHNElBHvoms0CEOcTECCM7mdcWDTUouHYNDR9h5W10e9S3HnJMc8T0YS6zWd7
XBDLRz1K0KqrBLjvm02CFTugw2KzwagG3WtOhHP+4zpaGV9FoYT1BKg58E0UETQR
0FjgS+DPWoEoPEv8PyHdLMi1IxjEe57ESAV2vDPXuvm276Dl7ablg9exefHZ5qqq
hL7CyXQ0LtbAHsHB5bKMPqwmFHYsGUmMY9VFWKXq2C5WLssVH/svFWNG/O3ROk/+
N9zgR1DpvHDWaqngbOddajcaHViMeWG+E/q4jhwbVdoZJKF1GL0KxOc1h7Fy9jBI
WIjgSn9Qwi2xoYJKUyjMZq9o/vuPSg1zR+A1C/5VVAb62bN4O3xfXQyiLFNG+FwA
vtvJXN5draTfnKFcWTsJTyQVXVviG0ObtOw1zS7CckS6mOkBATSowNXIj3BRuBHV
4onbNshaqo6S3pq73/466SHLH4DBDa6C5RyQAbeL24dI1ZL93/m3ZrOErw21MK02
GuzuDVdiwOIBviUtLF8t5VmGPanae19MdTQ1kCpYG7Pvg2h4u1xXkBDNP9IAU/S1
WushGQd4LDtp/Mk6hUaCMjXZEFLPU0U1+P/o0b+ff2Y5AawNg21d1LyYRP1G3VzW
oWHmXRbddG+8qepOW8zhZ4pdrSWyvpdVbubCQzTqWLTKGD3GK4HPE3CNHYnP2fzF
tZdIvUgAnakGUz0KDy492rMcZgVXBYj4gVuRrPZ9USKg72oC6ZEArIgF8blzb6WU
CxTlJ6TpPbrenNaoZ/q0KMyDsUMCQO+xkYJ74WcLZB2+z2f0iaoEti4ZrbMBmtys
hEi76rNBoJ+GdGkjMRVPAbQDCwRv14CG35nERZ2CZpm+uH+uWegt3I05VvdljCnr
0IqqOECCVMbOCYh2fQ2Te4vApaWDXb6PssrjOSSoUR1EVZqkG6Doav6Mg4bNn0rw
JVKZY/W/LB5lZL6AV2D+2u3pdP+QnMqTx/DIzxsCcdiib558siTSIVDxZBH8/8bl
HOStVAodoTCl+9uKT/UhGCk+h2DCYjd0sIE8zPTjdKN/iflBmvvjz3LFvOeP7hLp
d5ulZXFrndDyt1b3Qb6rm6pR3gC724bOV4i6LU5jYKB9PdX9ErmqLhwsSqNcmjHE
T3z4Un0cen6SXQ3fa5cDCeU/pZGjjGtU7QWfML+g+XZSYPElpCTxv7fDcV1PzvfH
5evpE32f3/Iez4mllQENz/WjKNlNJZmyOg+BatObhchE20BkyRtuOzl0Hp8mmPqn
UvW9UkVkUX6440b/IFXPqM/JDoNK5RZPpeVrPNdYCGN4L3hacaRTJcWnRs62pXJH
Tjtg3oY1a9uIpL4fXRyYOkL64qmd+bD96cYaj5q3g1qJ3fXQVLdhxFFtQGVM8JHf
1r4wOjCWfhPjQaQyXd9rJATPb1jYqJlga/1lnTbS0u5p0+RYm11f1mt3V8tQIAuh
TDg+HDC3o7DNlyTe4hDlV2RzbQm2QbI2+/MvBw+3/Wi9kxOnHc0a2dvNAkilpd3a
Aj31o4HzBKiiGOgFxh7t2iSyd/AcoKfSz1fTfIK4lnZvJUTVX5cPRTytyD9Ld9uV
75IyRf8D+EVqXPJ5MVgLJnx5EgDhD96HzOTBhbwx2iKNQL+JsrQW1tiVEVmmX4hJ
Gw1FEUFrKrtfc79BvU3l7ceCUNSAc2byCLAhvGmxGEBCSJAdT4RelUrSbb8vG/6e
zrLmroGApfTQPZTRA7yFt8z2LlJzcJYoqChS/MlNrx1A1IqnE+NWh//EJhUbYcWy
fq2DsETYLgwdciWCeH+n2w6+8nSP992eWYZzicBWvQnkcu2oS2GbLP75AvaCT5hb
v7IhtzlWvAcoI2CJ5mUo3NI7Y+wX0Lje11J283fdjpT3JrwzRccEyG1YNhYyVAuu
hX2M5keYPm3fre0dJhgv5p4WDwHfMX4KH52LEzc/Di9l3NLAXwcUYeB+b4PIUIjT
kUQgXqRxzuadxkWwaTheA44sksxUDoX4HOvmCxZuG5dOTlPT306vwJXzckvzmH7n
3vv5nmBbvEOfiQcGBmYzvL/lRoo14gGwfNN6uaVR/wVmc/lPZnBWppEOWNBZe1zU
Z6MgT73f1ilADwzqcse5w3ICkNbzJTZS8gvoEIC5Qz7WuThHj+EpqgZoSr6mv+/K
lw7y/tFy3uucouXv8a2FdVC2LnVLZrhKT8xFD0wMrHRoUVn8mH2+CGWyXp1Irtyu
xy4B6rzZSnPYoJ3VIiuixD9HjjRsJDsQL5HrSgffl7N+M/u+0xZy/4ahtaH3VbsZ
VNoN0tbQlHhbpVRwVNtfS0O1ycTQbQZYsQkMT7nIuojvPYQc/LI8Iw4lHE/LUVXX
A4NbJYXgSmyp6BzEsLEDSdOlDG84zjCnKBElkd/pI0b0cex2X59QfLiTii7W7p8d
SUyLxSJ5Frc6ksqs0az9f4pKltpelw23ZbCkE9X4A9WuBfAvdWwpFArjeaL7IYIO
R8QiLEEJTiyvRed4o873qcK/Trv5iKjCwbBONtAGq6CKiSvllyhB9/xy/dcek6Iq
5h8Pht9XR6FkkGJf+DSMRBh4r68UN6nbD8Crwe3mFHCEU+wNA4DtfEcTDwjdb+If
XD4j/vty7qkq7XzrPSBCiFpKiDxXIuT+u6nJzzCGB/jt0EgHrOlcTPkKhmgf9k5K
2PRADGH/O6+KqJ8oPO9enX9VIGHPQDnORu0WrPD+R8jPyH+iNLLs1eEZCaVU5uOc
5sqK6db5Wy/tBUA8FHl1fKqrTXs0iiPQ1BNVshSbcc1Mm6c9dOi03QJrCizFkTsN
RU5nK+KTDsFKsSHJrn3oXxAuSSCODETPFkMWGnv4+575vq8xyURWvN9yG18hDglF
b9MJc6maMfeRpjEUgU+OI6qvD7x3eyUB3mE5gRDLIAUsAn7b3Dd0DTLKRuE+/gwg
QQ8BY0Qb85wk1e8gu7dX44s8igx0lJjoDwzwPmj2Yv/hJXWtA/ZdRFP8wXvjIpOU
zwvu+7gvY1nkTyWRZ5GwTgha+jSdKrrkpsSbCwvYDfHCVF00QPoAyJ/mq3IlV+d7
E+FhuG84N8VUlV0JO8t5LuSl+K2jsovMX6uoxKg0YKYczusKWLKUhMrE7G01+btr
sMCCmJmsGNUm2HMlB1X1HmaRzNbPO45D9kezqd9vlk4G2is9mFz+aanIICa94n+l
ldhVjFCUxjRk7J6+8VzoI1sAVkhUtbNENLt1qifr1LUF5MWFGVkWGEspYO4RqB6P
ephDwFagSShbSQaFDfTsMxG6kJxMtQyBalOuwA+Fv5E/8i/Iq/fdDwyTkWL1DLAW
pl9NJJV6V9nbvvRzewhFmqQAJSUqHKWgEsZccVg47h9mdMZteBBxobG3ZANdgYVS
q2/iqq0L1R+0mjjb0HE/VCYqvJZxoahC76IhV/W4xTYbYwsO7JQzm9rjpmTi/1Ur
itOIGs4syJDw/fd+EXsV5mgaGDUOqKMhdIYAYQOVmv5B349hEFEcjq0YxAFLvXoT
qFfHLTuN9aQOKE3av9JHH+Jyzjy8+w5PcQb8YJ8t1WdzKwkTm1iKKleFVRAUJipb
llDl/CegWZvbBNITiahY34mmC3zefWtfSDFSYwlx1CRM91upi7vU9sv0HSSpgx1e
rGyFiIa5coJm14/y3cMVl2Z1yoTkOut3Ss1xQ4m9qMVNarQsbvYb49nZXOM25Ndu
+D/3zFK9DFfKgHw+8bNSP5+Cp6xCZErHutl/404cF652aZMvDEzAkx8KXuO2wsQP
Al1yG26Ju1uEaq6eMl6HOD3613whu7Skc8N8h0JfbW55fsQ9SpYj12qiolUhqB66
wAL4Hm5ihskoKeTCBkKCnJ5i5hNyPhGkM4Wvq1o/TbD54hE4CsGCweh3CPd09LR4
5RmxZOBDe2ukLO9WnJ+PzqSZeIJ4KLfrompJ24t/EiqFJ//+Ynx32GqYYD1SlqHh
TivySgLPugBCe0JM64/FHiweXWRJrW9U8hyYw4teZMN9gRw1Fu+xLwjQy99S62oG
yBU/hhESpFfZFKBXW4ep/ZeGvYNybEkgC7aK1FqOz+YKeRAQPuWMQsapfwZtWrgU
Kl9gf2CArVxjs/zDQ6QOwLjz39mAFRiKzS6AAvyJaaLR7sLmXpqb84DoWGfrHPM4
IFk8W7fCNXE4euXH48i293jPKzgZKjpxvL2VDsVayUqwn9G0o8f+640E9nGnvnQ+
SVK/zK9kChsrgSlqo28yzTGUEnyzoZolWQgdfNqk+qFcz+3eglp50uUjGNxOdhYt
MjjAvNTVPnk/RJGPIcrVzqW7ZA7egMzBeYsSw1fhbW/O45Z2c4y1HR2hoWYv6Acf
tesvciVzhZ7+daOgX0wrQHZ6EYG+70d9s0j6KW0ROgVU0KGvmco4jJGQlnJnXMnN
cG374U7OMD7bei+R5M3m9/Kq7k8iF+bOsnFWsUaWVIzWrvGCpxEe9Nz7d0z87vk7
prwwo3TQoYg0pF3b0zDGVgyYeqNz6QuDyO1ztomBdk5N6sF4jpcthccGNVpAGVB8
vj8mDu4wC8NW+8bYfzCypdrX+4JIf1MfpEhR6a9DyYTyoXBI84KsCyBVl/KGrxmk
c/OznqbGja33j3F8BwP0+RtmqolS9lwy0T8MZMWLW7ZZx7XEH9tsLXdZWyO2pgP4
NEP53qDxGOWEI88VfJNxbYKS4CN8GBPzS+olOYykwhoDSoV0ppc2bjHzxC/rwdJE
NmfS44sUTM3oU/A8NlGPzfOpH/o+y3WaFYFc5CJ9jXPFZzgUlt3b6n9NW+9dFVrR
6oi/doUO5DdzoxYoDtJlF8SmcVV+MxTFzeDt/7XYCLE3M38GBVcYL1Cc/VVggSGU
fSbiESusJ4O6UM5rnpjnoTNp793gmlh51lL1xzmS/0okKO/5Mjr2++3hFCKUI5r9
YabYGjoFhW9THcGcVdgcQG5vHZ2vd09eUEVALGaGassddSUuvbLKZejG+5Z6DfC7
dmLtS7Fwphzcn1cGlH+XrJjYerwFkf6T26s9dJm4suz/h5FpGzizaBTVMDv2cAcG
+9+5/JCXToxLHcq8TvtSjTD43arek4TqNpb2mH11fdp/RPdMQf+I0g8PuznrPXeO
o5dPLFEijczFsETjMJDrA0Ao/TQNJbJG6kPZORJ3l4AGD3a79krnIiPxl0wheTti
QhtCYtoLjLZV9tc5VBSpd+L28OK4W6hcIcVmkQ8JSZnK6C/z1nuahtKNOVRDEnV1
7M4Rar3wR0j1mEqu1XMHQymP7ymjoBEPWsCykxYmuX5dxLjI5GdvuJNvWUZQehGc
HUJ4zL2TSHKijKl4TsDvaBi4OPF+1MldpFFjmQUiCqSMxBU3TqwKKSlotpVBDsYw
gZiVgegz94ilmmu9g4GrJPWwIp8kkixS7I7hX4kCK/GPFyavXl18R7iUbc0hC5uG
URzlMM4k2rtanZAzU8pfYbqPi7QLF/TyN66jbysWnzO3HISxCr5G+2MpLSKeVIMU
0RbrX6BaNp9N5LBeIlZzqoJaopG9gfJrgzwl8jIsLOPWXoPgmDXxI6ZZEUQhl8Wd
4RQyqPIjqf7nJ10VdmO7Knn9bAQAltPzraBWT+9xThe83Etw8XN2FeruYSsatWet
mrSoPAGdSm2CJ6f5Ecr6P4bUMZPJYOvY88FT/kz4D7guw/5OfiliYmjurCoW9eE/
wLTHXLaRTQ5xhDrOytjUjx33evlGX706Y9NH+nw2nShlUFxpOywS0w89twkDiuXn
fiH782LuD9RcVdrh/u2zRAOWyj9LzUTMOBGKqbgaOwZJNj7SI0i1DjrjfemIX4SF
fkT+ceBBoCx4sQ6PbQpIegBChP5vdmwi3Or+ZmI5Jljdr3YFRElq2HM2lEsMspSF
0a2uagYbRvVh/F+rrDBHHzGXzBm5x+oaWX5e5QDh2w8463ST+vSHXaKYYZYvK0jh
IarNLjsSFmYise7SpeLSABckWBMJQRK+MVciCm+2EwyRk7ksfR+5P6lfvOlcja+R
mHS0opAvYZySEoGT4iDjNwwCM1Hx6frdb5KgGIGPJHJVOOKzr22r08h+fH8xzHbp
XYrJ0Jt0qm6s3rPlmrv2ZlS1OjSlQN6vjtFBOsMmlssxD1pfnQcTM64rn6P9Z3LE
UJfqkpFN4sPo6ovtsNsayePx0f1GwdIdseaoTNpNlbgICID2tlb2r1MvEuEUzmOe
F1QYS7oePBlrk40FZ0mPA0Anf/DNSpeLXxQkBQovuZdu9gmr+uig99N60Es6wHwj
q5iz7NbmHSzCqoAfvntnCqCfFjrBzqWPMeW+bLHJo7zNc7mp+aN3khJZVsfowASr
mjNsY13+TONZiOBteQDmN+D6Y359TfeQpx0/sXIf4XCQg8aWJH7qmofXB29hQMwA
th+wC+Vvz3OYTMfuOQWcK8k6ChmPpD2QOx3AxoCb/ZwGbFq2Er9Rm61ncO/aGzKv
+hU7Sb66DSoZwFX9zrWQgGjTIiKBXZHPoQSf9wNlZMiyLA1gKUyO931mVO1LIcJ1
N6Q4cVcceSuC73u/An9TiW5sUMaUvA3og0ny+wATwt/5QPXda8cRc34vJPMlODpi
u0oIwSDcidh08ckuPhu8nvMDo7ghFuax9QNHcLCQPuzL2R1aQdJUxdqYfFsVjBzY
nPGAM4twFU3MOR/oORlFuBRupi8/UAwCEWoZ/og4/jnNMvA+9A6eD98Vm49dM/sO
n5/+6iw+lDklgeuDt+zcveOfyLjLt+30lgLrmVV3zYT6+bdgSM+HButDa946xmU9
GPW7KMCNcp8deMzNOexNHedYnsn3Qq+px1zf0Rshnvs2TMQpzJcOoZtv+hxxsInb
8vQ+DemDzWeXrGESaQQV3lWpjZxtsxQonaAh4UBBY/U4GgO9okd9BMQj5wOJKQTX
gL6oO0T2LeOLkYgoy98F8Ioh87UghlJpGce1kzUVaZR0axq5v53ikW4kNvhGyBfO
fkXdAplJDx3hxnfwWbIwOrvhOKScL4QDfFprp4z6PZAFnNyGtMWZOkraDOQIiJFC
6p4JLqBNh7oZeYRDA5lduT4Bi0UQ1Qa73ZB0LSKhgik+YLf1b/NjfP22pafQ8Nyp
4YQrjEYATRb13QtrworVh+90n9JJcipiT9zTUyE1YtPEj/39jEhT3bus2mGtT9Jp
/V3mc4oUzF759uMVo0sk0nN3LFtTEhq0TAH42ieic5HU0CrvP9ezF/PEwPrZXzRD
fSnKhGiHftERVOHoYnEApX8522V3HvUolgX7sbhDCJ/gWhR2ZdqCDqIkd/FQN6Ql
U1GWwa1StLu44i6ZRjqwjteAsMmgzgkZ41z4Z+4XsDEHjujdsMZCs+S3YK7f/r1R
eXqPK2URf698q6I7xmEs5AaWqwYJQWvt07k0jEfEe52afMZgEhfuyoCgoB81Lc9Z
b6Px/W9EodhdMv4wN7n6FIsh4qJ2TV2/zLsKq3MNLu38JVe7RA78mc4ZL7QtGzES
mU0rmiVM8g8udAmuH+fFDcOiIfpyIszWzFpESD1eLvF98EZez8zRe7TqLPYFxCKv
SWdMnXmeC+/+yM4fjFlVojtPjklmQI5/voTUlmwyHVtvwzeH4FgiJyqgWgHqOY6A
XiyRoOwzjVeJKn0vqcPGDzEqNMPDq7BPmCx9SR3gu5s5N98jY2rQCxsRh1Ve+ehz
doA0YNHGJFgCGzq+XMPP0Z59D9V+nIWPIwXGe0wC4X3BO05uqOc0+t+tbyEtZg+M
XfXpilLUJ6Qo8aTKkCRsE7dlYkFmSkNgYZE2ClrsgG2TBfxXr7l+zxC0BtJUkouw
s/o+LpsRzn5aOLStQWkKYrxMSClh3pxxmRAgFPNR8QR1wkII+riPjIPkty0tXVpL
iIE+uBrhYZHJDGwVujS6i6Xa24ApmRcIJ4U5vxnqO2aVGGOxNkYbbc6TP4xSKiYU
sOJ/6qM5Qw0GSk1o5SDjdbIuawaHWVOICLLX8I/F2V8XLUcZqlJVyJuv9vbNdMxk
MeIZt+HMBw9sjc10aR3oKwktd07jMrcVMXRjENc4WZL1aSNs5nhDFR6yJOuIlYIM
2rFxEwgX/SW0XEOO+AT43F+rBk6hvhiz92qHUk5nRtYmJh/Vx/f7IgCOX8UHSdGl
Zdc8s7LkIs46VjpIJecaYrdaaZoWX5xIK9iHWs+/McFS7UXsa2GvU4+N/djVDJ8T
1iqMbg04s+/BQr8QtBrLK77HuQYvdiIApnagQ99DbmNPttRmtwNUH3se2xGIouDD
Z9XsMgWf4/0bDo1xgc2fVlMKiuByE/MRMUia3fYupfyxUmUGL9wIKA24ogoOrvGk
/jSg3QhSJ768sGhxtsJb1PyuugYNlHRBweUYpfPGtJ+pFyw7A+NoS4NZWVL5LCwG
s2TzNxE09wKwwc0n3lxLh6h7g3GsXUQuxodpy33msyPhfIeT5+X6LFw0PIWmZRLG
w+WICox6SOJ/l0rlKL6gt3ACvHphko1g9iJfh0wiIaulX7a0w66zEsZCMadgrqLe
4wxSxFWqihbym42yRo1CgXrKWrXTTZNzqItTSWkM9BTKHfRkLhfJq9WcLl+AcqJC
cqoFtFQQfeCMpBkRwS/JZe6AQW9sJES047HQws5mmHhtJyKNYBArlTfqA6YpgvMN
qGNnPiPyYx+omkA1sgUSwAskyVhQ/z9nMgjaPtJnRJtHnJN1eCxwuh/OKHf8dB9W
IW+IY0pqguCFL0yCFAZSQI4tYNzCiRyW70M4SQ6CfzqMSYDs8KMDrvC+OGXNCpw9
O0KnojfQ9J+fSVLBQHOru4QXgZQ9uXqEH8kJtqODf6QCQ1qylFoVPhvOuGz6DUjF
iajwxuWrPzQ4/AJnbl3kanRme1tAsW5IBSBorHQX33f/w/DyD2uba4WYRTLh27cU
I2lNdXaYbOJP0G8xKfYHYB4mc85TgTyuV9Fp7HBL40zGXkc+Q/5MvZWHJ8cgPvDS
ld+dpg0siaKnct/lhgkrUXBcmBzToe+Wnnr4tKjNSA5XEVHf3Xsh+MPUBj5rlKWh
1EyNIvoDjrcjXWNSYJ7ruIun02kayN9tB1XJIkmpd6xW7wOeujrWswdOiz+0f9oY
YC3LAHheEvUI8v+X3ubtED5/Kf7wiqULQG55IBCoC3oXx/T3KV8PuqTxFyoANBbT
AkWexUkSC9wJNP6t3IWfxgVlx3BlUpG2D6AMBm+8rzebzM8yAszrdp0YrrD0GnnC
L0jsgM9tQZK2abfz+DQxc4072iF1/tXIaT4sH5zWZJ7Pz7ah4QzJi4qSceoxjT9B
j5lBNVkbdaoj0JdWlVdArApPlmuUMnJyfmSpxoakKnhlXJ6IMboqLjXTSV6IQ91h
NFyzBo4CFg5EBHvHmJx97ZqgRH/A/nnYS0b8hIvTOUi/HCoBDBt6tLmMeX6K3QAZ
Gtt0mZbmBZu+XOUeE4IQM5/MydkEPW2aogM5OD8taQRVELarYCyUwFjv9gWC2ceo
RA2D95HdaqZkPyP9o8b39IfOeorfOu1nYV/glB8sXm83PiuCOariPoH6Qs3Ms94T
dX9/zOhIJ7S0tWLTu18sc2Erdyt5QgMbja2dz2bHPfJL3dJSURMyIS6wSvexr66P
HttkSCFZXRKt9RHBzAy4OLCaEtu9RTyhHQGV4zZICWwkbbPqV17dbAq8qRakVWAt
wWqtrq/iZgpNwquN/L7g1WkkCaW/KqnT0UimYaDhWoIFmtWJdT0AJklYYEkUpoHC
qNQUUZnJZte6R9OlGFKf7uQQDBVBQrpinYMLq1V/SV9PonlMilupufXqV7RnnP8G
jpWNGojxqsFl/9Lh7ipNoj0Dq4cmKzq9GMkCAObpgamGm2Q4dsju0ZKFVmeUVOYa
ccq/7wD5hbTKd+dbq5NplevoGWFnk0EUtoEvOGrZQ0y+NQp7aZ/p/XR0EF+rhFwX
Ev1PmImQlEEjgJpYgILBR5gcP1Q0smfHz54KrN9s40DTB98Wn7Cm3cIpMrISOkxB
/Hu7QKPFXSUJsUadAILjsDwRhfMJXgcfaqKc31YBfa1isNjvwQQuIxUW0ccjBTmg
GKIq+V5dRIhocT9dvUC0i5XmDI9VCfy4bzHswzsdBxvz0LILpwRJa+hdgRPngCM8
7ZaeB1wYBO8Biyc5pSkbMv5GBj199aeT1Ee4Upjk1U4Q79hpPk5NvQUL8zoXd3yx
OTPxjN6iLJ6IcMvPnrrBWd79LTc0VW29QkdA0PtbeTpdVaIeR84AzrzvJ4JZnkiS
DsQUULiDltH62uIvkbJuspV19jEUgs+2ALvdhDdn7JfsZcyU/aUoP7Ibyr8AWODh
3AlGjLT3sTxjNLQv4+7mSQx1xgOublLobWd5CHbDd0ZEhIWJILw1aiyBBZmPn4DJ
GL6GrJp0vkmlXJHqyn4wvo7+r3OY/hYPwQ9cWav/gIkycf+5WTSDzn6baySIkNY+
22DHL/3tphoJdT2qavIWhK5+492kkV36T2iEL/wI1C7qqECC4s2DqCe9jjl9robR
E922e0crpMdZYziCK02vrgOLGWoAroWHL+8WK51dBeMNb/N+hFfTblpm6/psSiUm
70v/91PCSoZLUl8aKIg+xLJl/XU08KBm0dIu3c16wOa8YEVyAZV2dHaXjxkQuf8e
tdlAPOWBVyqffkARx4sd0jJjKeJtNFIDgWQMF22L9nEw5HsXlnaXGt2AtkT/YVF6
8vpi2tarhrok8qo4jXJXqs7s1+KjwzuY0F2hkrPvEFFXKNmgwoGGo/lH8R6jLFDs
UQ64GVCPq+sXxHRdewDLYr6rt6Mf79iAgAZ7u/Be0JWUQoPcFXZO/xLVJbOHEEFk
YbjXmYXNwlj8RtMheCaq+4H/H6iokyCwy+0KAH8MDRrlHAx7mHvGJUOIOqPQYGQW
R5JM1OWtwGB/Vojt/m5L7w2EZRxfvJ3nRAE5XiG5ArsoSrS39BCX6aYA0ZGPwj63
/p9wLwl9rUsgsYTT4aqdfk6GMVrMICmfpLq6TeYxid6ldKqVipIcTDL6fIr7yl+a
4m711JgZxpOdZXTuWohz3NmgL7APdUAmD/71usFlLKHPRnslFc8SfXrznrnLmma3
HfBuFyMsJ43EfKB/7i+NDcBQ+GO9/qkklTBb0ZY3Tu8A4hU8L8ec7R681+WSktHI
6JjE6Uu2EYK5s6r2AEuEgoBPH2iw6ZOGmHhcFquC8hmEqmbb43N2qQx28SLMd9PH
DGLCCAB5Vs8+ALTu/FeiReCFrWbWRLyx5JYl1E+tRWitzLZ50vEOgG+FbH4wQOR8
a8irN7I5lkQhED7k+wOxga3o51h0nYJqCR3/fn86SzZWyA+4WmOabyGWRTnQOX+V
64bwP4Ot8AQ/O6pNRbr5A0rm8VWqtY8aPewH2Qh0K0DMYfuQljS9zfnah33zf5t5
WzB0xV0qFN8Of/FkyCVO1VLkgtho5xA2stu/koslj8eYZl75exwvm+rxhUUX1KmP
qC9uTOA43nfshACIGmCDDI4w8IJI8mGBzumA9PRs92JBbPt6UgcbpGfA4Ar0GUWq
m7eY6lOQZ2WCZfrV1L561ICN7JJDBDQxmrSEHOdUiT8HOcHSTKi/EZcHmvO0jn6R
UQZvBrVBYjg9bR/VjWu2aZBy6bITp0YsoVMqFLtn5MJTiuk7rdwuSDfXfz1sStjB
QrlUGGdfSHczv/hooJlPWKC0qavQo290hkTASEzvgiIB1GZDSBm0K+LLxEdbyn4v
QXLtSBnNA6VUjs58QLMOk3hxAzFJoQnJ8J55GlntWs0QYRFMFvWCOnLEUaJVyrFp
UZbsDKHgVjaPk2iFU1K6Csc6ImC7/1q9anRzQBfuoVEzKXYYCzNvpq/Q9WIlD8Wp
jjmvNjJfhQ8CPQKSqcqPO6we4EClj3mZyjGR4+brvNzaOW6b8jYHea3ujJzliO6F
IUfPCZnk0bVY8C7PquIs0whvgmBC01o5H5ygdRR8327tj/EKkAeCCuuujLj+ZoEF
srMoUk0Q59jfooTbdMWjMX7qoERqmIUrtm2if0jvdT1yw++w/4Y4W27gJtviAHFl
Pl2MSojpK3rvPxV/9vAha8XSjxqZWhwx8gpbpBm3SDzdPEb2jSWm66ACV9ifQJdG
j0kiupti2+bVfPAgyVNyHnSxvSFSRmeideVEevB81s19Q7zMhoRlKReM2lbSko/C
sQM0EFJIZdv3VVEIzvjytdYJhjBAOkdekqTVWu2EffaQw9kUzems9EkRBLsEBIS1
5IPsFPPJraHhRYKJ/MmZeK3YicZyhLwz4j+dTauiJIAu4B+c1fOQxY7DsyOEEvq/
WKrx3YQ0f2ah8MEsyr593mmgxl6f4PoPekN9gMU9fCbjL3elZsv/NtMECdOCtDq5
at8fL32GXGdxDMNjk9lxxMiSAbAMVhA/WT5GzKwFswa0DTizUzj+Mpr2EFYxWyqu
INf9xN1JBlpfMMedTXv32sZxQOU28f86TatcbB9WhjeHWQIMQK6Z/80T+Zh/qqzO
tXU9/NgVPkU3ddqxX+l19eW7GC9xxs5VHDos5YJa6vr+7BEp2INc0Q9A3tI6dogj
CsdC3vDNCVKgl195p1twmZLiq9PeKxhn/hMptvEeaobAA/mrlgtUo3cszLNBvhYW
FlLjyE0V8bRTrK6ufCuzcjrDitab6oH0Md6XDXhxBc6Wy1rQIJnUuC8Y/07MfMDt
EwL8W/uf6sxXc1Bj9AXzD6DvIIyQJdF48qPB6mKklqm0volI4/7IimdQu7caGh96
QASjemvN5SNqCnm/0d3N7opeyykNKQsXgrZFNuzzBfWvRWx+euR1slIyXUS9tcIo
2Nnl7kLfryX0amHWJtryt8NNXwwgKYdJlu6TqU4oIfx/7L3pnfEIxUpKwJRpb/Uj
f5rKzcmCmzBDJE3Y/MDzkTcyrNYc6h1tpet5HV+EO3qr30P5LXcTF2Zn7GOIwIa+
NwlmfsGIE4ArCUdBd8p0nmEWPqVrxK0Cis4dfL6peL+JHvSd6PNxnEmFVENSnmp6
k+QNBzopq8wpwYr87xnL+yUBfx8BkaTuH+4tIcoL7xj3cKI34ptluVULCJonhyXj
7d0AGSMx/J+6VKuBkVUQduM4ZJd8uzGX5Yy8plWMTOwJ2EzG/7keKOaffYdtE28R
Xtihg+P7Mj/nxFk3JdSKQ16m5kkfQx1gc/zlWWmslE3PZxY4vlDP8fTJqak/27I1
4uQ1zD0AAH4q9Z8nIydOoChs1QqbVxcJU9pbX58XvCsDxZ3tH6fvv2avLV72sLye
BfbaxD3xuWKwgA6lvgsTL27GJubIIl/crMYyLE02IvLKyqhdQ7DoUFcHBnxi+UaM
4FDWs86IkBesQXGG9F+sAkTtOD0hgPVhsyJhMqgwiwRFEFg3DWs1REGPTJYdLZrV
Px5KbuMKoGo29mPp6jop+rmNILkt7mgEe9hAKtvZkAn+lNKvOVvKxha6ryOvxoMc
C/NkN5BqFoFb8CrkddpJjD7IujwTf2fu8uIyABP8ukuSDURpNMT9F8n99QkD03be
KouGLeSSkojAo47V+yuPTSkYP5THIs9bcdQMxP+rCXz78cKWjnjJzjYgXlKySEmr
0qybXVVldXY0PUxjAqx8BPCVQ2xCm3nbGJ3uEmz+v55qaW4v6V1Sv8HgSz3jvUHJ
DF0vkOk+QS2a5zgHNkkOZUqswcn0BPA9IVHNzEzLgkoXVhM/DzNxAmGta8lw7k73
+xODGrWyI1w3/QbV78wWbffEPdBEZRiE6PGVlsr7+vucOh4Wln8DRx4UWp4jInJA
dCxm2wguVqzD8F4lFjrfiXz2AdUo8N74H3Yu2ueflQH84+vp+7QnK3eSgPt+yqhC
1VKO2asi67x+o3QZ45cz7CH51kbp+7iHd/Yqldbqp9Krtv6h6xTCVf2G7XjRtsiJ
wFmGdM1ZzRTurc/41pSzVhGcaJ1LNy+K1UxDys3kVduhfZUmmQNFn8wAGvX2tQ/r
N8lEYtT/O5j03AXYidY2YlnbayxGLsBokAyaDa0mC147iNJcHE+zGZc1VK6q4aEZ
NZvo2o/QEygC+hzqKvDRg/40P5gCDMvqAjjE/D7/s+509e6YVz+jhSeUhA0wzTfN
Kgu8s5j5SuwsitnkrjH+F9/cNtM1y3JdxnwOfAQAcbBdMyX/IDSLfGi9dvj5oxCf
N2nneHn0M3RtuqYFm1sYoX4rwJ2yTmpxGMQNj3LlutiUJAOUh56rpI3vdgxOrFiP
kPGFzdIFNLF41GTfBWYZfHHHY3VXPJve3djWcfvB9heMR2K7NTrWi3x1wI2uJSG/
VROE4phF66CoeFqHceO45tfmf+NuyGY8niqoJoRV3YZ8vHNKS2lwjKq/sYwbBBEc
SR4c/UR34uWQukiKZDXVS1i4FMgmdlSpAUD1OxeiuJWBOlivHPaFYJc4IKUSPOC7
uqM0IRgQAUmK3nD2XgtCqDd3Q47RXFlyIqmgZOwfJRcQX2AmkieFn4BXsWMqVHro
G3+qZlcsGRXVb09gWlrIwJHcCLPJMU4Rz1+s/kU8jXaS9Dbt1gtaWHZcjG8bagan
t9PMjkQ+5AaOFD+TwZRlTlwmxdiakdqxw7IM0h4zMMNLSGrCMr1SNcTSun/AaZwk
ida+e+Vb+816Ba5ERpGwT36DWT1fjabYtqCrLQqWde5Uz/L2hNp3RW492e1T6o/+
SPoMUmIIlY/rQFhh4mkTVKuffR4BZ8E417pMXIFgDv0Z78F9ucjt/J9NtqYna0UR
p9smba0V/qv3yn9Mbtd1DkKH3aa9H+38T46C3XEyPSE0ptUulw3nFN3/FKP6Ov8b
gZ6K/IfTqhfNHfwwRhiW79eQdkmzjetYupRKrctWfucOr82sk8jaJcJFt2cStiMr
S/ItpbEUOWghEHGAJ2oezQ7KupQRNEGVq3UFG/4hQUtnWpuJTbnTTWK9mNtF8wUA
GPMU9NqdgRaqWQKf0uxSO62wLo4sRP/sABwyryZZYpbDZ6+N0yRaNFcCmS8SXX/C
KMz24zJreIWiq/DLqVIfon/FdqyEpD08ontaFhhUaDk9xBSgcyTD2Wa6wLHMuO9s
qANUPW1ql293yMBJqSo1fbr334M8hfdz1v9J7ORRoZAIdkWXl/z7HA7m/GfMvXxb
3EQDoFpnCI6V0sv2vnT4MSN4mZWwQc8XHDx/jWVQ/ziu8RhsWE4OTYKO2TS29/Gz
1e2q/DVO2pi21bJpjvAi01aipxXCOfonAhUAsiLx4uhCBjcFSY+jr88c8yS7AQ54
sUKgbLDE8WdrWwoFch5OBvsTuUnhwAsI+69eDViVGezlTLcAl2cYtn1fBROqHZjV
8ou68fhhCvPm/M7KZgE9QgE06kyFmLRWIlec/2NlXNuAygPHAfduTs0PtOzNQJzQ
Nl3PHgZWxlPr9Wz3MC7Mgs0aOGtOTa/nvtr6ShOQsWlsaOZIMH6iOjmx6tS6Vu9u
ANJWDe3m8/AFLbr22w+DmfpKmOcWDROSZ8CCI8MjPrFL6C914a67RboaHstT7339
19HtrnlZpy/Drr9tDgw6MJ0KQjIdAQjXGmXwf9FxVNoJaLOJCGv1eCyfCddOsElT
DCIn70bS9NxHS6IUggReJb3CSkdPVw5LWX8M9aNCJUKIceIYwucd9bwYXDec16Yo
JMk7XakHzsfPIGg+chb8MnKRWgCaBwBWGqUILsfLA8o73QczObTf8/7cRArgCL+Y
ROJy+yJHjshk3lgeGBkbUXBozlr4MOgn2PgkJ4ChAdrkzN71fU5NQ4Z4SJK5GR9/
Trwk5f/6JQz3DpMOBFfnxT1T808ZUMtj8FZzGPvsSFX9z0yckdku2ht0QQ7aeL9J
0BTpy7SSrNlBuuV220KmyltA4fIHJOYB91H7dIsq+fnlbnz7U7EEtRJFfCs+VD9g
uVJ9QfUeRcyUO+Q62w6Uq+V6eFFHvOyskWA2IazIEy6V5X7Dgc9S/uBQ4icQT/NJ
4oMd5t+M6aTf2o7xQvvqYgjis35tNL9fAwQDNT3+zDyWWAFPkbzsjscR/cMXoRL8
DB/BFW7RO/Xs77t54zxtGHu0OCGBYfmhBh7yhy4B84pnleVsE06O/OpX84w7ZYtk
gZMTiY0vZycoStCNIJxCwZej6aWPCuPk8oZvg6xqhUF+O8+227JrUAN/oPdv0IDN
VxzHzs6lTAba5+ZEqh5nG3kAXH+IozM2sW9acGiIpVpBQjnoKQxeh9thWovAEF0S
OMweu6sl5R/XGaUI/nbdQRFk5kF73fcukhn7xL5RLhhTaElLGitYbbyEcmneN9EX
qmDN8V1cidq24vUIyhOstC19X+N9bJ2263G5LjQ6dz2K1DyIU8Z3SZRhIIIm0dfD
ySyydvECvDykX6sjVE3yz9X6DPmq/L3mMzfw6MSLsWUMRC5xGIthUDnAaItuMI9w
+/59thSSSmLANHfQwHxI5zGGg6CvOKUUJ4McPnhyFSJ3W5dqSpDO764HZN8rq16e
3zusMr01q8l9NooIyIqyxriDFjYa0jz2m1Cd8WeuaEpukfX+S77RSnHc9NS2Tj3p
CiNvW5bYWJ3Asl/osMzZJDQFO36s+sWy7vmqhj78QzO6pOjOQs188ctmLjGbd+HN
5hpHOOj/0JTb/UcRTcQypewEm3WytspvvDmQfBZFtIg4d0ib9LQxwdqLXRdplN/U
WaBN5IyRAjzUchBRIvMsfMTKCWQiNsRpoVLzqspsr4QTkEQ4p6gW5zFYQlzQ6S3E
PwFgpcp6afa6/HqQL+e8wPNvjNM2M0skILVZJ1B5zo4zxdmihSwQKN3qnOTfiomB
AWIk9HNg/74RZ25yAybNbB3j7eaVbolqEBykMJt6TKn34Bo5Ps7etOgnWPeTnVH5
f2hZkWtjQFOZX+lfI9VtOzi1/R2LyIcJtNE3urxpQkRqzlUugtyRTRC/dUnL+ul1
bzD9NFr4DV5gazMQZFXpqyzWJk+Yg79Or3w9S9iBOf04NjfCusIk3+7/ghnW1Qw/
NjlO+AQsD/4QcKLOpvE7r7PJ4Tf91ID/ub6JLjgFWdTssd020mAvkeXNSGRrQvhv
MzOX4HTnFWCOEg6nSKzeWJe9hCdTqz5yZg2XSKIAhOOB4gXT5qFtKWVql8FprGRC
KN5g5/dSDhOABIHiF2QSwFNyw+N9TeR1QJUvbBa5/jdIYUtStqaorRo9SwO13dcG
1W06Ia20kN5304sBRmRMTIy8mk7DQ5zIhPUForXFTxeP3coXWWMORTmKGnGBIC3E
KtB2Jw7mYkhL83rVRY2n2pGez+ksAkwALeVVbB7ElgvLb5S+n9GZ0AYd+8yTnvQe
awSI0XEjgit748BHwTfY4Ju2Gvc+InbGiKN1eKoSokph95wPF87af+8t9gJ/ZurI
+kgI6YPSshs+ccq8hPl0aELhh1P8eie4wtTjNOQe8y7cLVD6Q5TTeaYMAzVjJDxs
a4B5JN/yIZckG8mLNJcMH3VCksHNuoCtmMRJA43zWR7gC9nt7qag294oivJDu/gV
kexdPDWNQf7KpshkY0tPLQzo6MCQXpkRqX0htIfPxyIg8YV7fVfdIhx/5Tkm8cp1
AFNqJBrigIdrIWCM4YNWu4g/qAGiPoPUGO1v/4rDbZMmxnegKsBqMRR+7N22vniC
4kKnxwQ6R/1snotbBIPouEsxyGpW3gDLtm/v0FKO/Rle4WM1rkoB1RDimuShe4o7
DVDeSdytxjSVm8aMqkGCUF8ZDmeLJ91wnzPrajzoP7tB1rfdOronUA9/TNFY8ulZ
wOU+WAEP8HHpWJoVSgOylIujG6mHb2D2I8vtwbcpqWRvQalQWsjVA4h/5TUE04Bl
/651n83VTZFthq0/l1O1SfW7j6WD796X8a0XIEU/b7Pk9soPsGXJI7C+et5VzZQv
Nlxuwz4Sj7/9qFTRv/gcN9G9dRssj1Wd14ywrikULOoAe8/Jy9bfE5dXamYN1z8a
MS3RM3WZtaa8mElqXFTmQp0Zfb4F+5kBaIQ5WPzLh6cBPbA5w3gWSD8U5kTicbEd
PRwaDzvEvCL4+0C5YfdCk6yPrBEWL2kK5hvClVRJ5k3mQOQQWaXB8Cq/GqMwl78m
wyngFPX746c9cxtyQ7yiR91PTTvwPoCJmkEk1roaIdsJyfJ08564AHVwxagux0Ot
JOhaVenBcxnnF/EAscNvm4W4OsnVynbuFsiRzC9xbH3owbf/04ISpfiQ2yQ3QHp+
gWwUgfbM8H2II5BT+jH2KquGf8nT9Axlh/+1Nioa3Jv6ruC5KL7y8TeCR4B73MZW
hV+jPWLqd7CmMdzIEFSJ6R2tYL+0xOYEfsYhuoevVgdE3w+0ViWbQOh/N6tlS6oz
RWW2539jI0h6AQazkNNecoorSSspzelCRjvrq01kaXKfo6vveOWeFV2TQN3Doona
eMKagOMSwFUoIjDh8YtmXbM6dG26gOhtcfkwZ5xFlky0qHZO+PcBqdxZawNoGp36
dNs5gTitVNnPjl2kWRjR6p7CKTmkc4uOqXoUk826V6OPB3T4FCAR6UXrKGnxO7fM
YjSQXxele7IdP6ZDC385Y8ornRPkiKKEDdKzjIDy+9ZgyHS2jH62jI1s3nlBSMj2
V6NyktVMUudvMjEuLw6LZ8+xif+dg2LU0lRsXbkQKU7OG7j7g2utGEcaX+GMKLwt
MLHLg0xdpW+0ojRixq35LsmMc6NTUenq+V8TpyNR2hpafRggeQX7nSt4EPsRsNL+
iDkwJCXex9kZo5922aZRAW2Zgz+sLGz0oOcSRZIvJ31lJyd+a0yr2wiJ1cjGxd5u
XBbFycNSMRhYy9uEqmuc27sIcihF/BRXBu4bcnxe6YM0Cj4Rp+pFjh0sK0AQINyh
Yhmitqms5wNQ2R0Nc44AHxPAlV5cx05wPaWQQaBrTmn1w8QT2enR1SOsC4T7uuyp
rQZJuFhd9GyyrS7oU9nyfF49eA9qJdTaDs8B6ERKRR2bIgghBankV0DDBk1sFyXO
1oaO0godPPhcPePRrcThEBTJB98gPJ8gGlNwoBgAtC1w6kKFKvNOYWQoDNQVhixr
WSGoMp74fjW/R/Wvw/OUaQu72AAsqrsFXAgk1v+I1N8lwx7c6BEmhQHjFPwGRZ10
zOGfgEq5Y5vZ1e3OwE7YMH5CvghcoOUV8ZiPXAqhq2AlCV25YMBJpOZ3kuJmYrgv
5li3kymgCUXO4mn0+f5fzodTYzsmgakt4MC1XrDALk3oJmAdSLDNDc+dXG2I/WDP
nMMqDYTdnOy7gT0N2hQiY/WsqDHRd0K7OxsVvMyXxADqSwev+fCcvuobXb6uqc+5
ykTxmeZEuJSK8K0IzEJOYdg/ixsLFiUBiqWPBWquBBjs+GTB+u6AWPDPjKHp6iQe
PqUYbyRSq2Fh/2vMm9AE0I1+mrdKM92Etg8y997mLU8FV/reNBDuZlGn2x4n3bZe
xKKBLqYsrKKGRcmN1yTmH1FmGJNvEkyuYgltN048UQ1FUNRAy3FM2qkDBhJ8MOmt
eh3j7qPFcswaP4T33HSNoL8yH4L0t/WBCcJTrTMc7Hi7HwZarjzMeqmbRk64eD/P
PcG80mG+j0JA9mW6TTOt6XG3z3Ht75gu/86bJy7scDiRBz0DDjhEJzY0JtAiEXFv
moljTpkAIW6l29KOKBJKXQfp8K3695jHVxW2I0muuDhGSqWi3Iufn/ujPlSypQjh
1opE/ozoQrUH1bqq8BU2lzkWWTUWz+lrBWX8Cf/BRIIDWI84xz/omgKeaccqTaLe
8Rq+ouavuyrYAuEmmJ2sFjcgOhbqNdE6xdlptQdaU4XzoZ40XBOAcVj7HtpTlfnR
7+At6YDhANlHWKioiy3uCeJj7ptJI4+M9islynQehpGfd7Z8Qc1Etlx2bDN9mIg9
IdtvjZtPWE0h4siZZzRJIwDncXbdsxbQoA6/dQzGb/g01Xgih/ck85jCbPPMRb3s
yJCrx//W7Rnpqi45ENCmmbZkNqgAG4RbsMkT4Dh8uabEIVy5oMe+9G/T2/d86qte
V+7yoZjgsnyIeP8Ss7sypDNzu6a0P+6wmiyGfr9xfgbQ2uQwb+/QDt5HiPUU1V4x
mKrvNIFpMLpFjbTiIgHF/bs2uMc3ffI/GBfnNaFDaOCb8TgLN4QJN9wfxOmLnHcz
q7YWTDX64ZrBURIErpFH3qH/wzbTkmKmABj390Kjfw+X+tZ298XK9hU3xF3XrZ+C
4UTEw4WR76bDN64924I5HPUf4HsP7/r40GAgkISharqQPvhrSi9HB83owyDRfkbL
PCZwkbxE2v1WCrvYsI9wEMpNc9BreyJKXtMZHyAcBm11+EcG4Bo6yq2abNgJdVwA
Ay7dVGaRS+whDIxvn94notGnUc0QPL9l7zlKUjeWN9Q7V9VqcyoWJh38tTCWGZWE
7DjaOP2TnZ/5YsnIDhlw1+ElO2l8jTVSThIM4/P1zDSs7e0upd/s8nJcPGFAgeeu
nJgN+lPAU6p4o1UvDe1ceGno9MCZbcQ0zah+4DDgjIN8Z/8h5BIRPi3pLbCL4fNa
pOFBAjqrWMifQBM6PRXwY02ZttQ8UjeKX71k8sJgGrf/zBRABdhOwPcIynPvCiRi
iHabDuxL71F9ZawE6U/BJf48OQakF/bc0LeN0L9OFCR9ghjs5Jmr/VmdnTQhWNep
N+rmMjJ0fOlQy1oOQZ1o8w3SoYjCdtgkHGWaC9rESd118ZqzdwqkFRrrj2BFSMcY
CqIShPAno6HgiHbX4qlqLax0EMm1SJfvCNNAnp9MUSpcSUcY/a+vZp1waFAZhzLy
xhMgY68FP3spWrz3SA9TjgnhMfgjp+5ZVQxFpKI9g2jfgDQijYd2erHGTUNm6Iw5
h/j6KUWT3NHRJC9RtyyBf/e1vzGGT9OS9pLtMmLFDekLoNKVYxPDpTVb3tEsD6So
YaEr9hmjU/qANkEVBT/nmk3FRw7nAeGskpuZi/jnEzEq+qyODLgZul9/FJIlFMWg
4vUZmAiRX0UD+qWAkgBJRX99+NPZXfJf+h2C2c57Ift3jqegoB6C+C01+rGjgRVy
iE1pnsEBKjO9gF2FwLB7QOV1k72XYRNLJuyqtiKyYqWB47kDxYhV8Rb49mFQhFn8
fCC8LFiALbqWdeqDPjl0EE2d+BzzI1BX8L/2Ue9vUp2/fthCnA041QZZquEzNZ6F
L2yJhbV8UwRYGGLf+WFKV4OZp4MgdgWRugWDFWwcMtQPOXtoB2arUTCGS0015WIF
fkoV8ANYKKtyu3Y/6ZsdQvZS7nVuZN8zSdyMo1pU2o54lCjXl6C3vzZIuCBAyNLa
ZlJGIUpUV0liwle5gi1LuG1LzaUlNjzb66tFJvGL6a9PVpkGRYRRPniGpQ8+xZaY
lmamkkBg8c06K4DvEuJ9YkGIXAS7/Imrr4EiNSACAmOmbTPg/DnkLzCV2g89zkDa
fKhAMBonr8HwbsI9P710IyoLXe3hQPD/Dx+w9jPbG+de+c/GkBc4A/AXKXsqJ/mK
/O0VURU6vkHzyvSlZA9EBePiUN3VxyMi6DK0Ri0AGfIqZ9O4aRljOEN4HNnMk57b
wIfydXT62n25KMimfuLfkO8Oiu7WN6GSwWbajsHTlFPFkVmyUgr1NLAGQed+ajuY
z0KlExQYlODtkCl3hf6XnmqzAFun4vUIaYe57r9q2EAQQv69LuMNPXSrv2L8przW
I3/Hlq7TECED1dcbakuxqzE5+4yQ6oOT5RkhrVSE79MQWLFro8AA9GK1vg8Kdisq
o+k9WwvlZ6ZF+/iArCObvFNjWUwoVXvJ3Xld/Pykp3U5exiH/u4s/fanVH0phZM3
vh8UKidzTJdVQz+iHue3i2tcKQLVVE9bvMIgjtsDFP6zXHJru6/b9D1X7Hz3MjSj
IhQSn9+6R3VkTo9S6t84ZA8T0Wf2pSBfIqLeP/1AZkd+MmGbGo4fxiJSm22ONneG
qMQ45dX9Y+SwUuCSg3i19J9PUC1Pa/AL43HgCOZ5gVHarMrtTr//7SGoRKY7JbQp
RxMBGPEk7MTXcaGefe6vmoKaHnPDAlFYn0CmKG1OKunmujZIoMZ5+cvI/BoAEoA1
7rbzNIhv48+qAaKtRWiq30et6MzSxUD3ROwQzEB35RenF4z3QV21FR0662uBp9uD
pGFp5Ww+ejNhRQ+xOqtIhuniOwigNfqg2/nLzM8sZnelJwng7vxPhRT+lzba4WXG
oFKFGkGgnV+hOKLivVyDXJnl0Wj9+F3paV9morhMr9fPL+UY1nUqkoBUR5I459wZ
TvdwCKJc0xFYEBJI0u1ayEkpwo7fs2wJbZo2eYQmT+gLf7ScfRoUG+awmiqfAnPI
GQ6rxu+2CzHdA5cpHKnrw0apxBBap827Cn1rWTTENLcobDTdGW9tVtNPmvZAs9Q1
XAL8vzOpBtHrS6wHA5CGiR28O5xlR9xRMExlMIo0t/N5XtSesAkVtm2n7xIuDi1d
bAguP55IuCFs45kTHZlBgpS3FMjuuouOXvSGvphxAvUlHT2kKUDBwxRMvWQH0QGs
9XvOIcyUpthxzP6S1iaAkER1E3j5MFf/jeyerZ6Z8pnIqi84263I+qziDP+DdTaX
S9CE92Cs8eIRm1DQjOyCdBQpSDqDv3Wg9TITc+vfQApUZF661hdaTK/Hzh8h1tlr
+2htOBo7vfiya5NhTWRVGG4BlDwoTqYn5TIa7gcRPXmLC6TkqgSVlHo1bRnRH2u2
yi5Hd0a/zFDU1NfXmE6xEEp9/5DE114m5SP6+/5ujXUnbYE3taAA5ythgE1PLkVc
d5Cz43DZpDgXZ+cWL+qy2cigV6FF11IbEirOjddGsUECNAy9ILy57CCDq92P5gFh
9H+RqpBR5O5i99qnFTOiMxZiqLSnBD5AHWgKBjlTucDuHnOkEOiysoLuu4ozp8MH
A0GxIcSMBTQgxwgP5ssX6TGXrMoP6pzYMXkWCKs3ckNZsBKADeOozDyd5hIKq19S
KtTrQI7UyixML57u1bvHbJhhkF3yqV9zDjqZ8yi8i4nL+ezF7NG0b5SQcqYO9VP7
kF/VxOUSftlQMm78kCTfAk6KCcRXC174l2kEKLfzHY/uPV1SvbiocmEONLpAmHrU
MT9DGj48K8zBiw76j27uQ0uGjrnYUjnWPJkDMupHhcxpVWh2/SJW+jDUF6Akgaft
xrG21+3Ab1cS5tUd02HRqfEu6OeRKTT6jclinyoJ+k6kdVLrWsb5tj9k0LU/dthf
1FX6YdhuD8UABhGzNGNhib4KLjB9vUSpIK8BvDfT4q2nDSGr1HXdwacbJ+UM8hol
PZqce+7vpsz4dgn4bFVqXRV75vk1s0Oe9g7y1NQ3BVl0igip1EhFZscRGMDMQmLG
HJozMtCcQSCFUCkRwBwBzB6dBNWTqgUsd2Nfl4X91ffOQKUsqx/IjdZd/ygMLwqH
tYkxyCSC5tdduF7wSPNvpCWxLchMw9EdXoZ1+hb/dwrDzNXKBsutgo60+F3mqmIh
F21bJ+CMj/1vIH0rZTnRF/g6sh6JcFDmntfxr6yHtWw/weKkm8cM2zgQrDiR31H+
ZqruK2jxooLIPWs/L0ZwZpIBWLvYnY6NdebUjQW51I1lgg9gnkYbOBBDF29Ex589
yg9I5wmILb0N0NYXaegPntapkfe+8S4IDJO4z7wNpuue/UuXbiJDCHIzg+ny4a5B
puqrT8dMaqiZqML1jWs1+MBxnlxEB6ts+8Gw4ik3Eyws0ttqVabhKnau7/jhE5pE
HaVHjWbDb7LTwCAVnLo/YKm5n3oVf8ZmsMwoVyKkINcij+lj/N+a/dv1CV8B7e3+
vmprgIPmAKUufwz7WtX7F60AiU6g7jj+YNLid4b1TbrbXSydwO2szKDryA0l0Ed1
4ExCVWmDyhBR7Wk8UWSBhrwmPC5FifoqRoLWMD+lQhUVs+0swJCoK3FLsG+GTWf3
vgZn5lN9mfqcad5tXQJzfs7+AEQB8AZWcdxGIcqJ/N/tU3Uxc8TuMZ6PyHGtkQPP
j6IT2+FSfyzJvBtmz+yuTjSmJ2BDZw0aH1HkMi0xDVnlg5evZpT+b5swnFRbfBeJ
S6kYRJHi4t3s/UksJMKQ2pe958c4Az0rgBkMG6ruxoHW7xnSPt6LblmS0c8Pagn1
2HYNJ0HF+/HytAaWI3ndqrmTCe1XyeTMWz2oRH3UpbtZcf5llZnvQu/j1vJ+80/y
LgZ+VwWe6sCa/nYRZ485jb2sxIfi9MLmGcUX9G7iKfikh9r2bC4lRGLOv1/7xfq9
9q4hpvaSb6leYYP8Ihaba9Dl+ZRhysxFcYVrjAVKi1oRpVhe+qbiK6kWKrOPkI/m
MZWohzAw+OYvclvydMYlTKs3QJe8NjpcZtCzqywqFDA0I1O3JL2qrFU9FUFzB18G
LvcBvrpt0twQY9VHvfqjovxQRZufy4w9cm5VHOWEKa9+hpQOQlbSbDjIWNAak2xG
EYvUTWNtyqhUwrKWWDE+LgwtxWwi+7fvtzFsvP0aIS2i+6OHQT402akEyo65ZbaS
xYbDBw9tLvARJ4Inh9SaCTGYu3Gc1HK6Pfqw18wJykAGtJlVwnMLCyy+vU1XHBTy
qoCh/9QWrJEovcNfCNTq0s0DMyEGva04bakk6aB/m7bvt5V0u73hrd2TRSXZbI1o
DT6txIsQfNQCInke/kNu8VaDoJKUd6H56Tvd+jUIC6uTQN55ePDZ1Y5kuyPqv3Xc
yz5W7lZaEaVOLfgwdT+aC8jkzWZKbPPw610kgWBqN7/XJvW3wvDAnebWESkCwopu
aChoVVLf1m6LvqHOxhXn05L8mzosIgbH6vfpd/Q+/5fHpcdYaj3J++SvHk05LpKn
arrb/3MH9Fm2Y23laE3EPHznvSieEKU7q5fIW84o4beNgbH/geaIJtpoa3pKg+ve
176zs7ic4+mrlRbtMKIu4D0MOlP206ThzIH+vWezM3MZyEyNNh5y+3NJaDSt/S9R
y36u/i0AEivcqj5uAGkuqj0PsG6sin6HdVPJ44e9xFfspq2W9I+ZvK1I2tUl5pzf
3W2jDcyUAkGWBb1OF6xvlNvpCb47f5NHSYthblANrUb7OWClbCH/7RoJhMk15OO6
/X4h/YlYTXBaHCKx43wGv22BJB7RUB7EPAkOrLv/ZHo4lW5Z3OtYgsKhLRQ+JKP8
UQhgjRLL4OlGoQIpPpT86x9a8m3hkJ1qy013Ol9j+EHN2nOb8M36bjFR2bYzzFwR
dJF0B5U0tM59nmhb9m9BbKnJParZKNYEnBuxm2KXqE10cy4kSDfpdjiXtndI15j6
SmogjysXR8mpnAyGJwguqLiWDGWN0QO593zDIfHrOAlD9eC3+Rwlg3hLm5ZiHlP3
D31QbwAiuWpU8f3Fx5MaNq1qhJiABMyUJLxD6KX8orscbRToXkllRjzLj8027RcT
3ieH2/+kx5Z0yhBXfzD5U/Q6GDJQf3XPlBkFw4LjTjN76y6WdJz/kk75t6qOKcpF
fO77rymIjy+qsiPPMURcTk6EO0cU/VebDv7pEsxroxQPpSm4jRI9Q4BEhEGn9FU7
iM+UFBJnaNfCHVDZ7t8nxRRMVeozx8tb18iR0VGweE/QNvaYz9prR64/eKnRhjCe
NZKUH5fJfkcfixGVEam18v8ZcqBIU4yPxkpB6aSnJqN6MgDCnxF59iOSZDAY/8g+
bfo9MmGh9t39yCK25237pbPR1Mv81z/rnx0VSMTyl4ASbWDmybLfPpY+Zwj3oy4W
f4SHggK+Q8FanSeTQ/siALnsCcolsyMcQb9d7n/yz/qgvjZBE6qvYEuVJviH5Ftt
4Jx1D7Rq1T0SGu+jfFhDv8dE21++k4t8ofGCCLwXwUM569n87ZiEIBd9vayh6aqb
M+GsarzGi/K8S/gfQ8BqObb00lSSoGih34yHCjsUgCeCe4K7u4HYyjkz5W+RglPJ
+mwgP+/AoTDALOmw8waeLTd6KwLvGfO9y1a9JmL1/U/e/hPC4TCHW5T78WlecSB1
pOk0ozYQal0ZSx1A1oS2TRQtZu9knctaCOKTw0YP1d03gsFRq+q3s2p7HCFeS4qx
k7WMQwMEH04OK10D3n98pG8TzOs0K9hMsCrNQofPka/YAQTCz2unRqPnJig7uAyG
4b74LDnPfE5LwLuVb849CFnFFCYqahFWixu2WgPjcqFmWuzUrCiaMvLoDqIMISTP
Ekn8dvDinXmq7w5eDpUSIPmU3IsgcOaplL9FMEPmvMbKLsTqvqX2hLe2CPTjVeji
ej1WrnRm7TH2eroVfN68xATnl7SIlx4sgC8XCmfUY2IpyXoXBA7kQVK16KYYvNL+
MYW1t2+YU4a7+b+SnoFIG4fpa23mtZhCFFGJA0Ipmu1R2dWhlMVpsdjF21mP+pfs
9noU2SvDyMjwNk/5QeAvRRnFbQF0ONhrSnAu4wZa5v5OqIigQc8+vCV4gzOCm9Uh
gzV7IDyHRiwrWKSllLV0StMk9RADFryQPfmz0r7re/XtGFrDTo/zO55WzW27PiLO
K7//t5r7kdmfbQGSoKi77SphMFyiBtup+q9UblHYPEf4GTFnh5LxefvLNMJ+b4+p
wRnq9KPh8hko/LEHw+uaVjJeImfIg9ncw3NlrGyl+6RGwwzhpKd1CwzU1HXoQX1D
W4aa4G3n5s6Ex0LYZQbBY0C+xXp8WoLs8phdN280oaTBg1HjiiHY1PXcIgCSqe7z
VbPXM+chPCrmFXKzc+NgEsLOpb9tlgRpzwAgG94FT/AExfFDph+0EaRPorUllwU0
JKc+xv9Gr94b9A7y/UFqqVGos0V1+gPZWXmts+0bY3PdTuRQbYNl1n7+9N7ttIqt
oY8ZHaCX5oeHK0SQ1VNpnQZTKfm3NeRhCpC0aIVWq26XDmV4g5HTdfnNOWIq2PWS
tqNZTs1nkvevLRmTwwriD/nmxdwwQfSJT9Ni/jAZEyvCAkvlTI0TK2Jj2ajzJqac
5CRYkXEFZyth9MKlMp1H1UVe8PJ4CrQMx7cwlkZvTh7KKa/VfHjQwDn6ENbfu4SZ
NsmIEGqXLclKBH3aXZFeg0oZPiU6KmhgO/pDarROohbRmlqPSdQ8/0jEOVgABpbJ
7SgCsmcImqrA0ehlBNS80LxtMzvq/6N1S/41ezQoIPuWLJLcM/HATnBtVBiWM57o
wrw4ePRjRvyk0DsIJ7SlT6tXXMaFuCAMCiKZOcOAvFkogKVV6a7zwZG+l869b5Py
F2KOO0Y8hoZewqYlifMCjtabk7WGdDSiatDrx0lffNkgmplIiYk3x9d3WctTOGap
mH3eIiz4mQcOI9oykt7yHObznp8enHpW/q4mv0pCXR3qCBHvPDbUeZzFLMwEhHWg
88M3YTf5jmuhJZlFokdZYHxqEe8yK0CMV/Hdjrr8Xz3C4RyT9kFY0CKWoCmQyxfy
85ovqrN9KLuLnOf6c5Pipoyuh5N7+Ab7u4dzk4xVdl1BqUVW196L3rsrJpxzNs2a
Ct0Xg3WjS4m6W5Omh2gf9uceojUhJMHFNN5vWnlhoNyxC3s/XuG5/aIxycs+RiLg
qlW0l4ZAItgKrkpJ6PN1HoEKiNQ3IOCOju9maCvvRImDtu2KFQK7OXz8/LLI9pq7
TCwbiQbJLtR2xzwfqZcpHj3j4nt1ME/P6Caaw1hQydQvRmqbG5OtYaqLoBS4cMbq
rzpEw7wiTIi+mppMHIxYjxjgfLqSq3fnvd24EMxzdAqMc8Rk4CBOoe1iU8+TzXyZ
vJ+wtuZhXxMsuqPnXP5XCDFzpbeQnJK4BAPFP5ITqmUar8U8KES8v+7v4FITH7rC
d9GJoXSUijuNjSt9ImOlOi2WoAeM0xsbNUBoEfYeNiR6iM3l1nFRzwIsAxzYxlHi
fWdSTkvSkh+0LxPc6feyN6ONoUCAS5dJo5HWf6K1+qOFt+44m0SvFXALyY/s24LK
YW1j9xs+sZejyedMRf4F5T5UbUHMtYxymhfbKAw/N5m26hp6t8An2RWNjQSKiZo7
z8nquHlQmaKlHgswRWMhiDcuGgq+5FRPuGT0WrzsT0SKFWt8zyTFOaITchvYZxEw
XEkvXaL8SGYkMNnnOCur0cSWECzcXkRnk+daH9YiCahyp4u9+6xeEJoUiZoJfzfK
xovtusJour3Py6QYBH3QotMo2hgfRwJHx+9ToCiSsBLmaUCETo2MIVVrqZAnXle5
QpkRERnecpcFyRzPSzcMLmtH0z4rmHixeLuqiEKa3dlAjEw/RnsAJmNXZWfS7ARp
z2N0QiUCiyX+9lhcmEGouGTZsprU3p2xeoYGeirpCbu2R2BPZMuaTE0VC6zgIEdZ
dVYgC6CoFJxBdDCtWz9+v/YqX9OF0qUTFmHEoRB3fRc5DxmLr3Sqomjy3qIllXwh
ugmApYiSu8M0/tJjwEq2DDH9q0bK7c0CrzzwA2Y7R/1e2vvh2iJYLESIwR9LbPgH
Gy/HEzr87hnym7n6PtS2EExaRyfbiyBBZV0sQWFnQUPszsdDpoG5waLVO+FClWF3
+KlZzdoNOYRTF7wsUBVh7dy3FThchQyljzsSBhLo1wRvyN+1jxSz85bkunQqeUGV
mWQMPJ6X18Zb6TuOajq1YaBoXOsj5XxKA8q/m74IzTt497csth1gTjxRZbz3RcoD
/VYB+Idb1FQgwFfC2tXrpXN0gPOrVWe8YKiX9J4MUc+QW58qpw7jX2DidGd8BYuy
d+wu4T5v/PA0/b8CSHRhgol0d3yJyKHbUFf4dPk6rq/y93GiDUp99H8tsDAAT9J8
rKgxw8AkvpuIlQ3oj4DHRrO6itoyzM36sb1tZTOL5e0V6xl0m3Upaott35ENnHyk
rzvhRn5FFC+N6UEDrD540ycs95ZyUNKV8vfEzErmq8q4NDuQPjUqze3eM7FiNn2I
qgzer/gigeWcVOx3ICnfQGMCBwlE8QBwMfdyltQRAqMJFl0ychW+QNvJdnskUOEy
7UZp3gh5jJEt5iqKIIiw8igjWsUOaqTLwMhC7MTU/pohtdwvSajHNbr23fvVugme
yg6rkkDvbhtTX64JDmXLmiz657l572ClYMsRZY7+dedgRNl9BRS1srlaVlNajBTB
7UULQJYNdO8jnwNFW6KLuXtNRUQNcugS/C8FG4AEX7HuaLuZc+YNGxQQMxYtYbmT
Wp3KqJrE2z08YOyfbFprJhRA7N2JiWb8JSSyzgdh6XABqfJUrJ9ZotcaJZ+I9p54
rcszluWl556D3PoHi22qxi/Kcbrgd1c25HFlG6W6h0G2OwnbN2ul9/YYJml6rWbN
eYpFGDkkKux7T4Aq1qCQ8iZVeAzk2OCYbFulKiIVvTlfCQoadsl+5cnLBerY+FLf
sCdqefkhj8GWE1sI9AnvvZs69F5H8KI0/fFEUQaUxgWd7ENcHpKUlWZODW0epfKB
mpCvLj1ujuAhXxzxgTs2u4LWnknUUIsuhn6TAAcXR5Xhjw3hKhV8DMTEnV9EbAO2
lNpmyQ/EgqbjPybyTMPb/uwzniR/lCY1WFbgv2TKUAYxIJ/l8DosvduW3qvnmflL
lCA2iUylKDlK/wUKR/IuOwY+wobAbMeR3DzMKUGL6suSij8kM7ZEpK/7992MEeyq
RLblqwuDilCsvqn/5fH6skoUaJ5vOE5Uso750zSace2MAGEqkXAj6lBhEbVcQbFZ
J/mmMnnoL6nNqHzPZiXhVHrShBycJyXLIWDwCSymG4QEKiKqzNef0AJW9etAXffz
FC+9VIG7YqYEPxbeon4L0at1Vuv86UDizq6Wpz0xjYAgIIxoKsQ7leJm8nENNUBO
dWOYvp8Cp72q+aLgw6F8DblNLUtQTFqvtOfQZVI+Be1Qe+IazNj7ttta63RE+EgL
fHB2f9+j7+82V6XgWFKHRxS7p1Db6kcmjt15tZWlMlyAlloPdI9dhLddhmE1rnTa
u/WElS66K/VzfoQ6S0VsjphokU/RDky0NqxX4cuJ2B6XrA5Vw3W4i96mn74o/e/w
2k3fADBvv4v2XnqQfFrvbGLXkPF8MX638ObRD3L9DzXg98rcDGfllUh2+VEMAJH1
E/k46HtH9Iu9OjCGAOuqtGvDgyVEdcnc5eTs44QMJBEO5azBhhXhsBa7nIcz6CZO
5JgZoBbXGqcYivc6e8tL7eb+paIBywwcbPl1t/wqOWA2Wi5zqyI2XLPJ1+cWZ6VP
3V7ajmKaH2UlgvxoIfndQdA5z67Es5P0ybcgtgVwT62Dv3WtgI4olLQwYIZ0SROY
VTvnFWk8kjCWdV7oOyhnhEHGk/tleed7dtBei4XFFqPgfmeNhUa4G68KA24xZ4U3
jXE2D+Q0mbteoXxcETMODIve60Oi3GBWUQU+ieiU9+o7eIa9n99kfycDFcgX66Ov
l7j2dkUuY9iM0h3snb89kmn15MkihKSe/cDDcSGtgy2ygQKjoUcFBGtUq8HaiYSl
5EoT0HNJfM6DWP/12jMpvQ7pjw5GWlIK9Zf+p7xJJwo4JYOYJ6QWa66IwNh5cS/2
F9yi9B+v/s9NYN9qbDDB2+tYdI+SkiF62pqMtd486axe3t7eXPcaJ1NkFefusfyv
JFvTZb6zgdKj2X/xsTK6JnWKHN4io8d+/1O2WuAdOTn/ZrSgJYL7FNZ7mGrMdGHf
ZF0FgNsBRz3U4dDYMfIdlmZZM75xYmW7jJubNaSYyotbeVJAbn2TdulogyFOw0jD
8FUJnEl/PB0VmLFhBnxSfMTklpsjEdmCk2Q6RXnPlcaKbaNehY1YU/68NNLFaO5z
Fs7LyOsGJnmZpbG031wTkpYvXR8EIaBL8K8hY7iZo8utbQuY3Q8nu5K+Lvmx9YDa
xAMvpjGC1Vsc+CIp7ST4isO5agrFYtbhkrArSbgmoL7QxsM8D9XHWn2YmB47zP+z
ZrEmlGrtq4nacbbGvFot8E7BLDhm7txEyQVjJ06xuoPcl74IqBbSVTiBV23Her1+
T637oRVaeL2izvijAic52fe1MjdePYIV052zxA3EQycwBCvdZTGHXmCNbckMe7GF
2oss8FkpDDAGmFkIQnsm2YwIA0pDEkmXp6a9LE1PV/q8vHs4jbgzVa04S7Et4KJu
f4StWsA11+s4XWAg/q1pKojGX42l+M3CpiZj5zew4g0HdT0NNSrcKYmVj2DzLYOi
ecLwesNAdYEhnfVrd+zbucyAW3eciuPC8P0Vt3RpZi6GFwHw1Lk7quppi7lYj2pS
1A67pfqRablzmJ2lrAuw3AXJ8rGJ15GWEUUVKfMuVxBz7kOjlS+8rZAv/ZM9tfk0
kWFuvbP+GaMPKbobt6fythZWw2jJ3y/XZHtcLxDl/TfzFLe/xjKPeCKPM3A1TKiM
ruD3JaSzKpPbDcE0doGxkWI1MdWdgSEy9OYDbjfd9FmJD8P6lAF38Klglap2UiY7
wEQlAg86D2fMZ2FVqCBGnS55NwVUHWJMXU9rud8J+G5c+sCygpDc0Ag7n02Sixgd
N8iA1rAh9kDIY1uBBc/7MLLZNsA30XEdhUuwdt2jaWUsL9yeWubINuGMprotcIx4
UfKXOpC/bruCL/nOyhFOR3h8lzMxiUsmvdDK5dVLLqU4PPkfXak23gZ9MPknNAgW
fVpkJFcx9knXLn8bIcwr+RfJ7apC1tJuX+G4wHAFukYoK+CdkJhSFnwLH/0G6fwu
8Ci8HSTyO2mH1d4LiFFx1YE0Jy7bK56ksBU7AI2oFV44h29oVe43su7S1rAHady/
wCcaJ8A89V1SLBYrM7/OMwQ7SP4eL76ivu0eJa1O0dgaG2624SQha5Te+BfVHJo5
I6Q1RcqVKmj0FVQ1rHqbIphMAkkfU7/f8Ya1+3uIEsNoznGZKfnfmZ51ophZVLe7
uyq9fegNl8voShP4Ik+fvsZwf/1mlXl2tDYF3KTfT5VjkjPKcPwGT/ij2Ib7vg4p
hZe898NOcj5cmXj3ftEDL59o+vel2W5p8hnlHY+qLhHjokiwFd5thXbXCZb3d/5d
MIHS1kJJq+1RaG+WZWIEcRfQ4I23xGEH49caB6pAI/lvaCHFvLvdca6bdgCuGPC7
ARQ5Ynrsmjt7XroMBhG1fOb//0qi8kRfU4U+AGuJLmde5Ooj2d2AAQ/IRI/vgTZl
Jd833dhkzokIW66EIaWZbHjgyX6XoSCVFv6ALTzKu3nTDYTRCWQnsrhYvMwThdNd
gCWXY87eJOQsyZZNqsf/dtyBDIIhgInC7T9bUOId0PxUncrRSKiK8B3dj0yMtlU0
lnNqb8EOgLsWot26J+Ddd5amlYWuK6nS48uqJrI7aXZyndwVO7GcTH9CVZxQD24x
iIzt7etMxZeP+WirVhE3/DCmANMSFtLu7czh+2xl1uvui2CMDDCLxwSb6s6YTreB
NMkeMuSKFr4G52x5HkXXG4bVil8EgfGYxwl5rI3w2Iou4Rn/8KTrdj918vF7ag6b
Ds2sSanOxiWNOMjfqZ0z2oFmePPD5VcxJBvA8MZQyakh9oGlqqjmPu0XWvMe6iCl
BiETWMHmTwqnuPNG2knkqo+ONosWDqKg7SEKm1xp27cqvlCttFwI40V5AZ1BaVpE
BnJZatlHn1TTI/yyosoYBewqgt3h62uAyYqi8iNUfGS6m70ls/SzoMY1e5A2w0fT
i+n27Vx9IcA5zDSM4iG7elGMO6aHaBmC69bNoOiA5SmPL7OlYv6rjQic6JzQddEr
xLaduNI03ihWUdzDdDLWKsO/1FrfYaKVl1cIBimqDsPTATG6hUBplyqOwKsOxoP+
s7OclL8yo5NYJ3CSdL/8SdJdrlg+F4yGEqPuVR39JxmoxtffvyW5c8M6x/GaZjMK
gMVxTb32wPhVEtm/6VUo6XMRAipTpETA/l6JVbcOCJ0nFuUr6m7byh0jYbown18Q
iGUEaSpuTFXLIyIedCXCqzH8dTszjuytF0EuuC7ys1EC+9+B/JCtw83I18QTkes1
iMrjtPwM2EC73LJsDW+lwfen9LQgLl1UrV5mcq9EW8qFHkmdPTVNhZvk+wKIvMxq
NZc0rBQTWTMHbHVGrpGLm1WxTGHEq1mjnr6WQA0iJcbTFtyup9GzyE9uzFSZBx6x
SasMdQsysCKj7rbt1fsRsnS5iKDRWOJu6IMcknW8zql9axaPLrV0a8IXudNGa7Jo
pOvmYsghEpB4RlKVCWqsQ5CDKOUcpB2SzTPniu2Xx387AttH9/ANk7CBvTzMAywn
ToPgU4kr5wFGlUtQXQ6HZ8h5RzVN/Q7tfOs1nuMPlph5Lwax7Qjs+YTr4FfX2Uom
mjj8TgpeyfdT/hYO6DTKw88bTdvKyNZLO7W8XzqtrXM+a3ukFfvJHsAGGV+9UgPa
NjWx62WrtI5qZu22H53YOhgG/WaJizaiC/DvBj7r9S/tq4WulfdZE8aeJj2ouu6I
kwFIq8KWhGD0z/sYeaOR7d1BG9TQo3Zsc1Ui8FTuE9mioQVVgVDmPB7t+NNSEO88
ptHO7gcV8lxzaSyXAb7Sk7L1ANVlX1AftlLld8hARWw5bQ+HcRj2XAAFF1iKM66Q
qJzGDvvUMmgCkawGxRzH4zbLxdAu7v69FvccRMCwwhM3rq37ejnf5tsV6pBKnlY6
c9mZx3WZii1GivQ/ehwh28NNIAKaKzUh+wbMeBD76oRcB/gI5tDx0mHaPpiYPiFS
wsXgAp34+PwDkGzw7W8Pc6KICQrE1HKffKiatZKtHXewm/C8nbiPbzAzksrnPRuP
bVKBCi/xJKj/6oDguCkY6BoDNVJFGtQJUeywqJIypnLYFLkKasjmjZCONMAwgxi3
JKEND6dPtc9lCB8p4qtSBKrGtKExYysK3VZo4905o0tNIr9hElhQBi1saG+oXqmK
2s8ikeqqYBWLNX70hJZaiBY3260w0T9KHwzSB1Av4gsZy8UlDmeqJIQannkRgHl/
i1pAT8Mclb2cFppOYeA2UHGiYQbj2TpEHzoa6b489AzGFZAoklmJ6U/oqFT2EmiZ
abJpG1SoiGZ3+1Gv5xt2eZs7RCBLOpwrUldFW/T1AOuxqrVIaex7r1muEm7hS5Q/
iZDNMrVsBSIINc3p7qwQkJQLUpmSspk0N1ixtjpnuR5S/XiMz9ALA6HWI8/79HMx
hW490jGNTCuAySWaELhGIhe7JOmtCCZ8NzFhBMqqqb6l880DKo9Li89LYbiVQKud
yXUtli7cdTVRv6MnuNXBootVvlMFju6X2aqNmpuiJTbjxuDwa/UikU34XR/mNIFB
8OIHanzbk7ILdWgjjuz/wXORY0vLUQqusVMmZC1YCqX169VcJQ5ewPAjYJH9f2UG
u1UJgzeRb+yJs6+VY6iomI1c4XmIkjU9BqYlvhIkbVZAJgAmOC69zyRVGoAXyc6V
+vgWQIIANQvQnMu0vGYkfJwikpw42uEhdCX4TWWIwBqkXFtBv1DIKSa0KHE9oNkA
bVlJlWrj8VHOp2YoTIOrZrv0azSlGYWG8UizIUo+YNucurBBk1AlGajXw1qAMAeu
jzUGksV/x1NHtTR+bnp9nQOBTnuDtXRC6wzImTyDTzcfVEXOcWW7A7JKqjynCT9S
k/ak8n8qGoxfQu7UJbcRYyYBmNcdSbVr35MHEgPxpRTGBN6rvZzNUyJiTI9ZyiTx
p0WPyOPeWzVLTWWpbgCskcGcEcQ5uNPKTRF7wUTdYQYR/UhpfTQvJ0yI1nkulArI
dyArNs5RmVJ/TWZhn8kafKEdz2gh9QBlyVkqSSkLUfwYk+Dpag8mA7ezGwmMjzs7
U4QmjHCaM2QcjG/Pww1CDHtZc2f6GdV7+4eIgXveZeQeXeAUqAk7gee61NVCeMwz
O8aj3iP8TS1zyC/hOYBq5bl2k796PrPgVXZRgPDdFaibELcpBuP9Njb9BIMq7Ore
mlur9PoykpQwF04GcUJRwS5oS7w7YcOghOq4H8qRNUyDtu7vFJFnncmaupYUr1Yr
gFWbOiKqumrdrq7xfKx18DtJjyVxN86RO//hRj/AZLPe3nzSR4YyaAQGO4l4RbXX
gGvdF4WrqkH+YYDf4eKDBEWRHd2fX2ulNG/7kkqsGcxNoVl+9SNdGuFVT6HlHkgt
ojTGPJ27Sy5p/2PRCLh7GB+SnN5dE9GSlx4O99LWAlAseVGEDCVzyVDNCJDls3+T
7GLBORC6WK9oG4uscLN2xzGSP9F1b0SUoWHiHLvU9L2J/2R1+YW6JYMM6ClyWMjD
edqt0A9mVprO7Nvl/WI8Kym+BdaRj0hcBXQBID9zCji7qtq0OFIA+sZCZW1klNlV
IGWZCXpC8bye04V11uS1FiqkgO7drV5hO7vqQxTxM+Gpjj6RZ7Qpjl359d3ebORg
CuYtxo7Zi3vz/pwInykGAfNOex98a3xyroLjqiV0NRD74iv3PoFIUKR+QLwK3bBo
vzV316NdeuqBm1gyxbswbVYsb7bGvdfnjL+vzDKXM3ueeqgw7ozVEEau3tHVehKq
ETiqnqFhhN2+9nApx5+k+0hx+pHGNJxZfz2zyZQrJnYP2uk2K8kBhjzt8Kjzw9b2
B2RGv8Om0Ub+aTrnlBw/XBayqPLNzR/Z2CXwbIT9D5nmLsdQ1yJqzH/DB83vijO5
J/ICDHEW3mxbmGtTyXgutn9gRpZ1RuJgOmoQ1fupNCwy3CXOaG7Z7YHnVkJPi9p/
SlVHxaMelBiCAm2S+x3Gzw1lCteWzOwzvJ+CGxNvhOIJhmbZALx+upB4QnRtwWUE
O21xLCi6puDYZ77QlQh45R/HMUGATXCmPli1VOEAIMK1ShtAS/VTed1yKsc24cUa
r3BU1Kc/VyaR7Y1XfQlf6YIf+ZvvgtcDHUwChCAD9StGjqpRKD+uMXpUa9lZK3xn
c9sBLWp82IRS2ZuG2IeKWgdEnbtkz/uiLLwFhQc8X33R/47l0QkIXIFEpAaBlsRo
ioi+ScqPLShk1y/+uBKHYprvf//jMRSPEEDnqKb9/+NKk414Vd5g17m52WdjWdP/
2rOVa0CAuJgzUnDJoKmx17GeKj3V3YV02ByhpF7xZ1/n1XQZgkID3wWn/pZ1HS08
YHOy1qJLVjIE09le1vwWlQYX5i2SlPlZcJfBPwJk8xvvXhDkiVCwoRMxLTfC7eFz
NPX04pFjDuCFMakYdirt5zd9rJAYELtgrLtt+FFvpsVeH7LMnS0smO08ogvNo/SX
zgYKAGX4ktnayVIYNzE/7khc2VtVdRgJkoKmB3saFOJ9xWteM6EiEsQsq1dMxSPV
DiQppLpnvcNmkYMGvg9NEPJUfHQ/mnvZdPzcm25nmgoj/Yx/jEjuDJ1RPFiciHA+
7ZeTa1n5+2Sn0PshUCByZtGbt1MUOUQhXdg2BrInyrcQKwESTZxBVyFTYUFNlCa8
V7qxhndOSZd+652Knx8yaJzGckYsWaWrw2MH5NTYCIOJx5gq1msvEHK91+UQFDLW
hVHUA5L2EzN0lwQpgGJdsZnOhTBwLtMlBK78l0ygw0/sRfO1OdJsunVuvEthOzAI
xmSC5LTLlG5z3/jDHCb9mDVo3ppw120hTF3zv0hTh0SvWYNQ0ENxnj5YuWf37jq2
j7t4N1As1HYpPKpsrrL0QVPGqKgKWQ67oGj7BKZN3L+WMvExz73ewXKzyesmdgyg
kBvWcwWDK8qGb8IN+CKN4xoFIzQKqBcF7FlPp+XUNfaItpHygv/cLg9Obnt6HOzx
v5ry1ueupKVUA0skycqcFCqs9Wk+v9YsTDZpaRDdftpBJ/3cKcq2c3Flhyu2YUXi
2IxZEeG4j3Z24J3DBLfd8M4L46j0Cd89nEbpI/udr3AMyd+zV7teS0KUXLBROw6D
7YYRTmYw7esaoBXichpLCS8caKQNQAuRgSi/ekop5QhjygKv4E0gPRS+4ClxjKFf
Dapq8QQui8ulaOYVOHYRoLmmL8nTDRiyPX/vytlcowtjzO1IV1HpXCppr+1/e9D2
s3eA5vTXSWuwWnqRsf/6p3NR0PYIxANHZMa4K4PeHiL0npt2tJoV12l7xB/JMpcH
9+2Fj9C7JsUX8hKmib0gdYwxz5OFhVSvH94fQI0dPgqeZ0kfU4J4y/rGFq83869C
PYpofeOCVM64JWRph34PaFh4N5kbfFVLkPqLTWmQEPPtNhVTwAzx5mcHCOOA9Aoz
fJkyOvCmdNburC4kLLak2kONUnK45Mlz3Cd1El3OtMsd6i17H0hCW0jSVI1C8WGa
Zhwqe509d0aZ/LRFlxp0f8J5nUVfZtSUOuHpsIfYmp0s/P6nCACfkf+2mrjI+aBe
vk8e0FAzboY3m+GRZ0r+LJYvGQp9MFzlpAilEToPEKhfts78FsTNXJzKTewYBq4z
Sw2hgy4Hlq3uon0FD0mE3+Q3xtP4HoFyoJqdub720KiyHSJDI+QizwLfUK9NH3Y4
dk+ltucMLiSJ//2Yety9susTjjpGcFqDcZKiXTL4bjtfielcymy5lVYou9xrbTe5
1W8DLYylffPjn39JRjELo58j72IDqmE4iysu0YJBFuMipk9yAayEgfNjSImajC+W
Cep45eWYag0daIUiYFHhrTwMgUpGMzjWtEENggGqi1dpt//LbIIWLJqBIfWnk+Fh
F7gNhVHJe21XUDqUVCKE5EnxvIJZ91QS5IHNcqX3Gxon71PoEaTh89EbXmWBPZqc
qddEXLE4X88SdrFLfDNqzU9aAaek9aO3VeUVAohI+zGUIWL+noN9zIOEbsf5nqTt
5Af0WswvGh44rtQTsIqTiuk7iydoWa2uCioJxkZyRZC/gvSbA1zhU4p51A3mVOpa
x5VcBrtMB8mNv8pdMOB/kVoqMeWs/9/B2mIHyt0em/oTa1NyCHhCp/0ozX7dMU8I
gwPGIGf1Hg042sLVLBzHcMlj1qV4cS4bfiuGT+AL20Py3F73iNx8bFefFFbWcypT
7T05K8L9N1RfEsUHet1T3fJ33rHQ5xycjqQZ6MA8M14yOp9kWAYlxfa1hTOR/EDw
JOqAty1KcftTrYK1mW8VT9lMfKZynAODDxJ6U3tEfFeCT79V6vCsyl4NKZe+P7s5
6onzKgNNG9s/wVHZ9I3NLukpQIcAurgmlWTZnGHqYuRwEzWrL6bxvQUTBpakHCia
y9Yq2jVLcCJV+8aXf9fhHDX3efhhvZMnQ2wRQ8CEF8525U84nMx9k3/wM0uTeppn
8wvye/qK5n2VI1BUZO7HFWC0+VGxJF+6BJbTbTc2ezB2gCaTZkYCKqVVtr7YHa3P
ETDqbkuiYoVrRLwmmRQ9cPMY6isRkh1M3bgICgJ6S6BA/tjwLm76hSFz3OkWURFJ
GDXaStYYIDux/PJtq0mDYnxl3QB37vKpgzCyDPierA7WKohKx4zBB/Za9iPQyXhQ
g/jMxeBtA/hFrfRtLgCDNwwSVhfPC0ZTKh83DOx2+dCARPq41K7TINK0hBvQTRpe
9xhENPG/9mMFTKFlinSDBiUa1xPjIoiBUWAwetcHTay/gavADzrvpTW9C2baUD0F
PzAgJpN0z1LKIGNKmZKrSv+wDvDNEH0STFQv2jlAA5KPmIhftXsUfuXAZWAdlUBr
l1SbMb5Cd1vOMVnGL251kocFnKRgjGV2g6aegpUcIWxFslILxAsNFQnrlPCACk4D
Co3BFOtqyhm0O4BI7miOnG3wcO1Xu81oOtuGyNBHPlXRLWXSsSJEcfGJgVsAOD71
Mj6Y42Jsc49AY+zhaxORyL/nfQo3Vk3ITnKxDBa5+wmPcms6TZama+eSjLMNR50A
KDrGSM9a5a3ZpSsh7d26ixhh4Vg5rj0+xAshqdDyEB0uJG3sjwxkZfm122thyr6Q
KbGufOLVoBdmE+Xt7Yt9+T53BtuGD0lMfMNkwUyTGEH7KuW9Mqp21Hvx/D5/+QYA
APoiiYtjQA4xRF1R5oIWonb/qHJWFnK5W7T1fBUzWupBNldOSXB4f4RDrj2pWvEz
vshisqr0vmQFt+IlW9TzNv/F0rTo8YLQ0c7XXp6fumz9OyJ3WWQZFZEXYCY03dXy
9rmTG4MBJZWY+3OMlCpwTH49xF+revY3sfRwlrEEWlSEYXsRPWAoDR0fL+Cu1coA
CPyG93+j43+nIGOyy8Dp6fQKCrmwzb0+e3Sur8CIWTpggZR1N41u0tMDiHg6nP7k
eDJKYPNtIvnHg811yVJMpLRLeYviFCD+esQt3OyUCMxdvtpZ7RlaJr9TeLIOdY8p
MkXGIs+seiWEYTPeA+cwn0mO8lMpWqhdMFvk6yeTXYEYM8F9sS1+j6xikqSt+oYH
qOWlWX4zll0c9SZMX5vmrxLPv+xwyDX9cZk8vCsDJBFho0WUmrvdkRk+ULSHFI84
wSMfNrh7Rbpusg+t44MOKlzoxop3KG1/M8jv7kldAW6ZBj726VzC6PDdGazq+37K
sXQjzk7Ghm0lgQxqGR2OgQXZIDb+jp9VdyX0E2xMHxyG+6K6muiNasRDgejorLeB
uqsQd+7HJlH9/z8/zpsKc6RsOzrjfw3kWsDR7AY1DKRrxgZyq+MIsMk7dKhLvcTW
zvouPk98l8n2pwSaYPD05e9gtM5YAksKf+LP8P1Yo6wpMt3VXwFP3KwU0wowxkUk
GGNpxOH7tLZm13K5Ibma4SKiOskbBo+o/J1FUGqLREHwFdp9SsusiK/yEVQEtDPd
iegTGw3V0xXc2WeVT7mit0m3/N4AqDNgtsBoJw+NxpaunYKoLDGzgMKZjPgDQPNA
qUhx2IGk6anJ+JiaW5MgVezOcPKEdJAtnrtAuDlJtOVa/qRmNKatiy8Jc4mEAxju
NY8+M+tcU4BuhvflKZLH0NRsJYfIJKjeL21r+AOr8kfXCVOXsDHw+tzWOxcmY0lp
xmT+lGwkzNC4+meozB/ZZdmuVTvEPow3czXHj6zLqhLAcBt8z02c1gdoJ+MrAVTT
OHaDFp4zByua5NXcP2dNx7cyMEHfZJBdqOAaCT+y0UWUnjEF9f1HCjUcMP7z2DPA
5SKVNnE7n3QiVv9aqnPv3BsLpe/GN0mQ0Ud+nVlyp3/eqiw+qRjLkUYHtYiIftBx
n8gVTYcAukWHV9a60ZiWYgRC2KCYUY698S5vdxNvaqO/nhIzPoTxzHS0oSaxJJ5A
X8yt89d5u97M4eMJnAbbdUxYuvEzDBa1mdJVmRigaB00o/5YbHrgSW7MlXCn8OEX
5v4ybVLYZAnhczhUpc6y/2SAug7OovHefYsNmwU5BYqsqLuaRUjHyZrswzG29z4/
9E9QCRxBJxjp/2orukpGziStIJXQklT0vOZekQxmmCSL6XbwfcpB9wogQA6IVDd6
shBXyB1dlnHvn7PPbx4F3dgDRPLf4MHnm8kIaMooALLkXLp0dF+TyqAIUuZzxXrl
j92obPtmfnitNS8oeHPnazkouwGJxO5ZvukoWXqO0yIT5/xcC9jDHNAY9zsHgKQb
zpGyAr0Ce9EQMdj7tXX0vrZmgBIIv8Y8ZVcIH7xb5JilSVXsFsXrriN4FYjJTUcO
+Ps0H1w6VLhPOX+7AqnUdR/KeJ8FB4sN7wk3w4N+slY1NJYzELTdp5vyd4yekhsL
uB00pmiq18TILW3wu6vBdP1Q9LjcjI5OQdMqq2IYgLDxlfFL/q7HQ+KKmQCzIIaL
+ZQtXb5/U4jTZqr2goGZrs2VZQGSTNsiBlSRhF3VgH6veL5prqWBsBBwoHc76BKu
uBdyxeoys6P2XFx+e8AFkcHNuCI/Pjh2xX07LijZ9AR0Rpj84hqr0ggJSxHU8VQC
MoIqu3xPzKecH1m5Sj5hCdxn1niDBElawPLdocDrRFkw5qA4ZZEMavrvVAoMqf4v
2dWkz9wjvY5DmDRrdcGJ7ohkm1ukTlWyw1TSIsmutuaGcoCshk7ZzXMVORckoShF
0jPSNP8y9c+Ty+xcAt3hZE+TClig0Aou/kiiVWvAcQlGPs8E89YGm+2yZL3WTVtv
2jMzTwMATvWH4XZX5vsv77QxQcKfoBMVZThGABVRax9nhrycfq2ZW8d0D8kEms7u
wgDysi0b7G8g8bYf0f9c3um96CkPKavjSjkLnOgaM+C6zNE1nA8S9B8TAz7N03TE
BL1xGp2Htl2btsfYXE78Z+q031f/nL6OL7jvP9UccKU0LBFkb6rJMirrJpw8yqeC
LHyikL1kXkEjpaaMBM9DUgoteAUW2fVgYJHFanu9PU1MC0/xI3AC/QT2nN/JG6RG
OkGp8G7o0CjFSzWGzzegNfamm1B3nyblGv5HNcsj7EPApWPxVgGBdH9MlFf5RA1N
Ebr8D0OeT1TjN45/1kM+58oYQf3mlY1Ekx6AmuKIcJ7exEN3XQa8udJhhHrzsrTA
hLbQwVjIX75mrQvjtKT7h5nUXnpMrRGfr4JC8Mlg4AFV2Z26Dyq2Wg2AN1jr94NZ
U5gzfF4HZqYh6PzYAiE1GYZrofWRRnmImvkIRb8kCtA+DzoetnuJ/zySBBfKFX4d
mYT7ztMFO/MZwZI5Fo/Qo+Tdd+CeG36BXL6TdcQIsEgEvaqIdgI6XwuEDaD7bvZH
SfEtOqlP4T99HTSpfCVqbrFacLJQd8Ss2CcrOzwmfay7HqAk3AcTMl3LUEmqwAvz
EXdFNHA9gmERydcJLHi1mrOcyp2T+aKmayWZcp+FY4DJk3vnn3ma0MQbNXeYgICm
sf9fa2jHnDpwrR9trnTzD0fNKTA+zwEzGd0ZAHtLCTBHo0Zw8JlnLVzScR5crKBN
7kNQHIEkHsUKbgt78f9qB4fYH1CGxwY3xoJ0ZZ/yBpr+T2CWYMr3NMrhiVdbLw4b
fCM0Nocw3wkgnlnt2FIXLSZz4ex2iX8Y3Kl3xa1UMrAziWCGOqjKlMYYUUQ4Ir+Z
3MUo13XCHRNKbWhzOKD8jqhg2Up0QvNGJ6v3GtwePiBGYa5RtcMic7aq7F9vqqoo
YURFuDQ8f65ZK+Rp9zk8bqcBeiVENycoe5rDu4Hmdr1z+0BV7B7bd62Xgu5aEmi2
TwSReX9tNj4c1PBTkl/OrTHRBFY0k5dhVr6OeHwbtigfrQubLLIu9RAOjOkoPjT3
1Viro15M4RImLLE1N0mewHD4rFelIVkSmehNsSDWzf2fP+JYcOwv4BJWitAS7u38
vxoJFGDRvHjjK/RBzC0Wc1GmI7JQWL77yVbpg7jpt7MnD9YOV9YimSpC6nCME5Pc
5PR0P424U+xNJiN9H96eREpsrDWsQcV2FfplCqrKE2fqE8gsZaYXdDnuro9tIhU0
cmGX4KeWS6Xj0i6+tHfzVFtBc1SMzOm9WXsgfmXxiHy4sjV9TdN7742FoFNT3nvP
9TNPXNtBpa5zwQU28g0QuiIya+URkpXOkaFJpYDfXHC3hb4fbvyAIsZlhsxiuNKX
gsSqadzKDaScQ8Rd+lQYlqRwKPvGEiP6o+SprmyDA2KTf5YiE4DmT8D8E4qeqAfE
bXRjbYCXhIsJjnCylZ70uX6Rgsx3df+IzGklWEpelz5wNlP91CJMxJBoWQqkrZoC
S0X0y13CkA9R6UwqWa6Lgx8ItXC/PldJwljujXI/YWc9Cpq/J01UJL+rD12jDN83
q8snAEWZbxACXhmoYMWPsXgqhoDPWzc+e6QUu1uwqUHSkBHc7jNq64JDApGBBX1M
4aFUdhrgBjneqDgGfHNQ+szq2dH7e9CfwllLbU55WF3p/ZVnaPHPSgouexlb6P1J
Xw5528QqoNhzUMpMJ/FFnPY7M5Q32KFlY4k+s8b2jaDrqRooQ9/jyzhdDZfvOS1m
Effja66JJCSOrnbBFZCY1NHV6bDgD9PwpZ4fHttmc0XCNC5H49h0HwQoFXDd1pEc
Naa3GWFMluYVHDS7X02tYeiY6VFYgLgJD8ehqh++yWCuj00WqCmuUIprlaxM4ei8
+37O99S8y1JU9hZnhqTHXpJe9XwxvVRn63ICG6ku+mbCtXab23UF5pLHyixNZJ4u
p6JFA+MyKMNLyaV2fTs6QK8GYYtQbyjPV8eeJX2OgQBDwS0jL7RwVKPM0FHRqFQd
0eB6cOYCNMSsxSf+BL11D/sUbYtIyt94q2HOgW69qSU8KuFOlQEj9O9deVfLpgCG
dMaaHJMqlX4KsBiGzEvHIRlRdgrw7pjF42Pfx6ZAXoKZhcci/mwuPsEjyzcFicR/
lxICDgdFu79iLtZJ445EKwZZ4vwTYlv6BTiOrLUMMd/+4c700m8Vjse6xtVAK9KK
I/Qn7IRZi91vg0x6ehVWzA80SLFLItoQOo4JF8R1B3hY13Re+ClwIWjUUR8fqoxK
AZaqS97Kuco2VSAbk6t4lGGvANmhyJjppASxCEVgZjgLYGMGQQU8v3F5TB+ix1xk
kvnin8PkOMQjQHyhoM8nibmFABgIoBVYGwGI1/C42bpMj0sz5zjCqOab4heXvPr0
Ignvum71DJx7HFFfCKuBHKQCI4T1yl9x+htuPJ/oC0JWbYDuFFuzx8VQZDtj3yS1
ncsCCYN0wLlGgNmHvMvJpk6DAzhnikwNf7x2oz6DSKgLlBWpit+u7SzL9d22cHT8
N+dvpSLKZJC44gvKn2kaiRI6MmXCKaHr0N9xWIU6BTRYejSE0l/Pmxuz3gP96nOj
F+U2PGWTi728gbCNDN29PTUsLBlAGBlg5x36biXFbaJLXxVzog9qfel7mH73BJlR
ruZ/Sh+nwNk23QGcalQcaZ2HKi/SJjlrG7IADW1BKGtWImy5V2HfA0KISlZbHsyg
M4Ngg4ZB9ASE4dAkkCEloFM/Dy5Rb0ddt6Zw/7vCvVsGzhToYu713Sub4vTSQMpD
rQ5yK8GRUwLatv1RAgQJtwjsQSuWE163sfDrkxhsrZ1X+++tn/xi3y+OawEcGmph
AAgZStIlM28daRUWpa4bRUG9rJtEk/Hu+tM7xQt09bc4Vf4Jnw/psyPdNKfv6Cr0
nfZXi00IoTktLsdTwzkCb7lZxEccqwwT8eUpcIS5W4fMBBMJJ0/NZ9kHlEAeAx6E
J/qfKEASq6ze356WovxBXdZCZ09GHCQGt2uj50LcljMPPmzbHd333awYEvAzuS45
5QlqKyzvVPNdcngSbw6JyjVD4AdByGZxvllfBV4tbfsld9mnDyxJ7ud0wV8hAacy
bVXJSbSxqOho5NR5XgmqO38W2iTYB5ZwAggv3OYpUwbj86wyunwbGkJlbxRjLhYJ
YLuGjTQioLIH6b6qf/+vzIJJuJdHMmxEF/JdyE4xVFFFMewvfr1S6sg5fKrN6juZ
/RZZvJiX7s/avmiJWBBO8QoQYTTBWo10OuawWUK9X9Dg/2BeCihIAlYI9bbFL25C
LlX/fU5NTitbeJ7zU5rGONK1SoAElpCVPcXU6HB7RwHk/pF4r1yBhvVV8ytT/mdh
us6qHhZdCw7iOIcRXg2U1lrXwShEE84uVFvK//N/V8RakbZk7tW9qyFfkRQJGAJL
Grq+qGHpm/uS3pZ/UN5ECGY+Ck0cAjfCq6eSd3ZiXw4CJy5qhLcQwb+WlCKhe4Nh
MymJ/nyL1+a42a0JYbXkJ3krmeelpbeR1hzXkXRCcLcAxowEKlr+9vk4oqTYyqv3
/YPoaMlfjMdY0d5kOIOVwGBkt8p8SENXYj/Pvey2VbaTtCYPPHD/205mUHV/6k8r
hwcrJWY08o5VvdXrB0kZKnRmjcQtCBYGd0xevGpWOddAHMUNlT0pGlheIsPQugh3
ACfk12ufnRvFyFQb0daG/mGWWhRzgP5ljc2wlT5kkBr07cHFz2tpngrxUwT/GRxb
fE6lhQLWwq4EP7u8lIABk5MtLnnP0gC0OWDvR4vhvWbwh7M9pQ2PAtajd8oRGB/W
bq8oWQDMD5I6K8zLJH1vFa7Pixf2+0I9ZNF37jxCAD7qkG5wLXMUx/LNwpEhDisj
WqKCbPIluXX7JftauyUL0+bG4nithg3WzsC88U18uCOaPVwo+5Dg5QW+MsUL9qYD
GK2cvrXtu5HX2Dm2mQSBzTVyIHweFGs1iV/qqvJGYrB5DMRrzEK8i0writFVj+yx
LaI+si+iwbDnRbHdjHsi9UvSaPr0SLOJYswoOvKW0GjXh4KxO5y9GDI1cFpslne7
ZhOk6RZ3ssP29j0mGRapATDuZXZk8btzcGLndlOYZo8vvmvUe1c99dnGhFtbnnuA
5Bbe0oLTOT8x8VwYbR6Lr9c/ag05cvI68Si5BYg71IIxN4OSUw7QzV6TT+++tmDG
XwS63a+99bDyTS5BIFRRq7GZBgwqMU7LYHDheXEJHvd4f40Imx7UiaWEAduZmR5D
+QEB9plAYaCUmokukZPggwTsrKvJT/ZsYCvt0J6gaBPiuQf9R/CplHnrer4RVhJs
owgbjF+lc+jPiUdpCzP3oltpWgJUK2lswbfvUqVlP6045mQXIjEsJBHvXl2wJxyp
9Pc0ziGxzLZzH6/kXfyqhskIs5KlylqhWgzGt2Fn+IlH+qC/V4y2FhvlAtHDbQxq
RM5wzb7lvY3/7KgLR2Op/+g/cABXITRn4slQWK1az3v6IRBL/rmQW6zbSX710TNn
Vc49va1sn/Bq0bDPHDbdju/tfxtgCWNp7Hxq/vkOFI/oUhFy0g+CSiQcIV+v1b9v
kBD5lPXXZGH/9cpBDCq6UE9w7Uv99uAERRy2kOtF7VOrTxyFN1siG134kzujj75l
itYrASwO+Xo6GMpA/+q83mASY7WkgIACkyUhr3WOBXFmk7uMtQxYkwIab5clz76h
UopBwLMxN0i63LAsi2QWaacbUo9nwFvPIyECHWHmaWu+26ri88caDRxF8xG1a3Mz
q5ba2UOvQc8+pHYuxJ9BXGxz0rHqRMelwqQsAbS+t60H9T0V+8xA5u0DF9A4p3yf
o/6VHObfwNklxsbZNeSw1BbxyIriVGXDbnDYT5WfyhB4M+CMqJfDGdO/Senu+0ko
NQgQQxTgD4IfH7XUnGI6OeBkFiGnOEoZ4UQ4ufXY3MARAyi0mDeIVxE/uJ537xIQ
6wVcDtXYCd8PBaU/Gq0+DetogrQI/3bzy51cUcQ+oun1iKBrMgyAvbn332eWChuA
CEOPwgMGBsvszJOjLcC2p8J80CaiOCwLJ56fbpRd/pJlII1CQGn2KgwU8G3u6frt
RzSj3zqzW0AvoRXE2vktvikTXmrhl1JMx7x3IMOf9IJGDq5KZF1Dzw/xus6lKKbH
C9cFpIjL+qrjrX94J5UBKpS7ptMcO/uZ6DEPuQ78yb0lb7jKbRNtuCwlu0C7ZiVL
SGeJvpzE5uaYgnqgQbQmGtT7vCCItAzMvs78ZzYtuAFU2R9NWybM2mGq3Bng5ypF
F6HQak3zP18wBsXtRLz2uNXFCsI0ps5Q6uzuOYcYkcG6s0mC5w5fb59LI0FFzlEj
zpZOmhF8KU9LPAYv3lq2tjB9N1G/sW/gqWl75KwRfooWNJpcRK+Hq1n1WzpJgwds
uhaHhSXln6GO43tdCTsvLsCYMCnOKicfQUHPGi944pnmrJCxR2fpfBO/pon8fQd5
frScqIWNwrogOqScasJ24hXAOacyhJ1SEdzIJLBGBMSQJgZvS7R1PTCb8YIqnFg5
TbWeEtMTSdPxmjOTeyq6Zx55igJ9xD3l6Pf4anVj10NtVumeLlj9WBPsFKZfMTBh
g/n76VfTGZ8ZUb7z3psiwvtLDaXrzQ+zvG8aZcjto1Pt6avN9o0KOL78LtESCqYX
fVWEQ02l13LFyE/bLU7BPuTMe1Gr5zQfbpfYRWfY8YcghB80/OYn28ni9GwKJSYq
62eclpWlteDdSfMXZTS3fb1YGbTen6Sg+D8yCAUD9MAR/PfUsybNMvCEIUyfN7Z/
K3T8k5N5EZGLAeVyqmpZgZWNL5zaKhJDOCj/LXweCclTwvqTWzOWqQg/8cRMHusQ
e/w7lFrkkkFCZfdoznHnmb22dU+44OLleYyyF2EuhahRyTbRweqhtE3xhaGUvUIV
5GyFrhdbxTiwZEc0dQ5vf+vf/DOqQBJfb0h9hS8MiG+tJgvFAkBuSa2+QFz98aC3
R6eOIS9k6npWvJ1mIqrpsLoQxfgMCGap/q+3JO2hKh/A4qYrjxkvVQE4fb6f9goS
YvEfoCc7XUcSlDOUHqKxsXSzVTLlom8hgc0p0rMAQCJTT8uEct+QHHQszLXfkeCB
bnB55KGFQLm0GLh/nTf2w148FXKgHKC8gL78AC7nnJ3hqRp/UbXEGtrSi/zwcI/A
zYNFwuyaCUe8TE0HjUg2O/vNdQfpF8eU8S8pieWghh9csJOOzIw8Qbacongy9IrE
c2rK+zRtPfMthC6JiRLEtnYHSDakUrPHazv3qJstRl0u4X+d+FbEAwXlZ/ltks3+
Lljr/0Cq9aVADqe1ePtc58KaLyNPPvnQ1KlR+HMYkN6ZToitbNXzTk/EPw6m33tH
8OrMI22LAiI/JPQuKCf4WfYda9npshgB0Y3Eg3iiRcj7XH6t7N7EomZkvDzVCyfe
dypQcHF56A3NCpx8enf/GihthPXJMlZh4vSh/IUCDt9gsl2vtxjh2AQhZYnQqPEg
FsXUqj725ruaGhLIedHB+JjXI7JwEITJV/pRjxh32Mm9x+60p2QDUTUfLdAbubBv
XzWt1oipt0CpQo99zwf6NA9bxPiY2dHFRJk147Fquta7dvXKwsWuiAbaIKC7uyxk
gTDR7ZcB70KvIew4UdASrDiMY0fixv7Pmpt+zFlDGkuykf2R++zOOjL5fPovHZtK
gg204bu+nls1vwxUkL/MpGDX9Wc88u3mM2wWl7t3kn3ka9NV0HelRjtto68xxDjY
fQf6Virwz9HS3vDiNz7vcVWqyF5582/VYHpm5dZDxvV1iw9EOSFsmeOrn8jaD8vW
V4iVpEF8iBpfg3EWsZ/tD6kVWvG0qKEDCuVfusRU04HtU2QuLebHrBuGVWsROGZE
uVAguyLtGR3396+tK/+lfQ==
`protect end_protected
