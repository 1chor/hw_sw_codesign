-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ZTCOYgNa532gzqvhfVTBZZxZT2TZosUff4bL60UnDswH7htxeC8BTcm9XaH7SfFf
PU6e8AWixACGCA99ebJFVk/lZ9uF9uLlKKEymzzCB7+OKs7tQmjXn9bkKCvQiqfz
dY8zNGOk4V/NYx7FM7xew7KlxRORiJB0QfYrHEEj4Yk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13082)

`protect DATA_BLOCK
M6lmKGBDdmnoJCLCU795ODDrAVfLK5KoC5IRCMCV1Qe5Ftyiu7NfPjW2KLq1u/k2
FcltoGaeApKr1zfmhu7YG5DUtQ2LEJhU3YvRD/yxcu9gJ8qQQ0/gCc39wqxEJV5M
l4SSRjQ6iZIcGhZBRbw9rIc4fBntjrmwHBa81vhswBAUErPK6wnODSUMi3bRlFiz
OZZEbNuAQfL3pyTYJbzf/d2MkWZjGZ71A1c98wHwLftGltfrGkV3bUg5C+JNBp5j
/192mofENCGYojh8BIZJe2ZGqruyD/4quhwfiGmk+cWPzmntjLHWPijWSnAjrv7S
T4kQoeR0NNkpFVVCuKojxAenOiJNl5enUWykKTOIPW1R9S7zDolOGoVx1e3uu+kN
st7/vxv9SHjR3CfbTMQfD3+golNl+Jo79armtwwxdZLPc87/yFolw1Tj1XzECYFA
dwr8JW2yDk4cq/Pc7ykMNNmO6y0O7Fubghiol2EUkRycBnarp3h2E4lYUxpMJSLj
TTOT6Nr93FsCnMPYNoT/Yik1PhS9sLL7fBfuYfb3TF8ke8FSBpczIuC9Vh/ZsAPy
H/R2leBrUvrvXgJB5TXmLHqEEuG/5gLltc2KbbKXyAOqiYigGqRguElwmTRXhkmK
6VfXe8OuInoa0IBwY8lXRNUuuk17p+PEin8akr3UkbAMecF080AtdK74XP5NcdnT
VtU5Vp6x3S3vo1JrDxO/h64xyi1fPaPeghxdoRisAUvObqmjo+YsXwV48Ue7ByYS
UcgtEmDmPgCrmnGT4tj8ubggwXXJUxRHbyayH/20J5r1TkIM3nC4CglHXFgAVvvE
383PY2+kZ3W9D/PYleOlZagOsKXt4a1b6hs9Raba81TD2JBA4juxTQf4kZocr7mm
yVpoTsPJalaaOfMm14s/DqOayUPqwWQh4XrHQxgpUw86Ig1QRWrRTTxH4tBC0xRC
6HmeV7EQhDvzpQTO+rEuxQUggnSBGr6Ctc1DTByKubjjwS1ZymyVlMVybcDGabk7
de3XsUbfG8um2JAgAvhcTHMt8PEvRFBPaKXsqlynZKyTC9sXhKre1XUiTeh6o06a
coIo0YNC+BodqkvXuG7ZX7QWI/Z2ryuHsBLOF5IgaC/QkarELTR7Yb0WD02WyjN0
1xd6z0inyHK1NxFgo7xaKc3+f9MX6WdeQlkcBnG8Q270qex30Brxp2smWVK7g0IB
TESYAvUD4YapI2m/+h4lOs4FjcqlB0gTAwoi087SUJb4XNYzvatuLTMUKmI3Tg0W
4ZLRyuU7unZkXhUrcYVoLPgY76sUUGJp5zoElq0NlE5UtFmrxfbRkxFnwdGdhPNa
4mFKvxMFCDR/62zegJjK6SHLGBhbROD6e4ozxjMNf/3JxotvsfKAQFbkqLZuxxZI
7orBdCxt5IR/X8Bd85rUP4GwxgjzrfJ2ZYLxMsB+5hH5SHqLNG/rgweIVaCgyws/
/I9V+FToNnTKR50cSZ/nMHWMK974uTy9mxw5CeJarsB7jvi+LMtQbsB6tR6KNQdv
Wl/pWmL48MnBP60vEvaFOOBzKI9nSBrtHQS8FIbKMmz2NQLvf7lE+XZhKBVQAZAJ
EgNio3mxdxl6jPBMFZkpgio0a6EA3pnWnArPy8ND0iyPVEof0pj5Qd0JQCvULTMR
rRTqw7VwNUe+zAQ5oEfLEq1QIy3bdlvbJNo0aFvzevBaAribArp5I7tiNQgi3VtX
vzsdjNOF4UtXJi5JJHdJ5R4rNHG3O24jtLHa3rnGHw60Y3a9duHtP7k6uUkNrYUU
HKX6psBjpcemuM57LHPeKUi0MD59kvsL8ghEPtqBrGM6nK89DeC/3CT5bTAqMxXU
lR1MZ09N+FCwK6Gqfl63sN+XI5xQ2ELTYsZZU1d5LMcBVP8C6dL3QCeUYDh12Eog
6WaCieCVmsyZq6waOZc2WxjZnUfiqQa34gyPg8dD+vT2yGlXJyx9TKxvw522fFz8
UAjCv5Xhsnj9vDD5ve8osbAPpjg/SfOmi1EvrRW8MIb355rLc+FWsxt+PQkvN/8S
VMksDB7GQ8ZWxCfHml7SWX8bsmRUi8CeUlz0+OxfeCsRlNxxR7zULS499wJRfxA3
2Sj2fr5CPdM6Y8nPQBjI1ookcQsupUp6hvB1gsCglUZJG/4lhHhz5on4GqJVStOj
wv91Nw0YLU21zr2xQiYJTjiuKQydnXLDH7kf/IUPq2M+upPwBXHj9bOLQR6VAaNG
5vhLODplsIaDBwaz/V78udROxUnpM9IENru8ZVeW53vTe9c0LxcuZp7gGXAzFUz8
Gfzr9uzaSa/FZrD8YFj9XWIANzlEgP3AD/OBzv/AqvFqBU2nlg741TjtcfyAxbO1
itW65iZ6WqzzvCRIv/ayl1MpVRugqj9hovd78k0kVejkzl9fQG5WgWRhR4oM1Mtw
VN0pbcL+13MvKD4FC48B7Q8pGMYPA+a2qcFe8PGopzCbRv7V1Ojxhogtv7i+AUgE
703BfLDLCVyoHsqyyF0WgAJAv/D1QqazY1SGo7oVW6Y5y8K0DWpKytmVyu+jlNi/
lJqffiAZpZFa+PkYq2P5lOWT4+C/JxZQgkUwS4mCntrlzh4geNluIq8bgl4uQ8bG
U7haMi/xGnf5BzoDut83cAN2fg68rNz4U3e4qlQQF9ZRnYXexZG5nEhjG0OOrw8O
DPX3PHToD9yQk50uuWehthhidpIC7e7jb4LgdHluK6fxZpngcCf8LxA+W70MUS2Q
79vDRmC+x7+P05924nhlvPyASyFd4VIRyRpwTri1yk6OgSF6m0EdlZYYWO0sOwjh
ibKf19+BAgn9a8NGLPVfkSfYrTEOFSfBKbX3Q3LabgGY7xS1tXCxbD8g1A+sYKeP
V2G2x14YfR6sOumC9jeR655F+LEzg+nS1kSle5FSvAyVf+X3PAW2kNIUPtkGmSUL
IsVWskIqbviPByuRjTE/5mSNydCz+z8/wLqCO7uLdbTKvlQBXYsJ7Xix8Jb1ZBMm
p2lBEdcaoT8RnqLRG9mMd30YxzZFdXk9hyKuRhorA3Dk3+CbLH+GlDvHrwUhu8Jz
PVUIpyMSt9ysiOWJuxZi5a/awFUfpO5ylz3gWRCbgLCtwyXjujvBha9MmvrAigDj
cOzj5nsVMlfse6OPIF7+feeMAIs+1XKQlbppf/VlXM4nRtJhUehArEndJYHqLVNI
fs/ORtO688D8+PnLPualmDAg2mj111cseeyalpEorrCsT5OhX6EX27gJ+3TO/IIL
QdUWB2GSunu6SmHG3GoJ5sU+G2Dj7226flw/dj+jJgdiTqTLdClOvnNTJxUG+NTN
pWIVx8Ib+Vx5nyG6uB5KPSnG8R8o6PnCwVl2vdlh4IOINHQeb2LyLqGGzZeJhRm9
8mCSdRketvEIidjz1+DMY31Suph/PNonN2QZxtZZFNivKOdxMSiRmH6fQs9PlJhL
xeI1n912lRPuZ/mcVzuhHeuFbSzOgfN0bNN+NyabKABAjhK+3TZ3iPX+hiKsPzqj
lJwA8bNmWaJ9E0tQVWv3rMKN2GolYPIqSE1Y+EQhJZDpBzynA0FgHF23fM0l2wLE
Czwk25nl5thrxV1vKiiG64KFUa1TQOPFwZS15dzMC+3KwEVvPDt9w9uQBCInqOI5
gxvvkkJeBBIf8fQug1UCKVFhmVzAx7oAye4ZYF7QBuMTg3DWlMQttoQjOj11ekVr
CzM6YW/uba9d1Hy8V+kP6/lPvbG/foE2V5fHDbylZ0T/maJIq1LC9dXtojTtF75C
tW5xSYxAUucIDpE23erNS2NppmC/zK0HJPMfrRjYG9yZR0xasdhmxpWykiUea2jY
bKPQC3lPELdO7Hvqvl/TLW0d3SgXjy1l4gR5m9WNHymdRqfDXYPmqEqsuCy3T6X/
JjgeAHSFKqk7WBZvpl2nwybm9ZChGWaIw8P+yYZ3q7f0waSiLM+oJFFaYFg4+23U
H8iajvTspCmkjm0DO9m6upn85MmfgWIyvImFPAZ5MVYJopJAewjHuCaeczkAUgLH
o0X8fUI797rKH9OHQOmeDSpBO4rF9B0UkwZT6j7Gqox9dqylFtciy78hAu1KXQI6
BHkp3A+UPPXMsCYEVwfePiUToy/vibkgZpZyAPu+RzGbDn1txF/XVCux/OkgDWNs
yKguJZ9HCm3xPaBwh4tJB74HpOo+vSU42oTdo3d1/X4QU57M06He2pEwR5eP5pKx
LnbPOeodYhhgvIfzmV7bBYXALJ9GEQ6xW2rrh+26+eIMf5hqohcYNDMZ2kkoWC3x
9nkwG13NaAfPfhohH5SWanisejY2fuohD/2mcilwzJu3annr/GO6RppbzoLOd2pE
B0Oidk81RpeSyxT1KAJqS2AVDjG4MwYlBn5CmcuJnohlY+mkjFcU/U/TQM7PiD7b
JPbeTNCIngHCF38AMXQK6nRzFGf42g04zcEkUUgcHIEjXaHchgFU/OhZY075j09N
9KZx1fd9ahXBzjTEHOcYgjxvMDskGYnaTqnD/OfRBjzZB2W/q5K7zUkea6XRL3Zt
BCyqIzjyEt4VLtzxBTRq494MyZzCi53khKvfPxsdgCnzP1rGeV858TGLLna9AW5V
09817Qoto0BvBHEP/aFlQi3IJXA3Nn6Bn9lVSjQpRZc8spbzgHcQHAx30cyktZqE
H9a84yZpo5yIURAjmJmP1yYva46JmRwUI5T9obBbeKpttWAb1qb2HwWbLExwZnjS
9NQTVMjUqBTCpEYSd2b2HNtl62g53pi4mMfjsMcTBzFiIta29gZzgvni84JozEQa
5D8ffaNs8F1BXsGkiHKlI6t/vD9hCpwj2Z8E9xHuVGopdmNw65AhZ0qHK7icsvCR
iymvNWncMG6tt4IuQS5zlEko6f77ums3okt5USP+VXqnFSRdiRqoYDtq6Gto9HMl
OSMbHEykDr/jvImDPycCHXTwU1qxMYT2cekIVyOWF9qFFHh9Eh3OXzV2qcJfw/QD
Q8NUmrj6BUfC4IUsQLrM6E5Pwe3pMfffcCVFrhTq2AekuNZgpq/wpaMVrPSNKU6U
tpj1VTw3trbPcCATn83bmnjalj+9dZ2zkGy7jgao6yUhCrhiBopEGS7jtStyCD+H
rCkq4NkC3xSvVYpmwoVWeOoLpuygfPTk60nStRbM92QuqfPb+zp4t7CPo0qqJkSk
J8rBTjEOH0KFPTPy2oQQYWR4i9i0gzz513eqjvwTU3vbekkPzsb7Kr6hYLLnzKY1
7KfGQ+V6054T+QeR3byOVOs9o0cJ5QHDyLHtuvxxlOkagRR+bFVoNwYq5IXP5Vuq
3SpFLiCWAH0cgkStZIFiRMAJKkWQPgz+95uOAkyZd99zvhCyWTI462FEMp4xF4bT
Bx8xkYphajUBXTyzj1dgJQSS1USnJNGDThFPjhYjA5Z1bCBky447AXlsNjvpDhMP
kxz4ZlQO6mXuJ0DhNI8NYXxz9tVIT2C7JBsKdUWjIy2k4CN/30ogkfz/5hfQn/ZV
oKyrge3AovIr2Nf7R1bmnvrUYTBE3zz4AiPxGQygCfMUouAJ/vWAys4I+5gU+rPo
VBvzWBfavlCSQcrNhQnWprUoU/FeRQHOYF9P9Ya3Xi+WJ9mOjT4Ar1ZoukLICb0O
/2Nli/agN3ROEhiaiiKlOb9egFAbXpT/Q+OEJEPggdb5zbWwvFPNs/AlkRmftfPV
Yuc+V0UT/SZL3B4tnmu1afaR0REgt3wYSGDzzhdThIo+gen72DLGepxC6J5+Od6s
lJCuM5vcljmahK524x5V7L9KeIjE/MH7zvNMs6gieHLJKwbNTgiXn44Yait3DXnR
QKqIIiceS0L1hitip3T6y/w75hVLRqfLTNAF6bZH5yrMEcqE7X5iKVGb0SbuVXVR
L/p5Q9r73Jn3pvpLThQydHbqbdrKiHh+TSU/S8/jSZbc8dPCwmN8qg40Uvpym1SN
gXKPZ5HVUO8rHJWdetdzLRhBuZ1Cz6Nh83+dXx3BYUo48qSqFAmTGvbu2afQum69
WziqOlEXi/Y0beKEpQ+0THsQ8mUnRUtsoBnW1ATbamUbz1NrAejrj2eFDsWy3aMv
wjGP5SCfT662nSGjN7o8GEBxNzOpGQ+xgO9kjTb/vwHu5lVH4/e9SmjXmd826345
h1u9HXNhXyFtclGxmOCYaoHn0skH5HWWlzLqVMKVEfnFW534d+I5xWQd6UaclaYW
4JRxe2b5AcgFyyKMcVFJc8NMlC0spV/SsAtC9lwR5sKInECd9uTyZr/KZm+07qun
z4V6cs4OUSsDnKUf1yeVpDINAG0d90eC0T5d8K6lqCDf10VvC5YoZX2xFz7r7NJ/
p5PgMP46Ne0tiap5KChDkXe0SJb9LNmeQPXIuTLDM7vTy1eOoh59/ps6AsUxbuHf
uIKoaw7/xXusJ2tKpJmnMasSArMapbf6p0Wwm1ZiA1dx0HJZglJpxE6SMoJUmwR/
XrFq6679ZSfyCeDZE9aeBvBA601Om8BnLiGWsBOpEkmmNnT3aRe+xoiuMaTmMiq9
8ffE8zXHpBYYusQ65RofjHbwyaHmXpjlNb+rqFWW7JIOQQeY12GihdPhPhzE9zMe
PaxcPXcHquGDwdcXUdp1XybeWLVvQe5bZbbfnAN7TeVGyDuGHhugXleKUW9MA+yR
guAoXhBAzAvHq2ittbGALV+MLP0ntgX04Iid8+JfZhynD/XhUnKF/Jw1E2x6zdpw
B7c7rN6DMXII3dLX7L+VNpyntd1nMYj3ztt8j6uvmN4IrcJVnaWWKWM42e8Vei+Q
NVQwpEgNOnpTjUHW4vOuCI9GZlR4R4CmtZ0n9Y9ErcDr/gJdur5rZ7iX2FTwg+8v
Q3BTJl7OkoBI2EaMMods5OV4J3E0NjHUAOOhVbzWvxdtx1AFohPKEseXAtU1F1vG
nGw6B10ynW4wYc9GtBM08uI1CvSRPxAl/dT6P/9ORNy7JnujEGXcRdDJsG+mbNsX
bC4l65KoMdVg5QTMNic6LkPK2uBxHSaWrJoBBTD4S1EJRamMEHi2sFn9yoMGgg1Y
AWyRKENjmdwQcKZBLP4DrDMI2nGaTRbva66rWLQ8dewj9a4sH84p91B3yKtmUw3u
0TBTnBLGouQWC49JIt6v1Ce26fB1rNjZ6p4xGQB4h+x0JJgc0EwWVjp3myqri3+J
gD0e/Wud1OT+xSVtzsr0TK0fxCFnSYZ372lJj2GskxbxTELUVYgNXW0DpzMoHWIs
Ehfn+IjM3DYGStgDRIvOS5JhX695zuEBTNtE6vdHhrm8x1qZ1hu1DFBMne8pNVus
aVL1vnq7oaCBYaCBTAlvwCnqykR3OVDmtspPuNN8SmE622Y72HeCT/M2ld4UWta3
uQBG85xYwueAB/CZA4Mhn132pw8a+vxGVqNBGHrg1HTEPXQwR/TJmUe+CC3SBarc
2UghI1nfcSTMSDx1BbXnWDCiGNXJBc5/PlLxVin29W1yrzKEqsuR/OZJWjYGV/Zu
tnK+rDNcU1CkGPcH7mbWX1ePYST36jgelxhvRtP+DorQ9Eq/Q684Ekr20a5xolYF
xW7Xt9zWj5LeCB7RYzEBDw1+3h3aAHfACZVkxAYV+p+Eld+wR3z+0UCUrsOHc5yi
a3w4yimQ0/RZONYJW+qi1uVV42Ka5F56/SEruB9mNvQeFGmlGuiBNz0g0cwE+rg9
yhE78Vw+ucHJPjhFTsUk79AiV/PQXS7bgTQrmQD5j3sDF/EM+pJf8gDeLmjMa2vA
U/REZYWUraO7RzQF5mD+N7/MN1yxv1JwklWpBR/+TqooAizS1ZptpsHBSucgIjJ0
+wbqcbdT7PmaNrGqXP6uqy/k8ey4eRHxkdmMl4cPgZidtLQ8AwBIqeLdnQPX2Jqz
+c5kaewCZzj8Te4C+l7bKJeoI4EzAhLYEtBT/wWjQJmICqnwfjnwU2HHPZLNlycj
ZkVCtSBBdhLqwIrrsQxxNxenxKxjb8DDqzcVbXAWlkrxzLnObKTuEiKEF8+0nOrH
eCFOghQEKh6i+x8n+Fl2dCZWleu5NxFUx0iJ4LwLwuRuM1dUObmEWoD8A9xUocga
ZpeK9WRSBQ7VU6BKzIcOjrzZ9qpVDvkvL92vFrUeRnrwXubf0OgTpKru4eHThHd1
qLyCInRMtVkCHLrxqQVIeIf6EyyeKUNcIClrJNd8e2zvVppTJMpfAi3+dq0f8Ksn
HYDIQDq1mk9EUjAMPkT3pkV7AyM/hTN85IAFV1o7uvfewBIXSjAJxhqFiUyVRdFc
MYPkjrhqaP97x42Jpto3vB3+Y6ogon16YYovwiLTK3mwgJOXuZBNn2v3UQlJgCvU
wHYBUfiOze0e1NdiqWYPlyoHfPE0QjgoQnjQv8YhhWR03Y7p0I0IUcyC3Ddq8dXh
a+wMc7vz4dbtaKM5Iujk6heSP02koSFXM7glg91iSauTb2UrNp5YZrtqgCdZJLrZ
kV0UxsytQjxMvr5XrKl6yBFb2vmTcJZ3nwQuv9gqhSWQksASTnW5J3UAblyW06tf
o+RIuENojGCQnozNvJcjtCEnxaKCQTBHrlpl/SOJUkLVr1JCS7rRAuGvZo+hW170
BPWAIYmP1b5FqAmqTBc/AGq9McVOBibTCQEL/8etbDFbmHPYBCeOcVqrK1Kr9S04
kVNhNqjpdaCQanQwq65o11bIwY9+LDgpdabmZ72A0vSaervzaqi2jSmUp/UxofcX
UJpw1MeFX3E4VETjA3/FU8pjz2fKW8uunQA4JiwEojFZ6L/i9lUB0AKoi+VquM5W
z3wiWIQ7MXUsXLj5GwtyPjGx92W48HWzR4T1QGmCTANTOrpwYmQQLuoWMjWQfNJK
wWHUAq62yLXYYGKxUUY6rxJ+4MwaQHdaVlQ72JegqfaoySDWrBu7lw+l7WOIzLVb
tuobC2+a4xoPxP5TL+nW+WJEl/FlcI/XGXeClR1XCnfZKBUaSbnjvOdaj/78Ax0o
LvMO/rLLoiYH6oIJargpsmAP5Vn5140XT24KjtUUYiXGAvDpt/zYLURZspuTr5hw
DpCVHXSxxr6h/Tg0zrg/3plIHUxDqTxxGBDFVCM48SoeN2DKlf66WaR1G1I/I2DD
VaPJ23DKnV5LK/qXhrRQCZvvBn2H2WlqF398C42MGDQ99R8jjQM8MBFkH3ENjQG6
bqSiyFY/JIi464tcDpu8uPI9cstqSCigKL5J4nP/8AV047/zTuTKqiklE4uCNYmd
0QMxLBRuWYOEPUjEcIJTBJOD3ulM2cLf2ioI3kVypl6rqIv/Aa1frT0xGlelSvde
y0CVk/E6+Dj8FxJ5iRsmndTPWGzXoUmhPt3GMs/eXsY6uZspVNQsbKhW9YUcY1kK
lMmwsTccsuNhyGUSLD2GL79PfHEqdlp0jHCZOsES44A81/p/8Rf71avwZ2TxBlPo
kH6MYxnVJ7/qXseYH+TwH1MsFfVDG4+OJQKNMdnwnZ5b0BycZ3BmGWyID/k1oExU
1Xa78DK6NbOlVu3gU/65NrpmzzHSHhPSlUb3EDa409hU5zXetzsvrNK7w6gE6vdf
iEj+imjx48L7bhMp5Ub+d8kSWEJaH8TXwCbWNdJePEjvzZoIMZGWA1867sIlFqYj
UgbN6Vymv7zRl/hFLUBCO0bD/K4R8i+CiTnBc0Wj5NvrPY6vo4guvfUc4ShqEqFX
Lo4x7YOoTBgXQgim0ciKSO6Mtp3yPLcBf1VRm1DIR2m4NExnDzCJivzuhc63cq0S
FpmdvFo9AEQuEO1ZHSIrGcOpI23vswKCWo7dYSiC8XWfR4DHfg7+9BdvrJz1BezK
CosH3ggDWkkh6EVDoJzcoA7Ynb6ZUB9HwHNLtoedQRqYukAkIriZUgDNOT02m8j5
MsoYloXuh4KvJa5WkeieQhWLoISYMF6id3QhrhwCmM/Vfi2fMKBjHLdh4+EfgGxV
VFPJSjSOtDfclA7lrB6ZLzAKcUZlleH+TReK7lE34aYutvFqx7SBJR8+0XYcvTAz
vVDQ8WHiTxcDvCr472X/+IZ0XpMN31jjzPsWh7aHJdKZeDKxzWtCWO+COgcBARmN
l2fNFvLq6U2v8wUCMwvhxfiDIAOF1GqOAG1ZzcBRDe4FVo4R1ACEoyZk7EiMXixK
7nvV1wXD1hpzUZkVpH/otsx8SPlV3N9V5N472WZZmA8W7JMweKfVfKAvQgBIFlXa
iWLb+rpTwh1sqr3/QJcpLI2Hs/JlKDbwU21kMsQgBctspFuokBbba0ZNn503glpO
K/WPH9VsbzPyfprLkzGViFiS86JPNIOEcUbnNJ1a39hWL3e8mbixDM4sxsMhxUbB
XzpiK0T067OSvyWgeAvcCn1k9JwhMGrer2ZB2Rwcvz3xgfcP5PALL0Ad+x7ty/sY
e+EY5pJG9cE2hrnyE8ePjTQMrtJalT5mAwrYg/aTzV9hJDZzZxzEqY94xPqAT/MK
X3k3SxwTiU1Jjcwt3mcwebPCK6gsjCYM/vYkFDSYnUyYU3in26pnVQemEpXUoYx3
Y/aeeVj9TAjaKFSIVVKKVla6kbXHlewuo6Tgse1bZuKh2WAsdnlOH9YvkOylk570
7fQ5Tra9eT2V3MHXBm0jpR77cselV5sejD8Zoi+gfzB2kpl29Sak21S/r66M0hUx
6sPo69RjPtiqNnCKbRbuEPxcbAUpylgYDcljcNlBBxUGIigDClZdnnIlHYFrCS5V
aJuXuGdXmm3j6ajB7uE+vbLtOjce9f0Ru/gKLU3V0H6wms+lUjOE4fIj2Q45Ul2P
dw26F+Z8w+i7frKNcl3581vghhToUo5LOztWNl/JrZ+W9AE8agEYYBLkZRcpl+Oj
B8WILkOZupc9fepn5z98Nkg66MAMP7mdLSjNgMd4or9wW/otRISvUNUw4STk2tRq
JWUB4XFDwcyK+Cvouosrmh9Us+OiGFK5Cc1H0VznpB7fk4yVzFeWkVZMp+xSHhvQ
ORpHOTbsV4RJq4FH2oHB9kDLOe4H7zPVxK9ROiuENCrGTDDCrxmHk01pAWYxaZey
WXmLP4C0Xi8t43OZAMfbdBiv4KV3dCbLnwMs85Tfh3xgUDzqY+1TFWwt4ah1WtS3
/ARzQ9Yv+5nX9LLOD+lcAM55tFHEJNhkXiG0127boR2u4AKV/7r9IemA1RomRyYu
nws34bguYJMKLTPyWRexSYIYrwTvtmIV6/vwOALoJOQYtFLK2Vyw+Ro7aTmyqGwq
Fbs7hhud3vj/Jce8w+SfStAmO6qryC76WaWqXhxfUTyHh/xeFm4ViYcIuIz8cnb1
MuldyMU7658/wLTI7Asv1WMjn7KRdf34cdaGEnLq38ZcBdDvAcwCFLlD33vx8fXS
7KN9+6M+KxEGsDNw0KSXAd3Y/3fRX6f5bII8T14VE6AccRJ3jQvk5krq4t0OdaJM
r+7TqowFczPQBu+WbOejFmq7KePenUqx5Vt57nz+Q4ZGyiy+FjKCZdKuzoFxjEJP
RyJNG0mSWgcykRjdLOdZ9hOjk+kmxeULKWek5WwVvqUMNZEV7Uo9ja8SCzVnduDN
eyTB2ImExTXFt5w4kj+DAJOxGdJCpRK19UHyutJ2uOnM7CCFbP0ZN4acM6Ghzod3
Xdna2RlZOBfcaYGdP4W7u5+8pf2OtvsLVU8wI/D/jx5eug28SU4QAxUGiRJylPeq
cFEp45MmVTVu/dRYVxhMhvGdAnwQRitFUQnpaM+ONn1hSPJypMEsNk3otY2KcWUr
N9Qq/KunoyXFQK695WhLsOGiIqm+ODwppDJHcIM7YkdpPLiadDg1qDYw9xXAbcvn
LN4+BYI72PhzB9DbesqqeuEuxrAeorQkJjm6DcYu/O0/SaYDsPd/YRby6tKHHxEC
dgwRBjF0JY/yG0l0GPjfzc3o20oNEtYyEZK1wJZRLI9//QZiw1O6byTF2jkTdTIW
WmXSNbroHdk6TSI0/G1QiUGQNgLkNYkL9/BFuDxofXRhAEMc6YkEoHoQccBeF1qi
ocmsAU+RiNDqCxQU7fbrPEqoIVcIuyjH+RZgRCXqQUlDNjwRHHJU3TEZ5aT3Oohu
XuIFKv3LyEihCmgKyDIlvkW+E1BzEza0wzJOnzP8SfouKeHQfOICjLfPO2TgHmCF
MtqNE5AIskTQeIeh4dyAmoMdVu7BmVr+LRcMSRv/IGgnl7OsOmJFX+w4QBgiANdw
AgKtzJBzmj8Qwt+O5hmuLaRGjIoTOMcz2YzI6qQOnCHuY9D9NTH19dziqfX2iPNi
uPXJuakmYEPoDX7UlHU4Jol0HRPz3XTBc1Qb0lm7HOz7OLvj6ebi6Ranj1iGo/02
hauzC3F6/R3BA9Yc0B50AOaCfzA1ybom7busuYre/oLLrTx49kZKMU8Wv0qYeP2e
3OnVgbRLMAO6IZHAumf14CF3BSElrhGNP/ecH1SW+X5JhUpgS8D9srcj/0DODFSB
IbmzuqhDJZ7a0/dEKPBhWPtFK3WXRGYEhqf4vFIc1loAiqdQoqQor6PfRfsl42M6
XtDkupFz4nyc6hwKNXqZEfWCI+wY/EFC27SBHezyuy9L/V6QbE6BSVTFCA2iBU7y
Nah9IZOuI6tLSbukh5b6wK0Jdi8kXO7abXR4pKIAmR0l5j+EuTFTCfXXo/1OXWs0
7aRgQ78POhTBQnSVUNhiKu5vHZMwOoWfL6dsifR+oq2mMnd07Md2JzNr4Zv8XMh+
jQ8OEYcf6p6b4/w+lli67BFy9xvbRjqxc0mrDC/8+zMa0E6XYRXXw1PRqytdByfx
IdMhzBjvF43qZOggjmv7fZjwwH+qOFRiIQFzmk+mupITV5Eb4hqtWSgnPXDfkcRv
HA1F34nn/yRwtFtm/OIhssE3eABcXyZ+/OzVfS4Rk41GDoOW4YR+ipZcH+/C9lFU
INWBWw1OOGwGF0HZnuU4jat9hvoc4U2ig9RuXx1ZxYbUcjnwvJi/pDgd1PDDPOGK
h430YccKGEf5AHdR8XP3zk1vvgdQAGfy4AGodd9n30Kz9F6INLVilxcLAZpVQqpO
e92idcFbxppqddXfeB8NpR9PnFRPC9xYTzZEjz1Bx4cunSXVb2wutN8i7ROrnR9M
eUZwldPOyvYvKrbeZh0S64KKlermZ/L0xDTVGVPVVxPLMU+dGCeXNP5KXVEOqnle
TlJgTNnVT/HQis2zgddQUyGLYQFRyRwDP8To7IVN9ko5bG6f8HFuAoP5N3plx37j
/r2hV3+WfGUUT1uhmhsHqUPVdXSpe0vNuKOI4TJIaU8VIY27pZIiXQpR8hZsVzuh
2cVPXhqO6+/GtQLx/GSU7u1kwH2X20gRqgAFOeaGqJL+vYxoatMiXWWq2xjc7vf1
JXPnmmzbT1d8+XUQGDl7QGemcDNet38WPDbaW7iV6h53A/J+rVI0Wxj/0e4GArc4
kFqOm4fH6BbfrElvwZdOGAGeHF3ZhmPeonffsZ3N5wIsugD7udo+vP1bSAuWGPmW
kIpQZHckXuX95+2evO7fuhM6YGYiPDXeDGKVoUo2fPyvf1EwjIP9NKWzSx8qxttu
54I8V83OfN7iR/UkQt3IV9ZF3T48PrtDYcZEmRg32Dl4kaeJALbm9nTmixJVja+B
OCTxIVOvtJ+N1Mngvkc7jo+jYddyfnIGG3oZ+Q6G1Mg1SXNN5+tbC45YN7WWzeqV
xKqqnfQyLBzEjUci+xpu6g13YuBFn6QLk/+FeEPqgodWhsn3Nvi9opYU7jVSoasA
rppSnOzt6F7SAdaWtL9sOSStX+UYVV499IZY0vhIkB0pGcDE10xdQsaHnnqznt3P
8sH1ONSmHhO3BNvzM+Cr7AyDZGgZt+MnRF497gtKIAzPwzyfP4jCMKpdpqQ9Hgc9
Ak6neHdeIXqLrLNK0LBkygy+A+cbhuVJ6BEKVeM+v4cpjcZCKBcqd3ANAJlibuFu
Q/4YaFXLDko6Zz41L/dS00tyzzeijaKtyWaZBJ074r3YgBoSSSs9VcYFzLdWWsCO
puWyauvsl10CPDC9rCrR+DGuKfSeoE3Jh/+OavGJUEQ/Z2O60G/NmuUQn0y7pGMk
zFBPFbMzopXYkRz50h6FcY4LkaMPPJUehQ4HNMiQDB3YWlcxbxynSqNdoR2WzWg0
K9hiQbx3TZ7YhwssifuO62vbQJ1JHf9J8hbseJexIKpW9YJY1gTsyVubmSdO/pGE
Yoh7NxXwd/eczSWDAWsW5POPk087qft8fO4xdoLScmfk5gnEr32Fxa9TR++0pVzt
1SFpxTlTS9qnossqRM5sJqrOM+5DHsmBzhdett6bhXbaDSKalq+ea7nAinCzgvJL
b14nePdf2f1A+oJct6Kywx+A0KUwhUZLo0f3aXbp0d7ED2iUUQ5XKKBZaikAxfsv
DftEp/zwYTy/guoQaLTtjN1r7W9pnGpdtceJAqDKd/EWcNW2++ijcqKcOQ9EbxV2
O5qggL6SHNDBtrf/3za2Nrc8t+SGffYAg6eYDql1bsFAnpDTb2uWPMzdf3v+GagL
7nmG9NHyZXn6xwp9N93JzKRj+a5JaOsHSUa2ohrlpk7NCPFp6++vHAh6DyovL6mD
OR8uwp5q55UABOoUI/QqyjDRR+rrF+esO+HJzidbZHau14+mfytc5s88fsTlBLwa
SrBK+bs78FJDMfu4UQXfVwehd3RIoOB3Rd1rVX4abp+fCmR6ATb/PIYVVsiFzy8C
2v12lNqDm6/h0BWmqun0g4VE9dPLKzqovIxHqw8UvMquTCdxK5rFK2VD4xy1nReK
y1DtV8p/6nAPfRsjY/b84dhNQ80ron0ZQghrmpNJ/KSUH8WnsS/gcKLitW348qnu
bqqYxBSj807nBOr8iSXnpOUdaxtypSeNRI5IZN3mW+gDepoO1QlHcvObGsgCexrc
5SeIwgOl/LColzBV9+KT5JCN3i4zF7rUcOFCJMtHbDg2s5Fh2D6SgGMhsE0auUTo
V07/J7t2slyQjdlVEALskM643lkG5ImPp18PtItmlwyjPOnqZSoJk57Mn0xO04E9
3yVhBNNpUzNKWKRFo4S/CanlVBxx0owVdvs0LxYX0ahc0+QxAff7TyZwLTYNuT60
f6FePYNHXYBQOtoQpGZz36gPDPWeOhZiTbPxaMjAWq6Bp969RqcdHSoPzwSLq55g
NMatkOoCvd6iTiFl6tCuNUbTeAgrNoOzHdeNNxJ9oye4KBiVA9LUSV6P2UVkY7Od
MCZ1nBr1Wjh+l2w+Fv/FKv+hCatD7WzvFJxcL2CCCiJYwJlju1fJCOdaOUbD83C8
2Z3bqekorVXNc6U8flQBCSDtljw8VTpPufxgZ750fQqbkIwZbLenrg6ocx/zvFmW
3gKKVJ5kvTvxIWXoDagHFTEMl06+7pxi1j+B7dFswBtGOeD1hVJGLlPs532ojQ3b
FKKMtO/BTE0YSS8oVaALar0wwcV4u6S51D0IepTGRGi7yKbO+2udUZFQB61s9j7K
m1gLkV+QiAQEAhEUwb9dytjy4vf+UNClawKbbIOMOGaXOYEKFkt8/4G4MmbjzNR3
72tUSVZsZzEx6MsGmjyj8Ew+0T6o3ZCfodLbpbrJ0XAGX1UNCjk/PuomDs6zSxEK
QHORNUHxTlmNx+79qtsbXS9ZUURBudeaT327dos3FFlQCNu7YQ0n1hyNvu1GURCM
vcYrN5cizJN0Zy23kJlprDo8YK5Kqe1nCDqhN+tPOgAjZI49ZCWmH+kBaEpvmHI4
b7mnyBEZ/75mMq/Ps1xhIddkNz6JyKngL7PAZQ4YLGtbR8xB6k0zPwb+bbXdpHIq
gLVYoLtMec73JtFbx6oCLxJ+LdY8sn5EaN7SClCXbkWiwYEQfSOUKv/aimzhSCgh
BFGFI0lEriL1mECL9+182q+twhb66lY9LMrZI+s6yodwNbJ4T6fy4YiAcFDuiiYy
X4tBCNmnQh1i2vEQb0+u8YKvfv4nnXkSKv/hnh2Rk+HDmiLXdHiWiHFpSYYs4VLE
5kKP6bBiEmi6rc7Gjg487BGHnXDLrSJDzo6s1HM5KoRM/eL4dv0LIHFsb/3NTePU
yZjxeIDMMArCJYQZloc3ui+8/GfgrB51Ji1YdPPht00MTbsKll9lHItS//IXSkyO
H4iIiT0xwJ0NLRISNzNofKNJxkMOKDrE8g3hOFOs1yM14KEu2RHD0P62UZhz8BSa
VGKEuWDrXgRALJ33NXUGqlc+1WvRleNVhZdyyDwx0OltfoCOQDfKqSjuudEXnZwT
qRwB0K7mjxpcv5O/tv3OJf3ddEsidK4QmuL5xQZR3e7W16weSOUMfGcLVh5Sf/Of
+6oyT3uST6I/SjnmBJDoEeie1Qym46Sxg0sV7A4onyfNc3eXijD16eE6bHbpulsf
rG1byi9HtmmpeVd1Pjv++GNg3YaRJosu+SkK3LJfN7CYLVAxzN49bNWOWNqT3Xfr
46VLdB/6JK6TNhUDzt8jKIcBIbR8FPBHd7QWQxH7BqFTjTfdR8ltDIMhcqKbEZZ6
VZ25tXtoMQLx360k0OHU5/tu6mDu6FLZPP/dDtCAxRkP4bcECQ+vxWY/f/NdvPy8
4dgdfpIfCBs8uispS2FcxlY3hMNu/Cs77PDefPI5hnCN9diXVIBzI5+VpUbeOqhF
2F3IGK4hdURgiOw02LUgj3a8ldYictsZXrGkfG65BBocJ+IpgbZOFdUa5VXwK/pD
pNxSeqRqygx9Oh2EB1vfKGYGQEkbpVQ6kZ8eona9gl+04OJG5ySv5mQHaLfPLfIH
oLwuFEBjX3IbRSEULeiWfqiI8KCnvkolWO3Npnf7zbau+2evHXEbT4LtNI/Mjybb
YX1ED2S64T53u5Ejype/heHC+S8kDqimSeT3PR64ls8Z6DUINSAhMY1QQla9UC4b
tX5psm+0q54TAcVNl8GJQdGCpOIhatYC6dU7eqz2qh5NzC3ptTtqcQkWDPtFTlTT
H7zD1SAmNHnq7sfYHrEVjt8pWywNS9y4XRZw8PquUg+WJ/9JkB3nN0eeb5gYxtXe
aI46GGMF3FNhl20Cx8pNK9biSnwHW6ASbbmGLhUJzPWWc3hm8iTcgxOrbuXw5Xuc
Hbmr2gyz7kwKk1NG57UGnLYW25h8tuenSpfGZFwSvzJ7mQZgzsynx62Uh+5lnVhq
yRsohgrZq0QcXR8nsEUwznKCf3/cJooLPtiMCRykv2v671vm9072gvKnQXNBuUIS
XEvxpRQUWZ7mdkE+UzNfNyHDllmofHsP/pvdw4p1UUe8nNzfiwDTZpJx42eUYV7v
ul4XwJilHShPHLCQG1i4DkD65UBdNj2dQA9PFvvbBufouemrhJ2Fq/U3Nv7wtLmh
YhQjMHtM6h0uVM+PnLrxfVzArvf6dJ+582yFtstUryFiDKboZOtgda28gcR0he9i
JJXN+EUVVGe7N5cg6EmJDR9gqYm00yk1+Rc1XufQP+O3nQIlRKvUJyD+QxdiBS2E
HjQYwBGjwAPT2tLEgqk3/Y5DzThY8i/pRFpnQbExdbs5IH04m9rkyRoL4DZxAD4t
`protect END_PROTECTED