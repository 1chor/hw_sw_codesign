-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
eriXYth4/yDuWh3dISzNU7JDxfmj33lzwXxxJM8isccD+n3DJwRfErzV2zKYb90H
g6HJ3oFS//iHi9JkwdPKCT1ytleJ+N85axopk1TImfP917qqh9hrHluMuoMFLa0t
AI7uI4LVvfs5oQ0GofUNy5JlwkeO55XA3YcwYBTTVfQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7517)

`protect DATA_BLOCK
W/WPj2SoWEHt50jbl0K5aCuCrQkfysS2g1uHaifYQsaYlihoJeXA1rBe4uYL/CMV
zdEkwL4gZIRcQq+ePrS8DuTzS/L6iILqgmnb91qMwjtYqeAtC0vVkoqqKpq5Aud6
dlLTAbSCDa4M4/ndfxiwvi1j9xKqcG771quzQfZCXhVphjzexlSlbQoRbCgkecxZ
WUc7WPs/PzAfclUich/Y7XLN9+p/XwgMOApZXqL5x0Q7dmCgeCOPDa8JLyD8+Une
2usSpW8oylnrGvfjuhEGLWLRzlGNEJ6fd5aDeyVnGGe9xZiZGPthadVkR9hTEjjh
RBaMtYSr2whOo0VzIiMz8PpvAKCj8FjN6fsczdsLmTdwatbl8uw2FcY/8kKHwR/7
T0FLqoIasoAwUeFo/wAD925cm5JbxUNN2v2f3AySWprGWsxDH4F7laQOw5DfVSft
iZxozvXsDzLUIHxw7ICBu6liC/0RYe/XwkTZW7IO8D+tkj6Pz/XyReWQa0WrszRX
Ft4Q8BCtf96Ui6IaVdmGn1hn4thdMyK7fQEAzPERvqEIQ8ZoZWLJ19BxSjfA8zsx
6tdGQT6u4FAYhGMTM3d3GLuyr0jEavyh2AbYBLlUvWc6fCd46msDUT1LXcOyj9Eb
r/CkPwYgz25VtqfzHuLdFb4uFT/BX0KYZdM+jt3KJwHATwXUanuxyOowe3hZ+mRf
JRVqhaAIVkybJugMku3/Fr241Fb9a/z1KNHPnrEEBK1wN4tMySFLiRLdt4uxXYPm
+ZawAvy1gof85V+YqRfy9udr62Ie0O+bxrIiAUePRRm9Fxni5ugCM8zf+QVj/7zj
ZcO9xrpPSWUK8GKkWEqMBQRlS42IIp8gVc7YOxgAk6WE7nlJybWhwY8efb2wS48b
t3YbLYXa8zZcADNeMEIgKdbthckHChtP/yu4DjlZUIqJdIklFvNNsLfvsHIbNmO+
j1gGpFrv0sl8V4x+l6KfEuA+pQjSsFaRoi//x9GzYXrz7QApyJ7upW+hqJfHSNEi
l3zvJOv/pHcozANvBqfzQLdztizeQYu2bmiOREEB6N0eAGBQuqQ/dlnTVWJB/YMF
Ozv06MRBQN4m1kC2GF91ps4pA3L8GqUfFv2mu7XNGkxGV7GOFo5dUyujfNT50X4L
eT/2iLSYTSNlq/vwv6FNG194DbDYqVXZv50FBmHgJRZpQlUQkDQ8ZmrjPWuoQXuo
pHK+5OFBciQErVRoXwdR+pHI20D4RfQ1Wiyn4KZ5DmXnGI6lZsAepkSwBl2z4aDU
DmUlvCETvrfx3+rZLz/DgFMKkshTDPnV1C+b0kscfZUSS1DnK8K1DxuqJt57XZvM
FOAA02nnq6xmh/2t48WFz3m3SqMdCJPRJMY5eYN5dSc/xZ/K4zvSGzOPAEGPT4H0
h6yIORXRtBiSG+tb4gJQHNer1Y0L/Rsogslk/TkTchko4JHdwntKqZMjLcmVVi9+
xyjlzgej0HRXRFA3uZym9QXBKIBDK6x/aCdu8iM39Blgc7xBHQg7vJ5Exclsw/j2
0zc3HzkXT611hJC90SqKaPtThgIVZ7Pa6FLp3XkocQ5MomEB5HYkfgHWQcks803f
NXY3sky6l+VCHFfSvvVlH2m5AfyZhdsjpc7C4JHDGr6Jc+cjxox+pWc20KpV94/b
h73bePKN9Xe/CwcwKlQQfZzAgBPtobsCmPmFUMV3+fXfWbJP3r/V1BOrXCMsRwkJ
PcuzEzJK05dmP2FYF2/jQmU2b4JD7QNkL/3JvbcN1C7XIkOFBJ487zjTUNqQjxU6
cjQ2ExVlS5d65yHpr3kkVfUtIXm4syImYaj20lhjAameHoCdpGpD/o8Vr3ufsDPg
hWGYzih9Z/ZWVb3y58Fdv1qAD8ocZ322sehPzacsGPA4JybC87AhsfYRSuceMFBQ
Olt88XMVBlpNR7BkBJ4l8M7/ZjFTnbQHobYdJtLsBpexnh8GeIz6LEyy/oepKtZS
uW7KETjc+K1b5GMAb2YGZYRXgIWb99xa1RMRUtg/I468g5JesHSx3VYCHi6wvAIr
lJWrS+B6eTBBGcQetvvHrRYstM3fkOM0LhxKY6KbOc/51odq+8K0L7tlzrHTTGVp
MI89rCLQCwPoLbE2xoLKV2ANWBTKVCwiuzxgVaqT/zxe0lPjOK8S5wfSttUTuQIY
JqB5ioaCTtMlnDo9fKwzKHYa+3oCa+KIWo7QjR+BiHJ2xxvfgNE5LGG/3ElQ4Dvu
wCZUNpwstnhm8FQTkSoYP6xNbROup6JymQaOthdcRPU/ybvrxaP08L0JzGAOry04
LshcCfbsIlE+6DvBs8zK2hNeOmeWAkQGzY73efs98X4Rs15XRWFiHD9HbWynif6E
VXNpsTcaEEx6YntDsE18yNAsQJxNgAPsPacHZiaVCjEU1dnDX2cIxIP3cBh/dlpg
1nXVvgF6t9lXDIXdSyFRxe7NCbhjoQ6TF37SCjD8GnP1MGTWRlGV90W0dgneFS6J
HZkftXv6RXDVKtyUR0zTGq31kH5qpDKVGWPvCQMXwwQct3Ml6oh+oyXWr9JrOo1X
/xOC4D/QR9aibLPG0dYcL1JgsCAfVoDNd7B+/rNCWFasckex8OnhCJOGoiwmI76Q
rn6qdjbl3Ehn69ZFIKnPp1i8B5oR8IKberpsEX+iI9RmkdCarQo15kB4ILqwMEHy
y/DUgaCmKSRq81pT3OTB9Wbg+95+7TDDxOpC+mP5LOcXc3TdhDPY9kVRgaZnn0ti
DPdpwDQxQ7e9avi3ZmH1dmnOMxwjzD9mBXtZn4r6ETdH/9HPzTHoUgISQVRAqU0U
lOVpltE7DXzC/Fu+DX/Jad1RTpfFtEwAVnVEtGC/pXHpvT4k43E5CdK658+4DgZK
yYjOldcSSlc80FUb40F+30H/LazA7SNEDhBbhYK9zbxNeV9ysbyJInbY8NPPnN9N
XC3emdu86SNGx4GP1nGmWpIWXXpDOXb255jLHuTUl/bAi8VpEZlFWY9LgBFVDNzC
Tj0p54HCp6MYFXd/ciKm+8Vmc+2qIuAMo+Ty7L2TuBg0qhU0hqbMHFBOz/Ed2f0o
fbZrtT2xJs9nzxbcDb+NjsuDNtUkckn3P3Ou99mQifQbZr0HGRtlD9Xq68NHJDCZ
p69gtewCneJrV1iIRF3CG8DbhObLhD9c1iE4xSlgIjDhETmxLACvyLUXfkogddlh
CBr5foww3skNBNM1iyGmJ1/kk6Km13133J2Gx8ymEyvfoIj+8WGZzKGiga2wujqu
z1tgdIvwaZCmk0Syp8vm1bO7yYG6PS+mmMbIEvlAiegTRRlp6sLimQF2Y02HcXSs
Up/qF1qKHus+VNESYWbGT7PpbwzSmU07h/7WEOOpa4vEoS5BuUYhB4t7eVP0od4X
hZStBKDpo8HksFP/ML6vE1eR9Hn3ASNtt9gaqshfOTQQqGISd7NIKltc7Lm/pa3S
aqreamgsVYuLivaY7OqVxuwjF2Z9oVZSR0O3OzrJVtQBNtJhM9+dCmnJxwiN8Apc
0OaYR7HJS3qKSmLkRmRPkHn5ajs1BK3KQXMpy3iVqFODtYlv+hbFBgqZ5x2pP+PZ
7+0S4iNh+D6Gzd4agdjgyyeUCboEqQJaHeL67rg0I9xkDvineQoxreh/nJ+bYmKC
gYY3VXsJ8oexF0LI+JWnrk3IyWHYpWzji6KTFeC3N12lJVxGsBIvksNr/je30WKw
+bASfSx25OsUuzZ1W0A6A498SJbxmgGsTs93zJRMU0AjNGxie9WKDOhEe4C3U+OJ
1McnqSqdn/NhaPuiWUHBvipPIVAMK/kAeV7nLW5u9B6YyegRuKrJIOPwxREJiobi
TZ/NGlPgNC98HwXowZyCc4iuDYmMsDscQcLVpaZacj0ZumdDBotua76mA1mQqHtu
wGKu7kpj+6ZElagI85SXo7COKXWBTqIrlfgdnj8s9UgZKr1YzTo/D13eGrlyVNd0
i9NHSelpEwk5J8S+kEjMhrUqhFFyA+Bo3ErWPLqmpC4cWkXwdjxrQUDZH3O5JSQa
6o15WDtCpdCxmhEyN4CjopVtExjkctFlK/m6fGmHzL/x8GRY/SWeiOJ87FbUwE/m
Ji2RoAop97fCddN7dfT+D7K6CxVgMZgpPvjQtInlNx0R49v3UiaydsJj68toMM0W
UjPkmnLuVARymOkNYn70kRDh375pDWQIF8UlNui4xf+nm8mj7aomcynO0wZApc5Q
YOoj9GbJKvh8Bh7kDTIOR0GrHW4Nn21+XNXo9FJqZfFZqXaRcIXsSxK/0WEcsi88
O7yIARDNFHOMi1BLuDsmFHh27/ZPdJTBTFVWoFQnh0LNoVMZV5IcbfiJbDy8wvam
m7SmrVbGUpzBrhKCZVuXIXoIluNYrIZlQkWrUO+3twr5Ng2Huxl3jZVzjXsdiGTQ
WcmXGiWXzBR8U/SvYIOnDLgDBd34VLJfvtKI/Gih7p74zSIQ8OvS0d2zJTZgQYo+
P4UyyXXVu8XIg/me8LyZrpNRxudfWcqRoML3BT63Zio6kfEKc6o4q1AMeHF52dgF
XXRncrgrAcPt4Ttk+4udac8vhTEZP7UX+39WWq34BJUVE0JjY2uxcFGK2/KE2Gj+
u1DnrLhwKsy0zVH7LYNCRSDrsm7vNCjiqj1CysLBL16dS/7g3XcR5UqMCvDM7G3o
Pc3DTNFyQISQcDYw/lPsIiKqH/4h9VTAiKQsYKZrbAoTJ907KUn9rfN9pH8gkzjD
VnbiZdbbALUUOdKcbpxYQskgSDBUSYXb5AHF7xedP8GBd2vSSSOa0VyceIHToSV4
MWWBRuNMO1gBRTyuuncnUfq3nEqPdlSxh36/yObVuUxpUg7EqLz97FAqpdhvjZmo
k5FQ57Z9EGzIIuCjgWnuHrv08PmUA3ZzCdgN+oLmMmv6cZwy3vrMDl3PxcMH3pR7
Wp0myQk4XZE3r+z8QBtIv9r8d8I6LixYxd92z4m0Z8Mlxo3vf9rcThvehNTljBaF
XFdZf/RIET8XgfR3xGpCOAOZq/5/BZueGwrN7MopP1TJEQK6j5YEQtOVmxcAoVO8
k4ZD45Yxd6Y9p79sPOUQ7JgDwegW7W4qSS6370PBThoczxrmnpo1dtNUmDsryeMd
QQK4teMoEjr9oIub1LJdN2feOoYedpE+/T43aSjl0fL6ef41r9z0VP0yIxy64WuF
Zf0vy9Q0SNv0NbSqHnTNCI2/4v92EQyvctybWfskxnPq8yLo+bt9230vQDGws2UE
GzZXL02dF+tsnQX1e+WQew5M9qXsgEuKxr4pezRWKSgM9lxcyXe06ivi6E0gHVvX
VwXd1buiK3tvb9aFW6ZdTekXzRzy7JtFJAX5UJUl4d5d63I1tHjYK2shpXO71lh2
T21pWzO+4+iSCstqCNcOlGaGo4nZmcHc8/7Zzwn0FlPgbz8U6bN2HQ+/5FVi9scB
x/4cPZcoAxdIfZ9H9eVSGFireaTUYuaFh4EkJigNZC6mugL3O78kWTOGlcwXxpIk
Ug6y6VUWCJ9ULK64ZuD/sroPh/iFPYO1Lw4agA4tmNaKk6djrDCGs5KqrhUHm7n1
Ong7+J4HHNxKmabVOOcMDWVDlYsi/wR9PAiyYrSpO+A8Zwf5NSsZOalpS703aJMp
TE1epFp7CX4X9DIJvwK5axAB0l6kCGKwYzPnK4Q07GEM/LdF982kC/Uli+DOX9pM
5vjfRcCewCr7pO0T6XDjrOR9gxtgrOg80LeIOIrDuFXGNSKjo02l9G5TIxEkuNnT
plFfeNPWEkojd89aGWKkDJb0VK5BGhpCUAuMyOkItkmLRDitX93OVt/128/WxOXi
fxmJfn7tFVYPpUT/m6Hs1tx7R9Nso0xzc2VdZ4spxa6t11SHyNkMqhQtHsj/jO8n
tSl85M70sTQ34ehhEWlIcG4CxkAYchLQ3kqQG1AcAd3QRljJUBasIPyqiiUuCrBZ
czOP1fH0P8sjGyKvJ6/VkkueyXqB8QbazlShJukV26nF9CiK+Y+Do/lJrZg+2aS+
uWDU0G0LHDTNQGQCxmGlw365OLITqLA+DGuOG0HjafKuUWgh8qLNnJbbK3SAI7rJ
9VgetUVvHe3L/2M2SvFe3jg8eJhjQZ1nzht9xHs59R/Twtyb94n4oBpps8/7UvKN
hLSiFit4tsGCwGUKUPnEqfDd0B2Xa7Cim/zzBNhrDoYI3IcRSAFXT/ypQrp82wWZ
uUM02CzzQUvb0gbVgLkWPM/xLhYe7xXIOTZlzFtfDlnCYkJwHQMnrFS/e9qXQcvw
AHB9Rg4gKnX3n2E86UXVjLLYrivjElBjAAK0xlahWO0NNlQAR5ThOqvOUxM5HSAO
qmrxYJVWS5nw/G4z5a+20xvpWQkdgDZ99NmtimOKEtrA3lFbyGULYUkN8aJC6KG5
1tPhQ/XiK9WuEBLL2L+/WtO7JuppzACIVP47gYyvJ435NQyRSVwWtyCRElV55wqX
9r3Ee3Ty3BjictbzJnbqwRYGYzZHOZqIDsPVOoqlPkjrEHlyDm2kheSYk89TLJ0F
gFdmhr6mSPv5Y9GOByndlCaJKPTO/AAE2KNqmvpfqE5x+Dtf5ArwU7JwM6BCIyJ6
L05ewWuxwD8cehtyqcgzlvWO4RwUc1gKwYkU31sG+zhj7UN7vs3FUsEuNZdB7Qmn
0JZ84Mr9LJQixUfP//6xfaBI1Tm9AGOl4m6OQJ1D+xwIqIoJbXD1cEseVzY0ozjN
hN5KlafMzlxEXF4Kog1SRouCvcjiz76XX144+w53TouOLXMPE6F3pLYFkAZgd8Rx
Ifhmmc3/a9BGiQ9k4Sjy2Vce1DvmQn0pUIyeZHpTKrcbtaKCBldtbzC1RXObZlnF
Aw5xFTNHyahJXIku+NsdMERdRIKsk4lnypOyOD0B9LoCWV5X6Xl9mD1qW3gSur7+
HpdmqTs5Z+HRLprxEjN3GZq+uz22lbXo71vQr6vM08Ac1hNZqU385VTAI3nRR92N
oVc99ndPcOx1dwzrGSC/hbi5yn8eAh/mpj14/2ARGk7KQ+uHdWxDlxJNg2aYh756
rZG/H6H5tezojOPuyQD+RCfIcKj+5zs9DuFGb1ICkpe73jO0ff4MNO6kOIdQcptf
mzrQ5BgA2XVwLgP4biQ7fONygnIm4yDColvNZAsRw7SksMrynNfAd/5a1wwTFF+m
ZLDz6X5d6pEHzj38w+JLQXAHfyk5ZZF/fmlNtu8JNf9T3N6LbsIonb1RU7gsciqs
i6DTLHroTihbwkXuiR9zw9lnqvHhyvEbko1Y3MBoGxJyFCxnaUz9w7BaEEkhRsvF
Wr63EGd/CZQCnr6BCgxk56Ejj4v1jrhXdP6pdb6cF4tnnGpyAcplO9in+GC8ALIe
/KoA5NQ/woFJQtigBJN0J5mTjQ2OyR5mvp3CCGCzZvjclDqxfquR/n9Kj5rfutVe
R+FvkAZAhpqAA5ZhFh63q43eOGS6g4D7Rw5vJSKAfZxI+nanxSc1LpnIS4R4jLh5
gZMCyIBhs1454OTpx1G6sqFHMTbe0viQq/36R+O77KLyxHf3s7201+Mn36EeJ2Yp
3KKQTYqrIyGmfZUpn/Ukr22Ipui8gt0YcIHDG1Mf3YVA7gMzA74cS0ZT/1H6B6dl
yJdrZxwS5mamZXe1U6QkOuFXM+5Q7K8W76L2E/hYTmf2B5wAGslb2qa47mq8crVS
FGoudK+IAAm+kUqnmNvdqL8F2+vmge3CULnVCNZ2/InmmtzvCasRkz1T0uVwmQAd
MNkXndmmlJrB1BNrZYCIlj6pcNv6zFwU8gkoKLjUgwhbLTFSYNNu3BfVLdclnIQT
7YTGgo+3ffRwRiqPXBw4loPKUemclpT0xZM1PohgDq1FQAfn5yy3RHj3dhRG/C+u
/Ey14itlejR8sbPBAiWnyXAHLuAugqqLl2t0wIzkxVF9zWx2JNJ8WalJuv+T8JY+
YfDY1m8uULQ5JA/T7U7UWRXBRL3k+v3QV8vQqxeEbASCnnPff1rBAxZCaXsqSsTW
hFK1RcfgjThECICW0DL/XQ528SAWyedQwTL9Xj5/jtxyPo6OLOXS57yDTOYxX0T7
mkkVgtlrOvY5ImrEKA9+ThoLQXVztbLaOo9f9bwqBYoSDWWAP/bXqD8DeWTypLLD
8R7NRAwEok6y+gJ6yuG6QTduAaVTsmvDFwv++IhxHEXDnDAyY22ynrA/Z2mr9vLz
7tkBfuS/yqPRvxlfzHIDYnsAAKIVtUBChIKOMyVvMK0MyUBHkTM9Gv/BkUG9FTFS
pmQogtNmxKnLqU30XqeaSFAb9fQJexkw0qPlAlFySz/Fki8aeoD6qDZWVqoFVbUM
rWsrd/ocwnDWVt9/bUaql+H1NVJ1acSzZexH78ZS4L6PRmC/bk3NvBytOnLPPZ6k
c1o44neal+DxnzYdSGiP3WxVe1goUsODGBFYH9iG24BPbqv3fk5im8qOO1LCNbw+
rowYjBDdttU6JX7Qjw6b/FwOdnh5Dvx55YlAGEluiUduOSccZ3w/zXVY4ne8A5BA
g5jTXYDMhuggZivhfph1rZedmfi0VAPoPbtZOplh1KkrAvNsdeBQ3grE+inKbJhP
De3CK37R/Gob4WQeuhPkBwr/vTL5FMibKLpx5EgGryq151W65gD+4K/0O6VR8Lqf
3wkTaS0NBGCYut8i478RDPr4t3uEUH6XXAnDSEdMVoFNxQqOcrRzMBQRxKK//igu
Nd7+cyTQ4wFmHgBm+IvI+JeH6dWm7+GgbUZlNQvKfPUXyBhyu2taE7RQV6KRv+Lu
EkhfGV2JrrsrkQN9svrN2W99kxB3ucJLxGypDHPBhA58EAvwf0gq4PG2Q26Pj1jo
QMkJXm8L8jhzalQY57VjNObl6S3FyiHR0QCGw/UbUhxDoGuQ3D0KVqA2ZjiHZ3Zd
Q2UKX8igyMCHdmn2BQbotaup6L/Lqj+91FacxeZTa1Qde8aMoevlGzHbAtHrC/z9
wVfuvKnynwhA2Sr1WVneOzyk7BbYxPyamXph2Xsjp5crNgeRZs6f143uuJJdG0zi
hCsyKjQL9hF3XTPFjK7NLrPk2R92fSlEaOwFQf5s3ykXGHY2YtKTOTSAD4Y5ZZbH
Q3btvTHFwoBC0RRYaLCMx/1d4KdkAygAMKQ47hIMh6FWldgcW8wzkJE6PVOQJfC6
K3VKYcDjD+stJ3JFvDkxRa+NXuWFbQn8YkxQNcFPz9784SunzKjzn/YJQiawG2iU
sI7ycMn8IT7V06AE74zDgevqTTVn9Jgt2c6etYywPPJvOEB/HLzw7ozoVB+0HnJr
byz3huT5zxkiBC9i4Ob5vlsUdUy3RCkZUl5PotPJzs1E+OTFOgwGytdMPtmh4Vdw
2gFviKQD4NHGUU9hK9eybtv1HypgxGU12mFqtvFpaLHQ9j0lVXx1ETYCknWaEQIZ
HVZRE2jnXZojM+C5P0hE7tY9yBpc478/hOG1ph7Ebl2SBg2tM51VOlBcBfippUXf
MIz1pp02vaBfiVmIJ757SSe7io4+1x699+ttx87GTDpAAZlGHQFFTfqwytJmN6bT
IHeUzgU65Qj0Uyc/cKn+qqLuDM+GnouDwHMi1bgR2e74U5xdSKCCgoSiD2tuhj+V
8UxL26CeiBY2+qKiRoFbZZhTnBqy4L3HtcwzoK+RB56/3qXg8PDQwzItb4R6lzkd
PMnUKuWuTDgVyIsHHaL3DxfDazp+wjB/Sccp6p74Zhe8CS84Qnzd/BTSkfGTvZ2C
R/5FtrS/cXa5JLXJ+HJX88IUbFY4EPZckHQS4/mgRzpDfEzEkzuXhxMwNR10vkXY
7LgJkRxIiIKMdZQxBx+WGjWXZmEZieB7MTKIEswDgNVR6+kvWCp11jfFZFfFAB5H
5JvsLNHUf3TIVwFalOmErlKBDm/hFhBItHqKxnoxSlNETX2RYIWuK4foFhn5o6pc
0FTvknX6O1475FaeGxPeQ5JKGQjhmok4+CsJ2U4MO5Cr5gtwWAc+OjJGnbVZUgZk
NAs1zlbpyFx5IHyr6sXWb2piUq5ra8LsH9ULHckGyiIvbDACDWE0maJRNYdGm8qq
`protect END_PROTECTED