-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
N6hzJuZjBJQKotRYmSy1EKo+Ty+5b0f5LLZfqJonh1o04Y6npybv5b8CHboml1UI
U79OlD0I8hq3VCbwefSRejN2rGavxJzaanYESM2wGByzBdOYAFmqHaINGgQld/Qk
a8ohNJSJObwtC15iCRkAXz6ABsTmaV1VONXTO3huVQMPPHNzIdZmFA==
--pragma protect end_key_block
--pragma protect digest_block
fyPlpdOxcSoGoLGuoIYJdXzWxbs=
--pragma protect end_digest_block
--pragma protect data_block
NPGkioGLwtEG3YeiS/yvzwwLPDK7gy7p9nED5p4j7pqyaSiYeizw4aeq2c3Sdmpv
EUy/APZEytVEzDmm9sYx+xp1eUb+hJOYF54hSuBFjx7VJ1G4VJNTjQMPXRNDXVCc
CaNpXbBnLJBilKGak6OkHSd+HZsyR/zvPP2My8qyu+1pH4exU02fsyosJT6buR2K
Aub7JN5264SwCmEsYxR1MkpOLzQmJxxoZyqhvsgYH+e/TSPUbXkhh9o/j6VwrAn9
maRkFcYLqUQhTXyBLv8XIDRlfgV79rJhwufNg2xYGcj9JDWsdsjscOd0NUEh2JC6
y0PPUCcd3CaMl3+MEz/fyo3hQN4ajQm/ZtpqZ9xWWR6e4nbA4aXcPae/K8PY5YJj
JSldEhS1SIEG5/ORnz2Hx3RLSXhdOHjkduJc3vGLnX6+/gNnnEQXPxAyk4r2Oxpy
2CDzGXpEbatKAKQ2rVBP/fpUXktTel6rmWRqlF07RQYa3mTeqrB5ffT/Tv0mcZwz
EqXicf5cmaEYSlmUqRyhG2/UfWEo6t8rT5MRKBpZrcA52J3J9ZnLlSwFLCBc2qDa
xSluTEuDdXkYu+wMJqOn0nukfbS1VW1kgfOxkQzFgd4BRq/S+VmT03eNDlM5xgsw
CV9fFytoXg4Owe1SDSIE2TlLJoqCW1guQ8giXlBV2IZB5A/F0VUtIT7SM/QohCUs
0dv5AzXt2hSsyHtrDN9tJlCKQcWiuHAaFK1Rlb1mjU0QkElHXTTX4AeCGZL3stO6
2IkrOLcfmNJ29hYSGbVh96ZVUA9G0MfuPGX37pcdPIN7lM2hHFI7S67EiDaJBxa0
cXy4lQ0QlRy4XNkp65a6CLE5G10DTR1HxeGsTWP14WZepTJYLs5zyc0F08U32iT9
xnwSLT7528ZgbZDcPR6AixkX32PNc6KxRhw8yncv1eGUsz3lME2TGeC5d0qzv4Ae
OfrKuj3K7ZyKeEYdxr2HjUWhsXV3V+HvfbWbe4e86+627v8Ae4IVA2aIyEglxzia
5SFZ4wOCJanNAHWyrFosuzt793lS5VRVUCx0vlYUjM/jkQcDWihAEXJSIdsvOeEE
e1k67OLkqNQGK72T9SGjzk6cucDt9bVmhjJCUDfpsVIJHexYq0z6aCByN5Sof9cq
f8pSVyhpAFfa9vHnE4G5w/lY+F8ywRb4XUOYzLSX/uvj8Z9SoIIhaiKGOCo76sZA
k1sURGfdDqXpUrFDxQ3IqOEgLjAWOAJWggVWdfZ3NAPTXFBtLW7YKvvKGewM/r6e
HsNxjG3X8iAgXGFMLWx6e4Pu5MSlmYg7HnWrqLBPkPHMppna+pgz1vJsYmcVUkSl
y2zlbgF7K6f/s1zJGD/TmqLyR6G+QgsoIHhTtASsQ2d6v6AtkjgOSoKlpsEVLgiw
kiMNmMorX7K94BjF9BDPDBQazAGilxjwWgqOpy1tk20byx1fa/N5nnzx57D6UQ80
PnEfJy1zzSEqfEQcOWVBYA/cfVyxHHaCDD+lj1+r2uw/y+2SVt8gUXS5IWI9jq4f
6AW2lbt92O6ZMX2XtUVJqVd0RT1hr12QvikBJGZI1uWemVwCSwiKJhsZwPKQ4jWN
tW9LHZgjp0M8BNgK0O/UxM8ub59Y+5bK7aDGkONUHw0epil+2AqRojZR0DDYz9HV
a9dGPspdTAflgOb9/SxsCn3azEXJ1LBvn4tX2shLrbWlfhH7zE4CjbBBIHZmOoO1
J+mP59mDi9+T/d4oFte8QkQTIhrGc+TzOIzzqgSCsTG8k3oB/j+rRKVPKVN6tCwr
MbMAQTcuWv+tub3mpmSzjrK6E96BYsqH5elBNVdJK7j2LV0CkG46SANjmmx87KiE
x7jWLIkAo3bWCpeXkCrUq31Gk7xJnlwy3SwM0PviVYQTb+G78gJVbVHMG1/a50B0
tJo+Kd81sKufZuO4D4fLUZuYL6BRd9VpRh6KUY7vNRO6a5+Zgz1HlC3HllOjsGWM
YdvWFCSKXpMpUuZ1sNNSLr/6OhZl5ymZGH0LVVeyNO8VSti3m6Qj/VqjIS2SWBQI
OJuRvR6xlF1llF4ov5HvGenelIwduEzki2Ty3ug9r7ufb5PsvF+l6KRRepT6uFhK
fuDsHLh0ZgBRp+Dpw45h7YLWnYTU8e6WT532TUNayzxnSL5ovJg7dPkYoPm4zBa/
Jb+qR9/MCySrNGatg2SUiFngk2zx2ptddcFrO7Gs1ndK136FrdbXYo6DGr9+faTb
AuqN3M8YFjsl+98BVf/3iB16WpGLmO7jBewSf4dfgv02teU7Ya+o7f/1Gt5YHqGu
Kjs3QBtXc8RpkXCIQmqw02bv4zXeJvJ9/uIZ4bjsgvWViqYscWP5/g9nWiOjQV9i
XhxQRBdghnQaiQ12/ycrPjh23xtmEzF/6fl0BbngRnMiiSK+yXuW6SuG3PZx8X1c
sfHfE/LI+wAEL2HALCqnmFb+MmoA27FojSERB9vldtB/RA3aWSSFdX3hykxZYGW1
RHJ44pw2XypK1/z77cdYhMTy4/gdoy1W5z/7Lv3Iw1bz2OfyPl1Hx5mVNZmuI1K3
th0a7XTk+ygfi8zl0fAXupWkZwwD6qQZrKT0AODLPGcujm/NpJnIHY7nRrDkpe71
x9DabbSWIo5QJtcwtQDlxJ8MzlBQ/XStdxRZo6DjluNfTRySlRaZK1CZi3Shk10I
ZHnHVTzZyz1zmLYso0b0I12NIgi4pSTJmZei98wl35Skpye+6LqO6muvWR7jpeWS
R7qEUNBvsKek0Wssy29RLImZ9EincVGvcFlftAdg3MKmKa0h1cOukbck2VYMdLic
/6tUX9HxxgZZIQbWoohF+9KkKWk/vMg/609A78jMOkPwd5onWUFTF27zoJTlbGsU
JXA7HVAuTXnbmqFAfYbbTnuCA03rZqWnSwXx9qALFgfeVR4h2exLg403/1UIT+tF
AuCovnT4A5LD5GYhPr/LLg6kMSI8NQg/29GGY90gzVEig7IdtkUDkG9yJ0P7D9Yc
21jtCL23YM9sG0wN19KUnhontkE9XGYvkSt6roIqsgh6gFxJuQwZxnqfkqfBtDe+
10LVDfrmRXLDtNCxgK0jMckQdkT2Ad3WxUMK9dbdxKHl5UASda+mUrP1lFQL8Z8x
UP7EFmrsw0PqiadVIURTQwbgZbvHKa2rB33VyxS6Xk0eqSLqxq9WXfGwcKS6e8l1
5mzDtmHgQ4PzDFtJLGfHIVEcseeBDdpbjqaZNv7hbl3ftoUIYt9lDa9Gg0YW66xV
VqfRDtBhQuEYrGttkGlKmOzS+k2Eeg2HQWzbKHjmSaSwR8QeFdTeT9eZW9WzVPD9
dTrG6epETMlqgJ4YxLb6d+aXJHi4B4HPk7rOQKrDpLfkuS2+8rsGQi9D+8kPyyxV
U7tZsBOnYvz+2xZC/pqZK+Kf2tVLLvT/GE1B8/4YCbYQZQkvrkS7EPUMVoPZ6AKp
q5OS+oXVqN0z2wnVyKDo98EZ/KYgvklprnRJS1D8bFy4F/Ux5NeR40Niz6Ce3Ppg
7R2G/5/G+Q7e4nvEQtGCJ8N2CubjBowD0g+/CkyMJUCnzte1yFc19O+eG1EBz7Wh
gMU+S+TkKZe9aeNZEW9cbWyBEE0st0yQObCdsvmeYlnh9pbA3IA+83QWdu1sHVNX
RQwwnzjEN31OCT1fke/yS6lJ5jwlJQlIrdtSi3EGqwhMk0awazNQLawmtgVmDOwE
SVdxNzMROJIhVHL+4iL3dXPrLrV/LEGC7FTUQD4uLlnZPje5vA5pIrK6NW20Pgle
pol/KkAVk2RdKSut/R56OFPjfoWLwh2U4an5F1qa5SjeoMPuurKYMIjUmJnjJkHX
AuMRb25sFfMHILke+VEYPNzeysZLcK0CL3bsv2OgFLPTpa4XRhPw+1l1EZumumY3
PbzWJUvxwkp5gNwBwmVk8hRszR8XciORSu7lUokOemb6BnO/aAlCjjnmBddDj0vX
m6btjRhWx3q/wnGM66b2n+vMhWy5ewVxn6ECPWF/WyeNQKbFE0cmHEjqVHA4gXss
iulp64CWYAafPM5cP4lvxEgy4o1tDspdie4JLcZNsg7MRu0K9aYw8v4/S0iwaTIU
76evw7vECxYywG2FTaQb/pOzkj0xhIOBc29iY78e/UhBfTIiwSCtA3h+qEpFveoB
WW5tXg5YyeJBwQ9eXiCpup7pP/XOOmQQ/ON15Px6maXJ82AwcvX2uV52nl4IvxfJ
cIXlL+OH4/6kzE6bxUiAh4ykKZ60C0A6avMwBqHNpbaOorBkyccLPnmVX0aMHtbp
MHnU9kAYh/kDiMsr6nXnWkPOJ0cv8//ffR7dkm2nGK/vPoY51zD2ns3zKgPJRE2H
XPxpwjOvbUm0CdLyzhQ6wdnB/VDCspcEvwIocnPeJpn0L+6cnIDf/rSeUsZw8l96
otEQ40hhItViaYc5I5d2I/hdgTz6EGdvQ4y6ULEUp68tYfSrzmAxuf1TwpI1bC3M
RuJJ5yeqnHYkzDeiZ5443S96yBoVeBsxYRqkC1HMqS3xuv3tMeOMWuWVFWmplTc8
wBzE+g4xUoCxCVbqwQQXz3M8I394rm8k5k//+ZCmzn12vJNN12zfoLKCTRxECY1I
IDoEeQOuBNZ+jg8hgAsQ7rWoBG3yBnx6I4mmRmeNDhOT0rj+V7iTNlo2qH1QSd31
vwpnAA0nSl4c70waJozKFTJmCLnMfpmm2wdvFUR45S+P4YnON0DqlVcqeFzfM4hB
KRm8Fb/TT+LDy9t9PF/GxqH8lOoCR+IYtmXiut3TEsJantO3CW6uZLF4H64Sfk75
AzTkzLvGiIX7hDps+CoHTbWPnSz9xsj2fBuRHC0RSg8F4XvbCbV0XUdz0fjzBFPV
RWBdMmLDMSfDWPzw07WrXtjeicWd0m9653JBCW+nMa1Kwkb4lp+L7D7U8AojkERy
2gc+S6LA7lDivTNPtG3LmllZGulVIkp6tAcPlbvYh4qCRqZOld3k7o7cC4jl7cZ+
kYIGwdGAnsnT1C2rbN5HGJBCvzAvS3Le1Az6XYGfxIiajzcSlWL+R5CAenqtRmDl
gBrNPJPREgLiG0VmAyGbR8R0EssLAU2svLbw6ypqvWkX3E4cMkYrnGiXgD6RARzq
Io5bqFDpdOWNBXwvOIbFb2OYbOUlP2iCj3/jBHc2Hv2nJ4on2QkeulrYJxA8o/Nw
9xhwGtsln+jFwYmp5Pw6cqK0vOKmFkE4MPunGiGr4E4dk+6P9gppMRvrXPUMBMX8
/bpUFOebyY8G1TEUdf+4fPoXGhyIZyct1bflUduPZqGlANvEflcVAhrkF2brVGQw
dsJ0SZfTDNnCIh7GNZ3VEFE/8GS+L17Uy5KIpL1b1y7cLk2DBEWhiQRoT3niVxVG
K7+gJP76UyeqVSm/pf7IdbcQKXTdqgSE02lEw1isqqKhVvj215i5l1sTRUHmPzv6
xM+fkKTEr2Kfe/IVcgCdpiPMNzll7g9BQOGvC9DwYvhtw0J9O11drRT1nxlseyRW
b4vLipMiyz0Izt4khK+Y6k8enhmt8DQIucKMIQPbSTa93ZSqx2M0IuYZBGqilxYt
bYKQ1VxKLP8JOjCOht05jf9P9/sCfkXja4pbya41CUZemysrAHzneDGLeuUGFdT1
zZZluKrTwMoIJMqRmrTQMPU0QPDkR8cpPd8sl6gFzfKIH0jWMS0piHxtuz3Kb7BF
8ELSQYzlnvV8SYEhsMvmMCSC74lXi5aZuLjttbqV+xe/RsosGUzmNTLSm64B/6yI
qYwbpBJmpLqhymw0WfGooP3z2Wm4sPDu1rRqrkfJpk9Ux3SqVhTvHz18xciKaWXx
Vx3kipqOOL369+t6jGvMIA3HKBDtq2eshj/bCmvrqib5QHmb62ej+BAyo+U1qaQF
ypCGjUr7rBzGK3ltz7ei23f8lKyaoeCDcDfc2psN1Os6EgHgRmZ0BPPqsyCRh741
39919IDOXHntfCIMv5fgpNW/jSpN638AqDlgV7CzyZMtaD4dJrq6Fg9Dm+/8VTk+
y6nk6vZqJEiNff9hA0JlCKnLhlbc7vaFMkJHeRiIuDQJG35P9pIr/P0y5hcGSVO7
VSCqDjcEu2Q4mEBQMACNpi2oiaO/uJ2Ehw9PSe03KYX5FDOQ9LJGJdLb6tr6IX5D
xMvk2EpXrJZkLxQ8G4P4drxfQkqpI0JtkH5+NvSKsR9PeKHeHwhERRkoYdDOSfyp
gUkY68BlhKNg0UIalVnETvcWOWY5YGAvyIdH/gQJCGy5NxxJws/Cn8Gk8KLKk+am
sMY5/uLxHrKiZyXhgs5Cf9RP8gSm5ZLwu/OkxHxaF01HE81OwNigqoWOxbS4/lI3
n52ruIQY9QIYFNWfiNumn6Ld8kskVMQYd4g3Bqj8pW0DGDiEH2febo+Mlcl+sgsn
ODsYmPGD5xgrjl1E1UCQ0bYpy6fI5e8fSMWmB5QMFOYwXmsr0wYIH6swOr7OYTx2
QlJmwXEj65FlxcEk4Fyid/Se31Ob3cGqxPt+jQdycMrFggktp96KKEy6AZpmqQ59
6Ayzn6+x5KEOcTlytGuLxu2PGuSIASdRDsZ/O0Thh1qSA+3QkmiQFFbdl3sulxCE
cDnCIlC2hbfwogSuqi8WzWHDrkfpP6Ypf5GdaXj4iH6e/6y3G5e6jHw90WbvC3D7
d5TkOURFrUAOEe092cFFnz3etxklzvIHTWSYNuKRnjEMiEWhhQaADKYN1UPefQkS
yXAtcW1VgR0eUdGGQIhh4eqsOsUtSumYkHEcwcj27WGBwTcsAMj5KhPe7UooW/US
hula+MmMk1mp64a8lrvWFnCDoLa13fonC4V+iKwNm9bsZipXrQXJop7G23w92br/
rRSCqnH3srshGr7ph3bjq7RCajx3EhWIjKp0yov7isKUjPmGyn25J+HS5FTuj+A5
cRV6FCtpFr2g/Et/ppp4d+RPIMBEp7UQIFRi5lE7TjOaSxakc5IEpZ8cbk98NK2A
R2w7pv+QMz/RH+I4cRgb00wlXOgCfOJDDtOn5sdPEbuHSi/o/iz7RagDv9md203o
sEbVG5U6B8AkL8enf4BvWzNOGyN4B1jYBmV7LHtrr08ZrAsXvHQEiEqU1LAZl1Qh
X8HtXgnJwtb1EN7zRp+dC40ngFChNbq8VftQrFw7BkgFFSWY6y8lglX6/aSrYdJi
eDcaa4vXA0O19HxNIAjw/eTwni1i9AjHKqqFFtFFuDzTJeDh4+3n4BBpzslbAf0C
0Zsxz/Y9nNh7FH12i1utcZEr2QNncDoixs2Of6Z/Yecd31Lbnp11kd27DOPpzzJg
UxtUWYb8mVrq15aw7VltWfsA5yCapINRAYqjKC3+0cJXIG/pQcvSNnhwDM00Yvl7
Gxye1g/UrTwOMFNQBGO4LY3EzwHQiYaYdCgRUhQSb0VY3oXjvcK9BnFUqzwLv7Uy
VDQuvdZKMc87ngEN8ywWjA5E0w7qNkpTS4WWwP1n3QpiYFBoXFFBDOIZeRsAe4lv
vOkQ9KvCbP2egxDyzd9I1YzOlq5Ij9hYTvMObKBuoKcIIm9dCBQW6Pgddpw6RUOy
fbwD6RZUSMw1qE31AbpOkVPRJCtRfaRBas7Zr7bE46q/F6jYboZ9vBNZNMCadVqr
G5jdzJfIvKJHHlMzHthvJNc/ahPTRPGnkufMSE0pyP/ZBq44dHDRTcH79vhVDd9o
W16Z4CbOV34F5+nTE6M+3GY9q2uu5xbJRoP1GQRU9wdohElzTJoATizXX06pylaS
gES979jpLAjGCSeVQ0pKwUqIJaWLMsjo8SZF2BWY+eTRYgvCS+/kXRoN6U3k4BCE
V8xh/8ooeicOOU4+XOR9TVNANRNpdrURrbQjsGr5WmfZbZYYgZT4sWSHEZTId84X
YUWwzVoHjubT3SmknwLiFXTSca4vAG/wz23CHkOD6IQDk5ZqpbkaqNaoz1tBToH0
W7hJg/XxPn9xv4PF3ca6sckeQiWpxcZEb4rjnjWyr0D0JqtsJl2YFoXpTbU21ocC
p0tIo6Ieqf/Y25EiWsN584fo4zoTWIldftEyZRZTDHkBnWaxE4Cz8TUNsL6B2z6I
ygwokSP/QtZkcHhVWpJAHt2E8T/9zFVSpxP3Bcmaoy/CaLBfKQHRYuZThYQHiwGa
22wvJlkBG8rjslzFFr8BmeTL5Syci4auDeAxRh2T9qjw4vQ0xno15F1VCOWfH+r3
Ic+2qE8iyeODfR7bCDi4Q1B3R8fYemOmGQwZ1tHA9UMcdvlgnXOONBYBx+BQq0aJ
nIyLiqYEZE5VVxzIovZjPdVTH9ybDlmoQ9w/wyCuMQ5DHcxrPK8yWVV3Nw9oye28
yxLpByEe5giW8upJDxJMr/thP/7BtmLrVaIW+RtC0VsrAchBPCVjseT6RR2hv8Af
xZOm7CIGHuZH8NVrRIwxTfSV8R5WeW7zWx1dh+CwnAjhIlGHwLacMSj1fMofSiEJ
Almkn80RHntYduQalgF+JHS9/2aJ0EejWrpWJF43UsgVz5NyLlvvXoSR9OtUukPv
hPOU7NkCMUkakwUCyGosMEDYY0AJmKVCpH8o6dIZ7UznhHYvuLl/rAwpRrPYf8xr
bjUlWqQmueQv7sCNTGMoa2wBSuY6CWmg85JnJvGe6tD7TyOqkZCoEBSfrB6VDYfr
dQqWa5SClRkvYZZFSzLUUZcUxJlWgD/GwPF0jYSDtmSCnqBzXYOC6YPu1TYfqPq3
2lk84yZCv3WBTl4xTL26R/EPXQ/FD4cANjVn6wcn5glkT0qngJpdQHF9EkwG1DQG
H15O1gi9E1m+bm0aYcUzECbRknD0gQcG+tDGEVwOEp7rIe9sZaAGSqd9UidAC15z
qFpUwPTYCtJfoTY6+8O90pkvmaQiBc0dkC6aspIZ8DF2LxYZinxMurDo05m4ILq7
5DcLXJE7pamxEwgH6Hg409G2Uz16bptBuJ0/h2X7TkCLhhf7ONvBk81FUZo1lrN8
EaawSYca2nnSo4pg76byQEN7pdhXpKTetLf/mKxYO2ZBn/n1uAqFE15b/l/3tA7S
wpzXqDfIA/w5k36xSqd+jmW6Hn2W7L2OTiWfCzww68PEbF35nycv4pT4ijYq6a4A
DxsYv6+JOFT34UuPsv4MetZB6orxV8Mt8t7C9p/ZFtMS7j1EvfTkhC7Ap37+C1W3
sjOVpdXEQSea9+ZibNQRDev/Kw9LSQ9geLU1QCSYYAr14A/mubX2ELbhEaJLeick
jSk/m9IFpZzluXXDjYN9U/milKizB4LlovQntM802VZrL7ene8dkyKL9IlXebQh3
em8ijQZCfY0w35DKDCrjo6OnCrN6rqYcNm8r3+ijkxVD9E6xfvH5kT6+s3vsQn9b
wnqLs4FxwlQFD1+HHB/CJrSXeEL+oWBOpKXGc+l7TlTnqb8Uy1t78ifSuZlCJhIA
hC7O7ckEZr2zJKWfdiRH7To3/sNRDVP4F+1s1I1HYsEzYdpHqBBFiBOqyDZBxRFs
KpGaehMVZSW0QfuswKROzoDOMbS03g7qJnGcYXc5N9rTpLLznHysB0ho5nxVE1Mr
ce4B8c7gKoXFP08OGqcnrTuASmNyAauGB0Qp0RcVOIfkxseF5gTJh/9OJyGAqiYd
YNTFpi+0vWSRIw1SgrDeOm1H6+aEitwLk0ZXRMoIiLVcDzCSIB0sDpbhjvqkgLuY
So1/cjPNjU0czwn09x3l5pg1QdvKXvcwd5z/5x4VhsbUx3U3j9zPMDfSSlK1cyTv
jGS+IrC3x4Q25MUy6qUHKHMshUmXn2V9+FEs9iGVnMa90ZBo7I9+WkJ4cMTobdwH
AdDojWOTYUejlL1H00MzPwJT1Up1qCcsMhIhYqY2VUAR1Uyl/g45EPAmqijzulE2
UKnwjQdqu2zOAx76xXLUPkDMVLqlyl2DGT8AiJ9j7SUFYGUg1MCDPVKLrqWF1zcg
D5/x8V/lZ293G+5k0H3LrGKdKTVAM+18sHJalp3Y6XsZW7T+MxG+gSn+j0Fds8VT
WNnqP5y4aZxorjYKNzlyGKnwCy/jwdJdRmJB1rI50bVKKB/C8iB6O7Zyn9mNk/ql
GjAhCPhdDGEqYUVrjZSeuScBR2JGRAWrJI+K4O42bPbf8af3Wk5x6Wi5elMnqc5C
s4WmZAkRRTjwDY3tjZ5tsJsipkRkirx/Ny++ZKuNpGxnI+WhzokuWrLPyzWBBiuV
Kop8y8Kwjn7ibovkgXMfJHc3paNfuhkK2IqLMOZYl19vnhFNIymbXcOY04n3AX2Y
rP9qhBs/hmSxsfQ5qS2zN/GLsNrkWb7USWn2PgUFE9g/C6rL92FXhSl++fLeRy39
tL6vGe1n63Kb68b8jJDA7axTHcX9zq7P90YGm5sIk1q6ahP0RMKSmhxtR/OF1A/N
FnPhSqV8TTHzbr7I70Q1AwXOMW6oNaQzvvVafJ/F/SAHeHlJiamAWpb4Pkn/owZu
ouEQo30BjfvPqknMf9oULOZPZPl1BLNyqYdWvBTpGGwLU8/w7y3c8yVCt7MCM6V8
FmW5+NCRtN0zs+BfLy+AwI2VIoRPk1aQQFEXvAJbpGOEnmSQkToGaeH9lP4E1P2O
UM6i7/FkmTyDLT2XljI2vzFz58deKUEiZwdd+uo53kWunB8q+Dy1xuHRsd4E5jay
HXlx3biqKMQa82d5fwUxgTnQQ0EjVQzh1aqNgYn57I5W+p222pwms/iAguQ8gY7T
jND70xmpEM6lZ0qjLkDTiE/Z7YK3BJbIVSb1Ge5TLq3+OQ8usU+iWAtg8nyfEvax
e43A2zKkyo/k99NLNw9hGct97mX52RnH9ORGbCmHnayuSFyr9mgt6iE/gmorNT8r
Rp2FU8W4z5iSOBBaM0KKRlEgBh0ChiDK0sKQRctPeHczkNgxmrvg1I40D82SsTUH
whEGtVHXu59QrWwWce2q1qwk/1DmsTOMOkLDbCQ6PLVXtkETwIMrvItNcBFAvZYE
uTAwuG17BzeD19p8vdk6x3Y7v2q9IXzCOKgjlw5J04VLaDD8LoSDDvvl9qsv8WYd
gW1X38B6NjVhz07G7EPISFVAxChg5GLV5WXQRy/hAYMN6CtThmtFiDc7rLsMf1/X
+mxs+wwTYugM77Fpo7dYLGxTsmr/uLoNzMYSpqi2TBTRY642uifdHx+hN7q03Woe
pLPyVgb3QYRBdg0Yk/izHNmZynwXltj+iIKBfwBq8qyJPfkdAZJXG/aX+gRG6+du
HhrquYt7AOO3EHFAN2Rnt05Iwa7qOD/edu0w6o96g+zmg8Jx2IXeAgmO6Ax82hNs
+NOYR6MzDmMFK/tJ+9GypB6TxEJPooY7X8JDSGwIyHkm4n5btcj5TpxQClrQn4n/
6DM2BAmOjVDsrVweHuI6PZUS9IyWwGRjtpO1lJnQ7QPZE6AfLZT+IV63j9tQ2dLI
zB5mjYPyyZoX3OqO/0liDzRQcDVT8H91YaWH/TE8YWKIpW/3rsbKSZSF+afQkgYk
uMn6NPvrmoY+doTKMhQpoLXJndGJSzaOcPAACR8cxXnBNhJ7WQJs9zRNy4eZyv7H
8PBxD4xugd93vuo4ifzatTq6NfPlz83yvwzLMNrqNA6C5430n1Xdo+W3GsYNiJBa
z6KymFgMgnE7ytmIKVZVZXOogffBfzrSbcfJXGY8Ddbdmo3MwlPwpnAUJZp/N/Ei
x2GKHID8d4DGPGJIqee7frr2DghohUq2nAkq80taav8ZGP/qmj8zxE5xEbnQc4jZ
kKFnMGwB3/cB5uXuLiMo93dai+lWSkIU/MrJnBvtIKYLH/c+8A4cDNF5tdMrL2bl
/VhW5lnRRuSJGBvAqfmo0hf/EK0VdUc+TyBUYYExrp5bnP4yB5NjrShwsOZXNAF6
jeAcGp8nu9b+Xr9qwmuouqqf87MzFlFP/jtiv9wcy9XJq3SdaNZktEA4EA19O17e
bHmMlmfLwmdGG0MQ7TB0OoJ0acd/EMD5HpDjRIHmaBb4FS2tmzlXPUiH+/CUeQ59
l/IBraHQ1w2vjF7KVIkyPOC+2Y3YUaltlD/fuqpywrCsh2ltEGo3JgtXxQzS759/
yq2Mvqiro3u4OJ0V6ymXnRqdwoZ6lfzIYFd8PpLXtkm5Iy/lIaufKS0bHZOc1bkV
3v2YMv8E5A5f8jA5ld8LQonJjMMPIeVXGbaDm2m4buiapQM9Z/nUBhKLKmBtQi9N
9tsn5n4mvjeiXvLToCG2CUXVib7I0ukfe4WQy+4C3o7Nx0wVC68/GDH4rovPUZug
AQsGcc9BhhyBpBsmxzeAoORlxhaYn+M/GIKkeoOJWMW5AZ7VJiOn6iZT5/1hj2zx
8FevsFWuk6xdFIt+YkXlXHYrLFpdq25ySX1l9eax3w+b8fx5cTUUJjW2nV+u/ChK
wieCFn7cAVGiSw6SyrAWumPiH1eyp1hVRLuCA0uJlil9HHj9IPVkBfdd6PhKp5vo
a9S6iVchu/+/bixXf0D7PC6I7tL9Ykx7AdJOeU9zvC38Xs2lbAf/O1jl15mwg4B5
W/cgzkERnF/f+S2PAopM2AVJ+jjJsYAJkuwCinRowBhNS62WXVPy7a0ZgXQTQA90
Zt/Bm1JpOs2u99WrbjvYEjAf7gzRqjWbZyOz8E+SEXC7EtL1eV5rpzXcflnnEAzZ
CvLPmny0BWra05UL50G/Tb+qmdSGw5Nf9NxVQQJUqtZ7ICc9g0RIVUxzm5GnmQeI
LIaQDSJguyX0I1fg8teid/Ov8meKUDu+S81bpr45T6BH5XHtdBFUZd8E528CJjMT
vDJ0v8QaeSOc7o+PafbumBUBuqdHSQhysJPDQt7YxIOz/ECfvEEBuYQKalOIG91g
6nm/rocToEEJGHgkWBFHSuQyjds5cg9lCUGemmfgBPQaAhZ14rEqLDbGELORV1Cx
Dc9hCjl1+rL306x/ACjR0dUr/9A3XaCUOBWM0yabfZfSo+mDxX1EDtcGNrb0mOPs
ubexLEhecEa8sr2cmd/pZjP/88EGnWm4aN13FpFXCNFKYSHI0yVICMPLfDqvrDKX
DZ1jQrcID1OgOj4cyldBc7TDkGVevqr3DYFcfYYcBJTPln9/VnIzRPZQtPxodDHZ
It26WP0vJmXC9jD2LjXxc3tg25qfUi9ltPqRqUY0mgO9t59Raq6iE883J8a44I++
gR6EEajKcWKqrZ6aoDW2i7OCqYXUlubR0UsD7epuJkUwV/5jv1rRIuqCCDTEqLfQ
XmEyB9eW+sQRAuEOUNEDOv8mNiI8DhLQNCp+4PhyK1AHaBdQh7XOKwAS4XAlSGbY
ayIPXIyu6py0NZgHM0zaaVAUFBU0r4WR4fxPOJW5sADTWHcewQUHZrcFsEXyaXhf
lUdyl2qRbrHTjw8vAHseRg1wi9HkAJW+X0TfqBVyqCZANcN6HLhIdQT/W+kdqOeJ
i+bQSi0GPcNGj5oJlQ5GfDRh8WkDf+hPngkAOz/GeeVtptQ5rSHX26gbeSVUcSeZ
Q+pjQi4RFTHdQpyETGyNfWlP81d+S5+DJ+5x1ZkRbnWXzAZc53x8oWDFrzqodFGW
1coNELssEd7DI3o0mtykX9lsYBjb6BrFH4k+OEu7tUDtU00+LS5xVgEJG//r/aMr
kDruGz7FX4BjdYSh/9gMujiojfQ3DtXtvtAJjUXOhSGBVUpJdz+S4bnXiMih7w+r
+0+bxjZ3P1aijmfZQnLwLvawJTAMBlWXquohXrlDPmekZ5oSWtQffyaDT76uwqQT
P51hMPGV3ms/ru91Tq4BoOe/wanc0nEGElPoQhsc2z32wf8Z7ErIHTZuSvfEjt7l
kJ0SYaBZaqOGMSa1v02QiejZtSGJYwyzSp5Gg90FdWadVKCvuw9GQsMm8SRNKTj3
u/980RTv4s5eqjocbU9LZr+hwooLmmQmZHJ6ycLfHPsTB32QiL8aJH/ItpI/0D6n
b/CN9M0veLcgEYSdnec+HGBDThHsCdOGgwL4j0kVx+NcBf7/lpUbDj/r9z7PnXfz
8hvLQ0n6Kv7xUDVu6Ugi/c7An+85HVKNZbbkGfpq879YLnL26WZPxe0FhGvYufj5
0Wq+TxQoFYR4I28L+UVIJhjGunTFnJNGgHidnzJBTTByFJtIc2GZVvhYdKQlFw6Z
W7uhz+AzX2cdJE3s6yoFeyN7cvruVZWBBXwFeJ3oTL7Q06tDhb0O59nWmHiBCeCX
q4s+zVLAhwpnqITZ5u+z4E8GEC1fhsOO07ajhJ2YwF8XIDTvcVn8XxVlbuATUoFm
E51Je7tuxCnBtgGLwRlxYRuu4i1lnmYLL+hdfY+10GsOHgf6+QWYW/1kedHfQ8rC
kzq5KvsQ2jGpkblz1XiLL2jwGNj/ed/zIGC7VR7PZFCTdj30IGL0R8PYrPrZZmJ7
dGKsaQPqbJAWIhVR1vk7S8+LZfqtGNUEQgsUGV//s9Im1isHpnaM4MH6XE4paNNJ
2hGbSXsalpDEKf5vzLwoHHNctiYUhB32QDzF1mAXrrfnbGIFRYi7Ym2MNm0C8BiZ
4h5DSpFbRZgV3M+4GYRw/NY+UADCPwJ7fVayiVg8MyPyWMY5NlvmqdUv4NaCRURz
yx6VaC9fjrH/inWbrFr/SEwuL8Ex/sh8ERoPlE0IhF8ZtK2uJRnSlciJhANtanj9
7irEAfrN/afVhKZBYjcVS/XIYTTo5XOz/EQS7nrFxcay7i1wg8TSn1hR2v/95exP
vJRrTBwx/c0fY7yB3t7WYdbrc4pdfnVQMtYvz9EbNfR31iuykjVrGzZ308MYZn6L
qLTizBKd/vXBr2TKTGxQFqXZ/NLTCHN8hPjBfWTNCIzU57cXTYNagx5O0tM0Xli1
yqObPnt7kLUX8UN15dkSFLJliWbueMKixIEqywXzoQ52X+vYOZ6T68PRJ2knlR4D
Vs7KUIRNAMLRBzpWNUWQNCiY6jwzNsOT9PFLHN3fAMiDKsb8OwgC5Amwlcp5e1m9
hpC99XDtV3lpFXTDVvZ7ygVi3v9mESdyfThvAp63s2xMlavvghZr1ioZILjoFPHd
lDgDBFwaNX8kFVpm0bM702TBZoS+weUW6Ejz8LZwh70nfOK/YT+3arH7heoW7Xll
ktZSUKJild7j9FfJB3LrWXL6sZnpD3bY2JqUIIIG9varix6tgTDn8RKSAHNx3PVp
rwIHtwEYLuocYI0c5+TP1XA17963pAFezzFk6P5OzyVZ12WHRVnvxSPz+VHka0IT
UqTrWXyQX4jpp8dygceicvbUS8RdZ1K0WUKtVkQKsV7tHXzedId5rWHf2AfmTaGC
Z0DtYV2+fhUKx1n+6rknIIrMBdr2GZdEjRyP1f2ZUdRxpaL+dKU3BCRB//Yd1D8o
oLOsFP08GUV8gJ50lHOQjeuQ7tjzpFUQBGnZAvywG0aI0ZVs72XLX5VwTIn/aFi2
4Pjg/q2DTA1ixrCVpBsKs3cFqbh1wVKuCyTz+if08ieMcbdiq2bUpTgJJ4qxZ4GU
6G1Wtt8uPaDILBM/LACNBLTz4FKi/FNX9CY5rTWgSB538U49Swcyvtkd3Xaj5NOh
A6l7kRdZ+SVjBYHS1VUZ+mKwaMlw2D11tkFXxF0g1ki0bvk8unha80tJHaweszaB
zC9JlGhxilyMJdXOa2N7U0UKYq/w/TTBmFmze0KOqST7NIBVx9k1UF42WUAw/VqO
HnSK3g27CGJSbIXGlvls18ZbXlcZ5vtiNMWyKzbq6rCmLCuUtM21vwVf/4tmuF4O
1hojlgNzwZeSpfhlXVLqw1PZNXZ5BNo7dwqAh5l+/g2sYXKqKLnkzX8zCbyCKaW0
odhk2C8qfjYZfYfNINMUEMW8PwEtfNRt048m+wAURcXglKNMVcpUGfjwx7KV/YoO
JE+w4aikjschPs2zG56eBPF/tc4UQKdFywSpunRIIuDRfS69lDFqCJXWMDSZlnB8
uCvoCTBJn6aArW/IsaCGTByzXqonpkum03D4JVOVaGFK7YZE9SxbVfMiLcKHoh7k
mYfq/YUIzod5D+qUbNCA7k8BqeSKmrI/sDZomGj1qsuGyu2gaUd8kqMFUko8ExBx
aPeOmdAtz/tYbmmoyeweVcyRCCbRLgAG/0/PuTKGD39BIyhO4wHoSlgd2k2EtmCv
Ndab8eZtRG7rhq39JxMKgWx8Hh2YdUUkCEoqYSo7TRSFUd3c9SCdtkJ577cSNVuC
SW3U9kMAZuKLG3aU4VdrFIVeAbwqBkqUhnisG72LiB7oOYK0xaiffZIouj/nJ7Ua
/3AC2cnAwrifSt9Mj3FdgRJ+XK9dLBVwfNN6xAh74kZzBupjD+ykA5Gk4IPrU17E
S6aXWXCLrnFvVhnMIpO2tNyFhoBAVA9IHr5/3QrhEgZcVljBj3cHDXZn4PRY/iM/
z+nmU/F9H1AUZrPRgSL1/2X3CnPrA5PlFF1tW9RRCMfpbNR08m9cOLsx+nyJvPU+
OopzxiBmtbprjbmlmXR3vgmr/ZaQyqYZb7nwXNslQG8Fsj6QFy/ou/bkhdEB4Wwy
GMpAP+D/3ytoCWIcYxRjgGrnXlhl/rrXHPMwEUWGysuVYiMyXsYboPm77tIglPTm
YMrSXpY9um3hk9SpveTLzDXmHYYDfjQ/HGpicgz8T03PuDpAP96WCoVU1s27X0C1
NxAkbNaP5pyzUn7bsnxLGEKrgic3tWKVolFjwV3eleDR31I4wwe8noRq6Q49L9D6
LaXR0U0bVQs2Yo6Gfw8cCkalqEfX+a13jFCSxcY6ZHXzlqABZOaRE5VIRRAhzh+f
CltLVFttDJZGPkJgyK7l5zjYAfr5EBUW6OoOPxs4aojR6cU/Rs3/WcutAtweAQZT
ZFAnDhU6obgbgRNHfDXicDn1DBQ0dKSC3sFkinkqTyea4lS0g4BKFbhrFO0qqvZy
urWU7MVF4pQG/lParJkzmlFUNYfqnLb8EbIxAVn5Z2fYisu0pe1jhaqdo1ZM7qga
MlBkfCQmlJaFqXbPO2x0HTbp4uSZJq+ov5TMZ4nWOYaGCadG9EOxBFQ1TLsHzv/V
bEo8zriuBfstm/tCQOOjUQHpIaMLQEOMw/+6ZLc8VAP1Q6W6Srcn23lFtpzrls0a
dV214jSrcr3ZAXFGLtkPMn9k8aczgSUv7QZwUHSywKsMBi5R0TVVbvndoad0iz/+
utMWuDY8qAk9g6G5Q3ZJEiu1DrFPLenkhaVjv3GAkyNmWfep5wEIg+nB+fMPU1sK
TiCRbHSGQM3GDUrFMKWLOx8D/QlvJxhBRzKHnYD/LJXa3RqF7likvDOnK0Q1l0Uf
hOZ3ONa7WXAiebzwQt5ugwGQTn4LUh+i6E34oH54n3m1iznm0v+5xMyBLLiYUMGV
KfhDu5uOr64rXa8bFWXiBkmQ7XSjgGVBQ3pWqnZ9/ZZhvLKDHyglODJO3pHW9tJ0
zLWFKPS9RdcspVgjl4fSGXCzGy1nq+kJzVUtEgVzp53tEcP1YCyeab1xe8uDi8UD
/LKmBuas7cNMhYDKYsxiBtRPlji3Q0k0FICM0KfsSEPk/p0hAoksIiuC6npjsp2N
WtboerepyNpDBGYn7WA8FlvnVy5o1vxgCVAudAOKhs4/Xz/hSDcQLxvflwxXGDH3
2eazDeg8pV00y9PRBnelQ+4dnmcM80YA1HgLETMaGfIt8+XPREQSRm0OXHPqb37R
RCldQy69KjTsbbOiXtnPXeuju2tx8KXF2dOKRjGsCYL9gX3PgmJ/rUHlqnviiBer
fbF7zDFN+WMD2oa1najFFa3RZgAHNesfJigpCJwHKsxmk6+MNqfGp5RhF0IPOzlz
+S3fvemomeauWkuFLTdb8HJtejxJ0wPjeSSjbsG4y9dvzNkiA2SLfse20nZmU8Dx
DlmojGGBqmiuSgmMCsqJtT3Rcq7hw6cj4rMUH2A+59mqxTCnT9EUT3+XlCs3xjGI
JrYncxq3f0VGtmL2L4+l+eAWmismFbZLIebLYU397SVz0WhF7x5qsWw9D7oDV4im
r2Fz6VWyWJvtBkSa67YA/JynOa0VljNf/mASW4lOYXgZMc7MDTtOs+a4X9J//ksz
s1ammiLOaWUBCu3Xpb+vQJX2KZTdpRoNe7qCd8WHGmBMLzbn9Uy/MqdbTJFnnLJF
DyCh6RXRwr7wGZiQCFnlMRgBk2YuEerlsPHgDwrf6sB3Er6a5MMnBrmHdIEuRAPt
oet7tfNlREkBJuxhWQAVQ+dv6ea9PNOP2Kd9u2LYo4NZA45AQFQffjt8iUX6FEUh
av8o0Wp7WpV34dDofVIgNfz60BIM9AVuorpxVtiIDqhAz/MlbQxoHiKMhFsCHlCE
u0KyvsUKEY6uqKNwdSZxBL5JLm/YxQR2DbNJqeDLDhpBzVsatZQIJr2gjzGsBSx3
iq1IzQlfZoLyd32MuXAV0FW2DcwF8+YwX+6PdZtB0ZtL0RYTcls8lOLdl4ob6iXU
tQ+ix3sRSrDtwXpQlE7TFgLWLJPFGqPb4lI1KKsUiKo8g6dkyb7SIwARq6/I3R3g
4HD0lnvQeUgd9JIXx4OCrK9XWS8ws1D/E8KPfkRNmuSpuO2nDj/SWjMTID7CQFqw
8kulSyyFisnDoOxzVPR7FLFfErWr1VVkzPc4u4AEX2hxWRAxK8MS2s9r3YRC/vEi
6IzF8gAAWgCxye9YE7MQb8RlYhT6v5CbI7nwv/3EgTmHUiIlZGQQNUq+kyHPMvOk
Rcig4LcPIqWgOh+0iTuLeguPhXkdjhEnHXOkVpp13kPy+MXKnPaD/vNm5UUwnNYP
xFJm0a3dr3KmsCIO9gDk5xRDvg6JAkJb7KhPcwkIvYkyngKBL8HGbq0k0KAnSicq
lxUcoBd9+vJXtTibAfpSVVmjOyeqKR4le3VHqVEuJm3jaN1AP7v9LwC2AcoWcY2e
zVDKFeWmsZdid5UKiLyRR0+9NiSVYoLKWsLDDw125WLzL0jf88BC0KrZcyV8vA1S
pPARZPFi6AjCNMYpAx39Ihi8MiSTHqLkWODTuIDdxt43jXBGzassLCPOTh/rWDyg
M1WipbgTGQhBiJOaaSGbXJeL2mZRhcSwaOilPGF1fq+QPiffDZNDayK1kt0lgHy5
6DWjV8RX7PELkSpY3U3V/WJkm20tqlnTRWeTkwTLO+pwp4tNoWJGUnjl6TEesjQ5
9BZvnbOTcf9vtMZ+12sqCXOEUNoYTgWNf1lLGfQfZT1pi3k7EfPeiQzD8D6RTQ/W
u1HQE2zL85ofcyc9AD1hhPctc8y4ABsQ45Zwcbvc/OFUmc4Mb/lJz/re55CskODB
CcnuspQlrtRMKAcmMv5D+hcpQ7xYf7ZM/vXADv+Ypdrn3xH6TZpfeullOLOYfeCe
VWQBWrIXrJc4nu9T6eQ2OAZEyQb0ENOO5zEDFsNYKWT6/eN7RLgOLyO73cSg3fzn
RsIN32VjSRZ92VHttucc/MdQIModnnDJF7p8fU5ce1zzvwI9Q+d7waSjCtL0u4pc
lcFs1uDp9VgERwH5/nh7iGpdBQDFO8oWFwXKkPGcMoApgygGUuWuTSQhS8RaliE0
g9910LnikptzuWcXWy19rjD6a36BcvHoz6LxM5MplkFAwW7X+YYqWFoyTg+iJ7DS
+GFY6fniGPv2C6nguusOfhRMypfjrX3vA6J2NT+SY+fS0BbyuxedCFkJtgIn5h2b
QIesVLo5VvP4kDyDvIyhzZr6NPRzT89knBTKRv+Q44DuH2C/BqFNt6oUcx/245Wa
EfI68AmX6S42b791s2Qj44qNb+9hzsyMEIaDQ1Saz6gwDZB65O8qRTJYXSnS3oOm
NRjQCzDJZXRUd7/E8gIgfeeTaTqQjPfwvPxvLy+/YeWkeMoOFy5VS6IQuLoOzCkG
T95TUd3J+zECijqByftTrIDrOnwhqBRj8DcTLxRwCLdH/GcH/a9HQkug/j54pfIU
E1RU5kzFkepQZ6ugsw6+7hRdtDjFKnc2k9Loo1LfuSq3sS99lE2MWFee+ykzpeIr
KhBYSDNOgh3YfcJMrJ0VxOVEsPAWNLF7ojtpXOWLEw3EGD/zoswnpyVGiGF4oD9Q
4+9HZ1U2VXfZIM8pY/dn6qhflnzDHFBI2FkUfB1a/c71MpuU9vVT5s0cQ9wBHvr4
eTiQl9smwFu3DO4oT8wXclMr1el1fD9nBfAn7/ab74QtxWIMW1pSGRXoRa7L6CSh
EzA4OdsrsOtXGa2bRuTejt6ROqvPu2kt8PoL/wb7KtPrHNOtU4zwryDsTJn5BKyA
l0apiWXmqpWteDJmdiseEDI3Q5pQr4t+V6NdGSOEPwGAYhq+Pj8/HyaDabmQcmMa
oKGunV/z2sKYDH5AlhZpMD1UgMtO/D26rgWK8sIDuul//zJtt/iY71vxx/BBVaaP
ViavUD7BXEb0Yb9zav2rkRRsna06SToZybeNAQj9Hv7r+bpLDJCQG1jXvV5NvY57
XV2DeVOTGDV8yqr09f+6uyJnNEaDf8x4Norpn8Fr0InTyCg7dpqiqCY2u1SMKeMW
DTaVK/UM8o8h3VUNbdNAo8qrDtP3aOpWtEVJ2xuWe5a0s+H4EwB3YgJ3EQjJkjaA
OH3MkF/Ks3ZTgyVK4491cRvtqpeUJJbTIgWs+RNCvitgZZm+Vjy6/Oe0oVcgKRXf
0tsO7B4JknniBN5+mhicFG8nkhmoDJlwerbABp5Z7d20jjLLbESADrVFdzDqZ2GC
mtyMahGFGP6aldm0Ln4TmdWYhquR4g+n2v/1TJyPW5o5wvgsOZ3zu9RsSf7fyKSz
LHHCsSiC0yKP2rZbgC6XP2WJvUbcFFT8GEXRqIprJkWQmO2yKZ1BLn+T3asdSdc5
08lwFq2Y6xsiZLJ+rPi9XeRzYVKs+bTbALZO14OUJzbnEJLCRm9NFlcscD0FT3iD
sV/nbV4Hgkrg8d4ltsqMuMQAj+OugO8B+Hfe0umHHu8LAUG1NCTFPzuceKvVeU8Z
2kcyu+onfPiavL3+gliZXaKIBbsH9XP5PiwO9kZ7xaHrKq5Qxtf4WFsLMNgvIpB+
dsLXimYZlA9UjOm0/6pslN7nawAgZKOtXOXIRj4MYODM5p06P0QROusa+Q3nmqfi
EVsDOVR+b00NXRlPWHkmXNuc2V3w63rVRNSHI/B7DlYy+802taff+uIXCP5RyChL
IhSrNbMEVyOafqjbNSFKJEFtYadAGirxOnhnMEOw610jG7/VMohoWBqgI+UN487V
LhhTJeEGZRjWtNk0xA/xLL15+9e/dJuJbvOoQnWbbMH/QdihXJ/PagXYQN6GsiO7
B4DSeZJJzIVav04QngXaptbhCAjhRWGDu6xY/oeKkJJP82VHJ9W9CwQ5pNpT17DK
/adPnz485lFPo9C5onnC8kX3I6zqnNhaChyJgfkoS5UNIhfTaNdqNn3qBikTKggW
3IeuEW0dKYcLzgDDqttos7uuIxVpL9bKwVtMzcDBGnoO0GuL+q3Hf6oDC9TY8gAa
Tevmx8qshcZuzBUimWHnkl4SdzuR+3cGuiMj0UHwT3s4Gh50QhTNSPUXRtDWFX9t
PQfC6QPk9SjMHuwXwO5d/7FP00o0qDhN6j4KzJ5+lFiEtt5FTxLUTRux16q99aJY
G5xTv3DmPynT5/mzCPuVActC0cABNoJ36HenjJ6U90gQJWZ6ZEuwECTJVmXC7+ix
D8HO1UopjzKQ9ijjykJaMThvPTD78nhfl4C3R1eO7AgPkRG/9wBphIPnJdTCHDvm
kLLnW8gDLkjsWpzR+1VKL6CqJE9Ta9606hfo9Et+/Ws1MGApVx4DGYJ4iE5B0LcG
UW5BReTTi8W4tX+YDtz8CAOH4xaa0zZm30hCHouGYwvVwrFfKUvaahlIskurriS8
Il4cDH6e2hnldsrZhyGqi1FsQmuJ6s4ZHQIGDKkPG4ztzcHpmGW8kk70pph4cneX
AHRHVh55pPsis061piqksKMG1uPDCuKd0Df16J8m3Do2RKj811Ttbv9cK3ZFF0VN
xSqYZUu5uD2zMcjBeTqoaAiK//ktQBfatoCgYSQR5GhEyjAZe9hu/zRwjRUNqGzA
J0YoeNvL6YxQS8ituMxDOPnmHftnQuJ6eCg3bVy0Rm2iurQj4rKWUxr3wssyyhlb
P4qXDKDY61PDmff3ZA1x/iLMkolHaz8Je28FslvtaelpQg0796vv8WvP3tHCjKZN
/WeTWDuolmZNrTYM/HuFROpxKZ1EOSKuMbaskZdSpobWx9EUemV2ivteUaNMJeHm
gz+KOHQzFk+wt06gGzEy1dp6EVHbu+NJQhL78no0UfL27G/7QQdvziIVMaPvE1zT
FTlhcb5zjvn0rLOlcqIEFSq415xUT11Prz2P7aT6YySC9jw5hPx/KSr2Iao09Ecv
T5twNQbM4aP6mxgo9bF9PM24/yh4AeLT549cWB/Zm+lRy8B/8VmCtaLk+frZOkGl
N9QfRFPBoN1JLdqyK/KIDz/UaOhfXEwvdIggfSNK340ZrgzshasPHlo+0Kn7nNCu
NjcS0L9pGpAT0ounCWmKS0sn1O5F18n0bvHKqW9z4CQ1xRygIP36CdHYDhAnVRd/
EMh7XhJpB5HhqJXLdlNb8/mROTYJxLqII7zEdvrYoXliXxEUmrknrX0tKq10UsJb
Itpl+P4RCgN530KuqdjmFcL9owyiQ+9HQ7sAAB5JaxhBG9MjtKfR/6E61OmPfrCm
ylSZ6k49SXkXvJFdQKpjSoioMoJokvQcOrvK7NT1du7xocifeYX2hB8EAAj4aqKg
h2hvmvFUKxqE0n138Yt1sgpbLxQxlhCBd8FU1UERm36izsgIDzelkUaiwBCm4Kut
N6drZi4rS9kcFQ8EVcRO9ecsCoUrU29RJg3KxruSL0dZoZZdT3cb9sQnRj7zgvmw
Y4PFbCfCF0mDIf5ENIcKTi3j8znWM62PFKDFe5cpY0bd3mfDdsrdH41a9kOx11tl
h2+8NbILbGZ7x/12uXoIVhAcT5j13BgTehZH8i5p2l0kUUjmuvgxk3nV56QftMBj
khD2oF6LvL41Jnn0hH2eLYPPk8l8LmC4Wm3TZQyGPlRKn7iR3BemsYRC2224vrb6
6x4AwcFh3YxB/zR6b+baM4wsimgi4RP2Nal1o9NnEQ6B5j+fQIBxSxBHyo8RVpAq
R22cuK2CAwcrm6Lk5r6pd1QV6iKQ8GGqnG+gZheIOJzPgXvxlc8p59fBRmXQy2g/
ankYccT7tXw+bYdFqcQjc1vHYvoaa4JlebZhriOUeFZ9P6nmMHII4NrkW7EQ5rJh
pczLC75UneGA88ET++ov8kqjdHtaV+LUOWw/VIgNtz+JNKmAuECB8jJOMbcMX3kY
VC5fHDaFIXq7Zm+HXMhUZ02Fs961HY75QlHFDjWUnBO7CFH01fTP7psD/SkjF1lm
1m1vSwJq0QMv9E37m/Ywz2FuwUhk5wwoyrWwZjG/IoL1ZP8nRpoF1ZmHxa+xdOEt
faVp8iaev7G8VruUseHikw8IR6UdQTRrHbj7AjSEqOffZ9hbC2rPjUDpkkWjrTzT
o0m6w/gv+QF39baaJwKjprus+9ESbhb2Z0VlDWsGOMlslinIJxM3KSMnnqFCQZP8
9powlGVJBa0lwKp2ZYF7EkDCI8PR4YA6EQb1dErrISnFPHSLhbHVwBdBOiO8jmhG
lxJhQhUBYKPRzqH7ncatr4EkpMP4DXr3TSbA0qhxGS/REmum8oYxMkZKqrY9ezdv
Ihh/UrVOdLaa0prfPSNr8tnnFsXVITNlJsiM8cojI8u9wM3DAeFC/eIy505pFHRV
T8JC4UF7W9ILMBAJvw65w4/wA8zUWnIeieAz/cc8gFQo95pk3hoOeUbu9zrDzAIp
AxSFqrhsIzPlZkyLR0re9HVWKw0+wxdUIvOw/z8O7eJBV1RGm6ysgJorKl5sfo9O
SaQXJgQ7TYsAYn8g/BHxj7wwGM/1YI3z8c+JDEDOsHyeKrPAlYrbwXjELyL3/cRY
LJoY0B/qzVPUcs6hKfSJT3rp37Obiwgi+vdPlxu9HsoKu271baRIzSwmVKNvbaFa
Phx6wxCfIj6+ci8wFAdLhH9m43xqPXSUensEWoBsDf1vWFDj6U4pGH1C7wgC0IH1
bpC3elXavP58OeviOGozDHO1hZgixGGjwGHE45XufmrhdFu83m6SA+O61VOJv0Oz
o6AnKpNxIyzw7B2SELfft3cqZKQ+YjuFHy2c0xEIrA1R6eNcwjt87nh6eruHtV78
OqIcjaa63sbzh8p7S5l9KHD04scouemTFGVV29PX6Kn37+SEu13LjQt+dBIdRIOo
EBobBwbbBwjwNJ/4eR6YtqL4D55pKEamkc3FzbIwFUCAQZitnvxZPl/mYucucIgB
CeBZB7sJ9RRLyshkCFYxx8wz6Q2+JLYNm9Sv3BWC87g222oPsP0mf9t+u4mWGO3H
B8bVIYX7yiCrN5EPexbjyEY+eanwhj3fp/74M3DLlNNlPnJgqmiunLlB1B2yD7gE
uikYMdqTd5OvCv3Zu31ziPsCCB1BmGV3AmSebdFyAMrStGDJT58sdyXGDPZeYsDW
BBh3mnaTInAJ8Gap4ZA5Z+xhzBmeVzhCk5rezAOe1y5fhhQnus1lBmqyxqzzpsFu
2PEMlYfeVpLSUYoCOMkvjK3wUxLCzfihBjWGhuxPXQ7w5Eg9X9urA5vxBSeO/nGN
IhsvFmx93z4Qnp2T2ujQoXs7qRus4IzTnjxtey5hYisw8M5Yc8niqshej1xl2fWO
XAf4Rt+LB0voxL/UaqPz7xRA5JmxI5hM+p69lG5qF/+u+fIxNf3+E2Lh/XbDeO6e
6cEnlovGQwd0dOnaX3DAhzmNMK1+nEaY8EM40xZ/bCvCFFqmi3jNurxudDrpjzPu
4HH+6vx2nHuR5fUYCpVI7SGc4Cu8OZAQTxu6+W3MIjXWCdcIjt2ayS7kokjN+4HB
ocg/TSdFECuw79Gr/+WnLAu43/MGpV64e7BlOr2LLdOGNcQvpBnK+xHixsZy2ZjQ
dO3U/Lq0ex+AKF35Gecj9wFjsUfFiDAuCrYChGoRbM5LqrrdJAtNdLxPuG2zCC+G
cS4Tb6fwwtDcz9Ih7Cgnasq2BH6O4Ju+HVDRz/Ljh+LHskZaBIKMoMFCI0NopYms
czr4JZuOBCdxILnVs6/x6yiPXhOf6UMkABHMgrFwQehO9Q0nqqzUbO1mUyNfVeCN
SlgNcbz/taBCPhgXWyfakoqqBKBaxIQ+aZOtg7aZZw/sCZwxAyrdB9thzWWHMHwh
5RYerYfz2DDfHsnDdRaMi0GgnRTBIP3RNy4yrzC6jtuGmjM7SUixNe1HbpNW1naI
4shfoxdb+lGBIEgFjhW4GBZAxDox3bBZrFkSco4+QX3omMW8mQt2Im0pdhkY0CB1
hEkVqHgQRqOV+z7P0hFB9eorjWuCyuK317Vd5f6X6+Rh6OrfWQKz/AZA1ZTHma6/
w0C/fYryyaXfgPuPDZ3FEWazGOOvAAezKfNdDYC2TxcIOX0/QLW94TmS5ytk/T0X
RAfNB0aYb0WG+N7nlrZ77FYWzfjq2LCCcklVVVTpY+jG0i5ZHC1+C/LO+RT+1dZW
rgHFypPWwmi28U46tw5+xPbCckyhG2xmjx8DGcjl1xRcvOyLetLLQs0iV5V5ZsVt
RrX7TnA7C6BKGtmrVlPASeAq7LKcHTlYTnJdzmIxuVNL9H32GCrTWI9hyJNo5Kst
RvH7CQanEKtn6VMstemecw6MSRJpwr+Uo1YFISoFSor3hSed4z2bQWtSxeoVVPW9
o7FUy8Ar3KIfUGyzc7LtxGjWZGdDLXGRCK/f2MFtDruP4/3b1THxTnKG2xlEK1px
z0h2Bz0Tiwi7VcV4RfkqhFzgh8hhMKW8J0ZnvNvtE8ZsTIjFO/RqDMCslXs9/Emq
GEyWCdoJ65ndPS2rvuTMkD04N/fi1bkUax5loDCuy5qf4VIHNbVCZG8szZc6rqkp
pXGfqks8GJhzs9XYUi5yB7jiBEY5nGUGZ1/ldJo+xhO63JJxELTVM6ebuZKfbvLJ
nbLDrLrcUGR+1Pyvh77DQpAkJSJrHSt4+x5PQDDwpH0igaYiZcKLtvIVg+MyYfNT
RkdA+Oz4YCujlEl+eVedEHes5U83ha++zR03eMv1hLRpjd3w+bjqajWBcG6rol5C
hTmdt4W1lbx1mIB3+n9BbIns1tNLj4cV3Hn9LUsU/NLDwovV5+01dGTooujWGctc
jKqEuspB1CYAJ562ed4XWQNscrmIVcf8Q9XNWrjaGrAk4V1RqONvZMfgneXdyCwG
MCioi7dDTUAMeLb/pXaeETSAQyj+esfT1k75qAZJu19mdOXdsctSthtsfJPw18ut
/fvFoiMS+MDa+vafRiu8VqpcXGHBMQeo9owRMqlZlA3ljH3EilvDQ5XgRHOp8RLm
fXAlW+gDscGVIayQFVnCJ+ygta0/sc3cJM6WBE0w4fMaiJkpa+ZIG2ydwDr8jh55
qFJataKS881wb/lYWzpiVUWe+I3u6TSPgLULJGOxv7LgB1e21ibDoBNLjWFALzPU
w4bXkFx9kd7StVhGGs//aFhFJTeciO+d3qFiRw1WVgGFjrxS+E5g8bWiT7ZJkzmm
9I4TLbEaqbaGW43FYsqHT0uFlqlpwuZFqsFM0o7otb3q03VCMSKY8BDQggyT5uS6
nnohar+0RSr4/AZFHhDIOJPEVW/TYHLN2dURunWLnMwPofGpF9UALT3PY1ra0mq8
F4hTyg+Ajd4frnJaqLZJq5Iv0ACIxtHbZt3HrJf89vcVlv7Qn/5okvMjV3bbaH8q
Z/Zdelii96QQrvfZwCTWNYmjUSFcxwxke0rQEpfU2/ChkhASXj81X637NfD+O6Nb
aWaDKKCC2iEr1nbWlSX+98ZB8jpu3b1qn9Gp7yEyx1M6WSoO2yt9FGUpdnlsEJ1c
OnURWtbd4Qux30udpz8kEVPWfKT3cQ1Kg30nKpgrUFPtSr+dcKTch8SVihtd5eZv
olfVU4mYGXOKyK/LWu8I5FtQVoTzc9YSq+RUmWeF1ngnvsnJ0FdkKKYqv5qNALai
6ShNmNBIxBt1X2mujvN5AsGuFNCGphtGVP+BEAS/rlNRMPQ5cp09k/tXuFyCq1IK
r4MEiyKOcjx7FQgPe1KV34BtNLf45tBmjD3nRRdL494nZCD45tGzToFLNJf5vYWS
6AdKGXwosHkESPzg43ThJJI4N4yDrtIDbVx0v+yvgAmZBrJXPtJZqKrZK90wuXYa
tsUk5hE4mfBr3axEccd1exNAgWeJsweNh2v4POd0Z7AjLDABwYKXqXmXBIfgHUbw
pCltRUD7XFGKRB7LtQwJtlA67UC7jCRA0a/UcjsvGqdjFfDWmaC65QxYUSsgdzD5
qst8Q8PTWyqX4Te/4A7hC+tmGh+UunPriNo05SCZTI3a/e75vT2UIkGSTDT3bM7o
wTqiGXZp4fPrOEfS9pcUcmmt1x+onDNRI9nTkz6b1LsMQczTSNoEM4AdIZ+gYozR
Pqr2RoSv95/vwKG4r4O1CdqKRN9PVjk+O1wUk2sGXOmwQOXfPDsSbFEYU5kxGhIm
D5ky+3qZimsEhcNhxFmfJ6dx1wcDGn4S+WCDQ3rbfsolibIjDO2MCMfrFpFwpvdG
b/H8E5Yv1947pj3r7r32j7R3WVvoYbsTgdefsWdpAQ9+yfqog6ujRVNCITfBicY+
9kWjx/8lmB9x9E21WWVLfLd/xitFYLdA5oRsrqwM67wfi6bIj36W90lbr/6QjVbS
Kk89kaNxpQwwZvrACyNoktqWubQMxCOMAecL3GY+2Dr8FC9z9abo5FQDLFdjLi6h
KJ88BdK8LYtDY1GuVr10Jlr2o+FqbOH3bsumKkiYGyeN/yxJ41P6mEHBBcypLlmx
ZsYuom+q4CwiGwD2/KmipSu75AFkxe6Bx0gEaYVWiTKnofhNXarDaSNlXFz28o8p
E1ixu1yX0sQ1odpIE9AtBwb8tCcWbHFChsOmRtFLyfgC2duZ3B6XhLAFYNSNhWAp
rleg7x1tzJ7/ZwOaz5dfK2NyhghQXMZeDALIBp6P7bmkFSFcg+tbn3yFa6Bw3Ssq
+/HOKhtUNACAWgSWcf4Al+KQ29YaqR6Xl7ehdM5FIV9lbiyKrH93bQEuuc7R9Etr
bD2JjdonZdCKTyT++EofTkRRIiNuCWvZQeSdZ15eJt7g2ieKZMJdydYcmIGuitTI
sxs7PIu3Atcb2KG3C0RaUaUSEeMkQ9+FE+CFxNct7Ud+3MZE/lMYxph1pe65xiOc
OvIsP7Wx/WpnLyjOFtSRAgEeckmdtetA1n0j5rdTHTwXzq7q9prWAHqrtdhYDqO2
qH3RqfM78jyPjeYeBPjotB0EX0syo5pZucL+lfLzG2ETCBn7tygb38bPREugTEsR
DrYYaup6F+VvcF2eqPrv35wTNihH59jhK4CLvGMJ0NeGVdqW68xbVdAS7pFJ2cfO
nAhkC5Ohxb1JolLzJ4XEzAjNWvMwOcwIFrcPCsL+IOfHBXMaZQyYnU8+K7U1DHpa
Ykk2OYW1WjKy4Cg4aYbDQmmCKAqPKaCwOW25TENuM1AXF+fVv7klLohZXwK7i2KD
X2Ixu6xCfj0lBI0CBLrazoNs4Zgub3/U0sustRYsK08uQWM7Hc/SQCmiK98lUMdE
QsaAogwV7m7qXXJTJrVC8niLXnmSCovOxZemglM9vQVRnyoV+lPAPFvZ2nHQZedJ
YsT6rQUVZzHtElgQco7o2nWnnAzqFj1J7WPmBSHthDU7I+aWKAhU/sy1Ev3zgi1K
XxTT2btriajX1ICccvM8elGHjP2BVZt517OkvANR7VMABd0wEoAP0wB5F9xtsrRp
5Ym/RB4h8KsbUPu47SGCklx3Uhh0YVvuqtoBYZSCHtiDlQYewij7WK0z+SSrn6KZ
qSCovkmhZLLz3vvnNhrdZyEPn4CLItGel4HI8KL04RYn8CovA5hVuaU1GrK2QaGu
GzdEaAylGQLniFnXhEhFMAEYwijPrngfOeav5ub3Cz5LLN0wJerTjsNPlK+BxGOG
Tkdzl2hqdg6gTm+gWaqcysYGlCKpR5yPMSf9xG19Mo7OXOEWcRFgB+3qaZ1PE+S1
elc5uHJnqr7GFooG7eQCYGZ3kSJHVV4vqJ0oGdz5xE5B5w8gsI5EMb9FnPoYsP6e
ALFlGI9cJa3DTfp2tinoqXfFalRCg1PFPXll3qkMEWh9aRtWiQKadGyyihKWHgxA
XfPoZt9/paQ/O27Nts0XHqRrU/4KJi3CnBEBFv0W11Favh2VFtMG8yOlY8LXWYeq
y/TLzVEHfcrVl65ooSVHaCoDnLNfMXeKUItcKr2VO88RbwFGcWNpz5E3FwlZw/OM
80JB/XsluDOhvXXRWMm+G+KZ+OkOeai35kNrKTeg7VIc4Drud7TTYslmIi+laOCt
Uu1MXQpfF59AAkVqzhShSjEuxK3YGekj4ydIANbuMu/pjRTY9lxjgJbuSvisG05/
fs9TxCfC2KRxBXOEXWRaAfXrO+7juU/wSb0i3r54iDfyuazMbqzb8a8IVquAcaa0
NeezTgm4bm0AW9egi6MCxeFm2DEusqZvPspFo/jEVxzq+DHKOkuBE5yz9W5Ew3BL
ijg7LPU1WBoLgvqbcdc8FQLi73g5N2HQXhuCBSyvA1CKGMqARK9gT3DSycdqxyHD
Vu9oOuDiFAx8/6OM4q2Hiq8LpT/pZijAVq/e+IJpQjljXb3br4gyAbyY0DHoURJi
4jpmX/Anypy2OFtY2iCsoT4jXkpM5XcmTDbGb5+ZuIcRCARcGNlchVQdihs403h5
Atk7TgUX1C+SffXM0i6Zr3RiUeina2x3DuzObdTigjox5ogY3A0yybfuYiGBtENA
ZWp8PKg87VJGu9QVb8IF5rzbLsYKznSjJf4I6repJb8OOTHMF3wGAH+/XSknmvj3
ZSDomTVN3II5s1kOG79xlmx8wvP38u0+zW4zYzA13IiqZFDIfABHd30i9fs8FA4u
eSly22yG93RqqE08/ee+MAjc03PqEVlwEJreRfhSoEkDVsP60t8kysM1et+KAMmK
Vo/UBg17hLdwrZGzxu9p5VT5Bd/lWQ04qdXZdIjMJQPMbindg8Mpqu+QjdFmFIFj
7DaGrvBm4Rp2dTAImdsHnuy4SUUq81Pm3DNJo9NQc5DHNL4J/CfqLjkkCVmA8EwX
x2uJoLoD2qDwhIw7WjdCPdHTUyDN9rdodgg3E2TZKbYJ/SbwYdLKKMVI4a95U44T
pTboga4SWlZExEv72GQ/8OL5NC6er7j4QBDEQSTuAXrYge58VB6DnDOVxiVJ1k7J
43iTBidMAifGO7JCEKinVLGAejNcZaFS15ejoVXzBJSui890ZSgPqvPYExZ+bM7D
4Mh3Uel2uX0QURN5qEBsdWcMDPejAoelONlzxV6c9VCH9hU6TmZ1l0tHcoTosYUI
cLtTqa/eRJ9Yq2qFGgFl0SI2OiUy2rreVWY+dOYxHJMuaGQoDOrdusZ/ywHJiGB7
Cixz7Kd1E89xOTIZmrjwQox6ae4QozcQXCv2OQf8RobDwI9l7x83vz1TOxADe7R6
180Kt2i8mGmd/qAI0CuynFPlM9BadNM8UT0YY1H/v6Ypx7LIwPjaTzyie56y6Kch
HyMnEdsJjJM0xTdGaiMix3Jmp8IVTbkKiKSMsCqsRFJaTpMIaZtuUbk4jWYzYoo4
wg/RuS1taOafTVD+y5IBQ2elK94SsWWTMKMY1FdOShrA1ztT3AqIycVF1gH6PIuL
6gA279uMMSijFL6KGgv0LbI7vREmbWrKMaYg2/bFxEhsea9A0wvVsw+zBI+1vEL7
9/ribbQL+3DrYjXKVe2RVMuF9pFy/f0FxlI+KmH5k7DRvN3XMlPCJQ+WHvx2qizR
c5STNGDKQgAGAcLqDfxdID8IEXKz7/lpT6lB/NbsjZdXmYl+AEVAYJBxc2Y6x0bE
SXhGC2uYOI2XuEDQmuIHx+hhkf85718IEzexec3p8+D3WXkdnR/rT6tTFC8JKhf0
4/6xGm3KIBT2KbA0GbW6dEJpge6/JnIxA7rQ2q8ZufiXPmPiy4EA8KK+r0wvjdXj
E2at1nKLanzsexk5rjG+8LeIB4+D/uqg42mbBRwzJH/wkmPxFkzt6XBXQg3Y8brP
9rOPD8LMEZMjeMIdLTYmlyBZFaOgmOP5O5LT7qwuYJ1jbVEaAYG/4botUGTP/ZEq
m9+nJYcwoKgrujWaDxgghLY8BxJp+CJLGoVMTFUV0+TU47/hj/YgzvQAasBA4Oa4
SMz675972aAxkv2d6LHz08azaQk5tlBFZI8+c85f1A2Ti2oxcUhiO1UjwfC00Ji8
DoEwN7VCm6w/lYLqld7qbgbWmCXNGHc5Qh8UP3RhhiOokrV/54/ESWZ3CfqxUFT8
Obk3UMO264BVYG58519khXFJxuS7vDfcEzRIdILIOa8mJgQQgdcuSxGji9I/96mo
ezkKgHQshTosIIk9qpJrga64x0LQ+/5ythATncJqqIEy1w5rU51s6/vtACxZ927Z
ElxkBMdbWboGaOkwySOXX4Eb5DyjQoFPYsTNpYDNZzlrF2UAXmzbc5iTouq+66kJ
pt3G116NYK5BGIiMubq8sojTZOqXwDD0x5JxqM4gZRtOe1m6NS4kodGtL0nXBsos
mDyICJ7+/iL31Udund+RLJB1OVpURlpzruPh91a6sx5Wfo3nurIX0e78SUSm9NAe
eE6hbfGclRZD/ZyA4ylykI6viQr+BHSnd3gUDcMYdr17SWxEbP2xC2wvRiEX87EU
xW1uc+GD0KGAeP4Kl7XNTl+C3VKj3UI1hBGoEYVNnh0Qc64/mO/bM2mm3U6GjsaI
5aHwI8KITIO+Oz/T3jUylblS2KShgrnna/RhLWRascSJaXDLY04/txqSdWQDsJv4
pg1zM+sadhQgROATWY74oL0hOsDOwWmmXArboiYx4hC8NKk3+Uax8lDUZ7UAmevX
hEbZF++LuMkFP/gRucR9Z7MuU/dzlFdzi23zUF6kvc0+95PGi2TjOMbA743V9vJX
Byy6kqPWMIlPMkAUtk4J4SbhJPjnZKudVE0GygtsZPrqzyJVUMSWcQPOGhnTz95k
aBFww5WUWQBnynhABZRXIB/u5FdnHwmXwc9Nu8L8nwdoT1VKwZbH8h+FLoIchYpG
hDHYLFDQM296CJ8Wj1tq/c9MPzVTHlqljAgn0DtVzjUCx9q27ksMVHevyuYMhkQy
02K5gL8riyydr5XemFsE0rFLVF/hyayfiBd4BytCKBGBa8TGhte6AhAUpCzg/Apa
zNLq2gDP0XEQv7KRnCK743iubyJDYmo/+nZeUsk0WXJ+DfacDPXWW4tzgvbL+M+h
/djWpCJApLfPGieKeP2moZCo4usPoZsi7qxCmxQYBf9rX6vRxl/r+zmiU++MU6Ks
BBgNzmeOdOtTf3Q2gP47C3I3+yEDoIUKNHKP2goXckJveTRUWJJrbrvr/pQfcoHJ
QGrlL7/X5pcv3LGRcoGcODa64gqMaqB8ETzDKbZBoTqPGi0cU0mOYojpMO95IsFh
6bwmA/zIHAspXJeu82Q/PdJ8HpofsoImzB/lwvkyrdDIocjhsKlxYODczDgN07YB
4M/PgEyh29HU835h7EFzunR8cJLxW/TVGrWpGtG6d5KygYrD3lj76Q8wWs8MzvRr
msMVmpbHz6uCkEs3iRccLmKEKxjAJTo6DUBhiiZRxFKSa3vx5UhZjJO15H/xe7Av
wbmfOwlA2w80pd0JyGGt9TbJZFE/m2q4LYbVhKCGQXLmeg9I8SxsK+x8023vhnmO
hRSBnUox5kp2Di+NN27moO62KQUeyNSB3gJgSvNs0hJvqG53KJnO0JGQizkirYNl
SZ9xkviW2wk3LaNeLlKwlNVnH5FJDOVi193alrmhkws7hny5xC6xYoBjL4il7Lfw
TeEKJo2JCwpKLsKx38d2GimC0V3TX0YAWpRUd8jY4bT5RG2pWBNyAQ6NRasrLlkH
JmgRC8HkvtDKJwsGzokq9I2/GyKtAKQE5yMlQlVLhVIb8q1PfKPFr4ERrv0c6RBt
DKH+Y3NHPYXXsqG3v7dK3pccav/s9YYAyU+HEpGC4X72cBk8hDK+r+mQH+Ug3tx0
3rVOGaQFkVb7sn7HS7Npvl0iO40ulxf+wFjpcmirNaYDFEBbYmDhTz0wHCW0QDey
P4I5oOFJXe7BPpU30kpY6w7CXH3bym+75qahMr4nQAHxqpPUQ2PndYLzQi3vYn1j
UiqrCNU8LJw3v9xAbOuNofMeJbsFW/82fG7NdRsjBp7RxX+m975FfHRYvQ5wvYl3
EjBVISXpShC3DpW0X2W2uZTpzzovHTqL0AqA6M6Xmowt7i1XC7UkfoCxxyFt0W+C
Pvs6jeNZQ4/vHzx3c/8H7iev4fhDZBzEqNQQbZHODcWsn6Q8coQaBHmTHRauIl4F
o9+wvClQm2G/d9Az3WzA990NCAIAArNI1qjbnGHj0Fc0fXoSvu8p25RYe2pK3bFv
bZy4vpQxvGMyoVZ88FMVu7fjCovda/o+6g0+3ypFzy6SNtrJnRtf3iRChiVs2JmQ
pSoE3lHz8mNzoJ9NxYAu9Me4eIJnWTj2VKc+WsZlvtdZoeE/KkgfHNB0cLUvugLV
36cLbRDBUZBCMuy+3two3h3OYHjseLGdcyLAxz/6EMJfXoUEVj+mBMzqx5yYm4K5
haD5eRP2MiBgNwPqHjFTh/q3wBxWEUdAakXMf0Q18dPKgh9ZIBSK7DBXRZYLyLnu
OwaNg08n7bXTrbFQi8dWIYMY2zyB8tXldr9wqEmMjAHR14p5X5CUSiO3W1rY5o4c
PcoFCCimOcRubri71TMBVxcX2/M+kjcpKrBSu0+Jfw975x8yFD8oqNI/r6RlDv7y
HBfg26UuKtxltn8zrGPLrN7mwjMnHw25R1hI4fiCi26MgpIIT6W4f4Tj1PFU7/Ty
i3cYIp09Ibi9KrjgcA4FTchrTRkuIET6OOgYS+vDnyPWR7DVpOMEm89wIc+OfUYT
CPOJ9GtuBQgYLR5s/UYrei8qb1nHKMIfTFHrZXFoSnyU9xc8sVQsxhjD1ShWL4iN
caQPXV3tSJH7a9QLeZMsh11YizN7hykkMFRwRUNkucYz1ZREE8vz6FVhwYgFRIkO
AdghYacXt+BohxU7fTyDEGqSabwrFi1MJGMDcKuGxc4x+ZXOPuw9AQ6ewofPdQ0e
xgu6W3QZGAlrONTL9U9wRDEXoa/tHxMndonj7dsOQTcRfWQ3IqOJdZas7xFoYlRF
WuTizAPX5l8LA8k+HfuEkthOHDrXHJPuvNFDIW7z+QB0T6QouqmLSWIxfc3zO0+4
1Chn6+lvh1nxYXQk39d6J3UsP9MN4D+LAWZVjNgS6FSNWPiwtWbxlvm9HKU7g8Wt
v7S3SI/D7bToRN18MYDVCXBL4QsAjvW3E5g8QvZvjY0uoLmL6aWhECKcLZLppGzl
539ggEn9xavIy6XTCAB4ffge7gBn/zz88Qa5AFgB29r2F57t90BnpQb6QnQ822dn
Sr+Iw/v4BommFYJbX506W8YAu72d9sBNVUIyNksyUHzgi5PsftEgEiVeTOG3DHVE
LdT2IuLOjOR1QFnyaZLIGvX7+V8Rtuyyis07LUCYye20QeUVsNHMeolq1VJktIYT
Laze9n9iFI4c0pZ+3OJ5h62c34nrP3UYwILgpzWYLpTIUuvFIdjCCUTZZhKj/B1J
NUMB35UttyGEF8SKlVD23yKy/WUratA3RIW/uwqD2hdPPGRs/66vfpXYNSdOuAiD
aXqd2CKlV9XxU2lcZYcsVetsJ875ocf2KnXk/Jw4mOUZkx+jq7cjLgAQEFrIAbiE
fcLbrTcIJDOmJ4xu67jrT6RBNVUnVdpdwfvGdYAM10GuARUkdvpOcWwtTxxqno5U
ukUXfLpzKK3CarkK9H7gbBqOfYx+z9otrL99eKyxFriRxjgKrLqea3YKLZFKbjPH
cDBDecBjzn2E+GIkFiDoq/Y5V+vypNcQ+kzDOM+j0dplVc3AH3EF8HpTgBUJqgQ6
lh5hBQfdPIBTdguyKhvOaTy+rWGxNEqiA7RwPQL3eLRJYwaiKNom4OqCI/jm2wqS
1BcWCVkgEwkTpAWxRchGoIO/isLMitT8He3Nsq1rX3Ne9H+jm/OznFa/8isbKTLK
DptOzAHKVi1fS9tsAbyd0+OL6AWknhR4WimnWyaO0GRjEAXs5FP8uHLB/x5UFcfC
usQcE+YkWDRnbbbZ2MQByIMH/oDlvj6GN+QBF/gNNTs89yvlcx28wJmnOkgy41dz
ZTJm/ibhg+5LRKF0kOyKkCv/YorWWjB7cl5mRvKyqx6cU7JTS6wD55Ae5Mq2+Sij
pEg2cOagXxIs/k1OWs/IgvNAzQG5LWd3QvwBThRLXWWcuveWQBrLDXS94y21+KrQ
USBkMO4Rj8UG1GpayjEsxrDxJodOCIN3O1ZWBbdiQfwKZDAiIFQT4M3ZjIJ5On3j
Ne2mDDwwIGB1D+5fE3CL7/zeyKeOt4X0DSeEA4nv8a83Fl86rLlA2RBiDLPNUyP7
0Ad8uPYgyU+ELYDZulkCx/jjRUOtEbjXv/VJbz2TqaCJJRXTHcYVZmmnvdYeCNJR
kNdBHcCIV7yo0eDcugbdU3UCpQ+Xpun2ZzCNqsKD1DqRhxyyGM8iB+bMxhnOlKYS
RafGT94twPAvjVPD4KD+4LkYV7W7a3PjpDppNnRIBCsW2mdfsPRGeTEkVzcIcYrq
MWSOhFCXJCWgdmKePdpbwXw96w3s9yY6wDJxK0HEK1Z11ckMYJEsQY/OVfUGrNyL
GI1kLBpS0xT6K7QBXDfvrSC8epk+4y1UEiUdV0BX4HCK2T0L3NhaMgK8O5hbuCFP
SCLdumu/uglehz0UmcaA9IoLRz0NbRmuO/1KN7DN3fQkYjbktbmioxobmGRQ4Lct
bGFh7mNUlW+JJvtvmf6iH2sFzSeohhICYGAuQWmrhjCHcN60AjEbCmuuOElDbLoO
ulSWfL4WxxhSYroQx1TV0sVzJ1hxkM2CILF4qsCERs3s1Np/IFw040I7wf0YOgzS
b0UweDvMONMvsnrmmENbHsEhtAWr3LH+nRn169ug0RZfgxpZWGN2mM67uaAnDaj0
RahSruVj3+ZHAgF83BI5eef5DN9+vgyqkEjBgfSKmSXKbZf+NttlxBzusTHs0MF3
WJgYz55YSYJWjL82Pu3B1qMP278lP8d54tBVk/Wgm4Bet2/kFydPxWtXj2mptLPZ
sw2cND6Qs2DjNKdpmXH2Dd8dD7aYUNarMkoQHEAX7Hfs7WkpHVb2VdY3uqj0EeMk
wno5ehCMf+GAHLItPE8yG+uAoyWqUh/FvO9TnuoBy3xrr3ZJf2TWdo3E2g8g/i3l
ivfo9zsOEDr7sjMainLUJI5F9hPgi9nwV1JRyxIatJrVA49ZLa9z36l5Nj1HQPqM
GhFyUQtboBYuiYRLmS2qfenb13FI5HWp4yh2xnxlIpFfbnNHcElo97nQHiigMoVa
EcXtVWD8hJvAYmK5d/gSoFsD6FhPZME7ZdIRoN4NWSCqR54IGEu6a4qZfGc9K1hk
rBROgYukY8bebwS/0CzrYF2IwFojb3IAWqJ8XBcQi3ukX5ykXdQvgcARjG/Lhc2G
1WwYVtCWrcuGiCYUT6pzWa/tMKZeYiS2qRouHS9RJr6WnUY+U5+f3TxdcTaxqS7b
6eu99BspNGyMOk2gwRsmt2Kz/6YEY7yGGcqD0qrVb6EgfPgThyfU0j5h4CxJ07UN
ZvO6ekzgk5XjZtrGOvPMultdU98XdRaMtBhln5pQ6ES+SsleO255lMIUVjgnh9XO
2wA2ZYW4cUhaxlxE/z8Tq8/6/mwqjimsFfpxyQd0YdbYkDMDAZKqRoqT+aEqtZTj
nK8fCwylE2NVxtdw5p40szacz18cPGXUPA6XvYeyaG+4WcSytb59az9SibatLDwQ
SWHRn5JGe7n4oOamvQ5+uoKu4IyMIAaX4T4vNN+ptUg4PO/fIGBYOglCql3NjxOa
EDvDR/KGHex6XlYPOCcEBglecpFllMhnyTJuJy4/Mf/TkOjY06Z+Kl3/VChFLrTf
mrfJUDbdpnLpwkyX4z0YgSeJg3EuA3LMZH6woSI0uQYZbDTzOueS0un6tJKkfs1+
eO4mSdQvgzsLAwy9PJArFcJjyLtREb+7554WXQiVA7kCRmOp8/4ylxXwAYfQ2Uqo
dA9Yv2dbGLB5eMSarbA0627rG2w6V8Sx+dtgSq/4Zeet+qXrvMSkEqf/Y5DPs3+L
CfdIBN34kY2q4Msih//7620zdOxWQLdnmSMItJkIt/SQVnFmu33Vc9ByXsL5IxWt
kOmhKqve6UEzAzWI6gfdg2+b7P398CRCsH2+XVbVRSxo5bjOsrbrCtwGfCCIMC1i
Y9F1o8ZcIqNtg5jprtvf+i9x08IK632ev1ZAy6+eTEKxmEvX8YX44mrbhHTq474h
WLOiGmBm6Kc7oCRzxJFJ9kWTLhrAGC15jGN3UMJ2kjLmzltITj1Mqd3/nDV3pCWJ
PEicPthemQse9CGPFpDakAB02DOkDNzcgYbiNSB1T4yzuBEeW+bmstRBFIIahp7i
pgPqEmcmUmE1BNwZX8Ed0DVtN/HklIOgNRSisdygxQCHD4kICV8h9GG7xLLDmA8Z
r3f9SblHfnVXLzgCnxJ8H3AacKyGrzZRp3LCb81fawMQ66ljfFpEO8Jn2DCNH4WE
LdnHHBq5I3maZ9PjbdTyGzJGft4Yq5ElAV+07Go//fZr/FKMrSKO7Z5lwjcbmwbQ
er7gRN67E23pUqvQyXGjc1tUam3pf5onZmgCHccdTWeHLGvSUF3YeVItod/FQTZ/
mKIqQASULewm2dFIRzspPaOljxoNs+6wrTIgMrNayhbob+S688KTJLJQZYg8E8bT
iuYI52wiDSD5AGCOOpd6E9Kocf5gDRP3pmHR7YVPIrl8ffC8NasfG0TUpMvDN7s4
Ppy0n6tL8ebOkNOmfnmfjYfuNwLIlgiz82v+atWbFozaMY3dDyzFPq2lsBn9DIgU
s9KIA9I1eyrajB3tNTG0mu0jCbzO3mN7Vz0ZAx4oQojb+aY56eIc9KePONvxaE3S
RhQYRvwYaJSX93CraSGX4aLIPaDfLM6jEDXQ7tR98EABlrg1cpHZFeKvwzC54zyg
as3MpOZkVH3UNaVcofXkT3TO1KZkPjpJrAt/K7Vu5hvbC4CRQfJjXjpExGUvtLkI
P2775WUFeTBo9FO9OdLmuElm1EF9x5O8xSb/uMAxBiiQ1Zq5Co35H9xx9CfYftpn
2KgBB0BpeGsy103ax38heTmiwX48C1EmKGVdvtCfMmA0DdUI4Af/6jVzqkLOQ4E/
GlOTaD6Khu3ZHwGJmvUW/SnI1Gpn8t40ZHFXWvBkIQ//1RTjmyL+3NyK2sXdw5ds
KP7z58dXAcMlMY2jG2lm0ZZpQjAmmdBPs0M9wndb1+B61vyb2lqwIlisoNzXaeIW
wcKvUcsoVfxqFX1qtcOKEi2LoJQq23hNoVSDim+MmRtQoGT5gLP2yQ5JHF8X4H0S
hZ9gWxEpJ3gEHs9ZceTNz26P4CfmD+fPS0PBgGbwmQOkAVDkUN9tooHeoMSWsNLK
ZZ9T65wrs4ckMCC5hA2q5lOyrr5ldeKJBIBLMY+w5b7OmxfiNM2mjUOqBT9xWGtP
Yw0HgU8o404TGNNRz2mWKuO94x7TXtUg72UGma5Hkm026upeSw+iHiudCA/8ZktU
6xhA2tG4XiRY+u9RBY4zjAbEeZdoifCzspCNgWditSZOwC8GsEn3wtloO1lVPfwp
2bC4Zhp0uGihAG6hhaAQpgux++0QzIgkKIOl0XfBBTgEAUjih9G1z70UQTgVCWRk
AzWbrvlitdzmayLGIuNeZBdKSb1Wd3uhAexPx0WYeyT7wvrl6+mXC9ehhdjO7Eei
Mb+HWwnHHcfEtKWx+jNYERf6SdteaNqvWF41lBA8wH2K5aLKG6OUBM/wGMJCl1ZT
L4zWZufix+bM310riJ4Lx5/CctIu6jvnvQ8X67CVaXZEhKRc6MPIZo+iqyFmXAxt
1gbY8QDrU9Y2YaMg43GmfKQ7LMW0khPphvJzVEWEw6ZJd7EWyGm0JpNsTHnPZrZb
UpllOkW9c60HcOZE4Ug4Rw2s6T0sLOtft9Qqfb7bs6ujhslkbBIWNQOfUIUcG0wb
vSd75WVP8ypd0lPKS3PqKVZfnQoAmkSMPhC+J2uPiJNmlTKLYMDp+XMPid/b+qj7
EKNd6vvwn3uu2YOYxSS3bSIxGEoGG8d7vgYzDpa0h3K2nceXwD5xOOO0mhifsJGp
DuRi/SmjZJhqbL/HNOLLfcJlXkQa6Dn97zuYwl3Va67LBuhZAEm+LKxc01/jWv+a
TB+2SCaKpxb+Kq/2yjO5EeZZHSDjg/Eg6H2cG1MUFkkiHLODFrpqPgfJZW512lxe
oAVUsDOSyUHE9cGE0Lb5VhRv3IZAPLb2DX9vUKC0pTZyjqlPlR2FlljhGpOnNgm+
Py6zp1iw4p5NYxmWyyXq0hdp2HHB9ZiFv6pIpp4zjhdEmoYsAQTRRXn1coh+DzyK
tvw8qeelvPHPOp2dSdTep4YezNfDjc5cu4nWkbJkAiT+98W+4P2ML0kBhdOrnc77
/OK++kZUiIuRoQQl6i6GR5Q+tXrc7nK1I/Mbv19IEm8/qo4guR+sPGAF7p87e60Q
5QWJ+0NzK51inPIkt4GB9dvIr0i6KGRuixvPMgX5xrHgHlgjj9APTzW7lhEQW73a
roztxQpJow5/a1zstbT+z9qn0AwB9wbl/agqlMH1R3DBOdPO1l8BTVYtx1xrgURB
Zhn+boteOeTI3hKF71CfOywcb0kvesbVNHSsCPS192UerFGHHqU+Mhj9AgYiGRQt
zxkNF7ZFv0QLEoalo5QeeP4SJKf1VqRyR3wYDc/1Vy9EypQUTBJTIW9tHdZ4vJ6V
u2a8vhFjXkAIMvbttgrkNb4iSA1oUtgZ7jBtwgCPngJaB1cL75VceYSrfmuxLOdc
xxWsMbTyquYrpvQ8K4CX5AvsFCe28Tu5TmZ/n4f/rR8sCaF+XxZ1mZ44zpT2g8cF
dnn9OjAycIl/iSbNuk4rfaJSJmLvqHhwwrAkjim9ggDBuupjguMNFW3Hi7Xw0J3B
3EnBwOFpgno7n+Dxl5xlDkdFahlNmdzVcrKGXiBNStoQhgHBxL152XwDrLZ3FBG4
ba83FmCMc3riEB8kHsTLfZj881+81DYnJMIOzom95ZDochlwFzakfIwfi0LpQgUD
v/YuKzKRM4Ml9h/VN6m1uutm7VX3/Qgc8AGNV8kybib285NAD8zagohhbLG81JTN
m6Un5ZDFb0HRNUiWR0vPy6mZm3kF0afwacbdTtltbK1jexUspXBRkm7WeU93YURp
QTPEcxIjjEAmoR/1mVWAL+Z5ma6AZV+eCQKUW+QOsZPTJmdEOVCPffVuAueNpXJ2
DtOPVIXVKHJPXbquVCx8Zoccpm7nEnUy3ij7Nw9r42ZfB2YjcFcSxR1jq+SEdlIM
Sa2zq1TYnp3rg5RNrywRtQ3hbzqQtJ3mT0+sEBBWxbPIzQTcI8QxDcyMYZobHbA+
5oM6mqh+hX2J4kJW/gaWNtgikMlujPX19jo+1PKepcympneyR+APnlXTvKav0y3Y
xuUHTXLM2W2YvmLxXvjnk+iaECe/c+Gg1n4PeiLU3NlqoWmA9eWG6M6zSpGevGN2
HUNUAf4ZwyjWphZ8U+FL9gnuQffYTIj/+kzDQ7rP9DX3j0lzzUXJgNFkFX1Xr8Be
y5Xs4aY/sfxJCQWKrM0DC8h7go5dWxXlZQl0OTcCPFVbWKvPWRtxvPLMBXW23o/l
FPmxcb2vMm6ZIp0Z6d7VxkGLa20quU3zIaUHiyKbnnycX4Dz0J/GtwGDxc1PM0O2
ufo5T87dgyQTVk9q+v3ULPrvOOEPIxtYvYcpN0clEoVgA5lEYXfTg3zrBvJOChM7
qVyc+Pmf15T3nx4mGJHsmpR1rx0YWjUwG1kp/pF3jpVPTqnBr6etexH/DGnAkLxS
qQ8TSQtpob5QkAkRlffzALc9OhGR29YtoI5AeGitQBory9kqhbv7oQ4Y42zi5JJ/
BcfjNETCXKjxMiXCHReE0uBngsqvJkl/NfhdxZJVR1urWS1tcBd/OvrztDHFfF8M
5cYPrzWuXjzbVgw/BN9bpVublRFFNpfU9tIUVg9jHqIbAi75TepbgTIGy2iKW1pw
MQQkM19U9q/FMEfX9tlb7uhJDIExze/99paa7oW3tJujtlsl2kqmAbPfgy98DIfI
U52nvcn9LE08ryEsigRsgmRSgYxLfCsd/9xVSxmVRRRnQLnf9EbUuH4YLP3FG7AZ
j41BIA+sN/vVbJ2Of54VK+vFe9QV8qrgs6UCTtFCe+xIqUh25l2ZnaRA6Y723ND3
PldNRMTHzZBfuL3Xm6mFFxTR+eDfHRKy+URxjxy1GIducX6yLNoJ54+/Ag3KM6w6
o7vO2Q9vxu4zhX9CNBCPbLApJ4gdoYyOOyJbddnquyUZaBDjVRTCVhd/yf3nWULc
oPosq6UZQZT/62TYuS5i7swDNDYaUaCgvANWcHRRxk3PHT4IA7KWJamskWYZl0Xc
lJP1Xsmp9XJhaSEk2+DARzkEZv95AjXfYZH/wtiSryLQCgFpc+Sj70JBi8rXC/S6
JpgWswUDCG2wxOLz8EXrCgpHRO2kpThTehY9VtP5DFF94JVR42uk+bJ0BvYt3hTN
3CYC9iQAuo00L2m4ma1/awm+M/4XzSfvEfe3fSvZT1z+6aPYQk/FaeXNWhWoRgAo
CJipQ4ZhvGCSoWBcoejdl2Awuh3EhDzEwf0ZY+/mJalEbTe48IdSwvolArsXS4bK
xDfQD7OAOEZOEfVyauY02lgSB4Yn2xDL3mdoOni1RBptz5GvchbTjPRDma4aiCHv
KtYmpwAXFcqR4li0THh/C/yNbcBgAkRItWoCeM7ZtPXel4A6uXXQwx87f2H65ze6
ZoDkEuj5htB9hlnl85ldIyLMT8+nljjUBgvQJh7fOWHsWBXgMcIxOSzx/c/tJ8BI
c7rWQC/8IC8b/RL9sCGQbhj8ERx35UTw9ckmtRhAoDzlx/bY7F8QR3rC6luaXxJ5
8I7V+pUr/vjgifrHutyzSOP+xtkJrlmUj6lWYF1w7W5NcRrJNhg5r+aQHamISWak
968km7Ji2JgAOQdCy+ouL0JfL0ZETbD1aTqBno1XJi20fEn2ljFopT3aKW0+1lbb
tWxTHrVaIfglNEU8JWz0q0begD7Yzwy0FkujoU7Fj2ZBpnxq1kY1eb3a2WPFC24E
SxhZ3oyFKpP0536Diu1rrel2UHQfl9woJlwups7dUhOp3DfymE5zEQo9bn540Ugw
Ig155Rg1Ux5Hbg+oZUnO+/7Tofz4WP/x+MTr7cZbVByLdcEwZelFVfQRgLAZGZC2
nla+B77Lr9Vck752BX1bm5wf4rglhglLluHvmRvPyWystQ0TwZQo55YsEffbsGny
gvOfOBx16jIjG9VI/ONfmYvgejDHspZOWXcu3K9cyN2JTsZTPMFTu3ZWPI+0fjuI
ejkHXYuQsaxNBTpJbNk3+o5rrDAEnVXP8iiDnnligjaSK2LkBQ3BtnTKNFc4Lawe
mSKl9aZsTUtLUrskNyDDjk61u7MZi0ncBi1qIlJk0dS6X+i/5KNnPxTaoYJNCcBk
UlvOK/WnofYFsrAxKEZGkjVkcu9VWQL+sgUdtm/69NLVNG1mjftcqRPOuaJuXTD9
YkKlU/oRMK8qChktbGi/cnDevXTHprZtK5BNAcFINNQ94b/wfq7GTr+6UT3tp/4b
DC0Z0ziHR1uLxGHyLxhLB80YjmOSp+4tMTBQ03ddyMD7NsJ5GEqV+ybnVU9knDEh
GGIirQxgk3yR5bhM/Cw6kMFU1WnnDpZPFS2MLIVUSJStolg1juPGbKughuyckp//
ojouEG0IzXosxtedNrxzjRtkl/BtpoPHHlfIe5lyEdxooOCv4Peck9ozE89D/b6H
Z2wwnFqmcwsfgAuV8KJmvVy6cEF4YxApA8cAMuC4I37FFnU7jrhUFrBWh/mH45Wc
YAN9qzHsZddsZGBvAv8BnaHUj0ddAScZGOCZ26DbBJQv/HKOm449ev6oVBeZhMHd
QIPjQRoB0P0OiNlsI7xAZlZjJDaq/7vDURV2KjTjqjHY+VwZjvpo3gimOw81US88
jgv9S1Ihkqi2SuhMxuMUjNl6rDAvvUaI81tInwsm09W1RPYGOJ1xq2SygIFmLQRH
PSXi/VKO5Ldm97mUBEfG4e9LF1K69Xmlfe4gsJj9Ss+bHchtxFA0OKb29nZHfJKj
hJLebIJnVY3Ee9FAuNVH+FAlmi9zbkdxhg+PC+nno8l/DCBHaLIvSh0lXl6O3Q69
00+QGftlL9oD5T/vp7hDg5FgI/cjH7vyZCKAvh3yx3+7xwawJhMLpqvv4W7hBjKB
2JSBm2qmamMfD+k+XBZLqpCUEVtf6IYgonKpNgTa9zxLXgJD+UkERcoQGWfYyRa7
eIUWzJ1w8hOp8lRGxUUQWagU13EE/KwmAcO2nOnYtknjCNkqNRZCtE7WaykrnZqZ
HfZ/dOBeXazUNbmlioZG4isBffPZs05ZcMw2WcmnUGfS6aZF/9XAt3NR5u4Jz1au
YasjyhrEXGm3E8HoxoNkrzWDbFgp3GNjxDOI/RN24S2gk2YrvURFtKYGCVDYE0ve
eBM/5H/Vflv3tZKqV0RGDZmyEsjrOwT/1EZUJXBf+XLmSPAFh+PZOMsTdMPOT25g
6RgETdbkasTNeOoias7STZAXvCyPhkEdbOzb6EdqLYny6UERpNoXwGnhU4RRstcp
1xkRhBBU+GDj7KUdI/S9gAelLXT8MXY+T7Xi6pC5fm5bRQIA4jrcFoZZNIhbGkxt
4FTM0SyVUxTRYBghnEQTLdSQLwMQGPnrB7+/36WALURhEeKMOV/PZUj9LXc2OVMX
1uCnF6TZUHd7KyrnuelcU3W6SMSmjRx6URjNLXoR6sAXdduAHMO1DvW0tTJ5uWgm
FdE8mJQ9zHF+rIM8DwPly6AoS2wVtwSniIwX5hKr+HXYONwF6gbgxygmKbGYioo8
38yTsuZBvlGq7XWZKI31O9L0IXJ675GQZwxDByM3cyIrs/GemrBkMZ34j/y45MgR
6W+noC2K38Ei6XGMD1Lvn1bXzrPGqJNEIHh8nd4b8hUyclMKkSxj3cT0+sr8ryyt
C8u2bhEhp5W59O9gE/bxEPjAnayqs/a5PVcIRnf3NYYg1ccfp7jNViUwlWlzmzZF
Sj/vJckePCyM4uZfa7+MHKUyCiAh07G0QhYCSlILUcYQQxASeX4j4KxzASFCxUiS
iMJU/WRW+pQzR5Qnkey/03B/JrHGtvIufBmNPDJEgRSoj1+bMYEkZqyGK6v4MpIR
ndT4z6ZdlANnUdh6JomeloadHajEBsyKZnMiOiZPrxWQT3fDzmFLeViqcOA5B4Ml
qhd7GW6PLjq4ZB89LLb8LPf902d/yPeYSYs8G8R0FXUKJKlZyr5wZzftOeggpGeN
Zap2AlSsSUkz4vYjMq7S3jAmOP0LL0QP+35roKzM/eQ0x5pA+5kYEEfkgAiZvjGy
CdFV7db+sqExi8tMBoP/Dfxk1AOSjLRhIqTP7UEye3cA57pGRRQQBpvLbC3p+usO
DAOafOl/UYPP5X5IFn4+iPA68TQ0EQeN5rFxXqBrz2/8utCjLRxwQj+kxO1Z60Q4
OAGTkOSnwJw/Fn8QHRlOYM2iVPKqdyathmyM0Qrat5fSvXq3M8qMTR+n0xerm2/P
k07ayO+h/Y/xt26+dBjKUdK29Wgoq41W6LjW0/AyAr4wdzOYuXcL3Gs7kJXq+wm7
0kQps2cXcVwyFT88Gtrj767mxNfUAC7psUL8bDhDo/XNqfML2XsW/7tKx//2b/gd
vy90VX3QZQAHuxdky3gaAcRBxaC6wfbpVv8YpVAtQiCXjuYih5QOjEHScp2Fsg6L
5VReKsDuG8gyGfnBifa+gWMsx3/EQBGSw6gxtzfh7t08TpeC25UVYAzFlQ7oMyef
FSz9eNX+TIetewTkD1/dD/TqWipqNcg/zwoGqNegPs9q9CrIFaLZCnb1dezR51N/
CRAx7D3FnmCh/Qz2N1g2M9GQUefrQU5h2VgHEnXqPqfVkCK+96w8PVb/DiK6rMWA
+rG52KP53YbUUOMvxVkbR/Gtj8XhZWlV0ej2OV5m3kfBErqHlrEx08bw5BWl+Ze8
4hU8IuV7KecFJK2z+/uBlrS54aQoIvIRsXdSu8Vp0BqyAXCWGmOHBxUy0D5VxHbT
pGiiRk3c/QE2rJDpqxgWjHDpp3Nbh40Mt/xdFB6dc3QnWfg1soYEEZhslO5SkUs+
q5Zf3xdhPrP/hLfWjhP3sAjwA5+lSQTHYsKD/2MtmxOtI4O2OoB6ddnA3rW4lIK5
wz8ocfxTrBSUw5qEHrdvsSQKVOBHDFGpZosHHVJ5zzGi9A24MvPevbeS5reV/y1+
0Z3zVDdfT4S6WblJKzpEl5Ns+g7ef2gogdgfilooBsZ0+c5mU5x+oKimlOJk0xkx
yeIFQCTnEsLLQ1g7tdA1v69HwNK7fDQdwmWKi+yKxu3t0Pzxvv/oQJ4RR8yPGLF7
pGXeE2/Ri8VmncVZQBCQct6HGHyL1eqMKqwNeYWPvBYDXtY9WlGkDXHrDOECimDH
rdtsBZrfahluXRfSQtbjMtxL0dvJoo4DRIEBho+JBqZIo2s/mqL33YeWH+KcCKVi
LT1YV5VHGssKl5i4yKiIdRx67ViS80rZttW/uQdvkzv8CidcBPb+2ePMc618Zw4S
JzTCKdBrlrnLKfc9wLDiiSW/ciirK8jQx3BdbMKGpij9kNvbFOv0l90vyQqERQif
5XuT6QSNpUCqB/yCxMlQjRTJZRFIYgBtJP1MvKSOoOS3/FfdErnmuQNKDAYMU+Ax
opDcOAdOv4hBIp6Esqe2BaL1j6LeAvxqcXIann4NYvuS2y/U+78jTsmaHpQ55j/h
fpTb9oW0hj8grds4OdSDwak5QVWefXD0yUdKRO8qasG9Dzz+J65xv9W+RElzWB9f
SoUILPHApeLs8BXjTzRXrl4zpe91bi6hYeyYQ27SlHa7DGQvjKh6uVTYDKCTG7Nb
A0amylGFjcDBj0FALw0UugcxlhpOowLT7tfQ1ZIwkmZwDn8eHOf8S5w+p7bSUT4a
MroglhlDhtdIKAXFnhStdc8KkJ6cpur0PECmFcXrHhLMSyBApCSKXNKZpC+/dOmM
wnLWlAqOZT4Jft3YxeiimoDW65jGfoWT1+XvZUmbvYDHOwn3vnkkWzQYjd7jounp
Sctm6h4qEwMiYoWkNoGumw7yQmYsb6uTvFi7BfNavRGn84DtxWqMcGL7tiYAHXBT
SZ9LI3a9y2R//BTQhg8ZbJLqRhqxrZsQnrwLYJq65oiVrsZ/y3EkIESnrMyJjfPu
i8qpo1tE6FkPL2t117EuWHMEejr4hGRdaIB/4iBsZo/QNb2Te+enDkHjHXDkosHv
EtwFT+bnmXfrHVXtGe5Of29KkMnonJVmqWQdSqLd4/B0Og/+P03Qv7A6UA9WvdUy
Hnu0h7xlLUXz95BunX3VBUWh5KFgXOQlYzOpyu68tU0pED+MHMA3d9L/goe/dHig
SgLnOpFTv5QpVgB/ZA2fVjZ+A3MLsbPGY7JJU0a9TKD8iEwa9m3lfcIPtc1cTVzB
cf9ldosxJ2W8HXc//e71rzc5uTQGquSNIQQ71ot+bJQDIFUQhxUcBlpcFuPKPlCN
WKR+vkefwm7q+GxXKVhEyYfnw0R31W+K2atj/LHXF/CsTwIOLAsOlbAo+sqEs11d
g4fPUm6NHuOQmzmgdXQ+e3HlKYtaC/EDUI0sSxVRKR0Rmi+9rsAKmRHEGKlrgtHR
N2EGnDhpQr+lGXI4Zl0lDyK5YykWoYQXIiypFewWgzV8tAx9bzea0FVhsLHkjWAa
5pLS0YzwzF53ZOAKea7gptVUs2AEJz1deDPy+NUvsZQfZk4Pec8LVTGQbXt5/hgi
8bM+Lx5LoY0tTo/U8RmwY4Rp3tEUDe4SXbfbfexN9OCBmGrokAQ+9xQjI75JWAyX
EiyY2t0izc20G2puMIvfRwLzMVKgius0gcsxy63gddtVJ6ZK9K9YmIkmnDNMJF5B
0kRfJBTmIZ1tPFBiYOygsl8HxzS2zjKTqPkfuTYrIQ36wekkU0Ri94dGkGwdOnpf
PPDUq7pbIpH0AnZ+je9Qd4pR8V0QwEU4M42VQK59MTmnwtpKn93oeXZZIgdOyAOU
bXmgTuIMrDymM1zMuRiUwtNrq/rb4g+0NX8mJjF4GK71fTszCxzw76/j1/IpxOjI
o6P/jk7Aby8DG5nmZZghAwKj7fsnmOutNI3b1M4yDzDes45c0BIOPlRxBxJXkbwL
lMgyJEDRuvBNsAXbnWnuMgzwgodFzDiNnpYYBsPL8EyvnEnCCpKVcYwnsGRF7/4W
TGg2Hp9KK8zLaQIGIVHM1AUdTbnkJ+znKmsXIRqW98Mbv5sdje9+jS3b4LcvvB8a
ysV/g0/ASAKFYfzAYVV14tKveOZ20y1b+dJER4N76WWseV6hfATYWQQB8v2ATdFZ
6BDZC3UhKEsM3Yjkiu2kF/TrnLpqrroRf2TQ2e3cvwawbD3oaLpeva1en6+VrHMc
u97MAo89nRTYjJtxiItCaVCMAZ8BvgPrB1gCH3kwqIRozfPHe4BxOFpbE/yYNCNo
Of/iFrJosdhJ+QwylfTpidn+D0Pp5cOy9TC3KFYW/z+8vdnlnKrZ/P/5aRm7QtFT
KNrYlPQJ4RnkXJMme2KzuTsN+M3jr+x0n3Yj9h6UiPa6D4fBgzxkDZH9N8FB76h0
zcqSRk+iff8otzMZsaw6gQ+Ww9Do8JkURV3Fy0ARV/9qURet2QX5xE/IskecatTp
nCDsxNkGlEIcgM4HTdiKTfl1oKY4OLnYykwuUCHifUAM+7zfOXfaPjvrtKR3thNV
W/J5guH9ZxANF2WVPBoMiN+R4//WzFqi2Fv3XOhczBGKby1BOEk9s/kScNR5EtF9
WUgBd32EEgWuMYEZ06w+8r4qxh9zPcVMNkIVFGT/9fl75RLAjn+IJTvB575cYPUA
LKHVFwTSSXzeKr63PmvZU5irh+KaxiVz8Rf5gHh+weYyJucSE3Nx/VR5PsbJTMh4
SgkgxRN20piq9b+4ch9IxhEuOCvY12aTS9rbuNhopam7DMFx9E9m5nCuhSu0Tjdh
JvqGq0vrkZa8kgZZa6ObDKR7AAfv/NXRn5Yq0uA44a2tpneVbvBCFjeWgdhKrAFr
BZhGw6nbnmZT0PMTuIJp2uStNVEUbWDHaR9cxj2klw1jB4JlOnX3SEuanZzOPc2i
MIzWCQKY5pB17XaR7KAbEc0uD92sfrK4rjPxI+oeGKoBqWKWdPMwNN0Vzmgah69m
b0WpXZID2l4/CBwDf+HCjNj68vBVNVaPGc6WG2W9d9kO7ASYNZJuX26hlVvpzTXC
y/jV5/A3JUMLALDCMCY6JcfCgiZSKd2bwX8SAU2x9QHZlnPC+st6+wSOC7MQk2HD
p4wc+gL9jLBaSaKWUDUvMTTsUKaeI1p/SQGSbWlK4dRGoDQJjdID9EgkaJK5tfrr
nY1xeuq/UgUKflNFB6lkQ0sSXwYfaT2NstYY2DJLIYNFkGf/dbdlWsXIpxkDVI7G
o3PWx+4EZWxVjKWVGiNUFi2BWjtQS88aA5RIBcJARyIPX/kxGrvxFh/6e7pWF4w3
K03eL5Ykfiq49n17LH7Ig0I0qZW7NNv+vSXPKuudxZnriwSBo2qdks4hSf9uxKhs
Zdttnm3DWWk+ncf4FuW8g+XJywlXnLgRjqzOg5I/H0CXCUZEn0Amc+OsN09suijo
/TXT7bpg9T8QYs+ioUURvlX8YQuuVIYdv3tpy5GfIlYdz79iDyqoBLj6wrn93MZp
XAzYJzN/zQpXSukoiKRRnmkI1RwArtNKur6/IgpnmRZo4sEHgj4eFq9UjsPUj2ue
ytgv7xb5Y26g7Ivj2Hjl9ndBAV9L1TTx0NkGvlEJvy43Ct+wKCCjz9e/iqEJ5S6t
xyCj80kn5Y1ucOAmIZVYaojBuM+fN7/+sh4kbbwStSntHFGGRDc5/GOAbiLUkjZG
ObEri6YJYON1dk+8tjEuuailuagTnh7ToYWlYDy1nAVGaPjVHSdonVdmK1gw0+TL
cbzplAswD/XN1AlStRqLmTFhlLxvPTHyQzXgL5Sn8EOqXdOBpGMracKB0n+A6HLP
y2dut2zDFjtLrk+/tFHyieuZUR3O6K1AoUR/luCP/Ma0OSN0axPVY5sjrQ9o9/EO
hvG9+i83zYBIMNXDQJSZ2QZNRsmmHBtypZ1HTzlmc/Y5PxcDoTwhsnfWSq43hT9Y
W4+rIPVslbPjuQNk5fp6a+98OKST8L1bOk90z9CKK5Unc4X3/uF5oA4ZNcge11ht
1XXZS/pJRe4ui4uML2crC+r7m4GordhgCgz3QT3cPD3xiXmJ5MNjvZ2MW07Qswun
ZPWXTb82KjCx8c8EWIWbzWmSyGcwy2UAGr/9NbK8asIC3MDw7hqSx+Mh2ls3/jaQ
joNZusQ769WybEszFqftltmSbCFYleN496jmSluTuqnYPw4UEKYROUMLfn41oCzH
9oocwi+wGyVTObiTxuh22st34X7dV08BByjBSOBkyISdSTMPyp6mh+d9BZ/gPZUh
D2Ijekfn+198dTVMMmaOv2YbDP3NInqFT5DybpV2rgfvthgTxB1E+2EdL+p09tVC
jRBt7RqSsTtOwBBrCPOV8IBbKUVISTb0b2reMkcpvL1yx9w/Ez/aOayVryHi13of
KyKdt3BrRvbrFaz/7347CvFvw8fJatl1Qb8faTgqcaSFx+x24FPaiMojGFYgH/2z
oqxGrG3U/wMic3ygITrBI5PdergCt+vnmR5DHzvfteG+bx5n3N/bydKvLsMLzbke
A2DveDiLQFowXjGwDMdFlYewZsvNXmLF/fsihZAjEUk51SPLYEsbiTcf/x4LXHMJ
iqTQa0on3ZiNRvXeEoSQw+F8pn3MDceCSPfsDHasW7l+phZ1r/jLv+EmvcHS+aTM
JhJHNJ0QE71bT6fU5GdyO/VsTZ3usuw+fRmvsnopdQe7km42mYwvpAJj1G/VgiSo
qBROI4m4yTvRfSp3HXrUwQXoQDM/mT/QaNIV6EYWBcDJ7dI1j1Kg8hqeCZWEq/1n
BHL0SYc63+DCEj72l4WkTGEmzd1Cf+LcEH4vcLhzUrU3q1g19GrnEiZ4YcvZ+7CA
l14U3Bx+Utk6JtL53af37uNXd5LpYES1zX3qiUPv8pRg+qC27HX1c+xK752BBJsY
CUEZab4GCWvCDWJN1TV6hdXmDK4gZ2Z74lTqLMddYFxyV78isqLhg7Kf99J7Busw
7B4WqJi6GVWII02XOntnQfBXFHbeudHed5b/ErryY0HADO2JAWKxZhNEV4AqbdwN
5fmpA+oS5crKqmV80Gf2hTl1MMnzqf/isUYXM9k2A7H6fCE883g8k1L9FMBXDiqF
PL72qLLqvsul8lAhpOqi/3eEfFx875LEs449oUQs4z2nEG/QBYhL1p7NoktEiZug
WJ5+4VFD1iyb/IwjCP56GHjVJXHH4Wxl20xyAi8Y+EVwOHPFLv4igp9iTbG4SR5Q
3ihClWyKKBWR26fO7YZ10/XVAEk6+7QElC2PccSKAoNiqxavP/QJqXPG4lrV1VPv
DQfcqMEq4m4suHCj+g51ekT2QtEr/f3lTYpHCjMfpGN41J5piBVVME+Al417u8Ur
E8y5J8455Hv8BTSokADXfp5MbHGiIJuh64yKp47yliPMQXgynentKPqY5DTCfzSh
19m4W44DYXE6qjXxINhLSg1MoEXoCUhLyN4ghvPpju51xncg9OhUcQVFKGwE21Yj
/yoX4ChALEiUXUNN9dzRACYjB5PKixFK8ey6bjvpgzRfPza91xf3uu6I3XNFgJ7Q
gUV3ce0jhEW+68PKf8xhq0tXEaZIXgPXkp29IaBgEMsyX32VU25On0eed4bsKGjq
4gKAeb3c3C+uNjxY7dJY5lsBrO4jVFzcjIHJ4DjqeZkwxmAhaqH4WJxl1BH0NmNo
P+IqDwyckjy5yNhsmco0276i7quqNV7MovPBpIa6gthUCW1HvFewDUToKQ1OuTF0
l6n0Ptl4nX5Cs6Nfkv6F1HNBRUl9JonIqEY55fr2aJq8RSFj+LkcmJ63khVdYRlc
I3a9sdY/SJjuHRFOuSBIUZKUF3Mp3fGqH5I9La9lGo3T4do8jNK1sG/GhTh254gV
tCfQibFiuVqoaJVr1GWDsbXxxFRmi3M3e7rVNv5llhwK/+YSCGo2oDszEtC6+kGW
hSwlJ+EGJ2EQ+VgHna2BTQBwnY4AvfinjP8iCqVwjEOsAEyi+OtvvwywDf1EohFW
O9FoiwOi8Bzl3xUQB0oU1hlTfp/DHQO7z8nfPIHUlbuBAPU/jJ0bdx0fQiHLYnss
i53nYNE94VEXuA+mPVs4L6u0hCq2RIIJHd/soJmYdAOdOTShcZVxYjH2o0uOwHY0
VU7/A8lhe6gzw438lji3o4I7SGJcABwuToRa0+rzNuAF7DPdXlzcbZw8C4+qtQa+
ckKaqSLRNEpokZIUiFAAk/xfyBoEelWv/P+PjG88p4eH+AWfHkdNvoO2xP28XD6J
uo1kAS7Mtlj+LpI1oW1dl88TpdbjUPWr+EAqcKN/peC6HcxCnVC1pzu/heuzWVf3
jVb8cLLUg3RH6BP7c/k4J//Qr8yw7FkH3tsLRf3m2kGI8xi+5pMYCqonSzT0843s
ITwvereEwaJrHG3vxE/Hhbw83Fsh+RJMEkADaJ2l5Vqw6sIsuzbIjSr7+Gyw5f+G
RbAmAjuwrgBQJfwlB9QooR68zvXdbn920bAVGnE1p+yNmeKnPkboP9xC81HPvWBJ
He5+K021hX1p6oJUlXSZaKp4pcyaKDigkyRmujoL9DfFejmlxMWAYj2XZHyc5bhh
W+fUBHy/4lkWkkfW5P5j5vmnfuIHzu6M1mPe091Ed2LQvEnj8S6SJuNA0BHuwtaJ
ZLk/PXxiIxNNGrnYo6T2Ye+I2hzAza9bXPaR54t8ddj1VzFCdbaeBO28qUzy2+Nt
lbVFdznGi/dJWykLwz29J+bFrvFq0WMfMI5Yj5MgClyh3FWb4NAsLmp0zIU7p02T
dt5OX79LBdf0zxdj7VTmpN3loiLtYIPuq1MaDh9UV4sYkQdINE9vKOGzgZROJtkO
A203aFEfbYGgpmyjACaroDZ5EeUWAf0hGs2AYryc8e9ZAI/9CuCoNo+kOqcf0jdh
DO7r+xmIJ0lXCV/HOxBdwJumXlneIpJW22N3l4o9r5Tq8Ml+tCCbXyY52L5YQUBH
VJJ1h4JpW3WtqCQl9GgUluwdj6lL6ETqCb5IbHPuDL9YWmk3/Qq+Aqoc7wM1vMDz
JVbN0zk2C1m6hSvOpR9aRvzTmxpUISUtORFteIjDCvEhjuCxLb2SWg0U05IscUrY
GYl4UWtwWs539p1GW/uKFPWpdCsFN8KrcqgUtEA211ZJNApamlJ+Mvs1ilVxkbmq
ksMC8KdkwvOQLnl/HMEzcK7v0cX0GnfSPeGT8GYqtINMoepZTDJjhBJHCVmfclY1
MJUGxVae7eJKVP8sH592jdG44SIiNx0zU8vbSQSIMhyMunzeSEWoos+Tvum8p8af
9a3Gv7bedul2DNnPE0qLLVTPoR4xFjZ1iOso1RcL9uG5l4VF/DTsLfYWkhXM6vz1
zict6oZIO1D2bQHGAuoEiDFFx9IBTtSuwzIFHlVEUdAPpwHLirMpG6/u6/suAKQY
3Uluh1IhUTVOFg8ltp1d0A+ItQBAJrpjCZNf9I+3L687HFQFuPZdJN6ZCh5vW/hy
AKXcpMK1jklIJit3+aFuyCLnPEVCpJccgnHz9/3jEGINqSlIOLPWDpu/mTrWHpsG
5K7LZps3bMmxw0CHjU8PAKHrzxT6ESgWB9N8qFEXtxIfhPiQE2Ej1xr0ClZTCWGf
iGbq3CEYN8Yv+jOgbfQN262XKB92knRiIq8BeAOx2olY+4WwueRfyus1JmUO4ILi
egr8hxPueBhIiKFDkQ0XAEoxu2+NAFydnfPJ2dXzOzGkUgyzLMYS3E+1TrzyOXnP
Rg69kRKGRj/l+3sKZfzwZdkKn+f9CogEis5xbRgNDCeMhSDrAh2ieRTDJdPgMGqY
A7SiT4KkjEXsCMBqW9nnEqGVcznwCEK/iQmgGZgLrGy7vAXpQHSfx+aWDuXJvtoa
BP5bO4mlFf/DRVPiUTRm5Ja9s6/T0gWKD/1lobyfx3MyxxHflspDtvJmfhJen3A/
owEg5pB097a8IskZi0rC2ldrWOrwgMVscZGi/u/4HlhRRhvP1VH6KHVugUE1Zlxr
7n8btwPrQALkjOfhzO/eHJMxeKRjxUAWtYa4jCnuJkJKOjzoneJWXmqDgngUl9y6
WgCNiAQwQd3hpTznBapA4Lwm1Ya9rjmVId9bAF6yuxxbFeSKl7DWholnAk4nVSFj
RIOZPCuAyrO/CrWqQDSnL3lXdm/xyrfhAGdPKGNecSzdMs446WNlsgVA7G1MIErn
8K6k+soK9Ht4iYzxLrIxQ3Q3KXmnsf91L6zL5+FLSpHvNuiibrACLB4/F69cbXw0
k43F19R71ZJSKNklN89yB2ef1Y+fdjdMNPAhfFkwy5K+r0dmKpKMTvoybok0V+MF
lHWY9Emj7z4I4AfCIFMt5hDcK79lkhuaSBd0BX34Wfl6GYjITJU3lkTQFpvX8b+m
h9gieQ9AbxQQC3qWhGjzLdXNpIBmRLS31JRyv0v4eaFjP+0Vu/FhKtWeEcFkX/vS
zZeTJjNJK2aX2bwxe3/NY/E0fp5w+H3L9fxgTOTi47MWxwfCIvq8eSV62T6o1HIs
UG70/e5MK6BDEEF3G3rOS4bfA+Kw4S6HVg8ZUDauv77sJ6RjWE/v8nCF25phxbcQ
lGH+3ONd+HEPYixXYwziBt4bb45TcUUjaRRmHEvl0YiyStk0ZKnKWeO7nvfkP7a6
0YgptmJPk/t7TFC2MbI3VscwD9yYS87bURTGGzUb3wiABHR6C5ZIO0DVrFakH5c9
S28xWg5hlRZT+dC5kHFLIO1L3E91B7LA8wl/Mr3MrZep5scO3g9KK1ZtXurDhSEJ
6Ro7t0ps/pi4oKI3klpfOp7mnVFi5QC+Ku1ER/EEIUhtFJ1aSRe0QFeUsvrs9cIq
Pah6TNTdVuixl8d/eNJDw7HIU6WMxBrK04PmkLfyBJ03t4d+c8O1PZmP/zRqQjUK
qFtP57W0RUm4g2m9w8Mljx8loadmeJHZrm1MQOQFsChF3yayAr+oJvbVDUroQIua
wABSbqMo6k4rRpAc7gW5YdaZDk+CYvtmOlFKE/vs+xYpE8Ei05ASVIa3zVn0N2Q0
2s3iFyF4xLnQsncjIdMVgBc20/qyMaEbotoSb3h130KpNQqJcSnrcOPCIG8wdMHU
94L1j4+TCAppgkeJcUeGcKNIZzPHFZujwCRZXGSmTJvMYZQz2dF78xDI2qbkqo0R
yKm9ABGKAYs3j4eJGi5xWXwQhiGAnpvzjzEzJomNax9g3iq/tBxuM0rHwjlsuNIq
EAQaGdw5VCL/5b9baJYgxGjtMJslOrK5SONBBYfLItn0DBYT9ntO+79xNwukcLyW
RQpvo3vCunhriNBTQ1uRuiHh4ac2A6PSLdiGSQwk8877OXR67u8DS37R1za5aYbm
rywvTlQ9hc09Xl8dhcYT0DF28I93GWdKhNIef2yA7DtlBuJCKmhffdnng7gfHXsZ
ROVK4nOKcefxgZmoHp+ZPglXOqX7Yeaa9u2Kq4sgsv99jjEwiQou8aJSAEaYHX4P
g+iMhrafrc6OkD93ZE9mh6LDtUJVFBuJG+8+JVTa+9v0fkmedbHgs3mgLOwjF8/7
AZrzTmtFOap/rqiDybif9X8TQ0gpUKIbTmuITA/gmyb3H4/8HHlKKXmGCeZnAoSB
X79Ls6kZs8eQWNz235MuUJYMvXyXF/+wB59ySa6BEa9S7Q5Plk+EHK2HHhsdj+8y
+0ATDFC3jJ1PWozRhRHG79hthJnIeo5u+Hw78wGE0kQazFcp5gQRFT58/EdpGw9+
fox1WKCIK/P9FpHGExbMk8kVmOZ5kUwBwso/SZqOC42h2DDA48p9MaJmxTGc92Nw
43rWwmYgPBU39+XedlLiiogASrdesynCpLlV7NX1kNvU0//N+IvzXIMs7u9rqTBp
Fl13SP2L7jTE2m8ZbdZUIcnbXXDIoFhl84IWGubbjivnBZSPKXlMe25Rd9Fil1Tz
qfmk7yZyD0EhM/vrp0dc7xoO+5qjD5CJvDmKqlYIXFaqlZdSFbVP2AsmE/G5hp36
pyeCCpnhxNmAAZ/sDerD2X5JxStPFKchFQRBNVVH5xyU+hwxZgEPCKySmbKBMD00
/cdpN+pNOQ5AcCklwBSVRRrT9fDtmNMhuExMPQPqPRUTGmTZFOhPZtg4R9ZIz/2k
i7xpOUXMZ5QZZydHXWR5fsyu86rCOgKIzv2LPGo+2M+gSJ8UxkeOinrJL7akL+/v
rn79YgtDfo17+IlvoOOvGQrzXRi0tvRrTDNIDDDc0oK7qrPjV+/IemeXxN+0GTCL
0zbF+wCbeQu2HgMZ3S6frobpBEAnDNKYdlWBBxq9hVDxKiWTAvh1YuOcjDpUnvyx
UBnz7hp/ANL3k0/fY7nBBbqjt75FVyPXQnDPsXNFhfYjDmvsxSQHBCzQz5XevNXb
k06A5ANnaSvvT4VMRpnbWsSjn3gLpcdf0APXKEwumg8CGLa9nr20Gd8fVdmxLYtl
Dh5u9rLqiUNfGnJIKoV000zSPDri0bVyXf8a+Cp5+ZKjJdue2DtMWsYySY1Rafkd
eB3wNejWN8pillq28t8TkiIzjOI9hZwQ34Erium5GjMByB8L3mTY8IPtZFumcHKf
1Urxb7QSz5qJmTnof6stUekAX8LLvNYn3VL4Vj8spmbuK9cmglMjyysYMZc+zSrz
EhVZYRDqMhNMWFC5NBiXpPvk5gNXsU2ByA0MBMPbJd8YxmM6UTVK1v79YiHz6K05
EDRROKF1kVV7xP5B0uZ3hPfcYZsmXjZ5dFs1PefyckesoVJHd2yIdhTbGobLKLr6
e9UYjA5eoBAt6Wos4XkRL+qkrfxhAClFcLHeBI6f80xF0/8ni5WI+wZYbv1GcZgz
itoLN8p+BxJeNjKuaKMTTn1e/cA5yO23khm1oxnAfuLq+feF9jvToGAB6W8nGUXF
eGKr+SamlfdK4FHVvWVbM3eqeq0EedVUGm+EFZBg17cOnw+rn9fHss7fyyU/eMsF
Ek5B0BxzOFOTaJFtPcC7YSTvxEl9JBsfnm4UWbuD8wvz2pwhM7griUAQAKo+LMNn
ZrYNgjmSYqmR8UpKQIpgIzGnXKLwD1PYlz0XfyXrd+Gc/nV+8te6FhuEcFM4VppR
Ouo581PkSIAXeBN/+2L0E1dgx7pyINsqpsPITle5zxIgC1gXTlpm0D78qMxq6tTO
CT6fTOCFUF1MWqNckHyrGmMcO35xyLvwRq53l2dUKLxcagrQtwmhGvbQMkpiTDht
iZuuFK42tdaHdvoOvgdMAX/mJlzcKk6+Y4bYkaskuJfNVRF9uYpVCganVvBuYcA1
jd0nRyDuAYOtsbe3n9k4ZssYtymp154A/qwVgT4b7Gs/LcUR22pef/4RlLgWI2Le
TBvDtYhtd9nabgjqtNkh0ebaaG+MYr7J4gBSiaEXhOnLoOPA2ufp8dmpIvtGTu1y
FF7Pl5UwadKCu2Vcsr4NgkGO1u/DFryU+XNmx9zhcCnoCEA3k4xvkZgfIxap1Cx+
y+UOw1WjjPYKYhSGGjHkjbgaNFvNHl9iuWT1irmC5Y76g3jPgRfwau3XOa7LBivH
KPujr56iwoT4Dsh7CiRabFLnvANYMdo1R77iiCwOO3dnRjYLNlsErEB9kLcBQJhW
yYWPjeZOR0Ljv1mBuHo1W3mn6erxAALLidA3IlsZmGl0NEx59wSYshpcAlvx/4Zo
Pb9O7kOtkLad4JxH5PD4qL5LLP8TrReGtFQA38SzkgY7uQDqkXbEOU8hDpFAGcRX
Y3l0B3EJwir2qGh+X2K4Q5qoaewtf671iKqJ2wy8qimfYVLlBSlOqCaMNgGM8pI2
yocBkl1Jn36BKpXfqKEy1QqR4k8xZqAXZAoe2iyrB56HRjwj/98kp/QtrKlE7hFY
CWMuxsw+M1ZWfpSZRH3hXax39EGTXYwnj+4Adtyr0ylmwXtnFO889h2azVdmHI38
Np6qus8JT+Z7zVNdtxDY+aDJPL0rWld5lrBvTpMFI9m6g4g2hZG5psQKhEgZcfGR
r8wKOWRAxJKP9GK+A/ehatguEP9/vK2U7HV2fNKeFB+uHeeoIjhdvR5yr/Yct+me
gXpKVqaoIeO0Zo1vJSHZ1oWkQ5X7Ah/6BHKww7ZZERAvNRU0natk+Ol7NlWvc080
DeTmITzAt3V7FwQZtV7A1CYtl3uxkhhWpThCJh8sThXUrV8lc2QLke0v2JmkIq5a
LfB8HB2qI5BHoXczW9AzNuyA2KgY6FGCbuX/3qMkKRq3YgIy75tL9TUo8zCywFcS
9aW8z6ClFPp71AwCtJ1atbkPOaMwW4X1vocETpEbifWk4+JOR79LLS45/TnYijmG
Ftgg+qAmE5NMItPuJcGM9yBWrhytEf7+IDzTPzy9jSf0BVu42xOQkZeLlGcOvbr6
19LJacQIhghCl+A6YEx49UvPd3mAJ/2U10PyA3VcX4BZ+UOKrfaE2v+P17AJu+1j
KkWtW+L4LdWW6FL37HZZwvWJQsMAxr8YwpuGiM/yR6HYq+Gu93loW3L09oMDIfBk
IDsr5JWE+ELNIiW0UBRbE+u7TR04WZVtkAVnnA3EPHPWLnYZaSPW/RrxL1zB3C1v
MPc5TTnJFTZZa79KP/vcQh/qvm8zrHMomo00kR04WxGJxGd5I/fV17SckGvk/dsV
OPazmSYppXAw97g9LwNzTxM9OiKOBhX3pra19l/ketzAL5Mpcyh2Mj0W93NhiwJt
lJkrKoN0m6T3ImA/xgWxYq2NgCUxTMbhmAekQiWJnP6BzEuWYVjmyn04waSLN5Cq
5CPSLa9+x5Hfp9KY4o65dbKqpUP5FaCMKaFoZxpQ1n4aENLRyhYcVdUaJMW5D9rH
dbuHAFLr2u1JrLdm23Uc3jkyFeWASA17eLK5HXYgObeFceVJ5WK1VLE2uj6vRecs
520KLSx9UCQael/VFDOaEU80TYsnFjE5rQHRMst3wRXr2s9ua3BgmNUZuVE7C7lk
kFPjinY9nURb8aoe6i5y7LoGwQNIf17GErjjT4ZVLA3UMDn1go2l2qLSiPfMuF0R
JvjOACDiVIgSx8o7iIUSplEMG5clbW8LBVWqYwIaXkj5qS6FZjN2MFZrwdBmj605
QPJfFGvMAWxfW/QzyamloKBKynA/11tXqONeUFKhnURZM+hXW0QIC4b+u+PluwOt
bYtSC1ZP4fymQFWlGCgOI+QY4zKCjO+zlGuAQgQNQ577QfkKEEl3y+n4IF3rgp0y
LSfIIy0DvsUzzwwE0W1ZS1h9KikbCogSvt6po2AJoxXjd0lYplRtcqdvov7exA/C
KQn19QDQ4+oS9w/ZWt3V8GiWLE+70glBkwEZV9tN3GJVyA93bgNhEK/pz+sqSsYq
ErmKNYj7PBkyDJ9/CTkU94NPr0yBQTZe69G4MkVrEPwF86LZEXSGrYsc9R7EsCWJ
KwMWdR3JZxXulElMxZRVDl8kzblzYUzasZzdRUwTQx/KHMHDxXKUCoxQl+nOFpp6
uohjAmGmNJZ+50srCRdMg1HmXtO6Jg5CYFRJRN2xQb4D9wsOW7H8krsg3hL6KBm3
kBM8uwv5kYHq9kgB0VrcGRDRKopQCwV6vsHt6BgpXoUTXKkqiOgYVnreKt4KkZOf
Pep7Ur8iHajBRpskbhiXEl+Q3HTJ0b2S7i7arlydkiQYpi7ECV9bNteLcByo4QE0
X9XGNC5/rlOU8V7x6LcPFopBMHKk8c9tAQC8UfraPSacl5fNs1mK0czSU9keCKKC
nBdXFRSkfp99Efu2GbCbm9yWJ1pnedwrLlzw/heoHRuT4+URyBL8fyxLETqv8mJb
PlgXRLeasZLHDowF/r+XagvRnJtZPDuCyxRGk+pBx9odqVSi3gbeJQUqsUQnDcXo
FohqI9CWxp1XxVvUqnZlW0Cz5LT/gBRkgfk4ppM0btNlQ+wjQJu40aYdEv01nvIp
NGNkc+WLDvJ+syUO9cAk+CQVt9hi8vZp0tro08UMMMWFOxp+Pormeag/G3JozTJy
cV7FYAi1+rFE+BWSKyMA3gkB1bSZ1peOyfUjSKCAI5BVQTW9Ru2sw1KNHqw6YpOu
VQn5e6g2gGhIeryG3iGLBx2h6bBOekOFhh9vLu8bgNV8d3c4os2GX9tCXhJ4Tp80
Gkb/A9WOrAQ76flfIQeZaDRilcPZvUHbq+BwZ9NwGIUhT6Y6+k9ACanLORP5VGz5
E2Ky5qUCc17Cox9+5qc8OyUFBXag/wSBmHbHgCCELQhuL4sw/P7OJOk5I3mYeOGc
qodi4qD8B1rIcEJbPej2wejucozRt5W43El77mR72E1m6Hdwt9S9OrEdMYpisMQ/
Ni2bcb31nZCYNcxb5ujFny9D851HDN9e2iXjovkr/nThnQlvGLDEFY+3+NUxGzB/
X8a3/tOTPIekAjXTh58TvNN6OLHCAPETrkcFeNxcMoGT5oT4i6cM4orQgw6mv69K
xUubUXjYqewf5vbc/qbQ2A7OXgMbw5c+7Y5cy9Cku/bbMiuUIaOKbii+uRC5NGl9
X4mFciaKo23sabrj6p/U5APHtyJ5QobVB+IzY4KN5Uij6fE1z39VmL4SD4x2czrW
J/8G2k/EzQLcKrC28bosorZWfpvw1ZWGEd+LajOfkFAuWs4dsIQSl3Fo45mCyE1W
QsYSVjaUFEqw9vjVzeB7ii4VWxq4ec8sHiLjD8X5MdWfTwSy5Gp3FI3mBdC70etx
kfEtycifCylT3N1PQ8B6CE91QBGJYQTC8BdTtmBqnpUIiib0+tMXAE/P4ty5+S++
ftR36TSSH/QKrF78GnPdLr1A5znfno02BYGl7+DnHGxB8pIDcoFI4ffVMo0iHW4i
LUuyOQCPTv0Vh1aVNWWxWZGv9CU0cOxj2/5zpBO3lw2OQq6sYa3a1wlrLCZHsSTi
WXOKlnhyLnv3ihgtFDE/8KdzCE6lbcS5nYJ8YnByhlV6j+JxxuGb6UgLbuumoFmq
+EQb0zScGD/Z24iW+B7qDrgTa4LEduAz8qsqP7+S8yWbFNRio7FGlWzwZJXVBqs+
+m1yiA6UlZdc2Qlh0MCRByzQBBBfn+vlgWQgOhBGuRe6y/XNH/Nbl23tLBhD/8iE
LTw3gXCS69QWtUWFWZmGcHMhDjbhEjV6pJ1kogFro8y9KXii3kuJOx5ha7L/f7js
BHaGb05Flibn1Lc04xG7g9y9LPtiFT1VAtcaIdb8S1pI/Ji5ZOfH1a56hC28CO1P
LpMQ/09UNCROiS2dgoqwsz86FIp+PJ3PmpzyX39kRnPN2/dKN1SNDPZMjSEQurpW
IzDMmDrgxTyzeJ0r0XgcYOEjCJW0tXAP5GUCEgWgFc8CcQoFvC8Rx6YYMrbuWodL
BlX5PnPP2n+Ox6zaYwmaIVM2Vch3lOc7uh56aHRA8wi4FJretvdYZsQbkBLUlRzT
wsAQ3D/Xe/FNmSsSCSexzBJ8B2S0hn4xjrC1Tna/XDnPbpzEiUFcOLIEUWsaBqZ8
1lov800VB2OnUwnif99BdUjMb9qX2As4wDuVdpgPPFZHIocAhUzK9OJUZOV2xuYZ
unIIeVl1T/2vyA4ltrPSXYOLvpSH9IgNGVaENi+Pn4XV+rLxfPQUmPeyda/etkU3
+T20aUYZE9ZUF6jCBXdACjtJ1kifz+RjNn8P/EreA6IS7XdRXt8h04T1o64xHYDm
vu9Tkx9AqYqXsiSI/O3OGluJG33sHaM7koTNcXYoTT2pus+xEruSCq0JOgaer+ZZ
3ejgYKHVWEHaGaxvrBTqmmonT6GhoxN7uWy9wOnQdTA15EQ+vnmoFTQonF+GJYUC
wpTP4t9zexF/1taC5uTqP5mPrTKH7DN00EF3YhLZCZ6C5nuqmUoifVq8BBPCOjJL
35NhiBXTM7x63IWnLXDjCGsfwRL8VdcaMjZob0TDLCqqexPnfw6uPjCu7JvwSmys
jL2VlXF8gMUyNJnWddZpM9YWdcQCC2TPdbtXu94ReQmtoOPQ4tUS1pmztvcwFioy
qvHmFl8xJIdk2A7yEQ+47NlnSw78xmkQUubX7MkdCZ58eR6HUS1zHv+BAFL+eV/o
RgVAQg+9zpBohpY7FmPoJPrJqs0f2Rsjg8BwQ8r+4SBfYdm5BUIgMwq7rj0y+1Q0
/zkYxXEVIUI9yNeiJ+sLTtgg2htqn2y7Dtz8P8QDrA5Rhcc+H+4daT/F3s7vrJ+D
1/cWEpPt+J0dDjtWyKjhsP22PdXSLaefCoA/bqQ2rd7M9O11QFI/Rh0eYFCVmbB0
yAGVJ/m5sufAS+nJDAVOR3bKevWwBLgw+EACTB+ev/J24UjMB0a4GZlbK9Mq2/h8
14k2rnXxmOzNZgI0u5aeqSRajBZlsSxUmAeGyWrGTul48cLpn4R7lOIa00xGzKi8
4obA2ouVNKPyw/5JzxZhJleI/wjGwnwBJk2C3IKWyHEJ6+njv2BSJ+2Jr/tNiV1o
bZav5b3Z2tO0xupa2fmase9a8RNMByEoy9V7yBYwGMJcUIsbEFAXlv5I5p1gjUE5
xA5Ue8N7guZ6vtf1HQrvXAuGbwZf1/evj3POhhkXcqyizDiFU7qwpjYjzvz20VwA
PSMhsS0nmk+cONtlMXbEby5EyqW9UWNSxycT/FLsp7lCIazyGzqtajuPvhO4avGb
b5VSmvPVAzEFENTVZXcbLS6BJQwaoCXIxmwZbfvZo+pOpx2xh9HgEtvA2oYQ62ir
o+TKKYKEyybSWGW1w3DOoky9XSZbnDsPCTSZAnhcICcMaX3hPBurIjX+npoLkgBT
eLBYPusCq9gMH28tDPE+UGlugPQNfBJmkBY2wtyeYaqkepKyRnDigIlPU5UIrZSk
ByEEy6XUqzrav6IJ/a4iPvNsO+nwEptBrcBeJsFwyRWF6ThEVUnrLuDec2qW+oHM
m8ZgH6Eb4SZ1Uh9TOlOQqhKLEMP2qGZSFdJPJnJx5KIQyVBGd0UdCEcS+wmHDVxZ
a61sJMxx25At+7XhUeBFOc+3GKvhtfaFqvdSgUw83RQMKsDpM0bG5E8wPmG+dVZj
OZqn3bhmAQrQp3LX1IHQMdS1MQYGKnxIEK5tpTwtN5jx15PgEyEXOcrqH++zkd9Y
HcAqXhobuZVbk+GjfXJZV2sA6Qu18QInziYvraIbLLzFn7xmrebuYsb//LvP7lei
jYSleUYoXeXFY94S07TeLv0qwKP39ch9/kFjxPrYRFirtD+NGKdcMVsseKml+jZs
LIy/9+3xRwkdtHHEY3ZBMLdMK6kI5nfSkLLtj/o7zc+Bid7KX2ykdVybX4v1w/O+
zA72ZWPTV8CSmf/hRchL86N3ClWfgdX6XVGPx/TuBwR2oQzmxHo2NEu4v30iI4g9
l4hmNE7N95PIF02OY7xR98uGZhUhbt37SxbImvJTa9eX+tK+m00D/2yUVCcheF84
TZLK1BMNLdyoU9k3eGs9m4FzQ+4VIFpLagOo7e0CWxu1Pz3T5iUvG3Afacs2AoQF
Zdu8S8jgxiPG4bixw68ZMOUuBtTXFcdMybdgN3+8ubCt54nUFiOOvW1eY75MTQw1
qQgrlO2LlEbCbANWv62zR0HT6chtMl7GI0fJdZZOL1S7MCag5JYCljgLTYu+xRxp
oMXMUeza9kH1muJmetgOAx53ZzXdcljNaPxTl4o7zDI8ImiKBg+ZfstIkQGgUTCR
kxQlL0ebAhBVQendLKPTligZGPuV3i1FGLW8gSuXq9/SakkoOSCAhkV6y08DxDd7
SFnVkIjtRNJw803ocjz1CvW9nM05ZhMuK//0rQg0I1S+yaqk9OS/jH40N8k2jGua
Z22m5IGbpVzSvhnsAhfjS8UsCTaKApau7OfDzLrM+XuQaqQ0mT+gr8V6Pb7B67RI
SrVNwg0qUFFvih1FGMKP5MQJn+l7iQR3cY+Y/UtDQ2R4bEZv9ng82PGgTfIc0E2n
acbPRzd9Pgqp/W1EsSH76Xu2E5GAl5hOZVYWQTbXQhyQdatqZAb1LpvJpGzDfhsG
Ka4SDT6K67W0cJZnid3CT/uwvMIytnCTr8i2XmXt2BQeg9Z7wQ+Sur0asirfOGIU
xGT6Az2VMaEabPfbSXRyBFcp4o40UVWfZYKnIaFUT+ZvGtmLQMJH+IJwg8bsXqC4
BajBt9WbeyCwqZYZwBj2WjjeEiose694bDPNUEVbEsk/xD6TSm4eGnrMIr7Cja/V
f0TzNVtF8mltgSm2EC95hRbuK2yr19AOwluQ4atqXROTdlpXuNnn8kfO9H9exwwM
/Qf+DUclt2c0mxy7/P9/PDm6YDhjn8i+oLy6ImER6d4PAfj6xCdNLkkauJQODV0q
k6oq4hrhsyuaRLxgCRtZZ2hGGo0BtMfECA70tZDb8Pzslt5Vgq34WaBV/7drFYDw
DbSAkYEpROpacHEw1ASrBi73DjoUIIY4NulGJenz0S2Tj0cw6T0qQnJD0KZPPSWv
30JyGi/s6w4Jfz57HoPPVY1tDCIBE1vFSbcv6fqxDtxsqOVQGD443hd1Nd3EPKTO
D2y6oM1KufotgEwqSxAk+K2CDotLgGX/EqW1LW8FBs0XXoJbg3SKsWJ1Pq3jP1qf
ZiBh7FIslZA1KFB1346LDF8JKygIDx52w4HBrK8MsEk0GAhz+oqwLlM2DE09GIxv
OtBN3FRvZrct+Tih6dBnQiQxw2kSzQoTnsx1Lqw3C182ksTHSK+G4z1cat1whJlZ
92R6DaDhE0zYP1PjINnZeYWvPtIBqgbVCU3huiNR/4jSU/eqE7dU7Dc0ARgi6XZe
JCds+narS5vmDHn3jhk0vAgYWioqYl0cuhFZ5n+piuOmQAO+jX+0I2qNEfE/9QqX
KOwJeLDRK+g63+Hhc6BeTdowr5RMMRYva6CVLbpr/MoRe7JYh68UNt/RanVwHrie
ywt91Frs7ecb5kvp0IFB8uF2Ji8VOaWga5nBySm29fLRyH+Fgn9rtJ+bHwe/iMlL
30zPI26501Cx6JcUk5iAx4UbDa6pfl40uTyyMzHK+nIYoCbNa8CAUKc3uDkyroN7
TX8niLu0VRINfUrC7snwqK6g12DL2/+H9BUKcbL1bOF5ODAJmbh0v0k29UUWOHuw
Vczl7gcvTMnCBLm6gx9lyFtAOsWTCxqVjehd3tHx7lixcamtuaTtwPFp46exhESO
i3Zoe+MgNqbhF7UIBi13eAUyQItm0RSO8z+IWVTsQkPM9OLCr1YXOIiLtJqr5TG9
+UsXtCZ5YIZMRUwV5To3GAbfOILWAoxXWBcWbI36X3MKOnanH+ZsCoSR0NiD10LF
gCvh/ShogZVqEFEWJMgZM06zSKES91tvogZMoUiEUX3OcWy1vMZsqmRGQ/tEJ/nE
y/Hh2rI3KrePpm+lMJFnl/hKcqRzZ8bRLcZfmEcUd/Liq+PTAuHET+HFI2eqXaE0
PqlbQWnGU570kZHeV4Osm51bQDZyrRQJVnC+zOYuyg9RfC5KopBHSvJyh5UBGJuq
6jigkEotVdN8Dx1zXhvOSs2rCs2ZVaI41Cxqyxxw1YCcfbgd1f6xlHR9I7q+KQLO
dv/zO3MvXolq4j8nhJAkK+6BaBuPe/qCL55Cic3qKfuctdUAX0Jkz4m5vk51354f
XrzcS6vKJEQrvbDN9osIPisiKLTP55oihwS3xOIySD6lpAp4u/kCZ1QzVQqViZGk
ZpBQFA+PV4jDYXoE4qLFH2IVk/DeRjMdoY5Ao5+zUZ/kiSMNygR7f+xm4eo0Tvn8
/fQk3BI0SeH+pzAEDDOdDjT2COWO19R5QolzrRMB4J1HXpS4zd4B40y3uRXLbcUE
uJGOItBNQ7XEgOFOwDdZRAR7MBCJsnGcMEZHAqPG3qh1QBDwFzR1EGdEU9Yao1hz
MhWURUeRa6m+STY3EKpjZo9Bw080e9s36nxucrzosjrs0E1ZHrMWvHBAgrXuuU1A
bdbTfIczkPCPYdD0tqv35wjcxbckq5URim46imloWU7L6NyCRBtewkp0cHasPaea
cbOsGRoM3vnZB9kgJSEsUE1UZC0zoRPLnoe6Y/DFKKRrsXSLgeljdazS+rTrKo9D
IMhdLFmn09YYrcS15NAC8C+PkTJ9F7oF9It0tIWtdqDBhvA+lbFufSAq0qySnX9c
DJrXXBwnjbQ1981WI+uhPAV6q6GmftTaRNs5W8Ic1rD9aZti8J0AGIDSKfMPCSPQ
+vn3ePzKm5wC/mzPFmsQWG/yFj8ISrByse3rPkAlP1QxSMt8Q8LRytABtN6WMrQQ
/ro8XlsMgZh0iUaUw960L0xEX8FNhTK3kE+4QzzUZTjcDO7486TdDCfVOiZXIeA5
umJAjZQ+iERWY6MAEVHnHSYA6j0eg/pscevhltJTgfBpdptWgGVoRnbA5PbTx7mI
bIzB6ItWkBuGiShu0kqYIVJ3F3QFEsVnMX/Rwg+Ol8UqtGlNUwpyVUh1+slPkvXJ
5IKbsgxNDTy7QVxAxknQS7s1kXKtJ4wxkNkAOO/LF2gNvzmW6dT0GHJ7fePo25Aq
ULEhZSF3uth2QjE3HSF2fM93nWT0V+WbH/DkB+NuXSqg1mcT7u/pobrmjuLUZ8Rb
YZPjzh8WWtvc2LhkJIBAhNgmITr0101p5nYq8/vULElJ1CvTfZJK7Qu7T6zzzs/U
c1rTT9IcKXCav8caDzpJAeziOOkqkpPJOUY1UMKkksI87/bdU8t+84JmtHcJu3Mn
2BbWS1hgc3ldiUIWUIzsgGKLmznmMJi+VSdaGCDqw58eopGSg86/jlWbz6Tzcmmy
JL4vx8DJuLmsjVqL6v7GDibHRb3ve2xlrBlzekGMFnmHZphjckDV/cYG+WaXNuV+
uNFhsq8V1Ce+ogu4iWg91ba/7p9YPVTLbnIrh2PEofV+ZnuAD/jB6qnRzuXCyiAr
EfW+NB2/3kM3ALSl/yEAsZy9ddUPi+FmMLVKb6HXP5gIKo1l/cs1EyS7gV6g+YkW
IOqBwfyt3sYA9gApIs0Ea9+u/1Ne6Ckmbh4zjxmkq9q/ZisM25leEkbS2IzSTjdn
qjVFdbzYlRL7ROdedeKMhNKSos0vqs7BQzHFl0wqoSIjQd52dgnz1CA9Vw2zsPe5
kO4aaKk+IkWIhoku58cKPlcGM0hE5iB29/bq6yJo0vWyN1qMJLAITe0+tghzWvM1
7eI2L06QwRldRXaLsPMlmWRPUQgdMxIvPSJVKp//G4obvN/078zQapflWo0TaZAo
JHrjoNiRJ4gwccro0n3BAWOZQ9sx34eTf3d7O2JAF/W6ekWtcnOX1WpXbjj/XMOR
64K+lYF+dWjycz8gahHlhp13I9VivD0t3OvyVqNBBCV5PvHI7PKNw7fywwvc03qh
P8lq9ZAS42c8VRl1/kvmFLzXdj/Z1jcOgb9ECS4C49uhLdlk1ZBDQQbH2IUCXfvT
wk+ZfxC6EoaCsK2QSE6+0k4mD+rZs3EVr0JVYMNv7AzwxBMFfEzNJQUuXmyPf9tC
A2gSLQKBJ++LeRZ2V+JTWQeZgqI47LIqrHkZptM2+Su9piG9Bc8ix0gbzIrqfBla
L3hRwTSiI34BhOK9Vp46a4dAO3fQsHsqdkGaYivzceJEwJBbpaRtGW54igXh+pMX
QrNlDwXExMj7PEtkYPwjQAdwo53MNMcHnURUU/y2/u7v4bM33wrf89+aQiVC/wnk
bX4+4n+Aa4NX2v0Un8EvafWBBRFMkQCcI0BUgB6STH+usCHix/TSHupty3RBLeBC
+w3aXbxawyA5vIstINXETojtJKJ7g8V9eZ/I6ASTRqw1l9311ZF2zTMIYmG/Pd9B
18RnjLj49QZWKGfrx0vm2/KModSMAiWscDVa/Zn+kWWyskSysdmI2pmxfFqjb9AH
jTdkcKdMPTRILH3pHcxhS0UF+WNbPgkaii8V5+ZPmTrQIbzL2JnTishNr0r6cFV4
cX1pgtC+jHqFi7e473hoC+DpXjQ2mGow0hicEz8jfwfD81hLr+awxZm90SZKS6v2
zmrqh8JjQHbKl+oj9ifVA+k3rwNlRwOSrJqvCkDqexKziV5410GV3VD+lSfLUOIN
Yq/6Wm0Co5PEFIzGwGEJxL1EhduRRnNeNFSw0xOhJqBDIRQ3HW9IaLfWzeSsW7d/
rouuN1QjxI2Eki6biTnJImaI4B4mg5zYNouXqus/Mmf7jauIXEvG7DngzN8y4oul
lxOJ2ON1EOjr7iFmg0+k4uS0CE5D3r7PjxUiiLdgIFMV/nSIt5bYD81TquJDgnjD
dV4QLEu3pG2D+AmH7TrGscyXVxdoMH6z575YMhkmRglm6fDV7capJi58Fn5Degh+
CZfOTBzTx65lc3U1b2Ob2VBYA8OXmkl0rVioyg6KWD7D3y09/9E9t3saBejALNDV
RqKv+t1+YPakAZPKT9xFkELQctsbNgsjDzXU/08GIFkQ0Ac5/LOczO0YuDvFbxMp
iyOqHwYC1FeN6De+qiFplHxEq0P9OP47nAgD0kFn8eOXOTZFXFPEUrYY/QUK84wy
S9LmZlVECuiJvsMDaIEsxwto6Ndzfl0mizLtX8rMJK4OzmATQtNtDOqrZk+6V7Xz
C2jQ8EhWPicJIWlSK1jqsPLsTH8n945cQpsngSzrb2F3uZP5tJ8fgouktyzs8u+Y
+7mljvEZBkau5JYy2vEw1Eteo8OzM+K7eqGuefTHFpguojyz+GUEuRxGxYx/MMqp
WYH20p5E/IBOFYhOKr6yMi6ScX+vxASAG+eJTYINPnjBxe1dLY3aZrLh6SIlK+0r
oNLY1HEtfhVkWZeYCwIs9l0MMmzT/1OAz2x4QHkz+8IgPRLVSnHkfXEh5PV0TnvG
UwQuKIQ9Hkh2WYdt3yV1gUB8PUqLjL7zDUInXTre21WuS1N7nBD6ROcTC7DkhXeA
rxj1s+778mQmhKCNhAuEzdZQcGdigkIHOuCDaBwPfLnWhYI00zpQm76KGvCNFcTl
zpsfg0Fvl+RydVrwZcGwp6kEuGe+i7vCQRvdcQtPH7ZuEOHveDmS/JC2Lj4GC4rz
nh1ISu6D1quUMe2mM5qy+GSYwBO4PlEv1k6L5ekOv/Luxm0VF4QkQKRsLQ668idw
BJ+fwnS4vxKuEodzdBt1fc7NiCW3R6fqxp+3I7GO28+HMLgzO49NtVyumQ4VC6hp
ubctrnAFvD0tYBZ+MYX8Vt77OlcWfnyUUSetkgzMZsDWfZzOenQbF981F6Q6gK3X
ITzeIUz7SXjthxEJQ9L9c5tQzAxmQJAXggGPS0qXpp65KDjx5E/Zc/79etGtwjoE
HcoMm3lvceAKfv0oO61A8fXmsIaOWhpz7Gpnoi3Hp7xN8VCZ+OKas0KdyNg7qore
7qqRx3jfkeJL+bCbByzo3QXOmrtWR5hJVF3bnF6ElqBFJHKShKtJ1SCW6xfHEVJX
/ath4WydSGYSH8z1+BIQtGE/lF+0pxn47YwfamESMw2rCGXaALdGnwxD9gh6Q+9r
gH7Gwgv1rrd2JLd4jOtptoQNkticpGBsQ59sZuxMNzjw9eeu9NvjmSgtTOpmZBSS
lKdDw/ngz1z0WYtwhbqImV7l93wUcuGKD3xjVZpSXUwJfkCZchuL1J1Omihykd5X
PHzZ8j9ng4tPyyUsJON9UxQ69f1aLpcS6cDucKsEl4Uar/No6weJ34FfvM1torUA
XbRHBC/6yj3MR3JvDvAx2qF3yle5urPGCc9yevCt8Pl1u64F4IDeCe0NwGJGmLal
G0bbwTyMKhaL9jT6E7WK2uIkJwmiwG7KmxPjhIYP2fN6wBN3sHiRwQKjh0qPo8jh
7aB4kbhkuPHz2sNRdnm35r0N9fCAjN2VT0dkHtXO0scXwOX/L1QOBZOZoNQyrV9V
x1WnQGBBZ9XLU4QJIRkHZ1yIaXjwPOvVGY96XAcDs9bQV/SnS++kdyI8SbUTndJO
ggr4kAhHqCyPPhqAiyMlEP3luweLkrbbB48izsWLi8mJnJOSoJJ2/2mY1XnFXL2v
1aiWxxUW7gGStvkl286NeRzkRYOP5IZD/4lV7bmNH0DW4rLDbB4m2MYVJzDqMlcr
e5zIIk6HFpvXzWGtsUUL53WVB1S9XFw7jVWT0gamMCtd0YnwLzM1k/cG7VW9izNR
694m5+vEzEdn3fWIESgeCMJRQPVqU/UR7R/cp9ZIBTbqMnEIIzGg4t8bHiaJfWat
gWkHt4sb5tDnrQUafsL2yF0so4vDZAYQwiQn5dhG+lj0YtQ3qMs86M56R9bQgryB
dMRB/D1rXANX0nlvQ14GsvbqYNyEpTzh2mYjbvR984jnkDYW14L5nGorKN0BrhIS
zxDUvPMfpLipCZqcAWN7HpIJCqqLOmzuxCb2Cv+wCJ4GkLJfAMSHasUgtZbrExfH
K9Hlr5tfetOiY6bYvIZV/3KtN0S58ED3NyYFQrk/A5BtxNcT2LN+9nUBqvxe/2n6
oY8gaZWKZVcqUNnqjrfOVZqlyQMahuOjsXrNvMMG2lrpYWPpUqNxApnWXpOEd7LW
R8JnsFcA0MiPfcNlmewyygssFvLrwrgAg0i2mCSYO4U17ZicEZy0BNHttVnCGrQK
mgeuEwrhh3ib6Jflqx8AHNIKcrL3N1cxe0gglTk0qMRLa3cBdmU027UYgoxDdzxR
TqFcU7sB+/GLfVkHk5h9J3xy5Nd5J3n5ndXfOIENpiwg9T5EhI5PVerhqyn+Rrgy
NEfN/lctxhBB85+mUFlsDf3KARtGUs4uIbrbM2JAXa7t372Q0hNEY/EJMAhqoQyH
dxCgZnCAtAooFju98sX4J9Fi+eY6z8hPbDC6K5NJCw4XX4C3Ja6SEsHPgVyBXOPU
OY2eRu+v21qYT9uqi/Njr0k2KvsAY22t1SFrjQ5rP20gUIsS+U5V70PovBzl32CJ
VWib53snjOB9HPChgiCVsu6y9jUkMVA6BB95rjmaVJ4gyrCCl2LxkeDWSFdh9yiN
bJuaTIwWTyJGPRu1QVqT7Tk9tKr5aZpAmEogpctdYNiyR+kHnrRwCbMaMbxRX6PP
ZNqzjiYkGbpZuttrTZxbTHBDB0QpFEJxYoS9YUBTerA9zRt3OwsXz4D2NfN1Sa1R
t5G0gdsskgu/1XzKBLVyAObBl4dK34ZKSK2yt5PUtlqqV6x/Sk4s1Dayu54VrU0F
PphkWgczenNQxH7UCEGz19oxxqOEC/8lHm4+T/7xnsE4qEJPJ5KaP6oXA/sPBy6j
ob+BdEGrrwc3AOIrhmMAT6jo8DQ/jzCHplWWmn/QjE0kCE3iMMKBSPkslPzc0W1b
HnPXRkn4+19rwyUZy96LjNzdsafRI2aMrWLuH67mpZ3EAFt3nwTQhgBU3TCqefAn
cP4U0r36M82/GevKVILICBpcSnXPuEIJStIFvDwXU6Utfj9XwvtmuDGJ42gWsNK3
JBMZAA9W95d2n607mb8mGwDzvqEzJVqWhVR1aLBheYITiTJtyr5tXmZwiXWk9eWO
qN4VZEx/Fo0xlWjqC6Er+c8JS/AGTQ/8XWdhXLwIIfdJZDXk7Rrw32jqNGhElM1a
3OAGmYiPb5bBBaHUX0e6fIV6GRRh3Og6ZPkUSYiOZZ9KuABIjn7d2P0qPL8BZes1
YeUC1DIY211BBpjnEr0myYJ0LRzdviJxa2eIzPqF58TtKoBvd/aqujFQbPqeAezB
uyEgVYDaHuyJafrhJhHIUpqClySz5ZFY5HCtP5k5C95VScwrlgjMKIVv0+XfxyNx
pgzOR/pQ/hvPhMonhl/JRbzSqK3BaaGfHqZMCqWLPZSz4lUGJ8oplkK7a/cnvYb0
Pf2busemhEY8Miy+xwFyWsL7pm/bBT29ebBgO/E1qyei0vRBMjTzMEjBgSNQ9th/
plUXKG/vsLOxdOBMqVMWSKBHT5aaBlIQrYvX4udOQ9z6w0y4OwrJge23AlJmqT6z
ZSAnKLWFcfYjblxWzMhnNLdQQXpneFDDe7UbYYiBjP1lN7U5AOEvJG6gL5jmaNn9
vJwVRD0cpm8phnzQtNU30kzfaQUgOjIpPz9lVwy+KwMBTcAcQiTv+jTwkvpLUFMU
ePisu/0992mpujd0A4phLSmliam/ltj8eESyZhwKYsdP7JKmoFPv17b8+ZuOl3+u
WQnUxPeDlXtyjICSZenf+dXtMY+s9A2l/daaFfJqf74ZtI8wMtZpLN2d/8Kq0XWI
nDwNvD32/Nzxk1p2Qd394YCoYHaDmFHuVONyMptmMR7rSJlMO81tggSX/j1yZ6Rd
OsukiKcmvDKidB916aXwN0uD1qfJytmrDXml6e4nE8v+zokv/PqDkFoILHxPyCLK
7c8DikgxkQA+vKBZR7FlMIIf8leSgY1ERl6E71Tz/i8/Tby+p6ZtjIwdiVtAvxcC
v2BPmyvfQMHjto0JBzFgYcEgnrVqOMnWg4o+k3BoDbCK3Qj/yx0QDnpjgGzM791A
g/8BZRfgGw7+o3QSkr1giME2l2EexkjPncW9KmFgXT6wtE10dJm8F0YkcJD8fYFu
L5LTzj17G9JNfgd1zO3lIO//ocDhRiMhUNVsrOcjleJNotBbWFczrX21BWi6qxat
kCbzZX27SFMD4YFwWp+8W6G8Esm6qvvA537Wq/kOJbh/9PMfBXy4wvcDLBd39pfC
5AZnqEU+pPW8FUx6pi8/HXNlZmzR9Dj3eR0mmguYpY1W5IZOVc29hTlTUc9AbzJW
ZlrC3uAGLAPXfitED+jjZo/89urhq4lSKyFHNICt/p9jNuYvkB4OF5dMPkp24vii
hB5EASd5WIqRKaTS0RblI2fDgqyaAGIVbmvftM84jRD0Dp8zbEfVS0aeqfJoXG1s
0fzWt3lDrOrAnDxTckqPdLSTQ2GHqL118y1Be8oKOVT9qQVm/v/6HJIW5YEvNCp3
HUbXHSsnn2Zfj5l2XgweWnNAtH44TreQxHbI7G9qsmGDhMDYR9fWk8KjDFq1/U+8
+6043U0tPTu3U5jWzty6FOFAqbWQMFVbZA44Pq8gJoDk9BNzsZej/qDENhevk1fl
3gPSgGZvWB8mRKXVugQSIc5m9QjZ6cjimhf9enNpAivCvkZgELNAUEJM0rZPJQWs
HdgfWKtBIhLU6DvkPfM50dWmcYbqSTEnmHD569UFoXuhoGywqFmTMRZTtZ+G/OJ0
p+qFBhBR72VFvX4v2kAeeL/lng63qcttGOIyt2Rric+Ix6Z5sOFHb4aZHStDFpIC
g8S721bYoXxYyDWCZM5NLLEGjWjj50k6eZZ3sKZ5tK2u6nq9tncR+hSeRkLqGYXc
XlCopWYutMYdithWHyGrZo+ESx5z/1qa1qRcKD+D96Q7+PDc3ezwJvfkY3h7j82m
U3m74vmORDrL/415licLWAA3xH6ouFV6wxQ+/w0G4iDOuDc29qfJ5D1sbW1qEJbv
uHF3xYbLOJVaQmahFoZhQXUoJy4uX5LgrNhBIFUNZBNxmW3nxfc4TGx6prcb7mNI
6LOMXaEg+LpXRNhLum+iClDdJ6asO+M+fQWxl8RuEn6dcRVMn2rzJSlF1/Oh5jKF
/42fSz/zM6VnpB4IVppBBgjzG9B5HbezMjJCZN8Ho/6QUnAjzLlhbe0p93kGtCTD
ElyurCKysJ7CqWbbWzIzCWvi/Jb4C4mRmjOQQEz8CslggYY85VVvH9P2F2scz2+5
LyYY+rBhQGiAO6hrowx7UDiH/63EYBVgouS/vsn/ceyLIEXVCRTG9LQ2ZqIfBHZs
gFH7javYacL1QMrutN1ai99G3jxpPcgh6o7+VlzyYe85jeLro9o1mCqaT8KtbmC9
fgrTUro39OMeDrv+hZiU3RYekJ0fWBSBCNOwEGMsvR6mqN5POXHBl+AzzAh5BBVu
QgZ+DsUekIKuGzqfo4BcXgSQzdFUy6Y4ezStLWxWGvyxqxgORGpM7ldtiLSJKIFV
tDK4i/V5kOPLNufCeIwF4YZuwDMlyla/gOUyXJ8xlUdolTRLpxG16LB4OgQ4zY0f
75783rdHhfF+Zx5xHt8yCXGjQ2yAf5W8w/r+h8dWS/4UuOo7Ivl5C+uhgVqaIgEB
b6SfRpHfIhRRwPo6q4CoOnnd3xM/tcnZ2EzUHRsdKXWYErdebfbSwl8TsoPfeX/B
39y9cly7Mgo7H6aiy59o8vdJSFoPp1tsPLoGX+AHzFSgrm1CJuFqNHX2S7bL6V6N
cFDLMaGtOR1L3GELN+NG/00CZ3EbA/5o4kM7p8g7va5lkbQu/C9K2wqU7oJLKtsf
uTzbNjuajaDNNrON/s8vZbYdZBWWwn1yFBzKOD/m+ogRqNad+o72WkyJmiMIqJEN
nlCppPmp2B7rBN4DEYYy7Zg4l6w4BxujHi5ciQGMJwPkxBVPkDqpDcs23k43OIDv
9tOhU65zZhhF79jk4xI8NrqmUSJikzCC3I1yK2p2qKsYr6PspON6XsnSzfG8rMGJ
bLmiDfdb6AvZdc7BAwshzjIrz3b4p88ELIOQLfxr0SCloLVgzsTkcz8aIm2LFAeg
aWnc2s/XT7L+zCPA2IBcTC18S6QC5kPm0w1gOtmih7FCss1ad3Rv6lm+r0V8CjkP
UCLVAAwY9R+KTPmJ44ib7uzqeCU8tjHocmGzIq/lSfbQkcBW6m18Lys2Zs6E9D/C
mxswysxZ7Sfswn8w8HxRVunil0lGoKnHGVQFrc33PM6JUvylWZzrk6gAXhLXT07z
5gosOPTT3R2ahUGxAfVSt2FDp9UXdCeCfV3pSiWAbWJ+lNAZTmPD2ffJQj625kB4
dhy1gGEqjT6L5nBfvcne2uBKLI9toZmyYDO+/GkwIyhYvHa5gLMS9s6sQ/OM1xiK
0Kwi7kCiHa1bWHc+UQC3333luC+/ndvYSWyqNbv3nO6w+NXpMGTb7M221Q8vumoV
vgBfeumMvo9+UxfJYNHLBGOb4qFHQQZ8/U+5kHzyAI6W/TrN+R49xAqmt+ZIALY3
S9VfNjvX57GZTkychKwZb0JBTUF/I+ghuV9lYah/PTKX4wvU8UA0+zjGHU1lY6Ty
R5ZbIHY1xfhUxpXuCnoUIs3a/bQz8ZnXlZSCnEWyhRTJVFg1yXGKwaTD1iVaMwo2
3G6F3FB13Xd9AN4hJlem5OIk8vb7WBwY1KxVxywGH1KYxLpGUkHSuGjEK4/yn/dQ
MLED5Aaqlg+LnMgQ20AOQPVyNixLy0q99ZDxFq5hMi4PA3UVf7hl1C9meHoFgHHm
+c1Jj3k/YRFX5AL+w70u2B2Ogf/oKu/iDmJJyyOJroPTnS6fIicm0QFBTIVrB0li
rR/KX6UqrUpc5T37mthD9bY5i5naRormu5S+dIkrsaHLRFonxoJmgz2n9n45aXuN
/xwWbiqvyZHToQMQ/VjR0uTD85tdvP+BaoCPRrfvStaPPiAV+gvbLel4Uh3Baqw6
NkXDxsv9apR3Up1CPBkl23XTTt3Oqwwvp4VDkuBtIbdQ8gyIigVQuwsx/U9cHA29
Y/wiKg1/ArLwyDREaB1fgbKiQ+E3l+3mwxwDxuFi9iercZZ8zaOmYhpY+NXG8KoU
efvYxr22JdUTiyf+9adHV3QD9j7u0df54r9bFYHStM4RvNfiuVji1auQYQnw0/ru
7rsDdymk4TEmbD8UhS8sVBN1fR+nlu8FuOtQ5SiDU1VGsCHj62PciSPXDlcc0rA5
zLMZo4k+TKOKH8Nye7bVKpwAdD7nTENIcCc8VCxh+QQrQB1ZJfj/ewMRXeFjm4Xi
+8NNK+NqrAPqjzeOmVBsMQjZpQI2dxzlwTJ2uPYj8kD9GTSwFOLI27N48kmU0grb
jXmII0QbkG/nun50NErO+nBWieZV3NujR7YG5gAzKQCWPsXvVIBacE98q01wMt+Y
qqQrSXqEe12u8P4LoWm5brNveDyGLsRS5zRd1rLdglF0saRIus7+LphGxEFHUZwy
ZXu917IlAYHFn7HVU7YDbbS/lLrd0ivD81b4f8E3e84KRDziEpuRZwUMMqeokxv+
VT9T05z2udW1AVFSdmvQw1JVGIUhJJN02MTP5mwAZPKdUZeiFYQKhMRGxfcERRRd
rrYzfdtfB8YqLVB7PG7wvOiRumFTtKelX3+tBOlPP/ouVlLtc1o+dZ21dmeT8jnf
o3M4tvyC/oOt3vAmQqVXFfyZ0Q/qbGY0U3kVFMVA8mo1EcE4MxfZM2jw5X2DBHZb
Z2rj6XWiVo5h37ORm3gwnwjreE1QEAd0KQrTS/28L2MIOzXDf1b+Sry5PvsK9RLJ
IZyHEKDw0tCLzs/Y4unne9+kjEEQVCZR0aJv+VpmeNG50Jq6ey0CWHcGNUTgom+K
HjLFGjg6QlY/s4zj9G9wtPdEq8JhWQS/EMGC/aRxgyyN7lWCS4x8ocNfvRi5Kxt4
600Y6Q9aE0/rfqqpy4/nyL+4WTmr7GOn6lDF40NQVOguhaL22gNzkS7v/z23sk3A
49Fp/i2ESwTNUlKNGIHvcv3wNIeJH+EZs9XqqjXtayuxXbhvgRhRowCZbg8xrIBr
RmunYdvG8Ygkucup/FF2EPe/b3ElgEX38UTNCI9HxioFyg2CoGRiHxQMXp5xJ2J1
dncBGi3cepO8b2qJMqqBNVkAyRZGgxfZ/VIfIWxzjyiHkdd0A9EJk4VwzEkS8cqR
g63hGSgJKwbPGJVnRi3qWYf/XRyrkxqhiZVuFG1aTUf9RVcwUVKLSYe31TavFO9c
7dRAqyTJkk69iZZHDJQBJQjUrdGNGKT61sHQgr4T3kjPpyQmaeQCHo0TrNbxcTPN
9JcbqAEu8HkwEjVJ9nXN7xJGimDz8LGj24de4kwUcdBn9oJ/Er2fs0yaBCGHz1tp
3yQNTqf2DyxvpoWHoIeoJHqKpAk9cCyvxN8o+6P9mEey0TMJthjZ72bPmkQjWYkb
ApBZMSGpw7xBVhPfKjwHXJ0TTZh+DLx84eA4hYtbHHeE0Hfz/gkrlLL2/EFvruGq
cBIhO64XXiUiHaniUr/8+lvuDPOFe9kC8HFlKr4yu6OkSam+uDdlYF583gXJbBAw
Lbpk4yM0Ecir4X5ouGZDR+hNomviWV2wPg6UYlEpwsHL2TbVrTLpHP0KIHM9+0I/
dUk/UKjpM1hQnkrsqSB40hQiacGnWqt3wGmlPjMihiQRwUHe+RbN9ELkuLjkJQJo
I40xL7HlXS0nN+Vf4F4ytyOOP8ASh4xbOpLl/DOd3QH4Ahsaix7bKWGX67HCnyN4
5yYWV4jVoQdAL9fDW9aUDEnXnJBwJIzaDLpWIsuoAviv0MAARZHw2PeUcKv+4jwN
p3vZKX10LqRzdUJ+vqXZ1mif6gVw7LTADoGBmMJitIRRLw/NHhZXA8eRdtdILjYg
aru1VMHFz57tIBq8LhvymyHnmT5ZpVWtNK3+Ph36kCtRUJ2hhB8v1ghiaIJL9UaA
k4C7MQYg6yMNh0eneXYTEhZV4/sL0G8IiIzR+QUq+ds48w24sZCxgVpSr8xgzlt7
R9PDu7R9RDp8oj0y+PCrYLXM7+zeIhMnVOeOv6860x438St5w87LyS5mBMEAQ/TK
rMMz3dJHr99MdTGQ48lSHluP/8W3MMzyXcjyxmkrKLd1AoKPTEh0cS9PSnHcMkWY
W5CpHx1Vav1A/GHB2C1iTZTl8kjQ7O3YQhb3TRTXfIZFL1M2RFACbBIqjiyrJLC1
b5FjuqWzjwsNuLxWocMGaP44ZYjSMJ/Uh0iFIoIvTmgL+CJpXqerP1Yxh8p48D5B
7L9vD7dksmnHb3XICU9kIWEv5w5xEAIfgPowXFNrMcnPKrCClqBxDkMRFZ7jCj59
VGz/38FebGUBINpWOvr7M3nfpPNr8VZ/QVm0Kz8fTA4LFFV4z41K6T+sHZS2EMlR
rE458JcY+8Rsxk4GoIqFqvu9dj949ucZmVsVFrWlHmyaByTcUtmBB/oL4Eq+hUa0
DDirSKioUNav9LZaOQuMas0APSBzJSA2V7EAJNHMX7jdltMxN8gvgTUEF8+t0nLT
k8rH+QQHUvfHU+Ygutjyn3CjK/Das50h27WAz2h8homgnmaew4HFGw4GqdqEVqwz
ps7dr3EkzzhmGtte5B291G3HaaXBZ0R+5qju6+0ZRXhGLTQ9O1RRaaNItiRPTURl
mLjjUv18yR4yqszYNmcEWQ6UyrECN1knozDaCgHJ5O5KVIHx5gznX7SCBWiP9ZhJ
TZv+Jzk/+l3GIB7hdIVz62orNRA3DMHqqaPe7ectDpxUFO/oujGSma06s+ye+NO/
oJR/akH9RbL9tZAWpgHbfa7OmDr8motPC3eyxxEUgwj75JEZEHApy9lEQQRTWqqO
O5pBN1hn/FPMEhRdGlBRAcCI5OBtTounYWrUZSxTeG8lmg0P0y7x7h9gsNkEWDZ4
+ctbRGFeby291YCl2EniU17WvGDvonA2oEFbhrtv6uwrwR7kgBJMlYm2jYb9OKzm
8k5nB/HwUuiHKP08g7g44ROKlJGokX/t9IkmDK8g4MsP92BLt6s0bpC5HVVvOxpE
fahuUld6cPHJS80pSmuln7gYeCGLhppsn8mSOyYxL5xnlWmbwvQMPDf/XAx9y+f0
SrkJI7YpCGuOMGmQzBK3p6lcq8qvucfNAopzLNSIfAT1hBpsoELu0mW5iIEXbY/2
oeVJsiDnoveZ1U064O3M40qU38EjJUt4JEokCJ6jfB3F7lzqu/JxPyOqj0UeAMmR
hZt9Od7cIOA1ovsBz9uT62yeKKVupaHmj3wgXtWMXaB5f6utur6QoIi7LP0ZMdI3
8Rrhd45Ro95zhQNyG4ma2Xfr0k5GsDqL49d2rx19c96YTT46CxCwb905ugv4uxm5
tCqE01OJAnwQlnTVmKM14Jcnc63VzCa3hymw6pcbw20zBJ1qSk2b6qBrzOwHcPw2
+rKiThyb6aOUI1o29PedzubfjK7ijcR0R6IMVHYM+BWWzEQr5p+gajQH3Bl0yNxx
wwYtgj5IgOaiH6uk3NCCjb4hqWw1qKOyOFdEU1844rst9Z3J5UkHdVxGxrIg9GwS
IGviYZQ0GI3hwd02bjixL5n+aMyS1JFy/Wb5c47hCBw570BSnotW8ZX4D4GmuKqJ
OU+/c0zSoooniHT3tDztAgoBVo3vYGBEGczh7Wn3HwUey8K7H+BrfDl61MvAbgYM
bYtvyaB6ZCa/eEt/gPO2hOfjq5VreApvDcQkHcjqreYP4UwyptXLclue0Zjn+cxv
EDoEAKttf5nkvkvpsjLT6CFTAXb8Cb2ps06MDtSzhP6YVZSUiu0e+NRoEXgFINQP
ETzE0h8MIjVdftnzrSjoog34mHX6F4v5pIDMlu3uC3sAfNCW7RQJb758bp9lUQTK
A2NPLxpeXI+Hudd0v17BdBSXrbWNlBNzRbB2Vpv2UOTynfIqD11jsCoJPTEwmhWM
TlkRWWr42GIjHjr6M2qd3/VrVn4wpkcOdoBoA48EDG2LBhT0oPj08La1SeSmjmFY
9vNHYYPLFkZswePAwZwL4HLkyjIttAvz8lRopgIgpgguDvZMVJsq4y7i0RTpt4lE
Wg04j9RrHD1pzZYgYiupcrP1dCNsOq+rtQ4ExpH2vfvrtQky5O4AWQENr3dtbieX
vvKmP4szj001rskbRfLzFotD24UumsmmaeT7yzQYTVN5T8zIBEflwDQwDu0iZV7z
XReUahUwPRn4sdtQmZ5+1vfAsjwRKxlJH/vOBooqmtQHIq5rEKSbw+jhStOJYNsH
IM8P687JZ/YzqxLThsD1rS7D7UkJImTCGqxIPFPYhz627pS+MBDll4KwAOs4nysH
zgb45e+VoyyjszXwyKa5Os4Zsdd5deReeHm58jtIokJFIm13veAvDpXff2vCNjiq
YDCQyTGI9y9WJrEH34/JOvlYr6sjh+nRQ6hDuxyyLHy//knaFk6qeP8wQfICxJLq
e6R6BtW92A/oPU7RyHLUyfIQdS+lury4HoDdEzsBiG0tVOpWh1uBX1unoYRjiHOc
tJ9S2Of4uhWxlyH2T8kKFY+CUMGscLz5pKconRh6BzAg2/MAYF1At5OSYL+ol8XV
hKfTznpmsle8hmTAf5fZofN8w9DxIRXJ75erH2urOiYXnNA2RtX9+tPad7Z65Z0x
50AXxJZvKIEpUs3IFiiTIbfrA/1fjJA6utaQ5jCOeVuXRtuQIeoFrN9voOazQvz9
8Q0Pwlm/K3BRD9xrX0tGKC2cw/+aAdM+tzWRvcbRH2VFypuwzVlNsPXL9inDlY+f
BXO5uQyUdSOdba9eTtCc+Dmch9/pknxon6DFfakES4VUSywmFfAvTM0gMUEeh8C4
dLHIcRb5txDYhcQIGayeh5vX99IW2kHeWs3bJiQHP9yutOXoEHtxT18ON6qnNOp6
Ae3ArOhNdf3rHN/qOZB96+O/hO/qOmrW0R1wvBwIfLQ7awz3t5Vk5U/oVNWryUAB
4g+Ppi5hi+YVWemVa8hoaMVvI6GnIuc+rEFulOsgIFcfpGHOaDU3ouadDLhhgawG
XTZ1ZPvFxppIVgdiL5LeDSs/zrrXBlBVKL/smu0SStT+teGG/a0faBA+AIqVZzEu
e+FHDqGChyOuyPM1x17am+e494Uz/J6bbhQG5FrDHZhL8beoj2cN8Y4OfOG7zOJj
P1Ap6jx3Gb6cmNlxc1LQ4st5chIUVrT4C4Q4KE7INZU307xaMr57IVDt7WuWpjvx
rzX8ijAYNjMoT2zbUveBGgSprx8/bNBvocEqVa5Yq+IakSSGdGc6y+j/HtjMEFz5
5Ywt7d8v5Aaqd4CGiUZdoBezbaglmxP370rszlshh1YZso5jFjTIEy1cWA3lvcOC
ZEO5k4quvbsO7QsmK46iKHTCA1c9K5mw6fBSWKsO38y5VShhnq+gixZYNnS4ZASw
aewymAX4/eMUVCHfOvAhXLK6WuESwufowbx2SR8J4NXAMas2zh1wPajmOEH4qAUN
0S/nudhwV2RSakR/aTujJTpgB2dJC5IohklOy+u9p9MU83nKQuhi1qhS60Xtw4SQ
Chtej4DJRaO6mXnjtc3zNt+viiy5q+9AZXRA0dN9pKnfgi6uX2HuRlumX6uBU5O1
hneDvswMlI5HmvZCd37Bc0uUlVvagpjtgBqR4Cbj/Xy/3wOMBL+fS8qx3gOEHWLj
kTDjwSsZkcjJPLh14HWqX5VSTfQRYSFlGBkzJUdQTXbfEnLf/m2Jh7G+URpppQby
7N9BjNT9aep43kTs6BL4aGZ5GOz5UsVTSuMNmsWvENKkdLq2bebpPNB/cf4p3IHt
aoxgGWtbTM0fBGHF7QL6+ATclrY1EHTyj/SsQvPBKdRFzjZaGsF8UKWmrijanFZy
J048eR46NzjF/0ppPjnhnjEb0oA3aKLZrsNQd49zQpJBsxeY1SvHNELEidiWEa9M
MsqcLt+IGX24qFzqrPfgWxaMSMStjViZilKfXI0FHRVtajZFllMRO4/Ns0jD/NRh
o5jR+PSvIuXPXYjsS63jmGAy++9E2mti1vSy9jX7yp3vw0hhggLeW+68IDgY/Iy0
9HZQaaAvcIa5H5R7J4m3g0kY5CGcu24Glq7kTRjUYAi8r5RwdCAoJNmc3H6Ujfc+
a+12fC2AY1KTHNBsBaVTFxAPLs5ajCalv0zfMdj0fiH7HzTRdPsFs7SZvROyVdFh
Azw/NeEEWsplQG3DS6ncaOPatseFxw2lp6ufaWn7e1Rj+Jz/ctLmM6hvQciWZAfU
qj6wS37vDpvX/7B9YBB5ds+81GP7SD+Wbtx3huJXHnmVVfVAPfFbs8BMYw3Ox/mj
VXxFATuLPNL5/aKl8p20zjXTD5Y/13KgMkcw6fhrb+1CppE3knUxeJA9QaEVBNXA
SmCUGnJ00Wh3QrJ4aDjcdYyV1Ijz6TepgvgozKT3d+hXsXuEghlcVwagMz8Gd45i
tnIEGzdOZSaJ88exnoqbLBVlYqIFmBUgk8O/Kw/MNB9y+oe7n0FfKDBhdKAaJoRf
VTRuTGkyqFn93YMpbgysvsmCNDAnFQmhSshDMmHN07VamOMVziVSahpt8gDs1UP9
2Okwk6BzbM2E4U1D7+JQ5p5lWJkHogN+npaLGtotWJRBg+NtNINYKcqxmn8Cf2Tc
yiV+LLHfpm7MYJgG39QZHDoFu7fuo/tC3gJTwAPtUwn1rc85jenLZu7x7Lu8dbbD
LT0QcXIwzSFNn3x389gj3TcTag/EA8ve5OhFtLT1g5VOyD0UWrFR6bBLN7pECXnt
xYxj6aY+lv/5XYJ9lD/FZKplApmKowdnroW0TUIbUytVBw5NsfLylZP5bqCNG+yZ
RHQZZr1hGfBkJNpzwz9rvkMHy4DXSYo7JjyJ7N6lRL2Dz9tq8BfsT1/zI7lqa3bL
O1/Dj9FoydxizAj9hTU8LjKF3YIMDpRi/ns1Yn4Wzoc9b8cQAFyGseUDQIUqi51q
lm6n/y+P7tGYpAK8KTv90sCPa3kJYrQOeIdXcLoTJXvyS1GIQro42foPhjSZ6Yo0
rvpAOUtJjv4aSkkpzRnct4Yr38U29F+KmMUNVnUAVQLw11kS+uagFXMaPhWGztpC
xGuqxROpS9PZjCjwH3gRqN/iZNk9FjtjZ2Hn5Z81xhzYhuBvt++R4MEVlmPLyIXd
K6U/xUj/pYpXFcJbHk5UZM57IOP9ocm5IT4UxuulL9PwAPcj9RWO4sPrq0kDTu9i
ggedecM+X7mEwq+0LdSVePtU6qHTtXeTP++ZSgqkdf2cisdP1hKTVVcHnWukAEo7
mYTHwh1hAWuM7P0HEuonzof6ELYid5nCnwVSVZwWsCNUM0maYnA3QvQ8ZUBchDaX
ce6DD7vrm6G+KKI49TCMxmQpUIug/mLf6j6Qtx9B1/aIUKauecTFInFC2Xrzt/Vl
Hw74srycSSqld2xeHmMn8KpmhTdiQzQKXfkdPaUHay4se9eTJ1jUwjQcXJBpdaOs
0Hj9YgPeTpyJ0hqSD/Ijby8mW0LwcJZA9P6tya+pDFWxOGETa88IU53N0C6OS+nS
0LAVVKcf1I/iS5nvbLquKvPOxRwhPinT7QvJMPbcFl8/kvzpZLIOPYy2KQT/KiN9
y+9QLlLjWWy7OZksc3yR6vveMoDJ0NDQugh9m0GUufTzbZkT5Uhl7li3smhGyC1h
u6wR1iGi5gg6uD5mvi9yrltTohtV48Pg9CqjH+VEht0lQJY+YYkO+d6OQT/NkRPE
5AkFjiNsGNqrvkAjE8M4akSOPlQ5j7U7XWhl375ffXcCEQkGuevr+7t1UHk83s8z
MBq4NBfzD/KPzdpj/0+dVcdkN08zFGSZA/eZaJ1TlEEKnhm9ZFXfrrcuPj8vncHu
HnMvz9e/DKv2xk+wU26AsTLaChgWrrMJrB/W71FLYFJ7mIPAIa8yvAuxhhjopYtv
WuHXNBhLvkZMPoq+5K1THHdXghiYKnSy8LJfMd3mIDlyjPrHpKAnjns3Z8VoGj6S
hK4wJ6K3d0V2+OPrX8AYLePwojtofOQ6e+vH878dYuvdCSmr2WLH8FR01p2J9SOZ
ZpPm3aspqR12HAVINBdQVGBVRUPXJEVUPznxMRAKaAHmg1jkP6ag4/VKImEOsgU4
FKqe8/ngKIaE0dwXcRGbUuiPtjwzCGv0Gv0NYXPNXqUptbqQdRP7xbMZ6DuZMjlZ
Mbgy8Ketk4ncDOTYWv85KYDQzsLfxJOAe55+tgE0zvkOuF/Nbs4zLHwWf8S8L81x
MxsFKDRcAWdZqTnL9h7cctx4cisPmAoP+swAbUZqXGZKqs41lexOoluyGskBmXlJ
F3afOwRLouW7mmen09qiGwR+Hw/FFXXwjVHKcS54QoSWKd+ujj838eyTjFZbSjkw
GYgcYhT4bOhSd2JQt0Xe7ZsaCJ5DML/UE+A/JISPEQsLQOsL0NGzx5O8iK5cDDCI
Nliomut2C/hzN3A4S085Ndh7AFHWRLBCtzM/tevUwjUyhJ7IV6AqSvp8iiAEEBY5
RBlXQ8uqU9ZccT6neT24t5UCzUHU91xJLLz6Mm2mjpNRh1Ky+9gmNuy6CHq5Y8/x
fdz3hmzQPcr/tuRJDkfjlRdjwKKgJR6ObnldVvOXt9w6jnhmoEUapdkQOH8oAd27
71F2P0kwhUMrajKVvL0fUhW8aN8ZUGNnQ6oeN1c8Tez1aMGgm3WoeaSYlcmfsfM1
1QvzvSoz9nKZ7gwNEegUdLgbkqMVbSbvXFQqlMgaIx3lOWHCDKs260ctljlZUvsf
92OPy+1rGZkP8Jztc/TsGL00mKfeiLnLvkKvOHL7vE0z/IynJw0CbHgxMai5PcCf
oVLT2nVqU2cs2vNZ17yYsGLDdLXufCUwWGMPFfq7WwidWJFt7lRZRnK9KdyOh0sg
QNig+xHjkv8PhnuhJDlHQqvb+9S4kOmkKSZO7ZsL4sz8ADrmGm5b2cFTkaKaLluC
p9coR06UgyJ0KxU8zq0AUo7IgGzG65+qfBybl59lKFwBPtJN94pYJsIrTZ2J1Guh
xlbb1jY/2RYyncZeeyBBhzXxiMj2oPvxdLoHq4HE9irWDMw9cAGkRobfmVvyRwxv
PvKUUyV4OSOnYWhE54aacI3p9A6y8jIuA/rKdFPYfBQWGYNW0T7rvEGbe3E7RLyE
KqYcNUA6GD3BAfGwELULMaQQbbYinnUMwTn+9AiNk1X/OMw9ki0cvegQ2i2grYGn
jHbck1LwC5BMI/59ZlW/XT6sfL/4y1MKHoYtlQEmTkwbkl5cPpbzRWqCNi0OtxoF
0bocsG2h4s/zS4nVhP7M0OZCROXsUjrqzAFYhyeBWAGEIPt2aTDLpCyASZ3yEXBq
BACFBSLVQUyG+SARI6zXLKsrY4XEW8bKP94Cxt1TjdkqoUCjfcyH+fv1P1nR4HO0
ozr34qXlLGVfuVq9mlfZHYv08/9RvjSJNfyOd1w2BxM6h0Op0b1Xk81XYKHaT3kB
8vaSO8iuzZBADWWe5MaIZHDeJjPuZsJZ4J20M5lYvohGOjLw2gk33K988Bkq2MGX
duKA3+idStl3cNJid4CXcLs8N0XzTYYwn6ABKpHtZas/MaDytIxxBDh9kNyCELGL
DFrDuAuELzpuvYKgv0QvAUfzm4G+jCpf0q14OxBvuAHgsgtpgjbRRq9zuFsjsjwU
4YPgk/yUxJn/kLvKoWFNrVqwSnUIVHhuMLePQHKGohcNJTwHcvaS18a8Irfh1BTr
eejCjK7x9uSMky4UTV5pN8aMjhAJqqptN4cwEodzIeFCpntb7jZlEZLsWGxEgop8
PF8kacDYP4ss/nQtojEKRM0JMkF8tKBqA+m2oTnzI7En5V5ALG3OjdOfUdhKAr5Q
7+PansytWJVy4LurB+PyvaQVygR+ffl/zUDm/a2td60oVf7xzjQx0mGyUFq2qJtx
8O+0WBbxb8czIt/N7Ow+JDl5i2lLZAai67vJ+d9D53gf/OkhwORqW4MFEVo/PBms
i2KThK98Ni4k+zI73YagLcdVP6N4Ekg9jIQwbQBcr8g5pPnlAi30/u2rEWr2Mj3R
kmEBDxidJd3I63geZ9ZyBTp0bbtCfRky7LpIaYfZRxLPW5+55mVkaj7q8Hsda841
qmFslmOEHPvsl9bJL1NhJaaF/SzqqiLaE9c3e7+YA1uEyy0HlQ027Xrs7GEAHEMQ
j61JJnyKPjm5fFDxPA9LjAVAsDkrcNw0IYvtbqWtiLuPb9LhEp471CqFtIcBlS9P
/K5LEOZXtnKDcQse+IaSOOVFBCTBAbIvdtEu2X8bw0ResqrjXEp/f3e82rYhv+ez
Yyw+Fx2MaoMQsiFFDmH8OfA8fvVuxBpVCP6/SikiwQ7dxiS3MVBq0nn81tuvsxYK
zzT9reGE+BElKKEKjf5xIWMINOOKeE/XTJhUmfVgTFizD5js9RzIbImbl8BqpENj
2kKPIqKrqulEZKVzun+3qRHO0w6H2xiZCkHK2jEL8gyBne7NUW4IBGDj3pVfljpJ
/ENuzmRtkR6HmqKqlEvnQ/K7m/6Ctu8QKeG87BXuyeZZGmHTVUsd+xkQY432Cqtw
/TzlKPEBWQGJ+LQP4ErcyH73i70BYCfBnXHxh1U9Gp75VtVnVHkE3xq+O3XWsZxP
M1b3Zcd4lVqI2bSWU/EyxWmognTKFagdfSn1N42DOK2vFRogBkG03IrP+yurFiRj
XHLGIZr51sDliEbxrzOqVtaYM66K1BrOqIbrpjClCamWCzebe4+4j3Dx08AEzEE+
I2O1RcClIVUpZOwCdcYYbrU/JNTAbdZrabN/7E6+ntC1FC39j2cQaa5Dr5Ptft/X
Vo/ZUj5RYzpW8l9HkaseFrCE7+zha1hkWLrOIj2YXhV+F3nO88ETlw9nlye65dAL
D+ZVBYmszgBi4iYxvzfb6alZuYyNd70PCV4yvvBCPstyKTFYs7FJMuAA2DtUuzgN
QqExfz+Tu98D+kKQNhrHmhd9ZMbLoTot1NQXA9Q3BUQl4yjMnQNaWp6YqaB76CcA
MTC4LoTMFhAmurHx8zRiXectHZA0iOsHVq3f5h9qU4R2xUTmh47uzrtf6DU/HMb4
/NZmhUrRmiQPLmiOPbE5W4W/gEI3E0UkWGC/hlo4Wj9RpKiU0+DmuBEdpZ4V+U+z
24Dl5KU54erNJNWj7CijBr/59GjLdQUTpseh4R/241FlZOLbIeMxe30lLSsifeBz
yjM4gRuWyTIXZDBo7QOZIx868xsMNBtnCgLlQegVaunMFSGhK7gypybWYV/Ncec8
np+Ni7yiBhbAEvwN47k4Z+l6tPjcQE4xB6JtxhFf3ciYNZlcLll0CbOZ36dL49vV
jA6j9df9KK5AMpq0I0vtJ8eynUeLdGqVaA6aB7a5t2jkKEW7vWFThXAt50767BW0
GwniOGn5glISiB2i2Ayo5CLxYItMBcLiBoySkJl+JTTk2wlGIzHufp5lUWXTO25W
v04da4YQiE7ZWWdZFP4OBkmVL15U3pK3esR12iBgCegrzig97dIOoN4JbdcKT8UG
ErexKTwDF4Dv+nEx7e2Lu0LkQDI2MdW0O0S18RxFejKBasa45uh1uuzk6+CUzocs
qRRA4A+tjPtqw4qJjtKDg5yMbGqoGLoLe5TwbmrmVr9ZfTucvX7hMZXbQiKqojg4
t+ZGEw2pWMrhPhvOX6a9AOjI98J7be51Lfys6C1n9IUEwVdWw7wBBhpRumpTUqHI
Js3URz18aADFq8c5t1he4GN557xFmEM34OOqINx7D3afrvDdMbwCD70I7Wts+Qpr
JOIQsXuAVrA+dVcRP6CsZ7o1gMEu6Dq8F1XXjvRyBQWGRdcdoqGCeDHg5ZVZgtWc
8rZEJ+VZ1NbmB0venkWgidhwSyozcO/jT4zkhmVsa2LZETl3IF3WhoyWT7BNzRIr
KdKCx7PEZrbkg2s1gQYkKywly5tVz30Y0D9kN8Vk5aPpgCWOoeRC7Uk5/UF7mokI
1q5OdmtFCtZgOD0cM7wiRQ6L0SBRL2rgVkQcuRC2a3AJOlSLskpwIAaLU8rEqg1s
+Sjj6tqn5TDMjROYK9ov+IDeI3FeJUOQo6+j0megeVeUEYm33FpvjrQ8OXvNEmQ3
HgZyR1deAktMv/CjNktiIJsKzKnorwlJcuZPhmR7W7jTW31MeCgktXa2YppBXdCW
LaTr/D4/1B5sgKdshMvzTqrNO+igLHFwIviPUSimFJIycPJr+z9lX2b+lwIeQBd4
qfiDgnobsKrFqANScxdabfj1giXzdobySE0dJM75LZRj32ahKGUtLbOUSqFBrp9h
oUJCCwcyfuPwIQ9lsTuSiw3evt3VOH5vJ+CybpCk0fJlqcptyXnhyxOzdXbiZyYT
mY3tbHDFMKQIJ92LjFckJaAYFMZmD5gFVj+lkmG54Y68Y5eRBR/rE/5HBEeisBa6
W+JdcuF5j54G1eFmfpUHfjeY3C/bxxT3pXy5vvPRtYggKGjLcRpbISkGiBAaBWVH
c8I0i1qLovHTx+BpWshXDCZNkcwhgF2RtMO1UESXzhlDDJJBe96sVdg7BIy+s5zu
k6lis5CPqb3XWFZqxJ3ysFKMrQiN/rGi5uf4rTYa1g9O0MHL276Iqv5aHcU4aYD+
CFVkpHxwwgJET52VCxLX80QT9i8VpOOJnyRfizAQnMQjAH0sv6MDhhvv2rd2zSZH
4AFkPID52bpOLUqHq/CGz90ZDpUJKIeeEE452V0YWXvIm+MwLIfOMTuo8XCeIgdk
n6gvmTXV0LbQG0df9LKqUE/h7HGbPzRzVyJdb2NLWCCfdPR6W5in4rTWIDhrVhVg
d4RT+KDzgm75sSlCb6I6klxZ85C0T+KkC5w8gdgsAskCuqVE1h8re16WxXLsTPRB
KqQCNAuVpGEHh22unHDTqovuUtFZ5z9Yb/vj89q92KzaJrh7pFxDdNP2q7jQ78rG
vQPsHl4SOmQntsx9+OwO9cNaLbwZeuvyDYOmRo4/3DlOvki6gXGjoU0Hu/Oes5gH
WJRt6joRcExPY1ImgUJl6AGXgx2ct8JGdVENjUeH8H1Id/7rGW6h7DXeFM9L1RVi
HRUmhVza+xne9CH0eKtbGjrw2P+cMAUQhhMCgB5yyoaKLOK6I6/cGP/LrvfeF1jD
Bq/u9BejLayb5xS65ht+fV03R/Cmdd4MtpnZgJPCMsBRJrGoItzEJTWGW/llHBUS
fqlOJUhM4fJLby8mwpfbYkRZ8F339lTRoIyyK4C0ekwMJDR1EJqJNRmV7i7dX5ze
modnpHxaNyKLpfweYjm5nA3vD/YJEWEr1lRKt4xWHJdPQFo4/XZnDW1A4H2o+ycr
eAckyEKeiRloE9rUOylUyd2nKQf6VBfuCHy0S2U1eadNaGjYTj2waUDWunOzPzd1
dcd8wXLUlsqGhAvs2ojVleitQVKHOoBB9kBt+5R/6oLUzVTfOW6OWaTx877GRvD7
HSRXs459qZVJd7D2I5JRakp1QUv6+BGpEbh3QKyPOESQNicEtvYUM0mjwN330WXJ
PGFLejSmf+XfgBZGwdbB7fxiXFb5K3VDp9L3iew9OpH90kcHH6KKU+s8IoaViU93
dvCe+W2OcxaIRGEtQAq0uyQLzcxjyf2DzW0M/G+LObDKDVBvfhKx84NsdDQCt9AL
9CxYRaa6humToC2oBp09tmcmAwXVfcs+DcWbsk2C8XlrT4Wat0T0DEXaHUQLr6My
118NwnNbgGzAN4ioVEbXL/gmEECwMwfVrlt7ibF7OZ/42+R0f6CPPjbkvR28eqUo
dfo3nqWGeSlz889s6rhYtZBYV8mKXcj36Efy5pdKSIzS/g+kuCQRdU11/rW8qDwG
lAcuFzxwoPu93kxA93TaaWdlaOcVL8As2eTvvB9a5bcL5nXnbuWz5jpXVeHlxwQ6
XrvDi6cRvjcTFIkOUD+nIEwGDEx2QBA8pjptfl9UWaA+1GwVdeQKwmYtNDAZxRdf
H4C2d42gHL4kHU4SsCxTpRxMXmE8HPwuPT7ppC0xLp9R+EsFS4bs9dxZ96KA0BXo
A6r48lR9bI8CrraQ0dOrtJzCCdru9z9tFoSH4GRtiiMHrZGqdzM2Gjh45p+ihc05
wEnbKVXb1O8o9Zr6B9ZCplDO7i4ETLbPaeetsxTycg11kVbcMge2zNGWfZwPIhpF
C27ZJkrXT8ASvrjrYXHvWyizG7Ul6wbzRlW2iJ0H8MduQeoUiklPPPf+dM5ZgWnY
zxLWAPy8o3kGHHa1gP9Zu+hlgKmjvUsbUU7P5q+zVqQhWhp4ddXS5lQyfvQC/G3b
coLlfAFzl+rXcaepwsZqET7DGXzR32AnMFER3jUX/Aw8+cdH3Sm1O984G016MlYc
folFdoKa/m5eUannsmH9dKtAPvnJDUOnIQcob9q7J5At7X/IY7DcRNVgbXcAaV4X
FINHfH9pep99SHI/PE1FpExgKM7pgM5TTuFEfOlOP9DzGDzp+rRt6lCU4GvDPRzs
jKdA1HNj0TfUApI5Im2AFj9IrZVI7qbYndjZGXueouJipRXdMtvMN9zXWgqqVUdg
XlTxkT7ZXt0kt1Jo2Qb5+icY+WVovk6QLTIrYUfxhZeLjgLaV3OQho0DNHvOK9GA
TiKCgh0btIj81VMNWXpSGW0ZgqvQiy65fp4Af2XTqLpdwGP+G2Z+m9dsAkZSsdkV
c/CCzMGLB60ItYAUzBrSVxkTxQC06BG7h0Kw1dn5Z+d6MmC1ZwdVsc8AZgfuoUw6
PIMD9/oUmGzGFrSQcaz296pik+51TxhiwdaCMPKo+tURK7K3e9KLhuGN6EtOTTIO
zj5GHLkA1+o2q5ZrCmN2/AloYPKFQH8ZCUpGs10JQKWWjGCORF3VGNgiAesgZVPb
PSQVy7IL7paPy0u+pkCVyWkdmHZ4/kwokqxTCXodCwHiTLwXj/2VUV3uk+Yudxq1
J41kJNsdZ9pzWIEzcfFVXOL/ErIjjeZOzJMRzPJZYgpAmzEgJgInudKoTeEIl6So
v5Xtupo9cBVkRoAl41aUTnER/6Vl6tv8ymc3nUGfB0Dnvf8SonWhi5NGpNJgrrCu
0yQmbAoE5faY9q8Jjn7w7NR8Duf9Cdb7/5Sadfgd4vZ8EYTuzfXPfDYSk1bS5j/e
CTdi27nlvamvvivhzAv18vRMZgxe+ufgpjCg1F1qOEQpQ1UFXo7kjZgKt1bhPSiW
ClJczVor0xcyNDbCMMGNB9LrnqjHDz1rbYBCBWy4Qt43+Sd6Qh0AMaLoCpXEGbCg
yu1uwSQLjsMs6gIh++1U75aqVI24SE6rVFb6/SdezM89sjNM4UcXC+SnCkESB6qA
RQbyhz3cjzKmOdMbis7dXH7GThCgJWC6YnZu3qxCq1rgua8BzWHEbwcbfoBH2NRF
XtuyqochG/poHmNx5csSaMYgH7/k2XWSDi9zvTA8PSuzzzKG9cfkt2O2FQ9AqZpl
i24kFoDul7YKiJyqNkF4r3/uK7aEVk2CFOeVeh0QmT86XVcnqnC5UHUtF/WtoRa5
cDBcrAOeRWVVvIDBJyT877FuSRncruNeoIUMh5HKGxGi7UUBsCmJGTT4ahWtjtu7
cOyJ70z4KDSHeuYMtUCGATKf8a79f+FYJRBqASbil+ZVtRq67rDF1LZW2IPndeBq
K+C1WS6ssvl8IANW8BTAvRqx/JVpJLGLMu+HcjPfLHIqsaP8CWiFSypPjkPmvhdt
6arTPL7H92wcpBy7aMwEMCu5YD5VFNrduSXy6LCn6NYhSZunhDTVvxS4YKuADega
UM8kwvJ21B2c8VQ2YChPMeFzm9WzUl916Up5aZd9VmR/fXEOQ4xHJk9JSySfWpAt
6j76CIJeThFr72VvtLIrftdzO/quClVBrnLH+YhzpxPh+Q/FpXH6B3yJp0NsmUjI
K3RZC8XEWOjwQ3+NqqiMkf9pkatmXltISj7rFS1XrPUXVEMjki0UWyVHTsmsvnsP
VTs4CrUrc84u6xo+f/BiIoKqqMbu1fFQ41VD4SE/s4NzQY9FVdrwo4M2lvx+iF1l
Izzvcdax3QLejqR79YZ391khJO7ZLJWueKE/QDlThDI/6iqbq6PHI9m06ujySfj3
YHfxqCy+ef9PZwSrDQX8fgtvRg26kC8rVTbgecKj5nOBaQT9QnvnBomE4SxNGrqh
QCjZINlv6fz3TgCvAJfWylrSAsmjh6YyHQfchMqyHgGssJG+a64K1Ez4dqlGGo+F
/Yfpy74I3T4TtU4AqQZcZcuDBytzKwDoug7zu/c6Kyt5hTl+cspCOds17VeXHLkI
aoIg3SvEtIeG2HgtYpD1ydsHhj0UVG/hxHLjYlAAqNf8o4A5gh/h5h3GVF4RtMl6
TM0whQuQiZ+zYG6Cr13GmtRTbVFy0J6HFUcZW06AikkNnELei781AB9mP6N4VXfZ
viCAzRTphVbhiSipzPuO+MDhS6SHdx0BswH+bXJxdjnAkkp6qbMSlMiPb07wim//
25ZJQ9ilFRf0YveeDdFXDGQx1QLF8WzMeEYnHaVQuwt/qAAzwaQOdzCM9jaHrlYu
Ov+fb/SohRFJQTl6gbOCD2nc1ZnWvVPaGEpHDvXkGnkqzvWk/f3cDFWq2XRZmq9T
9xmjsnl8hr8XymAxcJIyPCxw2eauBOWihRLvVLkJLzj03BPZeYYlWDRl5BaKmr5G
ZCEtM7VJ3W3wNJO8tVLMaChZCJEtUxlLPUVFkTNwovjF6rI2zvaLwYQRubBPPa2r
oYK9Ny0Sb/XHAg090uU8OdM0FxsZSzspVkE3wxT8MbMzRMtRwJVuJDHSJN/9sgUz
jJmp2NK3tb85NnsfHHN7UvvjRUZ6KeEUminEHDeQQrFj7zyShYMyuYy1fb1RqaFl
A1uZL3L3pPvAF6FnXkOB7xAykiqD7mEXOPPS9ev1iclZgGoNwfdyKmSd0T4exhYq
At7y0rRkf/pvpam4rCL8y/NXGkSj/WZjfejMpqwFsXut6e+9wY2rUlHibqR9vLah
0WCtgOLg/l/Mz1QyaeCKJ5HTgnMAKMVAVS0s3ett0EmxXf6KE66HJVvuFu6c0hhc
yOQUz5PzHeOj7Joy4w6+KcdFwlU1S6Bjm70dyfTboaKxaoQ3J2cxTZeFhXhiXBLp
Xok0U+4iV08nDm+Kj1d4UD1xEh6Uee77dFTEkMlXXFf93gKupMtrb2kmOxrpx6hm
H6CQMm9Ra66RZgUN7G8k+spWkUEV+3HIb+fzzqZpLZER24HOD/0SyDpNw9A8tjcx
y6pw56YoegX2xUxUZU0YWLSBcFOwsnDzzMR7f1Aim9Epbx0uwZh3p0gncfFKvgzx
fMBz9yd74oX8jnxBssnj16HQG3qlYsYEpDt3SzJK6PM+bYEBziezE/0IbN9g9Qvo
5ld1ZkKg4JoXbdNrqVXKtvhGc8lRbPLYVmgm5P6OdgpRUS8MWn0PwqeaLTkqFlW5
Gb9DvvfBtPpaOOySUW9OTkN0zC/Mx067xuEAP48qiACchy9ZZtxoBNssb/2MxFS1
zHw+qOg9TtJ7ZsYknHxi23HCCqAvz5cFXs44pz76EJRd1q4fu0AzVVyhjW8aQxXR
3ySmeKXJHkRWteQ6FgwvUzUMKPlYwkxoiLt5H2UduLzlZIn+YZmxkZmbPurTeyCW
ryYxxpVbaWjGl1S+PacqADZZij3SNOd4mSbvKpMHIPeY32SRr9WjuWOslxYLQpaC
6Pfa9Wvh5VR6mGBQvvMosJyK/+boOUB40G8elEu4AWz2yim2sr/0xnznEXEauu32
fQiZXODzzVN9zvB4F+78JDLXNDej7hK9obuyz369QjJ8YGXCyWB3fA1BdwAjmyou
eJ2yflKj/6PC8oT9iEqq/54VCQsHZd/E2T4NHo94LXGERqXzZl1F0rTY+Hr9B9AI
w4IqqQ/IroDC6CZMPEDpXZZTK66ASFhulDXyqEc2J5JnzMyAxpvBZPA4K3lSE1EL
juooC9gJAA6WANJSCzY1p5sTeUyJRQR+l/GC8FDiqy6FHAKyl9w2C0MGwn0w+4BT
SY/7OpMbmiT8ROqk8Uqam9rP8WE7Tof7ewb8mc9D5/H+rUBCj4IzHN3hsdnx6ovH
fCKUm3o7VBcMtHXs5rwsoA1NrPAgkTVqHUdi8Z3IjsFBxIO//BPekexJqLSnVcf8
u4cn0mr7/WViWajKEGEWZRnRVf/OJVGa6f696oN/GatzbVSrOV33ponxhpsLfURH
io09nC55fWbpPexNJQWBsTX8rXe23lidCInjayrdpluFRARRkhpF5HQJIBOz0y+l
17UHRCA3W0KSgyK3AMTCpcAdNmW5WhGxXFGiwK2KZZXyNxAmffNeH0hj4NTLPbGa
iGPxbPWqVuRBoqB9eaYiYhdT0V3I1vQmj5WbY9JLn80c/piDtpdGeGe89RusW0mg
JRs08V3JMzVYqwMddPgZlOVFBemk+T8/tffiyFhbTqVjIBxfkhcHjb1+AzC7bJn1
eSeEZVZi9x6qsE8fBMuIKku+D1YKPDVJnGmLFqrvNLZCvceudO8e3t0Djb96621A
LFAq3YWq9O2TfwNt56lVjB0kUzFRphVrRJDcYq9GclDPWZQcMOJ9B1zQTrbsBV0v
9sIh311X0diBVhMYJKwWGYmNZIKsMOfpoBAOlO8G2pY0/wlq3v5AZ/qn6v4LZCnO
xFBXYnBaSxuhkY3ey+waNcu2OCPsocvh81nzyLsY0nNien8cBUlSic4Qxq2NX+Xb
SD+AhDcLxWnWxkJQbIO02+4FvTdRRq/9u8EEN2zUXfCNRazKViSdv/PcxICnOLSL
O0t/mh5cJk3zDz0NIgWPLJbboDpGJCiLR1aWwLRnjMSqNpvXbP7CuQgqsqCkeyoJ
8PYRtuIA3nQWGrJKAnhzA8g4wQu7vm1yDcvOxqLUCdSeldfrR6SbqTxO0N7BgV1C
3BYaV5T1/e0xJ8BPvOfqdvkbYd1+tKSv9bOSydHlWeDSHI+s6JDwK5kNGkfBKoFd
NM6koF5vlQ5Xi9vBq7Yir+2r+qoAy3FWC6z0bUHusO+aXHOb2P4fK3nwOmJzvY3q
ol9cNkQu8vZRZxC99mmSoxhjtleC1ZaLQ+eh694UlGnccsyPzb6Rv6KnslAd6ASP
mlsKuJUEvaEPUae0CMuF2/eDvr/MSK8xl7EiKdc70dgHhQDlYrJRwLEZjz2Ttit4
WyeM8fMzydB0DVuVqD3wq6GFCsdG630z34HAuZkHnmSkBReUOMhbKyzFtYzl+gLb
Z8g94dqUzSn3jzAuZWluVWYIrcVaZlgSlNnwXKF7wDjtW1FyM5MmJ9ltdwJWrxC+
Ff9O4dxUr9fb1RkPybeUmNvTBlsoQG44ENetC1QqgiYxWnUJCijdDZy7a45wX3PH
giJEK4g7IBqnqR2whwqc4FpTS330z7DPVvNwUDRFCsb3VViMfVjiA1VGU9+/Nyix
LeOj/ShXt+/evto75+cRTf3vvDP8OifPs2Ti08bX9HgOBWWSEQEbq9MHjs6e7z0E
13RXw3cazPTPW3mMbYwKC5JFTgR3Ae9zEiMIWZoXshiZIJjksCn3kyrEMCuJFLyl
jRGNCpHEc9sK6qH9Yh8xTFJgDxNC0sw3LhSEAR9z+3Y5V+Zk902juV77AF8qq+75
Ci0+aLSgyEwz8PP8ISx/ac6VhDLkkO+Bq7+nDoB7cBFP33KTk+mtP8h9Cbhg0U1v
OPD/+Ngnkoz6MeQZfrf0pu98abOBwCKnpf4LAcYm2o46gxU8I8EsVctlv6w8kLkM
zhtknyxAHhzYr6BGjTalulbn0QaEd6ghkc0Eby2I/wgDj6Y4Qr1C8m/DlE6+aZMJ
EHK0HPqtAYuicKlXhfS0pMk1EgzC6xp1KRyUXYrh6Ud+9DvAtLIvik0cNbsr4fsF
ml4LbQycBwAHWAGNtxb9Nt7N8LCLy8jAxDYqgR9o0ZbWYgP/AWHbCHgMmyYOthmZ
qGVN8mMmRYEEsH4rR7pqfsoEpXpDVL9jQpHdPhFUOS7mufGbCdUt0HXk1qe9dfsj
0kzlcWWBo+KQBp29tzQ9evXQHe+GT5nZ2kZNIoAjLux84D58+yd0Hr4hfwMAoD1y
bJmz1bzJk16gPJpxFJ6VYvspBKYOcLLj65aZYqCCWMTvbScdq0lBmUSwsp/XeqjU
ygfXe4LsrM9CvNeK4cce1kFqInQXDTOoYlj3DtTY3uIKWeVZrGAFfDUzNp3stVt4
Mcp8yqegzAaJip3QkN8Ht3770i9NBYkLCt6mxYrioujvHvOXFaebZL+YgjnEQGQz
4vgIpJ1dmFtvgtwu2KPrSYPaoTKDXMrH+cfATUmr4xzbi6cTDa+tbbm263e2THXm
YMV2ae1Mr380f4CLlljh2g==
--pragma protect end_data_block
--pragma protect digest_block
k+b0p8dHP4nlby+TFvQD32ZieE0=
--pragma protect end_digest_block
--pragma protect end_protected
