-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
PnWjQjIHu1Xz/2Tz2SxEr7NthySEEpqu1Wo+/ECsOtSFVWRDWGRjJGHpvacYfmPy
OHau9qi2i3wTRbqD3Pt5Nu7UnxGI1uuCZihuI4iMJgkHkKOBUOscc+5+whYfTmyI
9Mre7t+TMPsKrt6f+jc2v1Psw8NwHnT+4qjseJ1bCeE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4520)

`protect DATA_BLOCK
HUjT1AYUgMPVoEQx2lkSq0vy41haDDTHTgyxHioVf8meVjWp0qD2ZMPupK0Ks/Nm
pi9zaHlVSu6vNsMXoEU2A2C+tOwLzEOcyXsF633gOOA1mhUtd1+P//pxxSrTpRTt
Cs2e2godJmpzRtI7oe7EDptWpT92pJo3DMZVR1xnQY15b6sCIzCY9mh5b45zbW3g
X/sIQPDdkS3hNCTHOfNLxHH3Y+P4LT2tT7fK7lqxXd1Er823wncDSXaei0RDqKcy
7e/DPoCCpkptCctGlR67MzhxYO7OSWLP3SJaeyiqHYYP59sz5fnQD/OCayuBmw7w
3sqIWeTrhgItL7+RYlkpTsJPmABO+40ZBG5QpnJv+LwFP9bcY135nzYtyHKiwFyW
3HqJqdLUJv7Q6bidZtRYd4/ULBAq4Hin6G5WQFf0MZXz+FgkKcisp8/w0V5FP3PM
+3DyvCwd6qWjmKQCIuiGLNk1vw7L0wij0eBcXTBjJ1ovV9fdcd9u40qnOVEeawP/
Bv95GkHZA4D8Nyo9n7mNsGRnDWjBurSNJxKM26HDZG5qQAfKZfOGK9WTeAPTregD
DFJFOaVLPuFr/fmdaOKZK6Ga3gi2RPM/hr5jgPT3oVo61GyVnLQ3fjTugau9mMm6
35aF21/uBCVPbYRw2rN2hbwurEuGGTR6/KRRFDnQLH/xfUWd3JbnCubxDse+1nP+
L6CZme5HZAaimKePIMyYr6FvQPs/ALfD3M5jwr43AfH9rjvkkuPK3LskRRfJEOkX
NO2cvlp6STe8+Hvt7yQ0//Q4kL0k6i6iVZDC9P8kAj+tMjINcVXdE0fg1a1s1YNd
Hb19eq8DA2m7WiOfEO8aM95HGAawnmo3DYO9ZY2Ne56XMfW/X1clEm9QOj8mCtD6
oJj8Mxo7JCeP2hCPatOnJjlxUU1rj4jHHLe7LhVZfJ7zoMVETHlIKNSXaNrs4ZpD
jcN0gfnFTqz+6nKYdjCj65zRXRR56cE/p7W7OYUpOhePSLPfZbq3AIV1bT5QiVap
6dTU0miZdla5TMXMgaqSf5HpLvok1NcSQKaxCA+2kLTNVDZ0IaRetaaFAoWKmclh
qC5jHkqAlzF2sTYId5slkyte00GuWyNG06s/1u0+SDknogatIOW52OWSVpG7uvhD
90nJjvmUp8YCZ2vmCar5C8ukX7Fv1k5DX540eyhBaH7QNc1hVUgf3vGGPBgsBo8U
RA9rV3Uih9p3BuykE6+t32QyjAS4y//dp1XWdzZ0zr3G+s6mKscdVMFnzhMhLweW
hBIflz6T1pXazXda3mfZ/GFFuR34VwdxG2W6vKNfV27z4eVSfkEEHsx89t25TgcE
csvPB8ZZr4ae971pJ8jvMhdEhldZ2eDCz0msLSZrw/mNUJoDFRHT1CyfT6c8QykG
zHOuLBT0Tv9+o7ltmdZPtEqy9cEHgoIMst9lrPDkF3LHmLf913GgwFIiX1WarD02
wzsOpA3vafzuHaA6CIlMIv8ncNYlaV7xo1BzNImLtfvnatrRVZuCLHDB7TX8ZS+C
n0KmWBt/4aKuhFRgQPaxMtwu/Mht7RlF9y63W8UxiyHjG5KIk5+fgD7qtm6cbgUN
hSHfVH7UihHT3YtakCbBt62YxLIUxqywXyZuUECKNSNSGK+R4qnTOuzp3KAxEW5z
j7IuI2LxP6aCuTqx2bzV8XOuD/Y2ZwX6JS8K8jL7cSGZYy2WG/g0DYS8JQyOnovd
NRRQSs8K3QtiTyvgH06azpESzs4PPEC06V6O0MpV2piiRWf/z/fehw+wUZjRlXEC
MlLX0h2TZmTXp2N8N4fudm07IBuyyQN7fvXqEw8VgrgzZmkA0RLi7T2Nwk97cNbZ
ICcdQXGbKq4Homxghf4ZTJrRcFyOMgy9TB/vt1k5aSG+H0fFMCFyJ087pV8EIRvK
/W3LkavonBXesjbxSdr3iY9mATULxFxFRPMMNdd/zTIYsw3njiTDZarWUH6oaRV1
foS/IwSABEUi+72uts7eMMVXXqD/kBm4AZozOf2ua4ZCQS84N0qpLf20stoVtDjA
xSaBlzGQXko65EJ4hJqQgnZejKy0I66waAiaK/y0IoqzqEXio9kawXtvHkTAN1Zd
dfB9mKT2WCUs06eUG7pGH83N/docfKFHWsEI3UY7YcnGxvNsZxGPOi4TGEyYSeE4
slez9F/Qe5JHK33Q+TDCrpkNfLGXVhesorkbLxuRzAUvm8E84cnwQAfGMEULWgrN
hQCpSmzjc5x06Dx9NVgmc+UJTiiPeUJTFUhzUItKO8uOjDsVOkXjsAZB5phOnCSF
0EBkGDR7CMcBKom5LD3Sh0gIW6CvTpQpb6Rpypxn5g1qu0MvWxPmkv102EWsLWtb
A1CqeaIRbL7mJLc5VABRigwz7mRVVwhb07ZFxMc/HiYQ5Gq7hN1M7xf799NnAfS0
oA9zjNBgyyfgWBDsatvRm+nlTtL/EWL7/6WauDRH2jEg2quXNowyxGz5C37S/Yw9
qbUCw12Za9/7Mf2IVy6cHNKrTRCL0khe87/8sxUeVDFV1q2UnbDJmUSUWg0VhEoK
9fkcZyUlkdSKNPMyuVPnHTI1G5p+8ieO7KSRZntxh8W8XT1AMQGgdsouzKpUxUM5
ZLPlAgLRScXfKvDCH8hTizJ3/hp8Nm9NEJwc5V4uFUC+SbSg0GVkJtBnWYArib4d
CI9IdUkie3IrjQU8KZfeTMgVzZzGRLJe1DRd9rE8fPpvHlZf15hGHk8vsZjCewYG
VUYoPIL808fjPkgGoNqDwv7jJx5Aq43Dq8OraXJH6lQcn3gJBgKWCxIx2Ztcn0uM
phm2RMOUG1Ns14S+zuh+BJ9vwgCg3S0bBhxTW2r1cF7+RWvh3V1Zl9flJntz03IW
s1ALYKA8F39VDmA1Qd+0eTwX1sV8w7AdN7sDYaaLPCBuq9CfhiD9PlS90YLtLFHq
lHPq3xC+6eGhXC4sYbxq2g6/LgVpK0oUR0g75htk5FLGHcxFl/aAsrN2PvWu28fm
G8STaRE83C5E1XgZY1ROTo5OzdfiYqgAcBuPvzK4G3U0jGgP0+RhbmirL2Oncej8
T5QoKJy8TF0rMnsjHOiW+4z7NaZkXBw3fUHetCe7DFJkUnme1bmFGz9Yk3GQ3M5u
hImU1LcFNvjsfRWew63CisBYE8tNyxzsJqF5RFyo2BOh2iKk3llUvUWlgZLsmwU4
CiNRB+AvsMZEICSFoIKXlxtWIM7z190DvCIG/KG8skRelYSf0dzroHCRxuwjhoR7
dDTsDT84aagE9Haf7odg6G9n829CPIf461BvXaaTEFNGgSh0rf1MyFJDQ48QBc3r
4UGzt7H70KsUNXhqBOSpYbq9C1CDG+ptunCnoOCdDkvzaIa0Orj3SMbNheUE+Jji
rBETPJpEhT5k+Min6HwyMuJMR07kAd/PNPCzfqQQimVAaYkTHTLqPCve6uDvyNbX
lokIIaVo2TAbTUr3Zwn369rTYYSvHziEPWxbGiirkjujbYzhVDg5wJe1xe9L7vaj
V3Av9FL8DLw6OXzygefn+lG7JbRzlJ3rckNTOv/k+0d5HT+RJaueTWVIxgnR2CEr
CHPR7ZEPWREpBMsYo7ZBk7OiEN4j259hasR3xmSjP+A4O0dOhfMl1XrS+z2dPDIm
Dby5sfGoMkXYm6NfbmnpKBWKbGY8mJC9MxmdeXNtY6SxBuWLl97GGvE4Q9RdoVLa
/FTGwxLSdXH8Ng7K2Y6JTFkdWF/IeGHY5Z2955fVXC5nwF7w65wuAKkFw3hdfwGV
rkpp1qoDj+H8pMknYnvi1ejn4h8QuYSs/MVLdUgY71/fTVv20zPY4Umnzs1XlFGA
B9hPQQZFQppZOtE8TSwRfxZeJLOwun/afGVNM6yq/fpyi0+uA69KnrJHIfvELORA
DWkiEDbK9W624sMOPF38FuKA0PIkUbEWTFuJNgDr1+e31GmqNKoouPnqPpNiooYp
TID3AJg3aAs9dZubNU7I6gRP11YI5MNZLUW136T7zdHQWSz6lhsVVMRUbx1TZsvc
3q42wUnmUSDw478YnkFxA+gERwcOMyjS4pS/X8suPHvWiU96ElbYzDwOvQ6mfDgg
DZS8f1Hj+dNAOZBWWPA94xUm4MGr7p5ZzzdvVRp5guIdHuNCci591jvb3KUQlaBB
fnbhhEQncePdKlI72Ou4GsoxnEK+ii9GhgotbNnafI5o+wuFFtV/oylRJbnKyEL/
FHAy3CJJdJ3vf3Jhd7rp2OGLrczEPw2eIE/owHperUMnw5UXLR259RzlsU6tBYv6
gNah1IsofCJqRGk4ZnG+Q8jzRo1DI7qFHA0Vizg0ChJNhRDSfvYYTt6n066q+Hxc
WN6KsB3OLF04ef92sDWTc39GWifP2dUkFScfJzIPv0plMxYuqShhrY4RbGhG41X+
4IuQOVhMp8n/0MzdeGqx2HvDj4bzqCGMf5ILG94aA5Qf0vmGCAHKEdBynUY+l8t5
6y+a0jaIko0s42aj3Qq+B9f0ueLVtnkr7JbIDH9M1OBSXgmxCayC2Mpn7AOWQaW8
bYjBfTmje6LBosgX02EhkywusTvGMEg+OVKs6aUlTtWEYJN3Ac3dSxgyKmqIsDoK
uLZcUInan1kbWswGg94eL/LadSVZXcbE3Ajzri2HJ2KcXT1DPwkrRkhIvaQkL/e0
lrGtZlZD5g3FdHEbYL7eVs1t2b29pVVcvxy/ZNaZH2G25Y4HZ1Tz/F7j4gTGp3mA
mWfr074yZG7+BmHhfMhC0JvBl0qs79EwkFxvXremSNXtaH/JvLr/ottIU9li3fif
LYPDKGs33qtqbucLGtXPa/QLvBfxIKP0O+VQOR97BYvqNJe+WMYvaRJBakjD14Go
oku2JltDVZwl94oQSMubJrGdUV7aMsVmuHXIkdjZ9Bcmi4Yi4OMKJSiVqyu6U+Ec
/FjNI1fmTJrpukJLtHMCUlcXALn65b72QdxKJu4GFwIb6YJuQRqK4QwUcd0kivoc
yYPON9MGOQgs8q6HRyydWkC5oBD17pjkL8AsV0UzMaYua1uyVp1ptmJmgK5lE14Z
kT6lKv+CXsvQFWUBH0Xn+R90oSQZWEBEUCUvVpHZhSkaSRrNLkKlSPXlOk6NPms6
u9FcLGQ2nsw7FwxtUyIiLKUp46DQ/93MVX8YrH2VsrshiVn/DVMngC37ZWapTwjR
dyk+uz9wRXyu8GaPpnan0Krd8bOJn9r5VrIwnf//5GIQ+p/eOBkbyCtNQp5jp1Uq
qWo/jz+BhHoDO73uaHFY5d6u0VWmcZY+mhqiuUI/PnA/li+Zwt9Rfwj0AbpXYsJU
HQ3ihci5oBuLDrZwNy7eqfglJvxXCRXHc5rzqEmBh1m5Ha+Dz6CBKWvqcRVZkTdj
HBBHw/Mj2KG7jaO5jq/yuO3s1U5+4tdIO8qjWsuVB9zJAFmHRwTDTbCLW8yMBEKW
CgWNJwFG9ChyhbAorzVzBugAo9A24NPRke987iDvqGVqMq15jxnegxEquv8XiCeU
H4Ofm+JCPH2YRViD1PYInY1siPb3o3Gl30JvzJY6LodG/Hmao1NssWulvX+UpWZN
ejhI4mEmij9uBDr4tDiphoYvApxQJN4dJpnCIm9iRtPnZ4C1RzcmVQwRQCLhNzlW
wGD6vHOAB8OnkwSWTMIACmz+4p1Yq5HJ5r2C7bZpvlyvdumd+/UsnQvXnht9Uxto
lllRKe8svxKajRiHJewDTjQo+UgvIVHRzePmaWhC3OQNH2aDwoDh0+XPxYVMicqn
4vBu9xmi4j7KiFJ0lOL2P5oSXuMiN45oeSDqh2ktsXkXrWRvnlmkbMeE/jYg4ItL
ILVOSJ3zM7LAN/XB6u/kNlmCEQmalNgWHIeX9ttRXSp64uGj3sZhO/ohfSUK7doe
Npn63zf0Y5LIrDt1v79aKa7YE2E5jBjHjHrIadu9Zc0fHKHzHLBB4tDbvnyARln5
YhWTI2Uyd7PdYp5ZZCPZAFeqUQ5YQwcD2Z/Ic2wI37+oFpI/oV9PW95EimUDLpJ3
xfePe7EoV6gN61mZuZaxUZ4512U6bP5hWDXLNWt7n4w=
`protect END_PROTECTED