-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QVfK5fFq8aF74IGlkXh1g/emR7gOj9L0/wPR8rA96WQUbBh6TdE88ihvXM6a4nEq
/EH0eg/B8dEsWcWbGd+8pE/QI/sF48my1uIoIbbdag1u/tDfPAAUOHABC570b6f7
k4xHQBTwX3Za70Ymi4K5+z36e+GxF2sB9Y1m63tkeaM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 20766)

`protect DATA_BLOCK
kiRB8f687hGbcT0RqJZpD36zDGEEGad26XxPa1Kxi7/gWkygXZoVVopWVc8RMrIf
NMcN/eKBgXZbmh2hyt+JPj4RMDCj8aaGupIX0gR0k3paOOfx3usW66MvBnYR0K/7
8ORSpOckjNk1WgXg2plN8+eP8GlOQz/lNgAmSh2Q67s8fQTtMX7gmJv/4GGoYRFh
hAeZNb12MVn2R3mnwHvxGf/L08DmC/mE+/8jsR5RMNX06N8NaARKfmj8K/q1zdU/
/8h6oGovWvVu7uJ6ueAXRlD+1e5H9/dF7WzCNCNCrga2U6gLjAb9UGjL1dE0gmKN
dw79vlA8HL+cXpcIHfGXZekzjYJ4hueVTo7oCoLYRWyjes5r9LAFqSrgPMuIYQy9
0CGrAb0jzDICPxzVJlfdZAt/pmeevgTTc7po5iK9WxX5MRLgtCJvNfHwpfGC1FDx
tfZTrOpzwgcuLoI09JNbxOQmyC8IruF0+tGioFzMCZ1XCCrGp/fiHs/Apwr8Fu/t
o2mxx5AWYy5MgaWkGkDFd3BkLsVmsJeGRaOeJotALZ40sxjucIhWIpc+5xfCy6lo
CyyajvktqfeLY+XRyXBWMqeTa2WGwovG0UFTGFkp6qFc1My2+9l+Dhrratf3TZwL
QLGEMdFAWhlsx56v9WRb0MTH/B97BeUi0lhde/zV+5UGaq9mcH/NlXPsPwBUO69P
DlaUA76rM5fKTIkHqLhAxam5hkrO4P5vCK6V9uvAodVx7g7qoJ6LUakTlt4mqgkD
l0XhYesvtGVd1C45q2Z7VRZ0qQuhsIpqy0magzo70Xv8044ooQEsYNz10Tk7srsu
S2q8daB31xJaw0GewYhI6i4miJxDGQoz56V0pTIAcLQ9iujPh33/efF7q7hcF3v6
nysO/1hYHiB/gLatcVAihc6AJLm/BMRKlyxevhI/eVg3vrokCcvqtsaFAXUhvbbk
7ZtJRfYbnbv0Gzn8lbARbNVFC43dyLxToYaQhxIZqCjeekwyBGU8oRmRYxYqbZkT
xIdApmCeX4IOO/x+vEbzrMT/0/2uYpkX67zcNQrHEqzZEhoHFWa9zvTVMvc1bwav
R3QZ6MS1loRM0kh4vm0UD0AfiFczDIqcB/hzyPs9TY6zsD0na/nr9tODYDi79Zuf
rkH1LuoBYrpv+69qE06lEqI+gf7eU4yJOYvCuagMO5Ych8HW/XcQrDxHnkJCnWg9
9EzrHUNogCcmmKGrQ3sZw+kk3j6uIrR16x5x08P9C4xdpi1ixktnN6Q7/rbuQZds
0h1nTbsNm0D0No6tAUFiR8fiGL5RKDpVPrSF+dYhq/Jcc2D2nyOEc0r683Fyn8dH
fQmyxtZutDz3aoMYxxxPPqr/5wQt0GUTdi8XqJahmtCJSyBkkqWAa0YnfYAD7JZ7
FzCEkXV32r/9mr/CoaZU+XJtwvLlkk1o4G/dcqwSb8VoTwsRrkWtI8v4ZIl2l+6V
HecvRMHhvf/7fD92a3TVHoYGI8C4PmDMg4IYYyj+H1BFgn0R+dpTlhhVaxJTCnTc
4pTeC96nRhL4OxW1w1QtR2HvIhUHI5pP6FMsNPfHKXEtWpqO86pKRKpTcjYB0Gqo
ENHJZYOjlE86QBfun+pyvpG7+3ZJ5OW9GwBD9ySSuRRcgChSSlXZIJcbAMLc1gK8
eIlWXEkn9ZfDexSja+HgKNGuxPtoB+lMa3+AIUC4j83lp6Abm1dCmtedz5Cq52Sl
Q3EKn2wlxz66zrAD4t2zliF/Ivf2nnnVxcKVvvODrBOFDLlaS4mNOEetnJDakkm6
EPeagn7e+TuCcZkbnqavS3Sft9yXdsaCWOdB75oEXBHv228AZ05n3SPlXD7MPofH
kmplsjV2gYDiliRQOj1/tJsdg2ooTtFcZ0G71ufrpsBK3PXajxR9VYliydWwCuJl
sbyE/j20igFIZssIYxHGhrUQQgcBZ2lXKKiXVPsgVm8nnKS1oTqzlYaIDikBBA/d
hIEJYFv7W9jFmvEYC0E3RjQArWPSkgjEH3uA2fFYS9eVc/AhjXDlTEX2CxHh6n10
Ymak33qV3PH81tytxuL/49pEgKqJzojonXVKd6MebIksBpI356dg+r2gN6onu43d
RNkn0CafGWRm3aGHN3JQWijptakk9En7DxuNRcmk/D3wGtHY1b8uiKg13hh4WHRk
28qedn+eOIb4XyK846O8K/8SxBRgtQw28o2HJLX9JTyMflNy9d2FDxJHuq8bnMbL
nin6rJSQYtSlthZH7nD3g6goTgopX2TaBFJj9I3XI1af/YrehjmkGXal/Ybgzjk5
EZu3iEBXbo7u3LnOdOMFJ/vcs8ggqnAEOdQ66KCrZ3cNZ1rmd/BRRqzTIhiBAlrR
nwZKhfzMkoYsEBzcf4S1fMulwl/acJw3uHwbKVkR8b9dg+pbtjChImiQ/GyAedzt
1ek64C4y/Dq1vKO4cfzZn2ZrSu5usJi2tbImonC8eLECq4cHi3LkWkrtLJAal2z1
aFZQ2XK0baLngVXrSXSIiTTvK/U1IDoPcJ8bZwROh8/iyRLLPsMWF1qKpdxtp8ry
mTFcVddIfj+miVD8GvsSZYDxxvPr0QeUfoVhXaPLSnnTXgWVvkt+1raJ3jDBs4YY
fyPqytol1Zg80PyqEVVBXW1GW9ylLhdJR+KGP/GTwvMOYlQzcKmwO+oH12fzKdmC
IHWpiyr/Iae7zzDUJQimX3gUgqy5Y2EoOswRaQLUDLsC0Dwq281SZrC/YLzqE9JI
QrlVFCCmfrWLrhg0l9uTjnQeVhoxJRnelKyQxbWfmpwLZxO+HHteGx9n5WexDAuI
S6sj/5iAut/QBtwFMeuvq3P8RQIL7JRZfd35OhGUVDz9ro0bKPf62TtimCTVq6qG
+wocjRfW5sCSMpTkgq/kBYLUTiJ5SXRgOqRiFGjjV7rmOF1BJMJ6TTNj8+/C9/9c
hFwkqjnM/+6Jo+uzYUUUp+T9w/+WSvj0YFx6iSGfD8YGgjpP6NmSqKXwh0jTDtN+
zU0faiGuJfAeApW8OmFSBkgsyh5OdWzMGEIYE0sUMKLpI7CMNMdzWWLo71wnq9cY
7P5kT0yLJhrbqc8zKCYdJAZLlrdfxuLMcSArRNXxYentrHLF4SHDYxDwkz872uON
Dp9Wm47uhuWNeazlg6dR3GLorn1trVtMbV7dB8C1bHWAgeVKUtSJhHyoGisHkVjO
NBkSiDeqtxZtLGa5ellF1CMMv/aWP4YJB+Nok2d1DlOV2hDVKwoT9W710B67WuzJ
iRuWlZQoZAY9vkIZyEc7R5+xQEjHE5TmFzibhMGKZwPxStulnJ6yLqxCVdWNcR2q
PB0i48D2aLDCLyqdfjtjSuCiwxWWHunZZFGFq/yJILKKdwfi7tGzk180Nc8D2Ni2
+csW8F1+c7nfZmarulcxKfNOxIcISckxHAIYv7JGg4f+lmG9wObdtNKX/39Ior0V
OAqQlt0PMbgGwzAqdZisRMCPqBmWyL5tty4ISj2fdd8u9Wyb79q3d7ViACUXwxmD
njxVglluDBeyFlSWO5TktJwTdiovqikvhp1H7tqNFD8fBBu9zD7N331Bp0lCQDno
mH3DVooY0uLW4EB8+07Cs1A9+JXf4rq+2/YLhmDo+eb3QnOjyOfi8Onata567Sfv
IjKMXNN0OHrwnjYCMhzhnO5UwSWR9E8OVAi+k9HLYYs31IknXTP6IeM2e+7rtwJt
t04pYrQZ+0XTa4u9CCj1MYeZbqlq/4froehSuzReae3cYgMM/yHT8nrd12FiG804
4s4NOEnMldali2/dVEXOggPLYFDeJtubXNSfds7Mad5iTZlo1an/o9uokl8FSDKp
XOgLxI5W6p1nM88uE6KRVYzYF9gv2tr7G8w+ZVlmrPf33btprhVZ6A5QJnz2km6p
8h7xQPOA3Y8HiiAFEafZeeGSU0e5etv5gWQOevRTizdqSMIGB7yO0RNg6cYKgVvX
84pa9hWWQsskJ70cx1ifKYJ1mBpJbhbEbF2WDerrHFhHFA10sDhJnzXVOUMpXC3S
2n0duR5ZSnWRfiggAMVXIzRKUS/tTAIo+4TVZJii0K0f0nXJDgM5DNL4GIDmdUYM
YlPd0HZ14MWBFauHeeoAYw8z3gvwTx4oTM9SuPTQGBWXrt11GEFy0mvuE81Lil80
Gts8Mhqov8RRsEnYNH66Dmpd9d/R3KC1QOE7jsulmgd4ya7v0Ixob5MTZ3+UjS5W
wpytLhzTOlmtE0iALY+DhD7VmUTItPCQ0ghdzV3VYrPUoTD4djdBFnmS9WVQwfpI
u31CU+Sivr20ahvScBFq9mIi7SM7gQ3uptluw24aky8oKeCOykISIhTa4NfVHz+B
IcAV/7KtnXlsE5wqC7oWEIxV9PHZFH9mUklfWPK6iMoDS+Fe2yUQtmMU3vVfLAfx
KVgW/z5QQBLE8BQBdjCDkxpwLN1yIh7VEoVALRrPuAUoKZnxD0TOnmOtHQJIRlBN
2qvmxUDP/9bxI+cRBXTZz1HrANTjpCv1xJD8jyHl0MMupddKhOgm30cTSKdzBjZz
3sJLexyAnQUjoewpdnjhVRaa2/O/0pJR3svETtPZ5Yy80AmF5Mvhdl64jTIwCfUK
W4SrjDJ7YOGsijSiiKWPJWfcu/bYDAKhjwU+71fa4IG54jbLM3sPCKfW5GzEn/PL
2Z7/ibWq1E9dmQuT30yKS6JlTWpLkW/v5L7GJ96ex8j8uziImXmqqbP+NJGu3U1Q
lz5mu46MOet3ekyxiHF3KTStCGHj3uXs6x/UoBXraFEk/jGxm/8e4cBnivdLwz/a
km/6WIwTbG6nz6nMEYhX9YWOyF8GMrD+Of7IDy3stHvrgq642/INs8znZLg0Fv4Q
ZXr23dJNxfXyYsJ/KM3T8KXNTIiPjkJUr9+Xbbl6a41AcrzapPROYQC73bXfrxKN
syHCI1QKEIi/74WFas0ReM7LFD/l4Zq9I/X0vg+FQKrhxRn7BQ2io5n3lUw9P2wH
F6H0GiMAoVvYXeO5GTbXsMFIMyurhRtd7ofjoQXv2xmbaFu0YR4UVtC9i92orGSf
erfw7BFDOpGiaNH6rzP81nWzLuwftNCSgRlF2j/OzEN+ndhmMp5Bvp9g2z0aAIdy
cLmlEhpIDaBy12rGkZQBhdjfs7FI14afxv9xMvemgPK2g1eg3LSdGyLqhTFDQLdJ
JI810GzsCVe92xAf7ayyAqIrsRGsNVmEk8L3tN9wx0wHsDdjZlG5IuwAge/weCE1
INlK3/CYcWyBDc2kngtWl7cmjpZxP3fypAY5tx6Gx1Yfufzd76kuNqqa95+FVuTC
7fF/Svxc4Kabx7/k8u9865QGX5ONsboFkSzJbBiaQ1QgwE4wKu5evJF7zPZdGtJR
z+bhji1j84mtn12DSDbZ80WmPBRWi581hoaLbq7hvq85KwAIvaxnPwtOzOVr8rK4
eGNEJNOwHtzgeU46KtHQvMv3RCKYZvqQNXreljin0YzPn8f11tu2inr1fRFk1a01
/kjGAYXcjNtgexyj5BaDyPenNNuoA52DZ6pNH367BBKovMi9ye1szMwamvLFNsU8
k1+fA8KSnmA8+N1PIH1xPC5szTewo/2kJSiBo69oAq1xiceobLDRVj/e4fHCi35e
NQyaCvIRgmaPmW8NoGcpH7sjT/sXZeNukssS+tSQAC9OfvKG67xfIXgNeyp9IVy1
3gEx/Agf43+xGCvNR56TCK6AuVOJnyh/4snVJEF2pMWVpOwLYd7TRNM74Tf0QOBe
knCSfCEXsD6ybOFmMEvGYwQPsAQV9iw6GVp6DmePKffmYlGgh0YZCEAX0bqVGZC+
U3pkV+2ZzYQuInWdBzLJEQgjIYwFHwm2+/ZemuplOAVFkKgcY5LmTb7YxHzbZQ/7
6oiaB60q2A861i5LAQ1kE0LApDkoTTCJrMSDyvAA+/YLOuaxodGN74R7dFTJSzeR
Emy54znGNyraRiLsAvYx+Z/E3T4DpIyRkPyh+ZxYJQLE7ydBkS8F8qLurDFowefn
O+d7HhHW9I6VSmYXIdvArH0a6NlCDtKPOBv+j8LrnaPNluI4SxYziaSh/bXi43+6
Oz3Mbhj9NRz3+dWFy+wf5pQVCVqAoWMMAUgUxoZfWlmYydf3sxmRPhcEUhIFBprs
JiZbniDzk4BCZGvukGIGUQTKzzZKSyhiQp38N2SuOWKSH67f7VyM4HN4KEPTo8PE
5I4Tk14WaVbWE+l1sIUqqn4wcYDXyfpf/R6U3xoays3Rm7nTeD1qXm3ewBCetsCs
XwToTkgLV/cqCr+X0658QX21fXKJ+H0PyYvhhNXYYAFHAyra8uyus5QDFztO5w3b
pNAdWviQrsk+4pqzmNTTjHe2X5Zu6fdwonl6Ndflujrl9RNSEVneiynk7Yn8Q2oZ
VT9xGAWXTpqaJSZfhF/k+MNGKntnQUG5oAYPmfwA9jaBr2dQVMH5ypPvudxTlsBC
8XYhQd8kOxVmeP/RCljQUREiP7OnYx6xkSkWRwVVXmH1VtBW8IpQF22R+eYYKOF+
5+hFJIVzNNslzzujWxmNHteW0yFsvO2hwA8J2KcAAsD0GjtVuj02OyVvEis0AiIZ
FPiVlXXQVc2sRKNdDJaMRJAtyKRDDkTwdSFIqr6KGeuntMSbdxgMGGuVwoUW2uy1
3Hxgwv1g3uGVqEd+p0iy4DZnPxVFG0EIoN7XkyTXQvD9fq/LtuZhFqRio+lA/zRi
G6jBsQwfScV6jxo3MyH4ciu/tBvZg5BXg7Haud0dhqGsiyLJl4EZ7qAbnmgI+psq
HeM2FNcQtV2Wg88mgVqnSUVPaH0m5RYavKXLMLGFXt0KRRrhg0X1S5utUURE/u50
DcUA8cWU5vG0v1zh1rN62ym+GQoiG9SoeQO1toyXb2OTnzUmG/v7t4qzZ1l45y9w
Z7tj9kfJqj9reHxeMOM92uLqSFxFuEfYiQPBc0neRXC/RrnhPasB2WLuMcmIik0x
rjDeZC6uEei/fNGodP+7FdlnoHXFE9mqNGyF7Y1rlhKT2iP8tAUhiVMZnI6TK/9q
HbOM0L02mVU2zRFGoDZqwO32ERPEOcrENOwWB0KT9aRAyEb9M4lrkV7rLRNCqfWW
NUWG43DWRIyRhdL7mmPdvA+0tJcw6auQEjJXM62ij/fPrc7v3Vwpz3e8PtG4EDLX
wzj3B2xD3cNLMiTncXhyZc7kor1q3kGOjAiCRHlMdHWV5r16L4uX+MtQ6JF0hP1G
ffpcS7esyuqLXgJ4IfWP45xkLLe8LHwn9QvghrgvN+JSRRIeH8cC4ySWxT4AnZde
qE+b44kPfOY5fuAkCYky9OKLNRuCD38NGfNWWeHNzyhG65vUy61frBX3/L+2wJRK
8xeStLXNAXEIFFZsBoJgG5VlVTYyCs8r0kl7iEJEw+uqP55Ai/Oo+CHzSXmcwa39
wC8tjwIO0Jen9Inofk4Ja/0Qjqox7fY6x5dS6z99tZd2V9ZX9wVfT+ZcglKGqC4f
MxBFBkdTVNRmbLqoloQjVYvwhcmsIt4Xz77sHVTFAe++x7o5lHNuh7WJ52BYtDHp
Sk/b7tbpg9lwBO25pluaNAWmj9x6HPETVtq8Wa9CNUGreyWz56XIyyZptynTCY8t
SpHBK0cIm9jHn6is7DvC4XTht5deStpzmMD6G8d0jUIAOBTDHGeEE1RLw46bTC88
E4c3PbBD+r0vwSOAXCeWVzFLiGJQnv+wgzZyqwNfhAUwtlby+R+Yc3SNrqx3ULEp
PDYLOCawEt/K07K8DVyAdG8iCIVqqAiZETulCD4wRYlQjcXs1JzqGJCKaliVkwAD
Msjp8B8rAeNFIM1jO7NVrJclJRidriLxI/ZDQQJVZ+r1CSSy2Im4fZ4OvO5K3rcr
wZgE42cGa21WZ5AVTF98Ra7/EZVX2ixEIrUM2lzDU5RExo0uy9r9hu7EIqrZw4wp
M/J5VEx5Lzv3Hys2NQ7maLRwlncSmpRdXW/MHdmWyJYaU9HsbaUs8m/102HpAy4o
33KntnVh5izYY0FmMIfWGGVbEN1StwDOfKfkxxFWMvQtwKJ4kCWVkEU66HQrGQ7p
xUD4n06EuPSrh1ap1lWuPW/+aEVIXP+pM3+aRlM+++haTHXnmUwL/kvr8JxTmZLh
dj4G5ofmRGAw8jyNZBwDHVw8Sb7tA0irFDq/WuSoz6VICdUfmTI48b/QsaLDpW6/
Ma0FU86XkH7HaiRuHQ6j3ZLOmKLMuoSkhHKU29mtKn73zn+MfgwzkHTTytyiOA/R
0G1/it/rgSWUV1xMXWCCjvo3sM+Ys9ST4tQHhQTsE2cmxseIwAPHCxzVrg1vJuEp
opQd0PngdRXwmWnD7PZLNRZNCpOb9C5ICFiDPEm59Z/hJvEivOGH/kyY+o7QRcKf
+W0heLRuRXMb2dbdfnKQVcQuNlX20gPt7yblrDZTS2mQYPracrGVjUP5ksIqZvAS
ataiH/ePovG1C0gSlAv50XwZazzi31VETMCsvnc0UWuTx8wEd0wLWSjGV8AnAw4Z
M+vBuPsq+7WUgk+rIWApyW1Cu1tYMvQxCftaAWSbSVYjPnR6lXuHtEvtQnktc+7J
RYFfDRjbVQTkSRGev80MUbIUcUijGxSQx0MSk9Qkjtw5N4WoFBoZtS9U4slagL7+
nm0HKBXJQrITIjhEcuxJY/sLs57zT880PR7TZSFbyfgGMsLeMVkGKgtvN8uVF4Ci
sTh8WJAlZZiMqnZV2zvq3cGfxk/QfCgBdZrgGAMVe7Y/Ghfa0/Y3DkuEOEJ4xi/e
vpXHfV/uq3TPjmObiAJylRr+CXR9QO3bS4I/ur24YVt/2xay4rC/WuYZigDC8l52
PrYB3hL4Cz8wDTjOzSyZApDJWRCLCM8TB8wLO1URDrzGqQBGljvK/zwlwI9u3TLv
y8cLOXua+nb9b09eNnuSEJUEar9LSzEowIJrx+/dC5ibuEQKbZ5/LenTu4v/SH43
H40MTq6p1zTlNNmCDyWlcBhRlTM8efSTJ9mDL5HfEG4B80rdgTjZtZSu2tV2OEtc
pF8OpHpzPdVo6aC3HFDkIODlCEb+PjeRrztR2hAmpWSiyfiXZbkg+9QF7b7+s/7F
mI0pjCVzOBUNF/Qg0PPxpH3Kyuhj26fKmPaTYqdG+0tsI7tZZvLrVzXrFfE8sJsY
a7EZJeWrBNn3OndpLABlhH6cI2tFaJTw01WAMt8RZhlGa90ax7eY+uNpp52263aO
D87oYtMaB1ajtqWYTYW7TUA5kDDU2+5WpSeUmnCSpjNTCvdJZzX5X6ZxkqUPuhRm
bxNToA5XhVebDfVuZpxzpTFLaBtqjbdHNDSvnLoHmEUuLxvLD9O4bWD/BsjI4t29
zVWUEzFReCXoKzg5Qjm6c7rNsUCetuV2GM97nj59c7lZtAgaKEOhz17IW7TIChXx
GNkSU2c6jne4+3DKhWZv8ql2SEL3DtkTS9kxTLOyfaIRSkukg7clFB5m3GRTFNCg
4u0Fb1QvlS3NuRNoJuAbFjHE1WThfQ+nuiof0PnwKfOMPcpBqwWxmr9ZEFGCKaIi
40GNekMofxVKNCDJxI8VGvUzGMHop+3Kt9sgM9KfHYK4GgSuGqWGdvZyok7UdwBL
91cq3goXnVPK72JgFtudmfmFVB7OemVw4VagLShxp0dBZctpjDsLXnXMXX06Xry2
c1Xqu1kwqWxudLPcncCbpAqYKFKZZzC/0gsymrYJcQc0TQea+q53YKCc4TzN/36b
Kq2AoMGlBAoncG/MLwpNvwTR1jDfeNA2vYe3AxdkvCQU2LOYp+1ckK5qvSTrQBPR
X1s6baz9EgVfXi5rtqjo0YsJlKLvLbFi/7GfLT0CYGwbcq2Y0n5d+4Bb7MNN2Twu
MR6cQrMMWz1voWWqnPZtDHNB993dS3scYO31dZjBMEB1cgEVMcegrjBpuZkoNFDn
iusOwWz4xv7N4WBbZt6m+V/dNzK4EzZVm2d+Mo3bHOgZ+1cDA8oC3L2yz2og3Y+E
27BXFBBqXtptYDISzda97783KNuwCKs4rAIJvy14OAUTNEFOh0u7EmOQyJidzPUk
kAjTT1dbql6fuKVL6E+MVmz2Gu/2o0En5OAIncSQ8IjOJ33n7i5wMNFlnY1qJF5m
RIrC2mm2/GFU3AWVzcBFYecja92n9iieBDXF+GWlJlnu4X5xYHcw6Rp8XYAGc+/b
ql1kFhDR5Js2o0Uif6Tei/pEOrFWiWtlMPU7KOlbe2n6Xn+dqqGp/I1aUrz0H8oj
vnVZpkry41jBGXjUDmEvNAfEtJGuzc1lZsCkd1QmHkCQx3ApZ4sg40UEp5sYjosX
K6EXXquHfMaH4KGhu5lzKMsK5uJB0jHiuGwfeE3vdsfSnRGyn6E14oLlkSm6w9jC
itd2LQM6hSg8MvEriwX3e7As5Tr4H1c8QuuTx7pHvY4QmJi3ToJzVPW3d3ZAAPmY
yx/g7jKlTJmksyWwIMJTXSeQrKHKWtRIVXZaoHcu0XaCFCU28Fl0MjmRJqYtnq9u
klSAJWQ/q8MSrlrPa/M0uhzUCX4ibE0+L7TvixjOmZadgodeFd94K7FMh5B+Tc9y
m0aBHlkTxbTaAjpyExB0BB8JzVCcq3vVSRRQSwwWc3pBKG2K0oTIofyBqLPLZQdR
q+rWRkzWS61794YRYRT1XRsBvUUrIM03HjpjpGREoeOPD8OckYsnqINFRa7+lMVZ
hbfK2VrbM6HY7Y6hQO7EEPbMCFGiF/rsNWTqJk7zkKR7VZIcn9uz69t6mYeV8Nil
wXcoL2ZdIstWk6fuyJxcPaeemFPUv458tETv9tqW0tg4W0QZNIaUaFnfD7cnGJqw
F+RTZIV/iy+tpLOOgd2Oz8c1AbnvIMNIgpJ+HHl0AsdIDaZ47VxGI8WPtqliRW5F
Aey/Ny4pqkcN0LZ5YmAGfWnNbw1oEXGyBh0E7NXgZ/sTdcs68zuPUotc9R+xJtOw
hoIo69oErWChr6/VfYqwjuWNhik3SDaeRPS6j6i/7OCNjkPfYoDgh+Fp3l3TyTJ2
C9KLoO6sW5X9jA47zGyOu7bIOYrMS+tiuWW5/LADSTLFJRDQvd691JqcLnwzozw8
jsu8JcgXYJwQVc2BNH2a+si0QU3qKhCl2+78GmMviLexi/ydiwJpfmymtcyBZAgz
Ju8g05vWwYZ6ECEpjtX+/yeE0fsycv8yIhxaqkBBtfqA/nlhlUGFAbUbOcloJ3Nc
s8VMez8NbzvjfU2syCtFJWFawEOIy6JZgP0+nENd/d5HYYv4iegVYMSPnuFhC/TD
TR2nB3rkMtuTdhIgQesEoDmDC4ihQdnAw5VoInzp7EJtpONgORh0zXKSB7wWOZ/P
CDcYvjjkKAwxjPYh0xma9wH2nRKaEIs2N3rERznxeogGKbrAtmFKhu82h+R3U3sv
4C7wHnZY/RyXdQYs/IT5gnqxY7K28eAu9n1y9780IYDpWzVN+gPhkt500dlqk61L
LuVFdI3eL5F/2d0Fpq0wvpyK+twFIc3MsMT6aHGI0MlvSOd/bcZc0wqfsg0nOwE1
8BKKblrjJIfhWtprlzx4K3VMPk85I5uGIeLYj6j6koetpXoGpGwpppdnpbLkdrG6
bErRhPxJQFTD/yPqaPfLTsdzLaMg7LAoP3GRjXRYdblCDo1FOJvEkUXPaVQEIBF/
hZw7lIZa4J9B8ZfaAgyMYZDvCKsRMWeLTsnBmFXRDP+vLfbL0QeoCTsNZSS1FX0F
UmtoX2e8BB9GlDmVCw6V92dZ0JTdnfc0vas/sHiCxMPnGUolSisP23c/9okGyNg0
JuM6WH7F/dwJpdlT74UwzekrY81GOo5Zw698akln0dpJxqBLlYX5Pb0WcQmDl7/p
qSK+sl9FT4Ue3vs/BpqGqDfzyWBR9O+g2z26hRoAO/s11IaAPKCMKHWWA4tNRUEw
a43K5gxMoE6GG40bNe2OAty75J7rP+q0le5omA8BLGLjSdwRcg7qw0Lg1ZrNUirS
VllN69rAMF2g2P7UK+thkawcNE69E02EHaFBJZgHu6DeU2pawUG8Oytl864LbmSp
1q0kAiBuviSs8lxZbYETBXSvqlhbw8JGnY3UMOKqIn0wWLse4GNaAr3MElb3hZdN
KUkOMZJY4PEoAMUoI/w2Cd5EiKRNjow0SZNHqUKE53C3CKWHoPTd83iASkYARKUB
SvCr9h5gE8WGPwlujzjvsHDnGpp2oamb121QZTmih2HbBHuY2zjFBbfRb8n0S0FB
z/A56VweZUj+EVrXL7w5ovJ7JvqdJDkoB4pardc6SDeW8dQrHQjQlPoez8NIDZEI
4BcVyIOOA82QWom2Puh/nSuGhwhFNvCS6xBZQ/Gy/BV1ANeQtM3uuySqo2qp19W2
ttorYzHjtNjXaL+RW2g5N5nNAukrAQDaEQzEzyxn+ZaCr+hSt3ev87pHEEEEYVzc
UWjte0EsqKTBoG72K1xGCPvKxUTvbMczTnjLvHpKzEq5B/YYPbCQkeywTWBIkg2/
X/FwxnBzfu8He/1ZwinXxyF/rJglJrwlG0XhWfsysnfpP30ZtXAFdOU4ODQQHDKC
OUG51wDLtq4weV/OBsGdBj2fY54okkJfXSnlkpie0Kiq0KUntoN3i+3L8rqJvOLw
1DFB8BuEIUuRK6YGX7zCqeqI6Zp9tbm5bd/M9whsO3VI6cck2AXyWGnUTOED9qh3
HCDlVZ46J1CAftLv4v59/UR7jiAlUnvPIyrtbnbus8B6v0pQ69Eqz7dtC4INY/Ap
uqRzcaNfl0I9dCA41VFK64aNoOM5ru64bTJUidD1bEBEmRe6owqr6AHtlEg7hxpe
V2L9f6VWnzPFsRmiuRqCHXNDXtJUZ3M+DtyY4XxAebm1o24au7X3TTLZgFhx6o92
C2btkyhJZnPEIvO1qmsnMtz4n1vZnziqU9HfHXEa6zvtjBrqwcHdOqJcV2crx2ng
QZu+EWvdD0pfGjaykru7WlXa5wWHHvevugxujkn06dMdZplONvf2CCQcf98UAawy
mpqeT9SAHJxAiiMobFhMW+KwZX9S3+nLPmybgPRWIp6DJpt/Oehfb5wl5VS+fr7j
hVDsUreo2x/IusReX5k0H/gSUcB7pmkWBQFRC5Qg53LdhlKQy7ejwWvAXbE2P0b2
q7F++KkOlli/sMJmdS34BMA2BN3OlOYnNl0Mf7pouyN6T+WfkmP6KQ1XU/iDjIbw
QizauJo9eAB+RdTa2cx0OU+pH+IByonVPuOd86xpJRFXeeq5P0PIqOUe0vikdHny
Lniv5CpoiIi+3Dze3zhSoDqip01uHvImZi7aT/VrnJ6dTUbKSmX3+sRR06VKBbkS
j5QXkClTKHZSObdssHxubrCyd2Rr7UzZ7HrILEScPhBgeiJWea5SEO+rTPH4SbS9
NEUKC+cgyDL/5/bTmDhTk7h1XlxmMCu+PlGD6g+Mhzfad0jAemTuTJMJZJLrVu6h
QlMCOQruqRuFNIyCzvRL/mSfanMePGJE8BTr0BMksydixpf/vhRmWWQ25Yq5ySeD
xAvEcmjYrOFzBC0RpDomvWQ7BSrh3rk9HJ46qI30JDZjePrGSAYWtsMwW4x4yuJT
lsPO5EExUiQ97sVWXpguxDGgZU1PerwldbsnPftZT5KgKAcm/pvoGy/GwhatDx85
D8mfkEpE9BoL1hc+CF9ktPVeHCfYhBqsqcXhghKe7dsPPeAXMXhSQ6cgKk2DHTiW
RATslp4LYucurHubI5AjqZgpUIaBFgvmGwi4dhFhADueITY6FRyqtajFaYbYxM2Y
xOGIkd8G2IKmSTEX5R2hW9Z9bFH0MBToV1HKCHRLGkxNr2BQ8l+4k1BAnCIDphdd
cqB4id7D8D2M1RCo2r4bQYuYBx4KCR9ADN4NGE3/EOFWRiFCPbvq1PiGNqXO+aQ/
L5eyTI74bIhtqabKWbuoLG/ZQXt2IQZhv9mmW/fv5yqqNLRFKIQZjkqFi9AoDMIu
aZ0pNYWd6sAykTsnT2zX6BtKtRM2AL8Phm9i4UNVNGtMWXNGZBMORHSoaKOyUVuo
bOPzHn44uRJwOVk3HV030gyrolDZYaAhbWJf/pCMEXrR4IY2GB1C0SbhPctgQtE3
RXQw4Yrdl4nUiZaLwGi3/EG6+7HsX9FaOxr5Ycj3z3jJ5eP/R9sw5uftPMLk7oWz
Htc3kB31Qmp6gTNVoWp6NAaag4vJBjurRADFi6eIG+Qm04LU694AP9y+BD6z8oAy
Sp5hPQbnQwGnV129SUBuypmxllHmdRo4N1ecVIsD7n4FlHN4mWP2PyBoaRrEGtrB
o6AfZO+Atnr2RAcsVLN85vS2iYUaBE05sp6Qp03s1kW8d3pasxewpgQTQ3p4wF0L
xJ4OClPhEw/a6CjkuZMEQkFfhhK0taIE+h+ebaDxzW9m+hb/akoj0ChnNT7ognte
ZkYsVdZYZNCvYZ6cBHCQBOiTXQGsZtP/rxdDu1Px9rp8PkXccuK2RdP0mwXlnfuJ
2fH3CKB/KJQOv6i5bZW0M5Ppqop0fpMNp2csjsjKMpj/Clz3PCY4u+flVTXlamWL
pCkcNn+bi4cQdRHSkTYSOCHr3KqWeAoYv8yNYivLkWPT5KJWGmWBf/3JB6hr/3z7
TlG+wGvwgjktla0xy870MzVIzsTDLJzv5lNT+lBV45iU2wlV6RJuGwIdBzbHwB0J
TysdQTu0NBbKbsAYUBIXazie+cSBT2X6yhgGhFfHlakEkBDotdzcugrwnafNV41A
uf+fbfwNuujQzMLcNIA3UZ+z4WK38yqANtZt02XIbbAbLVc+SYOtgumY1ogXf87k
FJZgCIkhVruFwCad6jIJ7bbGFXmJuaSRnQDPiUXmn/VtPN9fGZ8bjTTQgLJWe7fu
Ii1ilbOfoZlMO+D2/MBjz6r76ZzCOTDchEHnGxVRqqa+S7+mXGf9jp7xsgrdNl3N
RGyOsBKmwpGi5znOo8CXS/LxaG/PT1CHQrsu1pWQUw6F8IEh+I1yK2B5ItPupqlA
8Wmrad27SJBcLWOfOoM8cM2LjQ8uSUWnxeLQm68PraOqOnjN0w8Bv1ApeU6BWrK6
nnDdCE7mnzaeJHfAo85oh/L7F/p2N8g1knqIUOjR0KmLLV9vQt+DZce1U4mmxoin
RcLXMlm4SvqwLEpF+Tj7i7QwWd5A5PdjBrfKtQ0v703sx/dN3FbAf+/RsnUKVuKP
Fhl4nmHeoAZzzXKBjRgYt5EFLONtLpPoPbxyai8CKiPAcRJ/jKq+e7XrxMaSRjoi
yomarF0Du9lAHTVtevNp0dULNkA0QmUabBcJc+hwp/S2GwFZ5JQeSX9JT2smtm/Y
jfnUy7brMryG89erbP+bmGgZKzc4Elnms2MxrIByyhkaJETJeQLvYEYDEQb6N9/t
iXgXSthhOIrolvMmP7qkZMHC1xy1TGznlObTMAKO7iBrP+xf/5kS6xtXVrkEqAB/
9nvO/x2LkqmyttXUrpj0mJ2G2sf60ZMIjeoy8d7CNV2AVngtolYAeISqcCpFCsq8
gfLJCBbVgyKDcFFsMy5+SSjLVS6EhXqkFvNg6esYHrB4Lc2isOEeb4BNWfag4y+p
l9sS/A+bquRpBPBEWWopoGqfjmuel/zMvuR9fGMzVkv/9KT8WuDoQVgtwDIiaTil
asJ86bTmNKWsOAVUUhvCa5TSpNRL9ELzofenH7qh902qhLhqqFUxW0qwSUcLGaFa
Frj0pyz1VqbfvL+LWj2BO3Md7tb3dPW5Iico75uZlhJ44zMT0dqJqq8l6prZTRnC
IVWsf7kllAYJ9GDQrKDXh6yE5qTvR6MXbSHzSlAtbscmC324wvJmFWerfCGi7uBa
G9KBKTzIc7EBmYB7sQ3F6asejT2SghHrEEC5zcNC9rCmiXrXSU6T0F6yr6Gk2Moz
qpfzA95EU579daDIQ9FHE7ighTph/T5XVi6dhTECXyYSRNjIIZ4hbuCoxGT5lqE7
chyE72LwFJTtjrtjXLB7LoUP7iKAOl7EKNdmQfhZX7Fus81QkbeyjeiCpYHIHTBd
joyPjURVz3UYwssDONKJI52zPN5V2beb7/iAgZiLXNWOhOaGt0rLpoAlZLX3ZkRg
RnyxXYnB9FS1ZvmmxGyOQjpnAlOWsiPi3fm1bBRvN8V1fjh62oO5HgRwmBjWShCG
kbBjpuK/IS61pVK0ILMPR1WtIkeOIQFtODoN0edsMB2aqZOdwgpcMvAkNGvHkJUh
5dXixxDXSJNjqEOfv6URwMkKSib6OhG8znN4Y1hM+7C5jaojZBzA1m4wou+rBJdo
lKeBxmh8C+zU9fTSCpLQUQjABo7KxAHFBWOLKtVSQ90/1Oxg1CDk6ZRQxNyD3Oni
0Hb2UWd+fI1Xe+pzSDc9Vmx7ev3KN4CpNROB2KXtYSdkx7EUYkHwoGDQASkMbJe2
0JsxB94uzwKw0B8ob8gxtXOSkiWUVmvlNgmAgoLng4x+BYsLJeoD2xVgpWcJYwtv
0h1yJuFdxO9CcRMGISrDywxzKqPRc3bTWkOnmfyyNIlSEznp7tUxhWlTET7GzN7J
VHKsJCz/2p50p2Hobuc1lsMiM0UA6J087KDJbdiPYrzATZTCxq2h9XQuvpEzM9E5
sOBohoPWUCxN83procqa2OVQtR4Db/3QzPLNRrfNDYjcC/Y82kdTMH0ucGZn4xO9
9Poz6zSlXdC7R+PndJtxhJrXLTy1pVXm/9tPeArAa4ojlmA0ymRtzGQ6GpQvjSUr
l/dbFO/mSDDUrw0DznZEihZtriwdZ53k67R87c4ekn4r+8vyWtjfGtG9Zc3v8kmY
GIGx5XCOJJGHHhGuR8nFtO0FjzSNHzmEZY0KZzkvzrtg0IAZdizsegxZzHknwt7/
0bK2bBiYxoOxdByds0TwpX+RkweygnhCi8USlfTTsjBMEum+j0n/w4K6ZLrq4TW3
MVTujIALmH+3+G1fE4yEYTFdreLbDbz9lv0l89OQQr9+emaebkOB1KPOvU/imj3M
IY9ZhldnxGvvoLV5Ux4F3ZlclCBNbs9CP+6F0P1c4CFDT4762yff7axlMJPyMLLH
ws/oC5D6H264R7EsmScIr74Zyq8SCwNPEZEH3Wm2/rRmB3+VFx6Q9yjlrbxjWzdU
0Gy3da55kTV+WBJ28/cU5nGLMPFY6s30OH0DL6wF3AXPZ9d+h7bvwG2TF0r5pzz9
UDLnhCCP0CNN6CfifbgwwHgxMM72xqmfLdDWAgsoODuk8ADvJ4JRsDJa9r+j9DHw
X5arn3q2Ch/+059s+P1yhznrp8IU/Eq/RG3CAyROQM8bD2K/g/7W+g/A78aO36Pa
zeE1Ip8HbvV9a5rKuj4bvKSWuwNlcsTJjItyjzAqXAcG5rNyT0bMmxIFWLiFVCQz
vGLR9zfEyQs8NZBRPAMDUDGGlFLRpuMKKfAlYeiGWQTP7k6id1tfbgnLKN/J9+vk
o83XxsiLqNofMDLUfn9DuefZUpaqZphP/34ZAK8WJSbqBLPimgrLssTpFnmn5u1b
TTvQGr/JNVjo6l8lyPc6k1Eq7ODXht5OQ6iFwopBYC68gIGzqMKBzg2yOv6wZFc2
DxXqCrMGsy2u+ilQlHrFx9r0UZ5uNDCbq1JzMNdZ9VUlVsmT2oS97vsQWP/dl1o7
Od3zoOEvSwPZpqfFvJM3h5XBhfHw7IdaUv2VEkYpHfHkm+56dfngAWvvjs7U9JzV
FP0ObYq8EopO7t8m+pmOqYR7w3MXqu6CLcRln0eS5ujcFlWCo/858ysYi9D2p/+M
ToMjNVfnIR0EZ5ujn66DV7u62ldBAbKEijanM5+ScOJh3qAsIRGj3Ifo0rSRxKKY
LWb9seQ4kq6DOzKaSKz6vQVwO7TLcG9HQsg5DUrHB43UBHPvEgKm7j1ahhUPHIt+
vdlfxvKmChrfrVBeF2ICch8FqSHd6OGWFGGzuSuTrhMG82MElNHDf1l0jgdhFlNh
r22NyU2FJar/R8RoJjOWUyiEkCXZdcdT5oWOri9zUzM9I5s0iDd3YDZWSdwsM4l0
yaLciOYTGmGzZ0ANDnER3uj0/LH/Cbtpqx8BZKidAS1lvWtOzZ69tSPVyIHpxLAu
s35gQuzV6jYjBM/1j0wZZVCkXEkHDyQGSjMGXLnevKtp3F6aYZCKCG+mcF0A6WNC
GEaO5FybjUgnjs2OG7vaHAiOs/9Gn9UMN4Gg4maXxG1iE4+09BYwHWTLR5BJARSl
OPRcwhUFxoySie/jldWG3eXvfNRyUSbrvRd4cwm5dRD58paPpQhJIT0U4J9iN6RK
9v4m7fMo+5X+DJQ7+NHhe9ErmhQozlF8lyl0jUQRtfzaaRpEHrmv035LkcZQ0X7+
zkjsan14yYrDUMLSWF84gXPnJijp6wM8UltpQvaWQHx00No7beaXtDP7fP94cxdt
h5ruTCN4QvvuBb4OjXo3J4utsGFLZ5NT7Ef5X4ZoiPVurYsNAgfn9jBr1S9/I142
XFLUVt8lVerp8omN1cjE840vnUWgsIwDyAZg//mSlyBrmXOSf1JKgX9PUHcJe7u2
io0gaGZvuJTMsrOs9G8ajWqHxT4Aow+OK2gURi3onKGBqXuH+qYJtJMrD7Lh+k7t
q1qWHqvtjYvkE6RdzjloXCwUnRvY2H2MJkgfG1JbkxJ1PSd9bKBn5lAYethWkw+e
TfyZQW25C12uDyBSAv8lroLozN7EfKqy2cN21OV8iaIvmpdDJzo7384h9KQ3Npjd
5/0Z5clJ5QpGzxfkJTs7xWvlcqLy3PsnspVtFAGqxemUJPpuzWgCUTWVsPlG6dql
TTvJeOyvFQyu67IcH3HXc6R1EogOcjlNDVlxZPKp6XUYSCLrvj+bZxE2XI1qXOka
aib0eNnkbb7lTQOCNoVoieQa0EBUjT5PhGEif7t/FC9y16a9mD+zTWlpujwWPik2
Xw+P5YJFF15DnVgLI0/ydKH6y+hiKfNfc3ShP3A6SLHd4vtfi5GsttE9iq71E+0p
L9Qj0sA3Y4s4WuE0CZgbEZaulf1rdM+w77FI8IiwS6nxGW72KXUilOzK0hJ1KE9x
JWNma3S79+ionlbuwH458oJuLqRcPnDh2WtprmD8DQON6c8GKsyIqvzt+wvZLHrQ
nfQimFBtxN/TO7VsEsI36XPvgUUdQqw6DyrK96/HgSMKOrC+/Ag+/Nlt/z5JTs+k
ZpL060zIMrFc60Ayd/juiQkYzbJIzBgfSLz9NJ2y+6fj0iWBcFWTOWFXhQXP5wai
28rn3EZcIoHLtMpeRGomJ6cQZAbofxqe6PyVJLLaOJa/NXlTDSLDBsLKigUVNH/p
x6Q+UUQQn9nEpA91jR7RQ2Vz0Uac0Y9cP0g6Wrf8BLF4gYJ6CXMZBlCTP1LYLzxj
1bJPHeOIUtnY8wM1nEJCvyu19iSU7gDf/ht1EF2VsCCpkPU2738l84pGmoyGYusT
PDJQyyOdCPtQrpgOg9jGIUCkQyf5ZsMwQ9VkNC7KNeVj0ZVz5rmC+Hii5SQrCj4w
dT8XoS6dC69HmoETjR6tozJLCpBminZcawntBNSwmy6uW3L0UDLXTEUGiDFNeXwx
SWQxbOOMERRaFdCN4Tb5yKbhOcBN/rOmMNfuKnQGeedLUlncJc60pb8aFSpy7DEL
llDen1+SUf9F7pvsixn3HlwBr2caqiorqA8d33xT7GhGgsJjsLesVsBqo2iKPIHp
Z6TDag9/Wtxc/6Ucz0TcmUPylGgNh5aYztBkXynvND3tS2ky2ANOIoqJU3xAQ9tr
Rl7aDAgm4RJIMuC5QTrOuLaYJMMDPGUHmwpAWO0CiQPi5IDjI5X1wjhxL/ud8Smv
S+9w5Amm6aP1uaax30DX+oqj4RES3AMYj3436RYPdYopPYUQbfIBGHL4l4jWO3w6
Czk9qdedsaH6IQWpnXvAernr+zOmV8htMW/YfK2fsDnJB2GZG9uRJzP4dKRpuQrN
IvqBicG4HkNjBfZcu7CnVs3gYlPxdOKe63hwM2Lxo/NAtPgC3w/2p3IOLlbgjmym
NAyWfDFHV7ybwbGbD8EX9A+TTtXuU+arNR4SF8sh49gGMveDEVDHXx/jQ39j5LF1
HZ6l+9eaSAKl4IY3J0FpnYghlP0PShsAiYx1mUPI+3W0pBRmhszVdXDNdj5iUPsI
3l+YBxoxtEbqVnpC54jF3qw2LdOWx0J6I+n4T+oKKQQu9EbgW7EyuuzF6/EyIiwc
P8GPp2V1bVY3mhmx4OXshQHSNT2xKIYoJRoy9T//bOWR+0UnWT5cVLSykpHlbWya
cdyQeX8j9/obRfcgzRlzYEALCqVkqvRdWfonOl2IxOXJeMYEFtRku9QFZbgFyhkZ
oO+lkdjCzRuYAud+IqZDKxfleHO8gOngFGl/xSTuclFfiDVW4oC63zAEoAWx+rBx
h5halrdCa7mAHfpcovab1xUqBwf4A8VCWMNPd9ml38U/9YzvZQvDTrBs0igwkQlF
67K9k30B/YRdy8985fWX52ZywqbBWGNqGh7iJaHZE6JpGxRHTMxCPMfHR9HjvVQs
8f/IuEb8oOH3X70Kdis0FVamOmEjueJ2g2laxitg4jmeA9EK65BdTa3Bw717AwEV
qTXg5rwRSwD/hc/EZ4zXrclG6/52UszWmRJjFk0GCMngBixGM5My0WCasqWuN+bM
0vAM1nGoaf5tjGE2IXFbibC23cIdr3qnuOfdyj1FNTWQcbx/KBr80beE1tbLyb4D
HLLgJ87PrEhSerZcu6BpDmYQ+mYgrL3xYkBC0dtrw2zZVYIhMM7VEu29Cf6E1GT2
IHgGfxihweQi1n1wN4Ga9O2P8FLGjWsdg0M4p9aj/POdC6sOUxnAMFzWKvCxgz2C
+Zu7bFxI20HxofkE2ZmKCaFeMgrgw6+xKktGpLcaSX0eOo0s6aXpoq8NpKqsTfD9
GndoxBB/s1MC/OHn1AAnLZ0Ms7tVJCOsa0ETpJZo8oagpIkadAiTfLYMoG8sKQX6
vy1xtkVlQ8l9BBRQRrwWEkO6lc4ZcatZt5RFAmWytukco8bpjNKzE422sABcC+Tn
bHZGVI97CuUu/twxmTvPJq3FcDE2Fi1REUVZpsO/JAyTU0j01qOCnNlNqGZJj+LV
VkTFEfNoXcLxRqF0k1eGKGjfwh/0ocCtoEX2j4x4WRY4F+jkuvCSputIbBfUjVCE
sSryNUVC7nWHPsdNDYNzSW/e7APBLf6MEeh/+OnwNcBfZAMbiyhs4MY8eg/ZeZsb
apune7ngIhZ2RIbgD7g5d185fQtZNeuvFR+0+oRUiy4Pm+QvFZacPZaVvdZjvvXD
3BdFCP6GmlS2h6OboFewORxt6N5ydnSNQ0NeZHoYR8BIB2LPVd6Xxc+ZuSsqdkRk
EEx20t5UbM4woCaC8HHoLENWe69NlSwiJfUtQ4er8QlCiy69ckGZ70zh9B1TqC0p
6SxGYbdZBHh6J1DgguT9xkxeVfB4OfVujClSlZ8Gvn5ROHtt3uE7LpeagugWCZ48
tCHCxUreHCiH9AEXq7QC66PzUS+KNHnYg1E7ggeBWyQrOWUhc0chw5A/TxkeonBj
qzZx+Mc75F4q/fV3H3dPO5pnhnopsBN9rh9aHcOyVr8bmYrkZxsKCP4tTVFqWecK
N7KgRNKHaqPOJpHikak+l4OUqJ8izz2xKmVqGjToyUUcbfz2daCZ81CQxlbyfbvK
4ttPQrpaerp2dYoER9d2mPl8k0TT+hxo/nGWyB4Yt0chSZPWS27BCKJ+E8zKk9xa
ZVm0KoXRtxx0TMeFron64UfZcwX3Z7k0vTsc0wizPmc5tCHRdc78IMVN5zqadoKi
XfmMBUAiOX2k5cWhUXrovehzUXtpsc0lLCPwa6YiVV/3X97vNd/+E3FMXH5iY2Jj
NcHAaiwKcvyTXs0r/8KUBhh+62qq9NnmBIPHPUyMsZGwKapqAOqIwrnmALzcP2tV
vI5JwiWijpMz/xL3b+cDt6oMCCrCCvYWuL4oVGHbcRsjmHlfjifssoOvW5CioE3n
xN96cv5cp7gRYCB2jIbBAtMq+SLVpkcj9PAHr/4DgWC/P2r/sYHstKPQG6+xzjYI
HitLCf06MVUVV+8VATUa1fYyAOPBmIAH2ewbGaNh2k5vxFVDWPotQgZTPxv4UBta
i0UTT4iPQaFovovzvueX62GvWZx2LFBkBz+sf5H0U+fJPXLNopuG8KdIV2HsmlVO
Wwn0Pkat0vojFejMnwGHn/WE8f6SUTOAfoSju08k08LI1Mrbrq+sLM1G7DX+7JFT
/D9frXrnsXUHXzgQzZiNrONF8Vvg1ZEBQl1ubCnUUiVI0z/7maJGkydvCDdtKAJK
Gkr2NgsIr6UwniQnwQxt1RU0Px/RldvaWq1L5OZrm4wdmrGDkhYVCef7zVYcg3nq
IjtB3+wm8X4edw56Xq2CosoVsHsETFHt343fdjZ2HruAUeJ98UBCte5nRC2d0P0x
XRprG9S8ckMOd5dM9HgEk2KkmA4pFMj+Xgv9dk+Am8yLHgHdKw6sj0yEPUQhkpaC
1hrgXgciMIpaxt6lrHCSSnWjCJKFHB+ey2a0tqQAnW5h4U4TqSUsrTqovJ3lh+VL
kXZOBD5y2/FFtdBeADlq9VdAiLyjN3ZRVCUYENp19Jzil1lEj7FUCAQCVmfDvV89
aX/4OYJh6vin3+msFl36+FhazAWgYkLKCggn0Ld54G4hOKKyC+jNjpaXuHbE8mPM
jmN4/nrfbRgoJta4ULOZmj4tSk1eBN4nx8ZTj2JIJ0SruuW2LuVNckC9qPTPp6Qc
TuDOQzAeZLLM/hGeQ8OZZV5Cfh7R6fJ16tWWgwuUZ2ywFL6Tr7kH8yUw02OPZLU+
gldDBAfo3cSrlfp4DhgtBgYBmo4DPK9/NWTeg/VZIQznfgF93DxhVf4qo49ThOaQ
/o1oF/Z70R5b5l9ack269dmVrHeq7fa+6HpsTVLVJEGPZ4KxV9sEP/2kfn6vTuw7
vDW4hSALfX8HPH8YCT6AMJubUzv7I6odivunyg/mxMrYsIFXhmAC919gWYFpR5ot
TlQt2Pr+tn7wWcxvfYwh5eQuo3pDTjNB70rY2/uEKkEBHi/CWLJPU+XCN66SEpmS
kWkVbMjxsUFr8L4CkorsqFnAMtLZ3Q9eHk9yDxz1tneZektk1YzGjJpgS9OId97G
qMJ2GvnU0Fo/cGjdrtbq3gmHqq/Rwh7BjFl5aREfyNQ2TGfcDsbPv+4jMzWn2dFU
XS9ciWgFrMNx5NNDWWEz5CZb6Syoo0l1xjFYwhOwrr6SEcSsAY60h/wDfqPjmWTF
M12aeg6mIT0U1drVUWdv+XbLbFnhssvs/0SpHKd9hU0dgEvjLrJHLyU7nuu52j+l
1aOIg1f2FDeGdq/RmmV+iHp5cX7WN0FuMBsqf6XL+8TStMtat8OO32M2j5WoVa03
wchcmd31CgBPOvyR5VKNVs9Ay1KHC2PshDu9glBDlH1N2E5qDP6FfvYV4n0TBKfi
Sx7fQnoOp1m3PnwhTImeUCsFQ86QKnw/jHIg/XuGWNB29Aip4PkH+sFt/CJRtCBa
VyG+ud9H2dm87HDR3CcVBTqfza3sPuV/r1ngSvpmHMRmXBPFjLoDRPmES0o8qLOs
O2zrKt8dW8lKO431OPOdd8jYBMSAUYlk89mpofrNxxqE795nY7IgvDHUsSDyLKU6
AoKtWnVt3p5yx2i7jyVT5wKm0HqimkIZNrOfjZQrUJ+mDygOWlxsrtGtLjLn906y
ZoOYrpQEcu0/vZv1z2GkGi+14gJzHfm4BKPFvDw34VFvSR8k/prNo71mzWcu0lkz
P/20omntDnaJD3hJKs3RijDfnWKuHHmYVE+fb4t2WG5eLwtsBzUulptW/gotpyP1
TaZv7C/1WoouW4bYjVY/pELGMsQ+gSODzT6nXSjTOypnNg4Vtsq+/F4XQ/WCiEN3
S7bGHStf/TlzRXJhY/NEIUd2Uop1XjPBgvsdAE2lY57V9n4p5/wHhGooAKBOXQF2
tevps/AGPao1db5t6lGTeEuIEuc7ReSXs28Uw4fKjhWIlbTK3xLdN+gnFwJ9OH9v
QubwM7/YxuscvZE2oCKN4cgTkXn83pfrsHBYmOke7oYLyUNHwsCQ/CBvwyWsyFnY
e3NLDOJap484aCdH7DYekPo1aCybDUDLh158PGikdxpxAHWZNb0mkF60BoQUIvno
7iuyEZlIxvA8pD6J5CcomrmMl+sX/Zqyy8alugGOQu8jeJ/46KHwiO4SjshQ83bt
rsPAngHR72JMQCUJ2DUPNiESjtB1Ur21y/JczxkMQ3VXAXIHCgBMjeME86h8m4RH
tHFdBcYMG+B9xGvGv4j8+ZGUPqJGS2Oy8bixOqo/+9RiwdJA2K/K7B1UUBSzsdis
mhQ7MemOFuSunZPNECnTLz2Za365HEhZSp2JecaZqKLOZIMASdY5azazFnc24Thm
+76+JERh0hkPwR4WdzGdNAK9QymEMdQogL0MyFy7tgDVG+O9n8qzJR+VEk4yAn+s
RKuPrLkFhuzOQTp7D27JmgiAS7TJ+SMK9AYCkNA5WyVjRaCjy1RArhVLtb5I0+/w
yZxHcdyma6DI8I2w9nj7URtCwax95xMQsLpXyFeItafnhc50yy1IvudXZJFe+LoX
miC8ATSxl3fkNmWY0+eZ9SQ/lHVapNDdohBO/7mVzePQUlXF2M2OJLOyL2Xw7Rei
8aJzLxdjVX2xOnwqyuLhHIB4caIAjecHv+mErnXR052rJSB4v7AscstnXj3iDFXj
Ja8qIEdwVJmVYYGdXayLT7GyLR8sWOyy4Z2K6uZ3kDhss452RJCfwHcNrmrUCzgi
NBEqTh4Lv1etl7HZj9T4hUWZtonyIii4zK3SOPhXCMFnbMQ340C7IWz9VqdQQZFf
CS1BjulPgNTsLjFpWEU9/e1iPWXfQ0k67enGurFvSjWSPxycgRb+aYhoXcjIeV44
9aUq80ArSICwMsK4jJfkbXZzD+Bzb6woss/lnBt55Sg/ZD8CTQGQsxJltXTBSKsc
ymNXx1ZbnpjM8aE1GK5U9xQrk3P9iWrEdm8QelMmMBBhfMTs+oI5in1OIENgq4aE
SFRRuYcyU6htKbbEmQNfo5togYlmRRfNvgKlTau0i9ZRDdZJG1F2mfJUjQF5Ndcd
AwAt/PFDF1ui/Jg45TZFB/Ikm9ShnKn070CZTga59+MKrI1SmS0ks9cS0+aOito1
SbzuB88YH0NbKBZ/gUa3Jh7fkGHxQDfu+U6PSj55C4zIpS/JO7woRoxHWpRWgoIe
CC3fl9jyyDMwhTdr5YoDBFmOtO51Qu4kHC0HyMQVUD12Z3ptmpftopfW8SVTO7Fc
zotUKG6az1GIvU5qNV0tfnUjZLa9cuDtnrRKF7NU8Hu+FB635byYahByjJ1hypyu
V/2G7c2oqJKuapHAKvc9b/l+0sQJm0/wbuO46JppJF5FTQKaTZFZFU2iVLUQDCK3
LMRK78mKi5OoL45nfQmmFBZ5XUKuQi7rvsv7OW/kkEkIfGRzmpBw7DH5jeWd5pL8
7xRa5lFB9TvZKpYjM3SzYCrZ1S3rcKzfidsX5bqsBNRJS5KZlNC3OPdJRjNCVEvZ
VDjYS6ieYiLFaKqttausv1sxUp9D934Eos+mvWuJ/Apr2Z5EEBrtzVHRvHZ9XjRt
8Rpk3kxpQScKDlBEm0QfSOWNs969BTgea5zOq+lYtF00QLXdqGpH5OIx/wV9LQ2/
iXSWmF73fiE1rLLRlX5tflsvXMeqC/l/OMv8BzFJHqiUH9Bt3WS1sw+24AbgrvoJ
j1hEM1wO4JxFrvfccgU8Hpl37od0igTdeOgDTBC1/DzwxH4I3AzzpQRU8D6+uot5
/D2Rzt1CtpPUla8p28H9CUIIuCBMU6V7ATY2gMMqVhbNBOHYp4qCl1QdNA2jNF0C
CL/E2Rwh6AEWHL13rzET4EZrFF5hqfe/q+Pq0Di0nFZR22onrw4pYz4Fdm7Np8Ly
ApPTzE6YAJmmWY/8xU8+oKZlvy20yMnWMnLBfuHN/53hh1S0ZzUEE7+Nx3qxWHCX
2+doqeAg9a843ggu4b8nuPtdy+wDK7H6hU/WeeotF72HYaGflbV06gp4X+uDd/Nr
Lrp95ZJ+uv9GVE1zutUOcNzd9FJNhiHtl9oiMs1O/5nBh/+nQKwE0EVqalwx3OTf
OXiI11TT3TF8WQcSH3KBGNH4PD8Z92rlSpzLlK8hop0oR+l2RhBmu/ss8jsT+BNv
K5bRJgSAcM5YZB5avKsWQp8LpMxNf4P5Ku+KKck1OLo7usCndUhCdDNqVk+G/I58
SjLivmMNFG0tBTclL2a0sJQKtNHk1SVY9x2NypPvuiPkxrHQ413DzVEiYfY0n0p/
+ZD9qkt/36j7kDJDJzbRAl/UczmmjuJmexAiDily4z5BMy9kqER3MAfOJQbuIIKb
j2uvm+KFkeg4FxBOI0Erio75ibUJRQYJ7VlK5BecId9xZ0PZ8zff+Lb+K6wj/jkA
kv0sd/zkbqh3M4geXuQWqzor5gZCz4XgDVUpyU6GPx4xpSjXsTjtO7OKeRW52Bx6
qi6PfLQ4t3Mh5eY4A995f0ZI29Zy8RSlaPeXtpoqtrV5I+GEY7e8IyoGk5f+wvWE
HTYLS9yEFE8Tg815GiGrOA7jzHEAgjXzG69PKfdKLgQ6Qrn2hZykW+/FwAR+19ar
TQ6VtT+4hnAfwDVtG0hrlrjQnS8kljBJePCNxz9hl7vg8fwczdP9ageMZL1RTwUG
KjI/PwdN3RvrT2WyNaRfXnWxprBMp6+v1LLAWptD/4gQlRHhQ3RU/l/i1+gao0dq
TtK/N9gqPFUfDrOXoExa++3JJPHAsojb/AWgNNDhom+6RdvOVWAGx2owyxWB58Nn
OlRwoTHOzpQD/FVFuu7koxFiQSIpfYCiD0Oq2E5e0Co5q91fvcWo7DIhrmRpdcm0
PNtprygGE2ZCWEBYEGKXf0JLuy0UkkgcyJTGwMANbKeTCpNCO7tDHKEV2MzdfUAQ
NgjocXvPJx6gvew8wnzzNSn4wRv001MByfpu+bt05CMke296eLj05cWQLw5bjwio
5YG0ab/JtBmrJM+pmgVM+edSOPfk3IrbnowjftHSPcwu4aS95hICK2Cto9t93xCw
wOT6G5rtXF2CUpajXiNizDBAo+U/QatQ5jRM/eWkVv3AOGEz5HOOY69v9Hbyi1Jw
SnBGAYedencs94LnVLh0496k1o+zV+y0j/6i8QCNq9X5gExGdxHJJM45Kucf4ma9
FwDcXXmEDxjAlS9idWqRKVXbs9EKZx1sL7aWy1F6Wgoe+UbiLZwEuA8DgbdKUgBA
K32mbkdRivWw9hwSi0P/mNHrBY5wjFMWxUJpL+U5/5xyY7pfUJwUFva0ZoXdjlMh
CDyGq9NmxamZ3mYlE4cKHL+o6OMAsmuIXnf2e13NRfgZu0bC7n5fgJoV4H20ymiy
bFjNqQpL5lp/1pAooLp+3dsrzscYOs/0XCBP8B5hnowH00HN0UdzD7CdtqPJg8PX
9nZFDwcukhQzkFtZp9Nx3m3QtlbR7JienuPHd07AfgtXEDLu8+mLor9cbhq4ZdJL
El7SgbllahR7iHiDMk25IRr66hs7WvRuE/GpRXgUyEewghjYzfAgf+tGhNaJXMY6
aZD6aHueA7ypuN0baku3LeQuEiVZQSC+iztScEc6OctDZ/+KZF/dgLTT1tgZz58u
yycMEk3Mcnav2vu1qUT4wy5spbEkK2V2LP7QFisXtW969q1Q0UdKkIul8rr3yVUs
`protect END_PROTECTED