-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
0iH8V3zarBYhUfSyQHOh1wZYIVnDp7Z+rE/3+qSuuG4FCvRQwX16WwbWqFftQo9Z
Ppqs8/8PyDVpKgXhBBA6cEhWbhwaFXRjcc0GV5i0KHyhqForTmy4MWWLE6DWvi0i
MTtHhkgFzpfaqxBJ7485ogzJOM3HSlE/rvdtuNeSN/A=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 29472)
`protect data_block
HsfXtKVmkXoKrHODls9/r4w3FwVSIoE4y4cA5AyiPMlqvE/GqnTKsSM7XGNhq03I
PfcnOp3YyAwzztbrN1/sk37B8tIB0xpV+V4oOuKfV/OjWYLmU/tOuNrM3HbPLVn5
who9V2cuRLDitQcXdDZMuZsHtyVenxBLNno22S4Vm0gdrRaLO1vpXaaGaSJy8YcQ
g8wdeaA1pLish2kPJyrVh0vXKxgbkWESPDz9T7OdPSHXB7bVorW/szRNVZHG/kDH
xqSoHAf9fAkjQtg06QG09pz9w2trSW45476diW0vJMokb0vd+YETLvoeZs73+zRz
wgE5yYPg3QzwuREws63LSDjY3B1rSA1Gorc8vuA+IsJ+mQMDYeSnnCl8pQiNqC0M
AHSOdow8k30mSYml775g/4cbXIM0g8Nt7pJI0oLpHiikjvzH49IX1FmwEzAtkfTU
1kVcOHrHYTD9UAnPeTlCVj813xkf1V5hD593WtAB7BBk+aPzdfx83RMjMIvNV+L7
t1rDe7h5C9gMGuxJn8/g4RG3FVpZ5F2aDeoiJn5uUwJ/lsHBIxOwHYRj9YshPLlt
TcBkIkiI9kY0x1VHxpT6XNe68B9Z6EoEHP9/Xx1CSZLarB9BV4Zd5/96ar2lKmQj
CqaICAevaaTc37IkqaRRHXnY8uzMI64rXQuLXDnDhfLyydpVYPzjNLdOKz+gw9zD
vtRLGyRAoR6INJ9MfOHefml0SR+2olRcfVJQvubRphPgeH0U/zwVfZxxq5R8xTbm
eZ3Z5LlolrLPd2gGMIUZ9oqvQfL1C2c65XbwSy1yNNMJ3rXySe1IBA3c2FyNyzlI
CKyBC6MWzC6lnD9tGP6OYLvaDIdxMzFyMQXOwFK+LB1AvLGrB5q7QHtjI1tP6MBD
fvDB8HfdjCrpG4bKkhBl+hDLU/ugHgaNJhgOnaNysYw/BNoX4T/tKtt4+0NVq1E3
qw7CBFOmczUhUefuRmDCT+g390WfUtwRtqv19KN1YO7dctqMbsQy2ktGzE5Ry1Ez
CHfsnQSb+eKAqIHqzWg4XAVzHiDjNUtp9WgNk+zytut8EdVhvgEjvvu6NgXzUYj+
VI4RjKpyTSRgFT8qld5GyvgQiyT9hNvVyfeMxKFQZYHDOhjKaduh0y5cg7IHftQE
YCKTzb3atXU+SWPuy/46QdpSPKYyXugHWHewmM0J+sW3F9Jy9k3EGfXSugiRV01u
f1J1aUldpsResh/yP+IeRxYXNSEm7N1Y8hPZG4gXntovxKYtblaHMP/ndcSXfQ9h
ZrI6gO+ZzCxS2hlG3+rfwOxIa3Mih//LXEVHhFmar+kHUX67o6DKfJgUqBNyx3Iy
ufhV17i0p9yyOGp4bNYofErnriqnsbo9FL4UwRKe44nOlppUNlbQxhqMYVaU2Jtj
yDk9l+EPt98RDANGkzTTcD61nSz6L1/VvDL76npn2UKTxpcnntf4GdGqEOKjY3Qt
+/AfG466Px+hyWRv6h+E4ISnrp5G8LDnQ/3UCrkipY9p6zCcx2Ng5cMY7twsJT+q
k56jQyAKHlz86iWGLgEbhLKrxX1eCu6+DQnXIiVrunaTYQcJmkNJZ+2zcpfttAwx
NhWnC2BxXbEOwbAAl9047PtnNf0rJnvfVZ5mb2TUkyvqr+Go3WX0SBMDdvjIXABP
uwTXZGDThvtjGzZPcDgKm5eutaeDcYeTTpRswp7skZYiiwxfvBvz0ltHdHtbilnR
d/lqTNXCXAY3P4s0wV0a4cj0abcD3amuk9CpHKA0FoOb6MeTRsWYFf0RFTyhFOgm
NnJVm0gq4Or9Dz0gzXt/t39v22lJH8ubzjMZdTMxLJfKXz8HT/YydUOdbcwfMPsx
mEQDaWuhAJDSicsmpFXO0Xzjk+xqDrEBwWI8aOkLTlvYxEkk6KQkn1S6S/3nOEbT
HID+xhDhspJksxoaXgg46VD6f+9YdBT79Pd3fyVKFb0XvrjlvvIt4teNcSrlGxUf
DTohlStwjjuV2XYB2OqvkNmYp5otL238kLFUL/zvruhWZmEakKGFQgT0P8AA5Pzm
WyLERrBfhYfzghxvQQjFWwaYP2AwqOUg2Wpf+9ULOMkRYChGJI33C7HV7oQTHals
pIV8fBasTcJ9B1kckEC1K3Cs6IJ4LKf1fo4PC8kXe1uTtTv3zxLrhZgQ+SINRarn
1kb/zZQXjvaFouAumWt9pFX+yYchw/LLA/4c4Mn8xETN0Wn5C7XVLYv1+R0xAM9Y
N/hhIkrWIaeQOX35ExFwYDbRL+cJib0hWmNNi+UI0T8nfZMRsQuOi9VCQYUaNCyL
0e/ZmfANcE6hA/Nr3c/xYQVmQSrYVgs9EmOLnZpzt17OVsi55+vXLWG285QNsaM9
gnWM+HJcexYg+nWyr/DUJUXESza6tuOHeCBQnIPV1TBjLKXo9vh3mGC1b8P3Icjd
xYh3+0WKkhgDWrv6V1Jfq7r2xb10T6wwDy2DXCPDD6HWEZUew4GjIyhur6Ny5i3r
k8vUKIuGXsOEDCLt27A0f5BZezufRFbUPJlZV8ojjaRREYycWyzOGX1hchGMSPH/
QxHz8GZUwoMQaZFWgT8oAqM+pjA4ZF9JvZ2U/t+AzHwY+BsOHOjtiaGmopqsuyEH
mDSSfcCdTIh2eDRpuyQ+q290cFwymoKKBSJRDkDe8fUtQVkdWwm+THXisUuNp6aO
eu740wNt388FS3ls2+6xvr1wq+8hNMSy1xVIWgEivrIYRStH+2xYz8bDn4Mv26Ci
un+m9MISFMuLyfOSK7KkoS8lcz8p+pBH6HGPyGfVDzrqsJvAngzycGofYMyhCwvC
zqgSVF2vvfDJNXcmLpw3xRwYWBbjHQChsmREoD3pZvHAJ1DZ6epJgbLqud+ujh82
AtRZDUJ3S5CK7JjOmyx+/EkF78gXhnKYx69Jun76it8MUmVC97Toyd545LUqp59s
+V4qg11Wr+dEl36AJzbB5LKH0QxCpwjbTaPZtC9SM03iqIbLx4vZEvEl9tGQENPO
ZzvuXh77uwANqOpNL4UV2PuyKhQelfY316m22WMswLFnGrVtpwgILloQC2W20Ba1
NMp2tygIwLnfp/4OgxttU1PmQt3fpIFeowxf7PLkK/5LhieghPcKrlvhtgOo0yhZ
A15+At210oTfqV4bG2R8rgTiGfXiCIV6OomqzWZENsknwryxlH+1Ro7zuQbPTv4w
xIIj5gvAYSvM3zgyRcDOVrumbFZ3hcfvzvDLPmd85lNquc01RVsbKE//arJ7DQ9j
Bn/W4PNjp6OyewRfsaF7y8YVJ611FNgBKVTb1u1UbMnk4SD24dVyIXvhozbseQMB
IhTEwi8Q6Of5ND38Hi6X2srNqduZ92XA1wbcNYDM5WzOlfM4rTGMmW/7g5cfJxnd
s03Wi3DiyDh+uI90Gb4DTDvu85xbi4mtTkpMANvM7ihvneb8wWapjEWXMgvcdUwE
cQA91pWk67dLpj7UOM2Y4R40xa+ZS4BJbfMc13gOLaB5O8YdRos54m2MuNRpXIWw
/HrivAe6bolShVL6Qr+tmg91Sopv+PrpVQDnO74Oh2WsAQVV+w95TViO3DsEOsun
PUfbyZIzS5/UeLA2p+ngQCrlUhHtB63i/aMdBfsEmz1r/bI+LxVWax6IXBcK0Oh4
bqyqZhuxNEWDuvty8hOvF6LSV7DbDsXfjFsw8zSas8RCmFDDL6ESrkt5cwHiXuin
+CX1EJm8BSR8uUa+okODeuKVpM6BhGc6ex4ripKDY2kMFIczIVYZyc7/so3YhISh
hPEQ5fKY3b3d62H3G2DqMTHwppGzKuX9+UVNrA3LO4uLYnC9aUSrHBj8ddnBaW2o
iSxmzh12qCe4IvbfaMElRttvjvSKsE4f/ARYnlrsC5rVy0qmle1GHfUyfFrxadpS
bXynvh8j8/xLYRJ33MzzbBi0tH8uxAkUZRBJktUGplKLQMfhyKQGnw6yLQQpSeLm
oteioq7UNKytEtLDwWwE3VtgQ2iUNt6JyKeIX2iZ6FZ7ODUGTWGWPA5JdxmrbAT0
UzvygLOq120BQsg+R/dZ/dcboIgUgHVbDO7ju9ermHfo/v0yqDzCXVvifmL5auqL
sdv9IHajnlTR+tC45+29kYLmfFvQkklNQB2u5DBHcAgjgfnqynzydK7EdTxzPDE9
se4RERIkzNco4+9VURSAjdqLY2GVibN5FMTt/s5kapqKpb5BksGG4uQBlv4jydu0
BCAr2vFhxtqcwaZujIVkjll3ZD46PIunAw98+ak4pLiPqGhcDEb3HaoJIlCOFjCO
KV5og28lqLrH3VPY0tXodJhUjBWP79vDE61vKWfiL1gVxIPyJtCrAscGvawVFEu2
hZNh55gYwnR03Y5WPAeiKMeEZtZTsdZl0thxRMOWYHUgGqUuoQTMmLtwu+NPZNf3
wDbAp1d060PR2Ubk4dtF8U+MrBfcs4MgBgsOjed1mL3WaxG6VtlYTnLPhLic+zkF
VpgHtAFr3h8lrvNv9Z9ZWmGhYRSkaQTcpAamUV5+2rLFt6fvNwMtL8MUroWOmGTU
jbhFaf9HnxsvvsVn9M7nqrOUK0mlVZLOKeDDxlPWlMcJOGd/cWDI/UMh808TdszN
l+2HQAOHbbz5Jo901VhQKdzuz+aYpAt4+AMIPT4Wxkx/FBBixhAydDoU+z+Unnaw
fU9LIqcQYBW402wJuQF+3ndPdv6FDDf6HVsY26n5apshpJWFGKk1DDw37K+mkeEO
70MJZhcvi2HkwurUpu3ssZkgnkQCAJISt/O8svs3Y9yCt57HDonfISsxjoOgmSx9
KHrU52TiTAk3g5O1JFZk7Zxxr2j8agOHn6BZtwqzzpY+vcx+bfdpK3P8qWdfLNJW
Wd6yU/dp1uoBqkC/9FU+9RMtBnyoX7ngtdSCZ1pxOGNaowjxJIMdg7SLn8go7qBG
34Lf7neeCBEXW9HMnlso6UQOedpp32DeSYf9MSFT3d/HipDQShxaH4IoxO1+OnL9
0C+h7R0cVJV9PcHeOv7k4S3UK8uqPwgcDIbQUAkRvOqfP4T+TX15fPag5UQw0FPl
OHNFSmu55sPu9Fk64XcG23A77FlSXeQk6n/+25n9W3SXnBrjjUb8boNXb3n8Jd3A
7i4Qhp0GgN2SLWywY9M83FkN9n7ls0qVxd7lmmXJ2nTNxGNGoI9r+eeLHplF1R/T
MUIlXqJaQ22XNH5rAkEQCFUDv/Xlf0eeKHqGSOpWZdTqApg8Z2wCD5fgDndMd0O/
8FcmaS8YRzrPWGwZZroOPmBtxocc+EsmloE1TdDEk9oVt85AHZ3X1w3V9zTU/SND
lfH14MGSOaKaTIqYjFamxJh3a8sLrl88BSXDpw2pR3qIEGbe/6y9zEx+Ys0OWW/j
IldVqD7f1wSskbWwbIhb0hcirKfewlXSvhtoe4lc5KkIavCZm2uYSslW5kFKQp6b
m+oLjTl36HCRdgV4EhBU9cIykosTcJoCMrRWCyWG4hVs6pzJzj1x7JuXilAVKqYE
8e8tAOotAXNJOczdTocsyAHTZxL5+z+V6BmnmbTYipeD24o99Cpi12O91ZuT+BTB
9Gef9OlqGBnJNluWc9yHOcK8Vr4YikneoSlaDlzVTqen2gNQwBdyL7PPMckjzySj
gPbE4NAJwpHQVAOD35a/XF6ZwNotuAn7Is0BZbu5ITCUlCLOzZbTJ+hRp0xA2z/v
7rO80+RZuD7PBpueWL4NRLlOajrdtNCM9086TZn+XTRS1yixvqWrNB0A3VHbX21r
jI8OweyH2NNvKp84yo+jXQz0IKCK+EM4CXDy1nb/bymhwWbfMjOthOmBxgLbKBsS
il7LkkJ3CjpkmIziywyMYnpNJ6ZrowKvTnyW9uA0/dQCxSgRyhvGvWMZlI7DqwhI
4OYkrmf9BS9uGqZAqXax+KB4ZOMIQ2mYLNb9JODf+v9hxWuGgyHnRF9E/ud/5bJX
54QawQvoN+X07+gX6Dpf+vMZd2HmTnq58lqKY2EhuQYqdfVOuFQsSXuA9Dc7Y7Ec
T2VBJ+AorFJRn3SckXu6L1dIHnB+fc6RA0j8X7bR++Jb2RhiWxZOz8xzTERe7goG
bSU6cIKGSc3jV+omVOERnmYqc8NP7jYjVGYm9mOTQiYM0p9lGgkYvYeJztBHzI7Z
j0gz9lwLY6gfK792hhpGveuWVl5obMRM1ljZSI+0mV4UcYOBqO95pBk41x3ovhmx
0n9U3PQSzIxmzRQhpgXAmUqZJkQpgWu8DyDJ9ptHClPEU+K9Sftb/0fd0mHAilTC
/KKZxhY7hK47Pvuhuxgw+nODY/OI8UlHS6zKOmsOgshZ9keVIIuyAOH0pfNRpoNA
FqPDgCJkFBTiD85xpyHFPVxdh26vbFcN42decYvQ/z7BdoqXp6dNYhvg3mdgin5W
bhkReOS8cgqeAVV95Ww+O9Q+l8sa+qQUgNtepii7YC+VqPzwDbV4CpWGwRB/jEac
utKgSjuMtsj602SMpiAwdaLcIYeHb7Ar8cWH1dgIts10TC5LEuTG9CzqsdLqg3xR
Oa5T3GjfBOLGljt24X87PLMyndGHJQmkVmUTxdpuc14Eww/ko1adGqziE7ElMq/c
J57GUkMY654OC9H7Ms9UqR+NXELL/G7RstLZeK9QRNMXImozlgKqJ93oSYVV+hWc
a1aLvADgp8MVbAV2943IKQlia1eYCCxg6ko7vpVy4TVRCLCdX/xPkmGKkMeltNcR
7DBjBtR1EfTL8t6r4LTgz4gWMeXyTEN+56UvNjxDviXeqhWfopJwa1q6v5Idv8Cv
ERUMHFSbA5PjRgq8S18b/mRFvRLDYcusA+EmQKYWIFZ4F7L734ov3SBEMI1mkF9Y
DUUKNe/EdYP3cTbssjn/IJjr981z2dr8yAScL4Qw3uwK9Tu1+H0U2MI2rdvXgKRZ
S03nb0LnyjzMkBpgh3IYaFo0mhNGV1CqWuPNnr+4pYnxfQp8iJlrfCbSmZnrqK3o
CZm5vqrKkrEylxFPIy6QZAdOJszmSixeo/fBB5XIunMtaUA0rzcz9zk4/Fohl+Zm
uhMuPcqo4W1UiU9ja9wuOgTYWP/xDK3pqbPFC3WN5UFij3XLzJqa/RANqbYlj3UB
Jum3+T1RBPreBjFMCCFrimUY/iL39xo4DnKDqD8i05qOVBkDdXWCXwHvCThjz8Xv
dA/zssklJAi/9YoUMGl4ZXPVekn3hS2QirQ788VZUYx3zuDvvp58UssmAj5R89hb
oA+ZQ6aNpvsWe16ecPxlvMyC5e8qXAMWBfaUTzAeoVIIn+BemBHOE42Na/IvMESO
qrfytpxD/H78E14MbSM3TjNpQ31XhzvP2zblItCEhZI5fu7tPLoxhfkagH1hebfP
HEy6MKigiJwsI7xdffvd5vs7hQ3soDzpWUUPt7xnS16d8xNr2Aljn2XTadX3+fP8
gCWHEpH4Ge0RYSwRiAHG2PkEdfuF8U+2qft4zsJ/T4CzbcaAy31YF0X1uyiAMHxk
auiHX5aM3cu04qvfZ47JgxUbRfqYM4CYapdhYiUSjR6MhE2d28s6FaAOF4jTLlQb
FxLYZx9B/XD+PN/3QjsmnFJ0UBB1h2eo5XK3wvijXjG56ZWKbA97Lu3sKZRQ124E
hHVuHSe5xyQEgUcS0tH0IOuoDvQxjmNNuALRs5WBE5bl1SM40/OkAVLvVrlcWHo+
BbKnyV9E4hwkRp+5YYTwQkUtI5Xs7TW3rAn31PxpObjK7iF0axhhppoDzRVHQI85
V0+VpnjoL0rwwSTdX0gkoBILKjMLQw/aOGC9puAlo0w8szzpsnOxO6u6D5ZqYC5K
rP3yAaa0j+/KH7/MpGuTHrHXqaSY2qXDdyMxNRacKd7933bn/9mhgBUMrKxeyOtU
+pHmLagXtqfls47E7sZSkOk35FZMWOp3IuVw5SC+5F47B4pJVMqL9sEtA5oSa8CI
260qM1TvOd8o4kuWUMI2ptACI1bWdOUAU8GqOsInk63t/QDd7ybv3Z1W7wLETdDQ
7MMhOSf0KOA57IsJ9rmRXMLDsE7q2WVairVlZg7Kou+UF+b6wSYXPwUaoPzJ0evU
rGrRqPG3mzZ3msseTcf0mxMS5OdDctiruUWz4Ec47V+3LHlG9l/5zfHam0EjP9wK
iu22pC8ZiWwvFRmydUJSeXSKrBP05BYnDu4ZJYkYjQB++w2k2fDkwDj7w05AI5ty
JWTV9OwzTg2I4y7iTKaZoy5kQ4d073gy9mmH8OJeLNhnuhiU8HphzSZ73rz0/l+Z
076V5Nvx1QmNUSXMcdEIL3b4QKtlDGF3x96ZAJUBCXDWXzOXcQZJF14YTP2jP5ch
nX10rmwfQ7rLu6oLFk62uJJHMJgIvi853SwVQ5r5eIVakaoKZuyMNDeZ7OpbSITZ
oyYIZy97KsTgKkR8BzuBT6eLcbCtAcPl+7T71zjbbw++J9+d5xPqhTfRt0oeVfF+
tCsgAGyQUymLQpED65GkS6xFL0hZ/VIplozWFmgx8CQcRB2tslzyQNHMfoUQK0L1
Gt/TN+A6P19kP8UL3yanuSnf61lCEsjrai9ASsy5LrwAvmVCLMsq5/yJX/tl2ehM
tdd18XMbHUDXOVVRVKNjuSjRIqGluF4MlaHFZl6Smh23DIe0D9kkaGdrhr2IDrN/
kMEbuS5AzPq2Qf5hLN8ymXb6pM17COE81cHPfd07rIjGMGwLmXXrqpRbKNp4JCVi
Uq/FYZqmr3Cj45M5QkEGzAcvy4qBEOu+ceHdI6LVmwTPvgPVIn6e6dBsVxLswWpT
x4DT4u93EJBH1rLxf4aoQusiZ28h8kL9lPHoQb/P2PZLSwIr+3wNUbt3JBZeQ9gt
Gq1NdbUmLOR5MnC/nia1aScPcWaXNzU1/i0ay8AhRN6+v3b8QFJD3qy73q2wvDym
5Tx6Hbp+hRREtYQy55zFDInvXwGGKcdXtocYQRcg1cGonflyBK8nk1R/Qwa+Ftls
cpJ5yMVPzXcjHCXLoovNNCVgW0xuZnYoIRDIcrATF78GLGKNKYqUVbArCUIPV5EI
RKidYeqErLGLqq+x4NVVTC8EuOgR+ahWQkhgZ/Jnpfso1tGN4vgKi5NS9Ib8zqPy
XV4QFRu8BO7EJXcj4kS430u7eT8w5oNQoGmHwhxKVopBiqbwFFnfVMLLCIwtvVej
jDRoqxNjvjetIr2nfT735fOYARJld6rhSGPaNnN6eUnrq/OQABxZ63clctvFD3ry
IfNbMHvzop+oCu+0NFAa2kw67gyY6EfvbrQbfnqhF0HAAwqka1PkvapZIA7AYPpg
diIaI7EMBsweTfVe6Nm6v/FPZ7eCkbdVTdOn3Yp8ABZYpFuiJEIpHbz6edV8OTfM
Rtv5jJWXR0PyEWTdTpyiu0fyr2WCGMazIy0KqNiS0/qHsaLw+S2Xpy70Txj8Pjm0
HjXePRITxo/EgZqWdp+TBbrtVVoqd9O5RE2van+0f/M743E67ZvWr1Omsy17WdFP
arxnjUBeAzbhdMF8awBaFsuv0uadF8FrNQF95V2SbxJYomTROgZ57gN7PMz8PGZ1
aI6IsIXNRpZb/349pQgPwjowSSanGpk20iuyz0wr1IGfYzsYPtrLdPb3PwUuxlWb
yFutyDose/6CoN5cBo0dA2Otno2bn4cZfIUq5LO/OTQKSy03tLx3rSXHvxJZZsro
cKbSsMwFvQ+srOljLfmysLLYE/TCcSOkDg/24ZdnIY6bXH94jJEQd0BlII+goeRb
XdXpt63tIXks2zaQRe4J0Ev6fMMjXLiygOsPylJ3HTNqZzk48gFGgPxEaOknFOZc
PPLc/gopU2NwWFx9ltOV72f6cVhHl4xFcCcNbMYJLttWyzEs3H9AdjhGjD9XdZlK
y9JbTyMm0sMRqhvc+9uh7TI7ibC3AXuG3D07DTVEgTjxq/P+RqZ2Zm66z/swMT7I
Pvc6RSDWmwpGHyjY0vtuqxezEa1ygv+aDiSauXGSfomXHVfTPU6Gyu8P3fzrqK6p
++vh4bHd+i0gkvU38hbSqq+2q+YKcIJrWO/U+POi0lxST8CpQlQBvkBXj5j7f7+a
a+ndsVGaN4ftzP/mktBwvzCBQXjsKjcofgvNGhHj9ipNNj+ddrGkrTLWWoMvaQRD
nYOrhBp+Gd0ae6YljhZsTkszQ4O/RKbqh8sFk/WXjTQwFxJWFrmm/EvPLq6Tp8Vz
J5XQ5cyRulZZBye3sKqVJUxoowVuRJUtlSuV4WS0oAZWPhzKJNl2jZ6+v0m28/pN
7y6iE90euUWPMRj16XeXqcFsrQkKwDuscrfIUnimEgvtirnwK0w+sp4xs3l7vzcL
m5oTREnZpaYtOd5gVwgvsUrOTe7SwHR9YJ+l7v+P/BW4p0lF3izjTOvlbY0Xx2lc
r9tgEhDoaLKV1Rr1dvh77gyCOX9fr/i4ED19lWPg45BUnRsjNzVmxtmMMyikn5zN
aexv8keWaDbdnUyb4DAqFlzTbD8WUjQqs0pHM4yLvCjXqaxjTyTb0lHDbZhhUwyu
A5mVitgrxXaiYJPHGa0dNfEPDt706bVXCiY12MFX1nZ49xGT17Dsfi/AJeCZf/Ns
5udg+X3X6yGXaM44UP1wOzqAhaC/zGpnoHFfHFiDUXSE5GHXQyE9lUohThHop1IN
4vs7IX2RvZRV7QRgvPM2KC+FcZj+cjI1juFpCsvl6pbDLalZ/FHgtdZaxcPJRVH1
DWXREPtna/V6Ty0Yehh8grOhj2BcykK7FeQCZNuG84nMVoiRT+a3nedHNLbQfl2+
nZguvnXQ+T9azg+uey8m+djLi8PvGcstPgnw7rjnxlWldqaWmToUZzwTXicVULrL
/fuFpS020F7Hs1iS7juwTToaZdwOpJj4DpRe7abSBRUcdX2FOSepx88C4Gb2dd/j
oBnDG5kokJd9uNt8rEOvYzJ7ue3FUOCwtBd0tvcwHGQIxNTlCy4le8ajIn1BkstR
D4PnA4pBwD6X3f8WwO62u69mzWYyHfos0P++pUwagrs0EUHCIr1s+YMoaMG/aZFR
CS2rRrrjwjHczniDHu9XNt4KmWPRZGKVXk8rvKJK+VXOltMwc+ENvI1h6IA5yEVR
/NJaxcGHSSBNPqRl41eKYqP4AnYR5oXQiwHW9l1B7RyuRgDjjDbJfIuM5M1zKTOX
CzzYrQFJfe6FDHLJVcdw/+YeP3FQfowSw1qxsGmzQYlrJmIEYZ0JwCyvd/RBPiZG
MJ7fyc19uzpxUg5S87Qzh0d17Zdm8uKyzvRZ5zF5oQ19L0im4+0gJOZt0KvCm/Mz
zrir71OCW89hAaHCI4E6vHKd33jjOdxYGubwhHbFn9uk3+y1p1YmVryvWBobjPoA
NwoL6Z4DX8/Qbhdu1PqBx3ewD+pYx7Sl1ZFxY3E16qCl1x4muCzYpKqWKEXxnHsx
p+WLHK68GArvuWetfDpVCI4pruvwV7HRC+fUNJ7wA/Zi4x9z/5xgNmGXPoHENZyt
UmUHFckuEeMTisIR0Yc5zV309Bc5BHal0ZqhVrqY4uTP8t84EhoNKZRK9LMCUzh+
KstjacMoR0VE2JvSkQmUxG2CZtEi1yPl080KWA5Xtai1xOS2RVAhHD5h8kIxbRg1
qBA0SAN5mVrGgUJ0apMmRFANSBxOoBitGel79HhLCuobH2qiD3gb8CakfQ80l4Qe
DeK1uzmaOlOZR60+LWVuiZ3u6kjPxttEL+Q600HZHtY0RvEO0rINnm5g44lrEvL7
/MqolTGTiAJiUWdYuX7ejYM3nNQpgLJJM+jBugPvsl14TuAVI9wp8T9DmlNoneIV
FVEoagpfFMZljbjAZKuRMzOQz8rh3XpwbYcD+3yFrAdF7jLoJCL3DfFy1vusmfCK
w6s36rm3wQj2ZoBuVI5FfMDqkaF3PSMuhnUe39fSMn0m6Vzqn46MO1cA20F8DqJK
pf2bqtO1vD7dpqoomz5O/PyNLBgnqnf3ysEbSAI65xaEjzy/pRZucRIZEBKs7JWp
g6BENdfhR3Yttjc8WYcO0IOqDkRoXsoRXyYW18skmXTa+7RNGXt61Sw8x6NL55G6
GsYAeMBB9hJvzZFuDSnDXz7s3LlgopweqnuonbrZRHcs1p+FNWu2JVcBU260rwhg
ZygT4wOBgmStKLqc9SJM/KLAT8aS4CSXg+3wVtwY+PgkiDb56I8POWCmb20i9Xjl
OTa5SLAX97vQMZZrY5Ynq69JVShTzQYe7lFDrLV0p3MD8PftvQcVvTa7GbzF7wwe
oEXEShftOr2lFkucAuuRImxdqPyismizr3XE8RShl3kv8wYm0YO+q0vJqz2mpV0/
nyV0jz8oL53n4M+fLSIIaHxKvGn6AflTLN9qBe1yzd3Et+5mozkHEl7k6/zO/+BV
JuzSi3BBWEWJlHMZ4nb8y4QiBaQUug0ZPeizrOoH5jnVHqYgTWb4oIxLiFeAGqMH
64l6oIpTME9YJlaCVOVHP0wKFHj6Osnv72lXDUXW73NdZ9h2Qe2k+LnWAXU7c+4t
fIFNc4+zIBYY6EXPwytNK/7hhijvGhdoldLqEj/I5MZpDHeIN0tp4WXaAuJHzbXR
LH5ZljgOhqUMmztCtDMEGrV+4xPeLTlZHvoVZxXBwE0oZ3rYyMI5u3B60ufqqegU
ap4rDtMCG7HRoZfZ8ZYxc1P1KI3C78oqmdVXYD4TI/ywYX5tMBUSH3mFM+lOskQU
YLerl3E/JdNFLvV+NY5mLyhS7H5zGnb6wwbrQ8Bb4QXPEdLl2osLCsA+S9qqFYZn
6eRc3JcHAEiNZstFVd3wNWEUbEOiRYEUuQYJ3KM2aA1q6wgXOE5f60nrdWIiGYYc
j/S/Uc/VRek6XNsfIwlXqHz7SNUqNZODAsLgIPb6pATuNFhv5BDHD7LxxVj0c5Nz
toEsr4ZTy4GYuf4iJst4pZE9Y4DI/x0ikWAMKm3R3vsyTLn9YmkjFuSO0NXcV5oo
k/z62iCjv1zxcECOlIu+VCdlaBqnRW2B6IQeu7QJn5ydwGR/A7u1j9xMsLYs2nW2
t697GNwWHp2u09RYyGxgG+AVnKGs1Y7M850x23Ix1VAlKQI+/OI+KHSyhmBElbaM
1MsnQr9QwBJQMD8A2c8pyXxR7aKk/pRKOkYNlxMKxxeXkIJjTIRRUJuS7RXtmoc7
z4a2vkUp2QfxoblZaviaufLjPUGrV38n2SaW7duStR/COl5LCo9937fT3wBvr3F3
LfcQ9P32bZITLHeXy2z1RcjtMtiygZULFNypLW/ToDJEMCLhcSYtUYzJtubYjeL5
8jfgjgf4GuXDB9DljGJlR3Ca34QbaVZYTxFsmvLjeIEv+m6hsyGmrMB29JwicjPH
WJDg/Jx4loIAdtRPcmrYKmDIHrGfA2rYm1CSnTNkQKL3aCfU8lkBAKOhaP7HCBoV
qCeC2q+c0sww4CL5L8c8ttNL/KDo/mvLkr+qfP+PIFnC3YXcmbOcM36mBmjOG4Ze
H6+Sgq2f6ZWXYQgfSAf2hI0u0x9oBxRtxBnpLheBoIfyE81TT4Lsuh3UHj+pxcCw
l+puXsZjxpqnX04J0Ww2yvFy8dlaMqcW6wnUXQ48kFTN3E+JuTwa+aIp7nN1rWoD
JilfQ5boLX87DAjM2qGyutAoB6GfmXUNyyTKBhe2QG1exWWfJnyIqASYh2q4wwJ9
fmKFEGqQ71yvfY5JkQPIvnFIRP/IRBvMJNnhoIei7Pg+aLBhJt5kK7RfNddlLZtD
xRrDfV4t110doV8AlixLLlSFels53CCdNafyv3rL8zsUz18j+lKoAl391dRUVTFn
5oDuVJvcK6DU6VSWc7EXYyU71R0Iyk62hTZpcpGqDn2I+Sc+Alioi9Cug4RDTzwm
dDv1C061Y5vytWdGgBjlwUyTg7zxXIuTux1rWG2W01f+e7SGFK0bhTbYZfwiVO/r
vj3r8xkJZLro0m3656KDqQBxkkg6E4b8BYoyc/MhnflrO0VY3lVlMKwCDrG+Oic5
8jGRBg8BuL9DE9P03Gcs6lJHotS5+fGCo+UayhvMXxV3Z7RzIC4pm7hcLoWuFYb3
a98ASTEPnofE8s4OSVhPGS0atqki2s/s4DzcyzdTUw6o7pP8np73ow0UfCBZItW+
LvcdwjSaFDd3q9kBxHpT7RjeQIRE/JcsGqHfY3zAPkoIFeIraEG8GB92/c/HB0xb
hy/S9BrsGZT6AqzPLTsy11j4QdryWg6w5YslAk9PuYprbO/5DzlWBY5uwczg7NOI
L1oFqSqyjBm+RSilBGqlCNiqEagm6+TUNNOmcTSRENZJk6oMBmTdRxHLNeGtAxF6
w1SHUFZS+IZLTzVQGAg4bFKgUV0LBCRo0ftnqw+AQgz95N2E2cvgPIMadAAeaEv1
sFTULx030pbVS71nos7vTcxkVa7OYkpxK7kWuOpjuZ2BmOXJGexaxyvWC/Mxdxis
l8oaqSue0NywFbn4hEsGkdpqucYBqDVBO9xJ3AFuY6irQMnlD4NqT9DxbNZJKhD/
7wdapU9X84gBaA6cwxy2VasSak3s3mf9C29TiavrCjdW8xgHdl6/r4tT1JlpODdj
A8N7qo9IzM9U/ML6t1JlxqWhHN7l3PgHa8acBWf1ChUGQOzszApFMjAM82mNXQrZ
68pk4TrRJEhFoDg1/MUXhGv5Ym/92UfDb+jHWDdziRehRx55VS9U2lsap3BeClMy
rZSByR8+5Z1OK3GN8B9+NDkw0j3wHiveYsBgaqUwm9ON2+xZ7yMZHlI9at673Ovz
87zpvIz4w7bMZb7e7eVth4GDPhb0ENiTh7DOqW7tS4ugP/r4Jgr2Z1Cpg1eQXjux
aUknyTWmmrn4+JekOodTq6gCxdNrggEz09tCCc9Pwud+U2ZZkK0xZ7AAb0vcVUoW
oa+MIiL8K7CvyoX1a/g9wtag9TZGvaGl92/dMmcR2cr7VUuWnlAIXdoNN8fzrH3y
nYY9dWbwOy7PItyW25LeE5BSIWdEW2u9lFIHIz9hEamqlU4R9zOoWcH4qlzXbAe5
EsH7r3bp03Vqdc+KoKdYLug7Tb9NBEOaEjFgMl6IKMonKDZrCvCdEb5sVrihWPXK
oVXY3ZO8OwBeOiDHapMrMIURgbj3T4l88oUKUzAAAC9ZfNAx3GLySZu0KH2JgojD
qk3qJqIktCRpDhDx3Bm8dTc3qZc1NNn0IpegBKBFZVV1oZ54Y7JjbPHcmrV5Ibht
Y2HKpL8HLhEI1hzhuCJWKe7VtzqTmzC/81Lq8VrXNm8/9Z/6G3GWcx5DhR/zC5f/
HmaxNgjhV8xx021E8bTYnR8LuO7TztgZKaUCaLwfRalyYNu8Y0A7s6sA9RS4zrKk
CoHNYdeplz1mVSguKjDhhQ6qE1ilWyfus4/K60lx73ux2sKgLoNqNRsqHkJqD9cj
0dTNJEJeNj4GXKZ8rRfF9xJOLhUUwHqpKHRlGpmrs5jt6oUmGxrcoLKDAnwcMdi5
FkfF4Krsc+L4bFB05zl0Sp2p2I1JNKPHJ+GrzthIROV2RUcbp+MJvfiu7xsEo8oV
smAtTLOuKI7WM/lrgxGFu0/uFgUflNFxospdX3JVeZz8Ma0OjGAkqF//594USht8
1KJn7+pvTos4EqUPH43v5NDb/j+CUyiWQnOS8wkWxUdsXM53/YeuCWJIV8rvloNw
ZFgLHiHypJqBx5CFTqSWhvab90xl8l64iTw3GEKGxCo6S9NC7B5lgFejHLGeP3+j
4iXfFu6X9WOV7FoReZSrseR5QtBDJ+29DLtM6Rj0//ovhkYc+1qL6TeRzqX3Wgky
E4UITROftgBSduEmA6zc7o4BSDZnuzTLFvEEQs/VLx3p0onr3RRP3ZFTcOYmjbbM
+yQZu4y3iqXR92mf7g75thuGB1pIsFJ0sIEUpmLsRX88SDczXqcBO5xOg2CtFK7l
v/tkxUkte+SYxoU3k+LaO/BqtHbmZL/KWSFB7Y3cD9hdpsovVFyM0XvkZS1zFFiw
rqw/5X4fXxvu5AmXhpylRC7bIodKQ4rUEhm3YToshV366nTiJfNb4bg43pHQTuP7
n8ksQTvjtm8IAp+YRlh4fszrUPQG8xyoFKNEaeSGOhv5vQeD2Mx/YynCEputYE08
jEobN/QBiMP5lrRRO5j5w2iYcz7cSHeedoevNU90i/w90MyyhrKS8kmQn199cOS7
nNzFfqpT+KoZUx6kC7oTdl/zZhZkfhwZryD4rlc+y8tX0M0hVoIDV6xsE1IP+uBK
XUBCvu+87Xn6H+X93GU17LCtA7P24hZd6Eal+3Kwn9ctgqvu234jRZaLVuG+gcG6
dMjHEByCn13SJ9kkyTHIwR+0Uk87H83m+519OuFufHpo87APq8fups9tv4mpjkZ3
J+lGGR/hfBgZX2kUWsvTwIop92d4cf1oHMUoyg5OJsNaE4SnnP4ED583Q01th044
uKWBaH+Z0qUsO8xcDTx4573bJrRPV6YQzzLhZfgR3+Jq9OtWeCZhUY9gLsFcNXkz
EVB/hvNg4LTQg05LjUjsiQX5c0i/niJcGCTb7eoRSbClknX2/WwTSFBdkNCY7s8G
AknPISk0GUCC03Cp2oCahi9XolAZget6BwXwLGA553O5q7vP6nByAv3IPy6aifmi
CDPU8pl/xwHpbhpoGIUV5lge6EexODy/6OgE7dLFg3MNzGcsDByVhKLQoxm+PXtF
ZZwp0cYUhFJZk8JyYA/FLBaWMuZLNJ1zXND38Chv0C0L/eh+QIOUs7teACfEaekW
/NFHFqEbaab95aoEu0DF9SFrSAAI08rHTxHiV4aR5zIPlntOhehK/wOFzYTxqGl5
3ZNPdPQClZ+jJHKVqfRbB5AbLtezZqkK1A/RjxNvRQQjVESekcqFC8/hF4awVTp2
B2UcqZqQaYizdkzATl36B7iapTyeTwRZwQUSQEQgct/0lI5mSwiycenBSVQ2q9XN
lVwP51HD7kWs3lWxWbZiv3gF4o0U0EwRcr0lcRuVxe/LGn923V7k3A1TcPZG76f7
xs+FsY3y3usRQj59lRAVozLviO8sFUxqYsp7n3GCXkJWTeui6CAZTRfeb2GVcCrL
7A93tmZltVq3jTrZjfN3Rac/qjZD1PTHCrxgkgX05TVPCA1vOHxbGMRoqYNxcN0m
K34bHLhX1EolpOvvnhtd0dwCxaCWKnDuf+mG7xFqAREJ8J2IVTgReug+2WW87+Ft
fN8Ztb5lhDch0Q64WvYyG6Ass6Ew3JKbVIvQzKs3tpqL1FDgmVQVm9aIhx+QPoQ8
r31Qs5fNjKDa4psUcMUSyLNweAtrPzHPmkcnvxr/S3XzSv3rJ9ER0F21y7A6oT5A
JxO7AAownLXCa0opG4sAkklwbqRkQqvlhCjg/UutbZv65K/POVDDtBwiSA8e7Z2E
rXdTWovZKhNNDRARHRfBx5ANldETrRUOXCXSFbZPArB9ckvfEZy/fq1IonWbBxue
t5jPhCYh3gpQ18Nu7uZqoLDLYAJOraiKgOv90k/khrILLLH9tx6gVgqqcM4HbVxU
YE8j120zTSYs7/sYhfCoyDQ8f5lfCaHfoaVXy0KR0g+l6rEySjC+Yu9DHifKUsZI
dwO1SoK0cM+utZ35fxxEJvZUz7NMoat9rcK4xkA+ml6T1jHXAkTmEMAShcde83e/
t6K2gbsZb7OZxJI62Nm0kjzZCzQsHe/eU/V6C72pMCo1pp/P8UVmkWI09NYinl8B
BHD+3/QockqXzssnFlYNVjnqW50oIekjUCR/SXjKYnN670dzUQSKAbt1VoHALe6f
LdQxsKa2YDaQ2GEaMkZHVrucFNsEpiYZdZM/B6p9iCLqUEBrbUpyIgxbosr1G1tK
IobIe5v3wHlz0DSLVGGxd9R8aIjQv9Lg+YahyXlcKU83OpjrGi9OCQbJU+H4Iwie
wqGxxvy9fBhlQW8PiTHNMNP1Fg97JoDsKxpTdtGDx2SH4i5I16oF0nSqtT9AjEod
1qYYPCm1SoaUfMlgC4c5YkW9ZejX5nUCPEbgJfIkjQuFRs4qHo4bNGc5Ys2JAtFQ
SIceu9WmS9BV0e+P30tsUl3UqzVODWaci0nlluFS3Y/GHyGeMYc9TF3Z9ubHdIbO
6b3LJnDPjmpT8bP69KWkmCJUtjawjyXUCOsSo4YnrwCVWNdpHhm9OYD1Wadsl7l6
OCYor2NkEKBOdlx2elczo7QEdyM0wpw4yw8s5vH9DDx8+Sb6BUIIt6jMY/4TKpD2
w7ik3i9F2pUf6CQCOwIIRsRBld3AAOOZU25rk5+n/g65qKnUtqRjl9fmKsd96KsF
wlPlm4229c95J19pq49+WSgWCfssL9UlfRIWK1+oJxEBTKqIZBFSWY5AToTR8JUZ
N4wtwyr2Fvrx7JbbNd5m3HKLFHdqHRE8nw3gpR30WcvUq3++nMONc/KriJruWk7c
SHMsv9O3LDNVdiGNBUHb8g+p8tADTNZa/2q2FKEB49sFn6Cu3ulVHWVsIEAkTHek
xg7nyFkid/V2hcyTmDhDHVB68V/dyzlEDo4soyocIeXJF+HSVWR+3dWRKCsmtAlV
DkX526KiC56JJUKpMMHvVvw5BqNG4rY6YKfb6Kmi+/bram0McbnsgSe7FNpvewyD
XuGTe22iuQvw35rFoQdrB29+p2R+Ndawb9XVFysQVfyHENxmi88RtOs2ZZkyl0F4
PQF3OD77pbj1ZgF0ESWMI+n4FUGtKQ709aZMNT1BWCAo844mcNHqy59ubZ0xe+fu
oAoVLFLHIcWnpDIhYj0BfVz/idHm47O7tWFp4+8oH70pqjJrzNjyVx1MqtXL+Hiw
09p3lIPUEgZaGyU2crSe9G8GR48aej0twwRF9RAyTPBI0AVlWRf+s+vMp4jvB8ZK
q6URiojwkpHCsiUfVjb4nNOT9iPaQirlEellH/IC9V/oKYlshUZQnlJ/eD6qRO4r
FGPiK/vrLy678jjDIDif6gPop3kZrqrOZLWEMXlki57+L6xllFartnX5+NsrxUX+
4E2kw1xRNeAW6apK2BH4w/LutYMnnMBdqTZwFKBJ6uvFpFlS9UVG+GsZORwyJK0g
4pqpHiJX+wQbpZDpibSi4Ud2kZJ71mnyY/gmBJtOlsbI3dly2FdcnV9dyM/ffcjO
hoqDxltImUxccf2V3Z8HC7pIwKUxg/uzdx2w6A2/gT+riMozOE717eZ+9NI+LEWx
mcZSSjDEEKyloQkPtnDr69CfFej/OuqVLum5o7Bvh/rdF0CDj4zEm++cBk3r41yN
zEr3Xmfxvr1lyPgwBivuyiG9pTLFDwVqJ5t57aIdKCDiX1F0+/+5aQLDipDPvf0m
/rHZwY32HL1M67nPrTYvbAGI5/KKVAyRm7+YqTYpjVS/pqX4cUuqXr1DoP9R/1en
jHv+c60ROeqmwVChbbSqrQdMkEHTWwaWs/nZIeTJCl8iFOG0Hlc0x5ft+GRRqFuB
HVz6Zai94vF8s51x7YVDG5xakV881G2sxCn0ot0udBo9wr0ILqPYNQk1vgbtLsZP
RL3WPAqy6PxqLpRD/i2LH5CYIVix2jtpLPgE3LtAyZbf0ld6eodBNNHxECAmyMWd
GLeOKrLXpumasXpOJk0L2cBU7MqRP7izrdIwb+9c8Ao310n6ZoI3ejkgKDMjLzmF
gTuY2gXBK4oXVVefULoirTWxLL92JJjzbFopF46uHG4Dhuf2NTq1Un7Y/rv/8xnC
TUiLTmJxs2a+BbicFxH3n0kS/F3QNff7yBEkHz4brooCb3fjeklvlMRQMeoqkW+1
2Oe5vRHveCVXqUGq6JtUQ3hZm73ikEv7tr9amzLyw64jylHkQYtl2VGYuA4y4tKY
JSA1blu+H7j2e+uM7+27DoKK2iVktUaz93fpJ68IWGCQhrnB1KibU85amPr9rWv4
MWaKlrTeZ73J7OtMFAVPbipDTFFmm3RDTFbEYpK/0qokPXBCVcrlft1w/87IjhPT
TVpTgOtKtVhq4Q0YmqS3TNBYTAdZx6B53aCLsGh3FfbMaSpc3ncgXhseDzJxObS+
XUnXpctXYLfU1PmKNr6HqZa8X8q2snhsDE58Xh0E4n/cAThEBLY81eJoHlHUphKk
zpa5cJNGtwqi+0qtQbmyWSjvQfbZ3cWWchsMltxITJYNHbP3yytRmM0m5UowBdw8
MnpygsLaiW5jcfqVSBGk7tyG79ZLI+uk95PhUO9uQhCBX7oJ2hr+90BQRtogmH7F
qS9sfjMl5LIHQ3P4XLxi+ys0BIVDVYclAhcvAF5kiTDzOEO48ZXVBj2iaZwHEE6o
Iaiah5h1Ay72Hi265+5eiQjmRjL9zyzJCfM5N/NvTSjXgjZ3LIUr54UaECoRvbXf
ly4TkWVjQgn2oZtYdjuxGtyhrxv66ycnbnNuJZOAJc6ORZ5rhpLb9Kzslc8MD2ts
jakEPHkj5A6Q39OJYC8K86G7ow7JvRVkB5hlxjGWyzzfFJ5qIoWRgj6upE0tWnpc
Bp74RthlZvgq0X3n13ETAYIIRYWGi+XCDNWM2+pKrtSIJGMoYN8aeQ5IsGZ+kU+J
Y2hNP6FvW++xRIONGgCV0WwnI4VXPlX+lw2IafZU4HurmuRPaVFsjTPACwqz8ynC
nPNKrbkV844llek8ioFb6+0cmxfRrbCIx1sQkGOMhaY7uZd2CIyqkT0qidyIkzfE
5S5+Ba4rcdoMRobcuVqoU1raLQzLXnPfR5uGcu8SKP3+gqzbtzzqV00irtWH1vp+
QVMlAmde0HHdmfO+xut8pzhQkhPfLT3PGANmYvcbDAMcE0LA95Vj7M7/An9CgVtL
D8kPJ+l45ua8XIvxZRFfuIm2xRf7wNvyuKGl2i8l/6vX95VreWtd1G9P0QR0sclm
+/alyGdGMAyySm6RrdGyskRoaihVxIFamwDmA+RDgEizEt3aeQkUS3BCcAVy5PZC
gtA+PPKF5O247XwVKaZINzRUqoX8a5RrV0hQhMf/rTqQ5NGCzGUvgKUChdlk4/3M
rtfK9uQAisptujPMNwyK6XrYLSikPUV/zAMHrmOLBacG2kwmbLFtn7jR7bF98xQf
O220U8JRXdY1uKX67yxHOj+IiWW5m/HIqAl8zPOQb4MO0a3X0rWI8X0HjQr8vv0m
MDrqFWuEc6jWChy+zMV1v7tKt1yYQJkgKVd0V6i7wnU1dmzNS5Bx10TnwO/g9fmq
NrQbDhsLnc5J7E9+dVQxbRPvfqZic1uDKYyRLbusGfuF0oRQBj7EXBw+Z16QnVcG
7fD0DDTS06LzOOPKB0V43mFHN6wXXe+vZV0iweLNx3w8sjcDE5OgcEd4MNlO0c1c
zOZGOJAY/4WNMUMkTXU1j+7CV/UrTos1j/4h2+Ctajdph60LJ0lCS8whWx5O8Sf/
mi9F1bG2ghOKfp53WaFBYlKG7yOcxBPlz+MMEMfeNVcwRT7pJv49J+zTJBaqDN6W
/TklHY3y05jjwGPHNULoLWz6SbYPcIPoyPyq4sSMiJu5izxBz50vXpqnt6xG66fF
t1ei2EGZXTjglM54VBWfzoVEbQgM4QEhqut9FvdHYYBhYf2xg3XkVu6cxsyX7i08
Xx8EVh59pFFRjkJOHDXa75Piw6PE8IhogktQ5+CSmBe/KcOt/AcbIeP1+UwzD5OL
tVVG9Jiga6mjIbGcPrCBfvSSlknifEEOenhyjAS/RvItVvHEgXzrx9YgPaGGNAWB
LxFzO8bfOoKZc24YxwJvbJq+G6VzJDOaOAR6BJv/d4mhtcszxJNkUnz1N/xjheBa
OdG09Fn2gD55yiBN69bUFZRfln+bE4JiBgB3wuS/JhgU3z6v8IRgDjRWtRDS9MwN
eSEmwkRkvmPmA/7cKGqWks8c6oLZutd/nJsHFcb2kHpQEWytWni0SjnEZsHx/dqP
vATvXJlcTK9AMgE/rWObHUIP4pvo8lqFpebKqkUGGGDWxKymlZr9IMIkshmPY/dP
lc80ABRLaqt6SllrTSUuwhWdYYPHU/fFKwJLzwQvYFaKNGBVm53kqCg4o3fJ8K1q
Ue8tA+elHYXVaHKZDbihrG4nA2cXk4R3c7JkbPg56EKF58JEEoKyr5PAQZHSEOBu
5MdOChM7LvmxcSGEMSW5CRUOKQGq1sRZD/NUjXgVSUNS5UrsCFf5KXxxIcIFpUuJ
Au9fCG5UHOw6W314vNHKrkVSMMeEq0mb2AmMqHHjWpuNm8b6gDK6LcfDPUGwq8q0
nCxd9Xrvg0DKmY5MI46yjgzx96p771LyThZqdMV/9yYP4Bqb5d0pEnmY3K6MDFPE
RyTo3CaFwYf6u07RgTEkeva5MJGDAYpI5luDJ2iUgxnfvg10HCBAosc7NUe2Hm1E
30epDvx/QV0j+lUMGgt8e7mLwoJ7DNrujsz7qJOEOluRBkG+YlhuFYblarCyvYgP
fFjS2C26B9Yqw+8uGkyJRPnqFe2u3WtgNpNjLfx8bHdd746ZVfTlSNynXQTX+/f2
wS4sbacKuSgc+lq/01+32fKRfLcRzXCO0xwF4pdMXLkbN/9/EE4Q6xQVe98Kj5nD
IEXYWa4WEkCgA53QsyCrm+lkZKkZ/7hvUXpdrJqiL0eW8JQhCeAhhm3Zl/nuh6KT
3PdiE4oozxMJnVBNUDKDZt3NRJmCARXxcmK+lYhM/mxTP2/Vte5DByQjVqu4SEV/
fFXHZ+mVv6gwoSGgEt0KYY/Jt44zvEXrV4irjrRZYoczw2ZFiztO0DI4eqEL2g7R
07umHQ6rE4xfE12uC/KqhTdt/AC8NTNeN7vpZA9B2mneSXw696+c5hU1WRVfxDaY
VnzaG091h5JPN4BNc3xk8uhoSoTm+IPEKQgssNV9+ok66+65sazeh2TXBlB9zy1K
LmnfjbZLMQ5aGDsnosKZiL4t4NPrclNhtDSmsivMpQlq8hYvVMscZIRbsxUXxyyH
RF2dNPamxkODRAGl4jit0Vm/BWyUD0PeI4r/hRwHvhceH5zlIUpg6LEa0q8JQkRe
s9pf7gXO7nHsfSNE+zOHKulLCGi2jQyo6mncaP2UZzecm6kFXhssGkkw/oxrPmek
9OW9U5nIFde7msvI5jhwmAvD1bfb/q+wOyvIltJcPKkQFITSoI2QcI9E4HVKw/qd
2tNdqCbovYorTnPGvKAgSHYsptTrunG/IB4ZL9PCTl6nT+um6AdOHMaIIDKQwtKZ
qgaOgsIas7d3AnZIKv5Cst2Vxlhe+OstoLCTW+guyG8T1iqfQZ6uHH4K3gQKLBeo
EdQVgz/l0+UVroPBZOeelZUFtk9vofB78FHrPM/bujWr+q5uY2irNdQb75xduUyH
zeGrHchw6jbXiJUpc5R+NqeLhd13eIGCjFkGtPFU0a3lsFW2+cmJU7Jt2CFjCTJW
97VsWIU3NV9KCleEpKNvSIlsagLMQKdmX/OYkReZe2bGgmDV8D/L+YPtIavrqaDe
+bJY8G5pchFPMcujTtjcPC3++vlE2Ob2FauaiFx9k996j+CXlojbt1wg7lhZoxK0
N2q4kaisg7vG9odp97KXa6yxtlAffA+u23+4001R2mEgYL18NnJn7Cyf+Th+PcE7
3Dh/stUfIyW3kMMYaA9ruwEa6zFFaLrTTBm0UA892r+E63vrlm+NURyUHq+0nRQM
nDicCT7+hnF6oPQQN4rBVQb4tsugH4BBfqxuThowHLJ7K5JEpwG5SvV0xGdcOV8P
MzbdxMUvTwLv8BKlQBGQhjjSHDkBoibB3qz39rZLV4IqdB1Q0mXF2E8WViCTvF+W
0JS+EOrs8LAv++yFvf44HobVJ2BCVxGxeqV6vE20OZdqgVKLLI9dorISsWuekv+J
FZKNXRsCuXf+jsakTgPYw6xsr+JahJ146/O5U3tEY9vYUysSbRkq+ttWABUMNRfi
ZBWctvlIyMxHkMuF3nehRjif4roiot+YuULIgi5Kq8fmUltEU7ojSQkVOC8fSckK
q94nRyT02BfLHpHR17/jZ3ScFGAnvZlj0AVfpxkzUMQp6uuTGq0MVp5AG70J54Xf
N9xG9M77WrzWY8DtX7rIQvSrqDQ12YwBaJtc0gi3E4wZwKU+iFK/zGomN5HicX2H
swZ2IRJgLa4EyqqEEzhM+9gEkfcDFzWu96RN5lUjVeczBzqkRWqbiUzrvpBa+Wxl
cDuOCZDS9hp9Gj9AtmVbBLXD/h45rSbwlhSyzmg12+FuFlzsDn3i5nyH76rzaqvw
roSwLXWVhD00y9BJb+KZUrSawm0KUjyO0eMTdpMak2qXhSrxK4HeQw95qPjb5orO
lv/PqmA9HLRKixzV7No8jlm69QnKObaLxFKc37BWtcPVXREK7zy2rDMrFdKMBr7N
IffGQmbUp5CEjMC0KT8kZQQ+hrS5tGfkwyipvUyYKQ6l52UTsOZK/OnOW7q8Iu6g
zxMCwadjRckdWZmX1qeyBnqwuVxQmhGQNgQeWTkv/Bg1ZYssk6KqaLk8WouAynNn
Jyv3t3V0Kvmw0e/Eau56Dg1niNlqXxleqC6xNoc/ZqbUiDMxRxUirHK3wwu0WWaH
ljD5La1OLsVzfqhh/xZhwJnD1eQVLYtBZ/JRrARdgR6nN5QUPochXTa5zOW4LWXH
8iWDuKRFQTmmAl/ZE85MiAII+WGfwf3oo7Tn7t9cKcEj9F5ZY8vtk3cjslC/EV3q
1bSCVcyMZZL3guI9MBdskhHyvpAMDPkOVK8yWwbUpZqW24QBvLlpHApTE5Ay55Re
tymDXa1S9KRg6ONwvkZDMkgHkFwlGseJCQgsA2+Vl7fWD4EBsVRmqo1LjJi+zRkM
RrtpqGi8ULVVGBOhiX6qEmmQr6LSeN0PePPaVRNP/el8PWcu8PrChL8a8rzwheHU
uIHa+mBWYIiMWsEFnPg1t3Vzs0Y6vnv/kDTcoQrekNwYoYPLtLu28p4sDmyAdA5g
Ae5NmsC+Igbzei+CtmkdyY2nI7TG35bDZXpy/PafHpsuSHsKgAspNG4Oe0T8UbIy
0R2ILeiqNwXSNAxSuqc/zmMz7zBgJBxWQVDhzp502pYe+qlbHeR+mlFW44FreDG1
1zvHTuZDFefLS0av9kgz9tMk0reXskb6Js4hRA/wIEY6r8bqh/kz2EDc9EYmaOGP
n+LSEPgwuWhLX4yL9nJGvGFl3gIHDnECfK2c8qTXR72/Hd3e5asgkzHRKArQgpD3
dXo6uxufx9hCcgy3cfSQJRjaeoeN9U0ZAvyIhBd10BY2ux2inQCSb05FsfUVjy4V
0lXov47nRf1192KbiA1lWPRobIDKkZEstt0EhrgYOSi823lhpI7wImzMWdZRnhKw
jTRaeQGogy2K6KShs8m3l1rGJsjie8uPtWQQn9QojCghyxbamVB6IwqVaeAK7NsS
fdA7QSLCWw/stiyeenfGTSST3xahQ4kr21QNfvPWUcOsxpBF82bZzADqLETlLicG
a57jAUa+gXyxULl18xcWexgITUhb2ozqJnNUFWrdpPwEC+dohGsbkWE6BPyCQqJ5
LPWyDWAWyPxjvO/l3Ykhu7aF8+hvLz5G/5b1var4Ngc4idPTIAaOTQSFVk5hKvuu
1kvUIrmTd1Mkny8vca9Z6tflH1SNYoT01GzZEM5ugJ5Yok18z05d6EOHT0oO5TLq
SC+0xMW2ccAnHpk9qC6dmlxC0gU34wGzXKkBm7Zt468VNAKmpXz7B3oeKpSDMANx
12teJZ1+UBlNips8gysIb2L8XLeOQSRz4byXdJRLf8Jokbda/2eDwY4WiqhdHTcH
Lcs6v+/Pgh4FDYJLCV8kEiHftQnRKU6qN7+C/T3zhoVqX1jV2l96CDBW8pyxrIMV
wYYsk40XVMEeo6l60f8ATViSdMN4HYLdk6OeWWq+b2fobZcz0V4vFbSPtpwtIRe+
0D/Jg2XZAEb0lDPIysjbSXDgKpgbbQZZRLH/R1BVQ2X+rBi5ypg9PDh58FZ4l44Q
AIJfcSWuU7G+u03jks2V6mcpinzsRK+BOxEBGm1qGs4P4UDTj2av2ElEjf1EnEjH
qxVQV7gkDFrKo8qjeTNTpbAC6/tzer8XgpfFb877+t+iXWMmVNjUjSLTgMgBeaDT
MadO043kiC6eALHXuBkPv1DFWfEWg1UHS3RIoM+oKlpNfsHO1P+yW4lTy4QLohIv
VmhW2tLIl49fjmqa8KmSH/bedRxWrDVrAlX6TTzRFkUM3NivjKt4MFjVF/I5Nl4j
gU+uSFWI76n1OPGvRzWQYZeiV09n+E+2LYbDUPuCkk7IHR1O4fhjNXSTP9UE+OUC
3/r095c3ZkG3K4+iiHyS6EhldiZ4mk6CGrrQOIoUIy9Y3ImGlKpugUTiG5/cuNvZ
faqeSt8q3ymcz2WblrTTON4ZqRyl1ayCOff44MpCcpEvMBj1jUBB23qQITpIfC5X
Zqzprz2zwMJVHazHMW4GJMKV7v5tvjjljqAZy+gPXyFAkbkTkIWknYhH/luJ5cKk
HpLFzUBAePexdP0YCKQAPEkGm4Q3R9RU1TFGM6yga7PiMUp8OaZNgpUQY7BacFY+
qlkA7VGSo7Bh1f5op23BP5xjSD5C9Z1l+HZi1FGLtGRau5zhcPL9OX2w+WuJN6jg
LvST6A+TyxT6jI1Xtq9IzcIJQBcIG+sjzsEHMeW14wGbM7Fwl2g1xHWszYlXU/Gt
S8YobmV7zilypkKABONrPnoj4E74pYl87LOgHpARMJeJShFc8GTbmxlz8QYDAQ7l
03SAp8xmX8r/FcihUxo8ckTdHfINiOUo4Q1QQcDcfnsAhwDlSFVz4of6piXhadkM
jzUMTpxgUw/MSt9pssNdfGYfje1mERdjUbarM7Y6eE1jtysVf9OUZ/GkcLECw0C+
awQrUAdc/rdWdfyu8bg/amzZzaaaPXf3kfATdg1lNGz8p8Ill8jeFo7Q1FVosE6q
i/bkwAp1x0MNgjcQkecBPExHY2t7tACMca7ckhuOyftWYpEtb67NWTtSosAAo/us
M0ZvYigo+UCkWkj/2gSBRQCwQPG9twATE3ANWpDKjeeAVtzAubUbmerOTM2KxrdF
UDaMbAfynp1XOm3J4F7Rc8kA9pAQS6z9aXprgGewOC6YJ/5U6V9TonRIQpvZdct/
cJC9vH5sRGblYFUvAnN0R55taxNL+Iax5muB97l7dqoiFmXL8Nn1iTr+PuNgDlth
m8ccAnEybAWdY2kexVH9wa5C7DOT6pa5XfTB3EVqBqT8OkMER9hVh6IzDJawt5fI
cKzgtVwKtMqcZHjqmCHW1OZm6R2TSvyEdZ8ArAieb6XOb21YxgCHZburpDhmjs/J
VPRa60mGgPywVmg8BzxVKCbvT1mZe10sTotgg06dzh5e9669lQlX0rq6ojnucnSJ
9OKzY8EcF1WYWhtMb71iaOPcmaqtPVSN+yO+CJoX2IwQldvaGWEuhOmmYYAJolAL
mDK2JKMTDff8TRgz1Oiy+pl/Kdwansvr5hC0jGIcDCrdJn6PDR9vIZKQkOZrka63
fxfHiZVd5A18+6ho9UT7T940//ESgxzLxw5SJxzRkDHdOtyXbHZRjDeSf+1z122+
41w56GG6uRopekjwTQEcfh04WviKfhdNl/sFsor+YFELoj1E9UwHHWnj9MDCiSs3
XD01c4myDvLnWii04tmGtYdv/25CMhrLtUYZY67xuNgcEonyXZgUGUODpQ2jlwci
lEi16vBSzJDwelJovBw9lAMrtEr2uAEFtlU0U8bzSwO1GGKZlS2+AzGJME9sY0EA
XWHnNG/Aj27UAWbS23Eae0+7vR25p1XFncNL5S54NhXiY+QZN6tZqBQsTXZF/ujF
CgLgh1p5hITTn1nP6AbwfEfejCpeFirHtt/nHkUnstbkFhpeXkqTMI6A9mXzEcyz
QdO9uAjgCao00TrxYD7JGeTZ4LRBOdovkwdfoVFmJrtlt8ppCmYJzO4Al1iWUYK4
bQpJb5xoGWcxYhxAtPisroP8URYM5j0PoGXO1notcPLawKspgDfAbF2mHS3yuOK3
JbNgFVE4q1/TZfJjbkdPluPAAKx3hsdbRdSO0uoPH1T0Us2mU77DqtbBzCG1YSz4
+VBi5IBFzyhxt44l50IwF0OK8lKbvd1Yj2B1F/z3ZiTfpsIjvWT14pOPQA0b18zR
OSQZW/P17pCE+D3fRfUsWehLiKAYqUo6Rf8eeMqjbJfeGcfTyIeykVDcynYG2wFA
vdANsCX9pWlbmgEcPcSQPfb8+hGwWHM6su7sPe8QqqkLZgoPyZ/cIuiXruIS84pY
xpd2yarZCoDDchzPwxu7mkuD6GPLIrtMWXswSke5MpFK7X3quSmIXoqc2Rd1BMoE
7rGlFJJ1skn6k38czu7orw/S5NNeOkTIXq5+0y6MTApEnYN9ks5kDJfpcyphLD3s
cu2DmKm3LKfwNyWfP6TK/12sGIXK2i+YsQIEuNfFAMubhvLszb1RH87YvfXa28MX
yTKb1IS1nHEp8jAQ2kH6lSmU3hfkEfj6mok5/CaEK48AZ7yqx71SWYDqkLzawRhT
8vGYahEpqL4l8S1wCSTBU0DjueY/GfZMfSzbFa+t9OylWgMKw/LwejbAxNxXkI7p
EqmznxU+RClVO6Y+zKuM87ZNxlfVielg2sJQf9aUodm/xj4aK/Z1nLon56QIWRjG
hNtfXOB1dQqGBsqRFyhHUFwOoNOJD4DBaDJBoqhCWitN9Xl/J2YNYIFRacH33XFW
hnlqbKalJg6E3Q1LHRiEOdZtpL16cpe8fS92OvpAIPtVDqIovm0SMniepjwhNRAJ
OPhdoqRFxBA5EmXLO01lRwXCDAxc9RjMyzT4m9970i9YQO5lrovLPweHk/CGVnMd
Gy1tj90XC6j54U4ZgCrmkqQfchr5ewNvzmUEMUDPf/u6v9VRdYpPJvz1b/epyp12
Dd/oMbujj+rjKzWYkvHK0TXD0TIRI1KWmTt2N1VFp3IzlU/JDfBMTt5hoyBr5G+E
IQPRHjVDtYYyJPgUc24kwujQpLPUvQkJfqDm4tP57LTySSBr9Mk2aglxJ13LUHiz
3BXL1Teo3qXI0jDQlPGZiNF7+tl3JgGy+Fv/uMyLG+q46rFHdTb7c3SPeA6EDI4J
nmwJGqPYnc26pCDTYoWu9xLhZocZIaMmZOoTsao65c2kCSqCIp/uEEyiG4PtEeOp
fmjdN6dvyoa2SgKeB7ButhP634w8rCGr4FJ6dEfRVAwb8OUrQ4sPqlIRhUekDCW9
S05voL9NHOmkG2dW5QppO0NWpRi/m2SkVIpHxmhnh5h/BLMeplo1earz29qdCWKy
T6NTtrK6db3mx0kl8Cy40XLyfXtOdlKAeXw7I6/gEBHBmTlXSEungnAt2HAsWngA
yE1eJzyJusMWrqBTDeuaNqQGI2aUYBv44KqiL9k67SIG3j2ZJA3QZBdAId9ryJnT
EOTWZ/PEYSyWrItfFQwFaJQ4No2q1JokYYu41bcA24PV3UK+nN/8JUkJgszH+XXg
4zn2XbkH3o4s8XFiyRn67XqtrR0fr6r8oWvtJH3OcnDDNAN+761YcvnBpGXCPHdv
Dqzl0wD32fm3o6+U2QeUszjO+HilRSxCK80+cgBm1VUDtCKjwQhFN/FgTqPJk5Ks
71Tkc+a51XbsHepAwAPl8VpbaZdB2cENSBnnk29J5rzj0xHY55xudcC/NCCpLVgb
tc0Fn4nzHJko4fZQuUVchjYhDZ6bNw2GSzwd1El0s575gmvSuZTQGuKBMwyLp/wg
K1p1O8waBdJYeWaXyBcKBvDItlOwDzL9fNsB9rYfC93M7YYxfSqBcFhKEFjCk3r3
gJ/3Hz2W4ThoNX57OdYL33n7jkxw7eYaxFDL3n/0MbMVHC58tQV5M508i/IA2KXd
cvZRqUfYkVl09NcRKpV3E0RIzUPQf6oIXQMPEmMi/mZwlOzWn16LYtM4LQGhNZDZ
jPw8HaAA9r8uiymwRvUNOmDA3NeaG5oOwJojMONWjwhdHQz43fvwC99qZN7eCM/u
2MrdTFATMZWCX28/YxbJBWa4fsqeH6vSFXxr5Y/9Ryd/j3mHo4CPEzf0CpDUDZdq
HkUVjfWnHqxJCKrF8+mX8wusF8URVkqYOigrpmNdtqQOoAEL/81Vpt58LRIE/frn
czpN/39OdERdgwK3Xh8QCxrW5vQhJD4Ttpq2iZFx5nquz0O+zUVqMU6cAg+ncfIx
sI5VIYyPYpjay6FMu2Wq7AeF0eGRkC4qG0l2AaVMmbxAl9XnkB5IZiet6cLjxHeC
SvVeZ+EJAsLhqkm+wy2DQ4EyoGu+M4g0KoP9vzya7g5/9R7j3969tHRggyLhXuEL
a6ick1jv+pkzBDGGZPKebWRIEc3y3VI+q6y4lZ4Unkazjftc3wCm/scVcYluMVrh
YKRo+VUuHgJ10RAmF7FucsMXy2ejccLdjeKeyRo3w1WMaCPuthyp+S4G+Q4ibZnP
JgnXiswrHGiQfwBhEIWO77UyrCe62cWux6d6LJV2uDFMQjn9rbMgDkB54b2ymU8Q
hpXX316sw2S/OAm5QpHcDn1rGPXqOrxAyJx2jusZFEDgP7ti1dZMsv0lFWtrPT1r
iMhj+SOWgv19VtD6cExVqfRvmer6Pdl5o5Fkl7aWzpvJ9Y8VOvYIZlbWHCIYgjzX
7ciShPgNII6aHilkRMa7mz722///p1hA+XB0dsxTWMwthFtypIHMyZJtN9d/soq3
GPO4+E4NziPn/NPfao6ZyCG8PzQXdHX5xBySIZy6wBn829uwEkh5GY9gAugsePP9
RaPcVMv3FIXPlfQb0sCKbu/gjssXAZZ+6FYEcrYGbJzlTYecuuqd+Sfn/PzR4Rnw
Rf43ikzu570cNJCUa49YlK/kaNAElh/7HwJASGiJuWhgfJ7+YDvYuT4M/BaBfRMo
P/q4rX42Gws2FaYRlSM0y7VZcmVzFlHpL8vMtkvt4vyCZYpzXMx4/t9aumgueGKy
ziQd9Dhicfkf2jUjMb+hLWJX6EjvA9w2YjPICuwRQPStF25ypxRd42KKVksgEVAf
1APGjvn13ZZqaZSX60ffHQUK9LU+xwsxls+OF5zIdSnXaTZPaeSC/j/M2Fvv9Rn0
t77ul9ly+yhFI+M+rOdwBuymrlE2LhUwPoP5fkmEnXRnIY9ZlAneyTOspPQ9DX2i
VsEOKPnqj+2DW6xI5WrubH8xu9O9MEW+n1OrfLkfAaqxIQb8YipyufM8t6/nyh9e
ezqZbJcd4hAtDV8UIk2uSr+CHoBfKKwcALuA9rKtyONZ2W0Iez1L/+RyvlYUNIRr
Gsh7j0XySCXc74qO2+FbjSCwydEMVqNmNDr64c8iAC0NtXCl/IHS9NAUnvVBsRxj
WHBzh6J2kUcyiHcFnTQaleXtiVMP9lXKX7+hCtBKy2HjzhbhedORsvNR3tLtR3Ok
7Led0B7Knsp/YRZ6KQ61dztAFGB4K5SLin21AOPCscBYnDRaRLvwQ15DUfggoSq3
Kl5M5lQmsSNwiCYDV5Uf9Rgd8MfeFWBU0ykgt2+UoQMJJxcYo2M0drg0nkixv4VY
4bzpw+9vQ1cBKCWqTi0g/Kl003OCs+U5JfmB1zD8WuqVmyoronqkMbP35gIudDaQ
lMDYRp7mgURcSLTvTzKZbtrDjMk25neeSmSPVTPIW4CCE2QVnP5aHJ/tjmp7cdcO
9dUBcSsIe13/otZMSJNS87Dv0tc+5WwMEs7QasDC6hZYWhPKRN+n3Do/fByj5zn0
f5taJpw40E9+FUo7OjsytqbWPh3sVTjW569Du1Y0hP16/YkHIyJq+2IT1lhcKNnQ
JOsz5j61/PA5DZSLKTLQl+bqhSBeIN27WBI/AZMNRAVdNXLTSDn75aNIW3my6ORP
WuE+FAXTy6MbD0xZwSmwF59Q/Aq44N92X4zT7ub/1P2bKUST4pfZJwMobynwDs8Q
ntxYMfIT4juDeCwYo6/+IR5S0Jqb0GT7ztjHofchRtZuWf+XZ+BN4fKqAOWbPt3a
20+PVZNQh399ogaFfw9wgXpskFWSssBgMYhBrVsahudgUGWf4YGTQhT+V+6S2Qcg
OGweL4zmLmlClTMnFtRs4k1TGNthnEJS8fmQ2DoH0sLo8YD6O50ODJ3/5ySM7eJw
FsP+Gx4UjCljFs2MFAvYHnTZjmLTXQY49VPMism9fC9V4fM24HLrVjVShPawZQ/L
siGmVFKoLBg8a7misrQ5AZyVByL9V8hDawXb2RQP03Tsao7NA9b9Q0GYBX8OVnlw
PVoSO5bGCbkHg82ccN1Hk1rq7AVNFj/YYCpX1cy87VCI56SJ9xtzRg0tFNVdN+aS
Zo0IlHqVyeKkxWcwuj5+CxGIhsJenjTzmrw2b84pFVhp3FNpzOJnwF2G2xHWvvh0
MFmlAgGiBKpHBQh+pGWS9h+CC7qGWE9LNSXL9kEUqlWGeSd2pcNV1Jjqn78xskSc
oh0EZuv8zM4rtniktpZSK7qXChq78P/8RgWSpDEsoji99lWMW4l/CWH46sy1ueOI
n2kVzwWbNgLrsxPZUtaf9YgpZgbe11PkBBvOdOl86RAE/VdbtI1Fj7e5BX4tLCfH
3yU6vWYdmi19/T2dcv8CodIFKN0Lp+clyzNKKTazwEsZ/Mj7LXzDpUcQE6uujz3Z
eZTeu9uygE854Zw/p7pGINpGfYEx1jr+SQmEl9G4J9j135ObCKuG2bNmmsEXSJWq
UdepooAX4zSnEKVjJOCygqLNDIeU0O9L34jP0x3A4gX73e+ABf1Hgfa8ncvgrFAQ
bpbhsGq7MnhyrR7ShOiFfz0iL9wWBUKZeDOppMjMqKYNOSN5Fr0OwXvnGALG6GMm
aUpj6Zb88czTQwa4L8UkJbjdKvtANLRQw47bdn5E0UMgbayP7YBudLzO5gKfUBWc
QgpVVzab3c1dQJwnDRCBJ8u7XVyFfVSK5k8EFAkM7TD0mVK4pm2VjIjxaX0XoApx
WHWCAy3W3Gqo3twEz8g6iAF9/o1hHWsT3vvmRrEoBSliuKQK0sJFGIkpnFwjaUSn
nAqlTB6XrSzbFQYC8JZnwLVkD5SAwZBV8wPgJ5chf6nPBHVOfhuUiZ9vfKI8046w
ykahBODruC/JNME3O1pWnv3BI0Oc2aa9oHtld+vMOeO3Li5fCiqKzV7GtrCsT4MK
Tng9ygT85szbvHa5hccLDescX1IfWjkLu4JHqLt5vsgn9M9Hq1MxIffXeI0UKdik
aICa2F2GLr/CuD4iEu3fFcHiCPKu2s1jwk2YoqpWyeDUnvbnIBfv/IVvyAuKF6DJ
zoJo39bm5qWntiF7vABxB941RkkcJCmDibWBu2ApPdheK6cUgqPukWO3ffNvSZwa
hbQy4caSmLvlkIuEUrM8DW2yx1FusPdZSBu+nkhJ07GmI/9Vfen7zlncWlkglQL0
YyazCelUzfrwIynuXAfiVJ8FIZnT4n2F4Nro/nSVRnnQklZ3QlunZJz9rM8sUwfl
yLVxmg9Uph/Ni/FMkvg9z1W0nQ4FwMWASQEqLnAFeZMntWQeMCGzM0Zb+HlRcLzN
RFUBfhsneVNZKnVK2CJQroAg/2QwdE9rrPWnWTu1W1BUNt2hB/YM4qjGMCchGnwg
rN3nWB6EgPxqXl9NsRKVjOJeZl4DlDbnvs3UwPK99UfbcViP4AHpXUrB0iL4z/0o
3k22sLmkhDwjNSzKHe+dkSWUniDPXiMTclEwjs20LcVXIAArMfPVroEojQaWgtmO
0mBEV+hU4foQSZGFvLrvofiRmT8ppm414jH+wuREsOI6CVS+/md9W91U4juKa2lD
cVHuBrGiocXl6gA3/xWf8O5EWvC53B9Gw0KD/XnNlRzAmUwL8KYtGdb8IIXd6XS+
UqvJI0kNdDTSy+I/FfsCVcNJSs0WBeYs9eQeq9fZGDuRzCCeQ4QPoaNYrEG0rYWd
O1gp7DHXUDTppzAwr2lgDtIdaUxuIue9DQ2rTiFJDoxXIElXUI4gmITuqIBBYC3j
aZwW11mSjhNcvpNz0L8Lu4jMd/ue4JdG1gpgtlPiymyQPY68XgMAkQg+p0qNowsD
4+yNZCnKcB1H+2kjuI9+wy9KJ90MOleMqJuHe0xWKo09JFKfKM1AlgVGp/cAeluR
IWLsOWspB5mYDcEifPtwU7Icd7VmDjO8/6Z7wB1MPn/4PZX1eDTlMXLNsCE9DrIh
s04EzIq6CncuJ47cZ4fwp6OKXrMTG26FqRmevOTtuuJKLLH4hUOjMMbu0dhWmOdx
Ze4HkmqGzytUO+iTzKCEAWLWXpuyq+/t6b+54vAuC8jtJ2bGRZUeh0oAY0OGXdh2
9xnCyndH8Xg7VHu2J9ObB/LHjhLWUWReq2Ddvoxh7gz7VgGylTQA1u5/DzNIWYBZ
V7qXf6fslSggepv4SjSCnqL4M6hO4plfHS4PySzm+35DjWhNWN8YK8TkLI203+jD
BlThvOw2vbkfzMlNvuB4AhnZWtRq4Z9pVx8x4OMKQgTmdoSy+FEUzwJyFNvzC+Ro
I1mKYYhM4sZwTZD70XmbBzOhc/U9iXs+Aoc4wfmzCEdo42T7rSQoYwER3S1YKg+1
SXVnsV9PU/+nAi2UPnHBOcbhyDcKcpfFuGSOgNQOY5ErziAPcl0xD2M4DRx9lOzw
r0V8Y2yyvmh8ssztab7jt+3Jae4/zi0LxyLKjJEVP6T8Wo4hhtRmQ0MwbKNYY16u
vcCS+9Vh9EyMlK4X4zCozZ+BAd6utG4GLKBqNdYX6AWFh3r34+e67M8ep3CJ4ZkN
9uMsobmz9x2ct6dsblaaaoeD8JAg10BklzCEMpbtu2eOlk6sdBLz75RaYjfo2UGQ
umSOn53V8jbK3Rb61Uiztj9/b6z6jdfuMdmaC3Jvt2rjrWw5TG3HJTfyAYUHX0ko
0ypeDXlNkcqwGvd+Gf0GhtbV17OQq2g72GpmcxkS33Lufb0CUqo77eN0Xs1vt+An
e8+BrHr4KZbuoyCaa6m+3bZoxSr7B9XnWanAkcvFEGDzKIg2nTTUb3xVhIOpfiOR
W61MO+5JaqeslwFtmjab72PHXURqZdfu0mFhK2fwbmjcrTq0jxyCZKy/kzGOJor+
152C/xZPCtsP88qaRS4HCc83u77JqEW9Is80zivnOwhFUoURJ0+/SvicPc6lOTtz
EZLgDCB3Ajz4fAQX9Gwl5j4CEWWfReDp7a36At9ebyTwcppkxo1dvmWNTMCxSlaR
J072LoKKkXHWxYCESYr+AzncKsLMwTzwrAg/xYYgIz5jgM0riFvIIjWawhsqWFgW
9OOZyHVoeltRz+glMJ413vzVAJTN95+WCqBzoe0gO4gTso0uG6qDAHGbdwrVbFwv
/d/zNB4qtM0Sin9IpYKBohzASQEAB8njJxHBUm8O2wxtBFIRo54hwwgQLtOGo4Uu
+0gBPuy7ZTfUgVyvrLzpByuh2tUx08rS/OxikChvpKYGmss62N8YN0rRe1yJllr0
QtaqBDZsT/VpOcztlk0T914P8q226M57dlUs77uXJcDlZojjy3i5sFfKqECDzRJ2
/CZJBzf1+4L2av3n3+NUJgy6N3gyEDnlEY0AH4XvCc9S6qenc/W/HvyGH8kUbeLs
87HjyHDQfZ9WRJ1yfcTjIwkL3RO/mslGsKsJgg3Ba2jOew7YkfusEJFUDIuhcmGb
K72vW8OoDgQx+AlMERhx3nNICXAef2OopEFSYO/JgsFS6E1adSa76L4S19jcYHLC
ZLWMF26n45XuGC7wM2OLDTm/qoN1Sk95Mo+3oe22PXm/iag2NVD61rXcCHw95d2C
HZV9ssLrmrpI7D0dHH9w7VGNg3mOs9GtsuyR/isi2MSvR1i7MYUciLQOySl8VjZR
7EaWXyORFSPbSzm1BQ6hKuiXn4IqbZxQRupRX86PS4rPAEgxr7RWWBIKHFAFEbv8
rDq8DmIqhlN0hG+v+hODQ3pbFTqze9N11jKSVfseGgNmJK9IYPrpHrAwWiwEY8ze
Ep/Tt9haexWwHLI+ZQeacKMfJtLheKJOPfh8DDKR57EUP9uSOc0GWprvJgAvkjrL
WeFgd08vntealua0XOAQWB5rR7f+OJHX50NoKSyM77L/Fz84ww37CY6Ghjl7Bzmx
4IxKL5ryPe7hjjbHVC/5ypc2PSVajGrPTsAK0w0vG28yzITn6+EN6bsp7pCcdj/U
HQg9AeKAzVjTHTLcepszM1CdKbTsb3htw4hZaRXKtouGoO/pxv88B6tK0OyIlL98
lsespJvXngusXrFI+HlmVRjqXQ6lRnFDOI0LON7d7SNtU+Bhz6ILY+OyQf4IMn5b
CTK9/hu/C2FYvd22HOMygZp7pFf/1BwPL5k94bd4yePROECkOCtEIS8f9W6doC7/
89X/k3LwlK1I70Zyyf1r169DFXH49xcCgxz6HGF8CHez2/FDIk6glIeA0/L/pCAx
KQsQAyP+dsWsKe2d4UL3k0BWgH1L+a/ST/VZCz1Nmrpcfh8wmpKNyAEm4eAHrofE
RQRuH8X0CfRLY1g3DMBzhsDx/r6fTXkib3o7OGOE7iLbuwtVIb1oBethc+1lkXBh
VepkJUFt7NFNF1RMx3yBl7vB2V6ADUQ0G3L2J4vP/gd5ko8k9R1U4Io/FaFykmPX
cgKOAGgM2k8SUt8qE3XN3BagGQClt7QbuJjuoDQcnUUCl+47B77wSm8UWOUU8BoS
Q8lhRViyNZ+uU3zh5zf5qFNiqeAJS8RiUZG8gvNtzg9SjEbkebDVLwkdqC8ZpGia
00Zu3QteS84Du5me+ub9zHm57lV6U6mkak1sOkVdcglYAglh8iOEwrlvWTMNdLqA
KsTz2HEhyGctaU00uGr6uU/AOouN+rA2bORnQNaDfKS3mxgZv6bBWD8p5biA0kBr
ZH0DSGLSQYNSfr5lbvvMsD29MaVYREDpLzUCLmMNTFQODYU0PQOVA94OxsJJgh9C
VWg7x1lpE4nc4XsA0MLN8Q+fInDRHP2aSkBGIB0tm2WnupAyZAWjrp6y8LR7QbMn
a9NXoWvIOQdCR2J5ERHHiHNpgzrlRgQsj+x9aNQ8zl72h1Wi+Yps0q8AS4tjPSzg
tW8mdgUmpOie4c/NsgFJIfRnGjJkuA3tmIyTMu9S6jKEjaoQ0ZGlv9s6qRhkIOXo
XufLfRPpj52mT/jOaH/CWVaXddzd0s8mbjjzmcwxbCU68gVegodZTEPYFXD0ABo+
2Cr3AIK6j19TlJaTwKSXLg8+Dp3kzRukdoaLw915Ji66Eu8n073FbCW4/DHMZPk8
NCsofCHQif1yeu3J9nYOl7I9JXtxz3LodiyITwE97eQoFH1bURrsxetGqq7KPVcT
KGsnYU82fDkXkYrBFDY2HWq3xjkq4C/vt1eZ6QTaFpVkAAJBfbShiyUta8A8c09X
VdqERIjfiZEUaC5RoMk+4q3L7v9HDG5jRd85NGMw8fx3m4vzrTp/7yp6JAN3AZtG
vxsC5qIAcowkeSPqBOBb23pm3PL9TKkNT3vObRiWd5vE3nfLgAM37FboyNTQPSdD
0SrQPQml5pK5C2gCgHK2KGgwUCNt6HLfy9K9RYNegfD4VNhlqQyQ4GYYtRj3geZ7
N/CSDqaumCOLbo8tx49nYWyYabsRmU1RGKTEKRhCVj401I8L1n1SJ7YQo0vIasxK
0+e4BdcpVrBxJR9EHFz6h3TDsUYl+v/0pa6Ngd7Rf9kH3XGge+Q6RAYhcsQBQIcv
kk0eCfrJxa6VI8ypdv3s7Du9OfA5UA/qWmDSLsZQM+TJeaJlnHIEjrWJTrSAQvWZ
CvkQylM1giu/PuIJA066W8Cg8obunnLIh+GBWvFIIxUO8bzh6gUvXghYpglsKaIT
9z6vIeP1wjuF97j19COmI2/udpo9kuzYKC2Djkm5MQuUPsXO6JqxN0qZ75TKs0bQ
kmcrjroypAF39FqyGWMiGjjxbVh5YQZzg2ZEbB3Uo8vljbVt+W4JeUFb1EM0juiT
YZsDM4Jjl9GYLT1NA9K+5VlymBm0iN+q8fMXaBDV9BiSepmuBrVkvweXl4Oj9zdG
a9oYmbJpa2fDPcptHcw3N6lDaeG2wvd6LVkVRPXNE6LosT9QGLRQrisB4I+q8NZX
YQuIKaII5yNyk/bdOCZ2vU7TXjyXwqDf6Nmkf8yL5RobDPLRdbeZqi5QqhknyPD7
iUcoOXcKnn6oB5FIKhPfJijNMRpqHFCLLg/1obiC61zIWsVk2ha5kaStC7yrifzg
jfPbcTUD45gjioSRrAXF95VkvneeLGtGEJo/aM8pwOtACBZCggqA3KrcsbHUsyVR
CYEd2NbGfz07D4tNj6vG+VL0TqMUiumLKDooVGzSDLzX5t6l9MCwlVgQ1RtOLtre
5zTcInEfk9NCszuEUzJRbHvcT+ps//qyAuusCQD4iuT1FF9v35E4h7gSnUw4Lilm
TZToagIo1TjoL68SCxkO5Vjl1U7Go4jM0ENTOuJmAS9GFQhI2pcIomAbAwx3UGCF
kRWWOiq2Gs7qnHxetwsJrBOWFXMY7JxNaA7/fFl+vT4UcA5pUZj7HP+D4TIPgbTp
4Gcm0NdlD+oH2RwXhYLJtyS4rHuNwu2nls2gK4Siuyk6prP7t9s8kQyhYRi4q8ft
mwxxI00XpCX1eX/MWmUjGW1HRCT99rrYzGFMw4UnKXe7qXn6/XQtFl0jfgxdHmZc
5occbIaXGPnWxZkn4Q/V2un+DAm+dj2CdpBpUNPxt68yV6RP0JTGGF0Vxwjwoxih
8+5/Pmr7YMOKy5eGHQX2XAdLmG6CZIDCYtPRMVkbOwc4PmGw/Y3FEUv3tXGTHkUS
9maK+lcVtALYX5mDqdWgxbLb18cN3TNA0X+uFp3/RYCFnpxF0u2FF8YdyJtCuRiN
rMeZOlmXyoElF2DJKr0jU5mf6aJZR3PvZtrugEp74RaIYSuwXMbcQ8HkA9DaF7Jl
0VXbnOYh+EEag0YCcgIGVjgHJff67Z31NSuFfXvt6d3pAb1gzZRUili1cYsGMha0
v9IKCI7qbSSv+EK+RAg5FAPB9gG2EU5xiMBwUd94p95V/qMjcQmQQhGFsY6QsQ73
9C8gRksbidl/tKt3MPI51LFmgP10pjf7x5gMiFiRkbjEl75DGaOjXPuXUqHu9mvh
dzDrUbawPaPpIJaNS+PhZDo1YG9i84o8e3REGdqSZVmZEm1GI/hkpC4xTeXvXURn
i66rRfL9hy8Gs5bK2LSfaKBIPV06MH87fjr3R1ZotRPR2nOPgn6efCFxQoSHGWaO
ow9Ku4bnOHAdFQJM3V9kpRUA3g+4yoMNqBQkeP7j7JvV9eQYLr/BHsTe29trvDJC
2Vb6doX5a6ishmPbJTXtwDrPKxtLa/ltwSbN8cHd852QvpzGQDAYOYOaNttAUqwW
360XgiZiaPhbp3RvgRfJFzBydqELtyRfo/8ct9hFSS7pDxTVIZVJO9zV3CZMGCtA
`protect end_protected
