-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
4VpXV0W0MKvae+laM/95d41kLooTpO6T3QSM+HDSlYIHDeHRZHYOi8fRGj/rbb5q
zFBcy59Pvj4A2eKaML7uAFjQrzXRmNjpi7qru1AtZFgNJEv/13sEd3Lb5oWnYDi/
d2vgpeZlGw8p4d/VkqpxUjl1688Ee2sgc+ueylmteFDjZ811/b25/w==
--pragma protect end_key_block
--pragma protect digest_block
pxoaxRfDpSSSGNXrEyUQ2FMykD8=
--pragma protect end_digest_block
--pragma protect data_block
dGu778KRD/K+OOrfoAYUD1pyecYywVKPgCmT3dC8EJQfUKx7yCFmEGhWuN3+IgfI
ISMsUHG7bvFeFv3gi+9yhoZ5nIYvMPCyjS833VIBa6umWNcdneVB7FljsfAlr5Sy
O4AIYhGIUmQDV+lEzGuTD4055ngdET2TW/VP0C5Wm5dGCR3YcdoQJCQv1ZzpFvmy
TYxVMGh+Dyi8NArhgHQRj5qUgl/SFVxiwiRvrTejrC3i96xUMNISyLi6CU0gDAs0
Rr+mZH2uovWpnrI8bBp5R2WDCZa+BE4R0wdOwnQs733zxUeQVU0UsshljRsu83aC
bHdetJpw32EKFIVy04fgyCmV7N9l5/3FcBB89GsPV/GTzmj49ZQtm28cpZvgwtZI
P6OVYKTwlcZqGGiM18sIVDANK0SkSb6zfumc++HFc9xLKyvGuvUnv9ogSgmZSole
lxDyO/Kf2oT/8ROupJ4mA4yoBNgNyBfqW+VhvRXzS4GMV0bXGy0ca7PY0dhLwd6S
4hStpQTzfMphvJqXZgy0KrynT0OIlG7lkkJUQ7LS43+R5Ja6QxUzaiLcXGg3pV2o
Uze0YBDPNIQ71hjcbsBNnQ8GpCQXZibQ5aYoYRU3rGc0YUqwcM30mPxIrQnR1/Hq
MbQ5/++2TfMpPBHuotRku+g4zOjJz2f8wod/9ZpJiHzAF9Q539VCW0+l8K4uND5Z
xoGMk9h86+1mzfRXkTFw1OJPfdfKwhWefSbMPZX0ZcUBWJKo2/9gBK/SMyVHAmPr
hc5EKuB5iQMkOKaw8LY8wtWAWu6jWuoL6aOWL0XEV2eBQapp4kMZKW1k6x2g13OF
PW+06V+C/i53/SGFqZemFGylBvQG5CEh+a95a1lRKRBEpViNrKSjk6jJ00oXKZ3E
DADgYtPTQuSeLJuzEZE9LO3Q8CAS3i/1weH2qPeK3nQhe/Mgk94erWOSYK3hA8Uc
jYP3N0mkntJtq9T6DQyRc6Qjc8eU4uIlcpfOR3jzKUzv5cAXY43qloXCrC2WNh5W
t0rEXX6jGy5eyfAyOdhW8bYYEwGIRu8AIEChPpohGGTelhngA5Bn0ZpZtsPypr3k
htf3T4vQpup4RgP6F8+HVqWB9lgcxNVFDfDDJc8zAex6r93GNO3/hXwhhPIaVMcz
+/x5fVewVmllVapmND4lpmMmqbTIg3d1cFzlr8F3P3g18vKB8sNEpz+jOMVPUfxT
V+U2wiT97hNp1oAwAfuAiS/MCus7tzP2uTrqtpFlQF/nX7h0pFF4a3QqbZWPmVvg
vgMVkJK11wxVxY52eKz+ruXdunk+q4ribsp08UrP81wZQLQrzcToglxA58RvfWcr
Wmn3h4ZVjQEh24bfTj7IlN8eF5K104lP5LIMgTRlhWZ1VHA+vOY5LMnL9mARUidz
7v5biz31SRj1fBNRxTde+Bhq56OLWI3T50uNKaThK0+w9HZKW6XsDkuFv0amkB5V
hLfK16UsAjMhx/9nYYU+wYa4Py0wfF+zNg6a2OJOLLbXbshUfyWAbgIPCPm+6iNS
QCVHccwDRpWQnpqOsLkmOWhGb31wFNYVLtByM1XJ/5kXZTfgzptLBfpnOVlIJhNG
xkEO0wqZEUxDi7n8tnhMnbw29/JKSWse3J8iR8lHgQChz4aappDQCjrmcBimpE1u
pZBTH0F4kopqwRSoRRQeElDxqhI5LB0FPHZ1/uePltsN+0SPl/eRa6H2p6EcAJih
j7WmwvuxAB0ClwHuhfzuiq/AnADolsk5sIO409bpBOv9Q31Yq9qJvAUBl7ZVbJhr
gGDszDmdp2GRE1IFEjmoYfmfVO3ydTcDr1u7r1Si8dZ5BCk08LDTxstbAZuScgJE
4Scg50afk4NQ1Fqji19KC0Np0WWsozPUW3lxS48saNqswJdmBpNU50OeAbI6F3ab
GLCDVSy4tEsd/I0FA3QnuOmoH3cl/LJsadDGTmPByGJ8qKiQ+CQAqZ3e6wQQZJ3m
KlHFn0mEbMGFFGEMUmMUYMCmIjz2IMteOYIFmSbCmr2+Ib/Fcwysrqo3BbfuZX0r
UEC/6ROX5MAvRrnbuVaLgB/OZY5HlUt0TO675FPwPW/Oi8ecMq/npPK/bM5RwKuo
Z9TsMGJAGZCVMU+gDsekVzyqrTLnfx+EClWyIq/4H+acnMbj7K3r3/TL1QOfqlSm
17OBQqu6AffqPe3WsTi7UsPVQms50xW9a3UdXH2dPlbIl0zkrJYdkxRyr3H8qn0b
swhaYaM8jVwTRkBA8Tcyc+zm3mXlVcSvi8fHz6US7eHFpf9fY832HZ28O66XnrI+
1zJT0oJTRRVEiNd3GKbCpqDz+o3St20GvdJemRVGGlCY6ADtUh67Tb4FsX1ZwDRL
o1sH3ATXsyotjf6ipaJuuvjalJSPxqQZa8IgrxcseKDtYI1lN6sdQ6DcqbypeeVx
9f0CIEGcY4x6lkVDwBltvi3YOJLsCRJPDX0mH7/3F2lFSYBhbCclOcFXIRMcv0A0
E27JZQfsm0JWs00HAXq+RKAAW9uV3g5Vot7e7wKArgwdXWK8juW56C+wgNnLc5hz
YkgMO4ywRfSxakfrfLTW7KuyXi8FBlyx32DcU3Ekx4Im0xbq354vB6bvwV1V5Y2I
kStBZmIen/yJx8NjRbes9u9aqNDYuKRuRzdRvq1bxQfa+HLWiBwyFrDvNTvFreaS
S5vWSL5PoSTznMy+Ek5nHF9J5NbYGHW3IMHRU8F+MB++fHLngz1VIZrE+qy6PxXz
1sSm1FR5sT3A7zAW3Kyullu0EN/R/rqsSvubOjuHaS4d8IdEPPzjEb4VzG1pqDZP
xAS0CfR/husPItK0S1ftk3PuJoHW3jztWTUYtYTYWa5rahYSoDXlrr5QvKh5bd1v
9XZTRxi0c7ZFulQb983t1gxlqrZJdLQ7Qetl9lebsHw7crawjOqf5L9OKzQ3uCmc
yXKZCpjCflMBJ4VEICyarrEC/UxZMSH3JPwFvhMYXpN6JfZvhNJ3RZRTYtkg2wUm
GMdvxEmN68q3XlqbOxLTmrDVN/VbxNSXp38tCcrbdztBwHKQrm/1EK54MyugGwty
MO8Ox1NWDDElxAHThq7XLPvr2SU/rbmBkkJ5S001WDp91KjD7LDaVLu7rOINz94x
/g8yioCwcLOIN7awjo35TkmvcRfDNQ95OePCRqWIJqY94mjumJTDBcgwXiuANAFA
qOecVa1DlXZHIy1aTrDCxEMts1KsXsNw58ldZRZ0iUpvTz9tqRLj4bYQMiw2J/pC
yQIvDiLPqpL8lb4hSAUkz9Ez1vbIqrpdFSwEGSC+1L9qOUUVlXvqbvIOr5sULk0d
8mlBj3xzIcblSL2skP7SqmXjJKqscmVJ461jvfeoGRL0vV++1ABRqwAN79ForDh1
xO7Dha5yzPveLpwdhfEgXfM1bAppMtW0BhaTmrhuXcjR3pMk7SUvJuM74XV0hHMX
YMXcuRobpYZAe4NQZgVlu6+56RW0OacTjKhtAELAaW//s0H6AblVfVYt7i6oHzYJ
42RBN8iEK5IZnA0tZOBfaOdLEZWMXOcRs6ci5k7xkBl2x6YeSTGr9OZzq6SK/xhK
sbp8IUVZXA+WOcOWEN9svh1QYfhDMwXQgWnRULoWngx4zDpVOKh5mbMcvpIVl6WR
fE2cDQeJEhK+44/nzpbNq/dQFnDsV6B9m2q/UPys8L6AGPxnEvqWM7AoAR9fITAV
Y511sg0ieexGywRqhhkQ3LcwCiMDMSNs1A1HwxUAGg0wR+w4gkIW3BMvqjv99Sv0
gJB+U0f8pgF14jt1XLEu6m5sV2sp68tDuqdlALLobY3V8xoEQlkqyhopvEx7EhKV
4eLKxR9ePfVsde2s3X0fjIOc39yCbM8mcopkFhwLGTABSwr23rotGgMhRw4XO7BA
nEb5Q4NysK675EkF1PHT56Coqkq05F4fKlf3DlAxNAb226Q0CF+UXGWQwigf1XLB
mHDzKkDztrtZbfEZ/megRaA8GHEcAipWGrHNd/PiPzv/I+eR/Tzo3NW6TfWB/dD9
Y68EYHpispM6mE0Kxxl+7ax63BtcXkf+Xf5AuH7p6P1NR5HAf39vo1wovzVpkLTG
BRABG8sFMbpcvIJOSa1VvaW1Vl0/W6Y5YIvEhn0VJrPWZQQQXg6LrXPuZJTDadqy
m9uOLgZ/k4EXOzQxicIsAQFcnQ51aJgghFIQLDVAvgWuANxUXEebKr3Bs3nttusg
N8RABM3QXSVx2VNIL1hNxqhN1y7Fcq1pGBHnOselb1Ai5OWOK6eFuZyUmIbQwuHD
snr/Pl6WolOEZhXSP7ouGIXNinkJKnYO1Fi29jNdcGvod64w08T/lbC2EJArH+H0
vl3YNSJ0AYlQ+8NVO+C/QMYJe4JaWeE6/weKVr43tQhOE4HYOfMaGJGbleWGVIQn
32I/gAQuJn93mLp4tBkymxd521TQyktwv8tUVGuD8M6CLU0Pp88Wwln2gSmGtnIq
930W8A1/ulPi3LlH1vqxJ0brkygpvGVZjS89Vy3ED0lpxyZZp66hlmOFpR5sQEt6
rlLQl+w/o5LsYMrG3K0JpETWvVylkcbVormncyTNRP2EaBx6hR5YIuBDslx2nxHm
UCMaJ1cWcxnihWmdFWEqBwjHzCuX9KYOL4AJ00UXQMqde+h0YwgyRjDXof+7a0pr
iq8oMh+WUDjKM8xzonw5kh8zy/J9OtitNsXxKE/8ty5/HvHmWDfjMlM4BdDitC0q
Iy4YtsJVnyQnhzY9t/ZyrkbC7IFZzYWkbh99wbox03q2JeTG686yWA89yqaVDnKm
x50pb8Kl9deF2wXuZ3K0cXYYZX4rG5JPiSUUYlTr1GZBNB1ixkSiKk79Bp0AkaHL
D3oOQiXeilLCg0aPge9lb4QscgQAgAP8r2MdXt2hDqxOAcjCbAabTAQmV12pkFZ5
GBqRUNznrAJv0eVFxhPT2MFkp30Bh/TewmthjIIF9M205x65Uwrt9SCiLMOmoIdu
1sST08fZuybtjY80zJvlfVgOYGC7nsulk/BEWUI9Mshkx2ZU6yDUwkvT0n96vsmG
Kdu2h2FWmH0Mvxd/lqdhCKTNZ9Ul5gPu1sMtleAZ1C8y5z7SlkZtUU56a7tEzqoj
HSj0OImQNUL2BxspMW6VIpbfb0dLVrDu9cJTaD3ClS5h4Ux3s9kKXaW2tke0MlRR
2MRB/pKDyz+Wliu+ZhQ/FsZ5pFV3ysGXb1Rm+NbZzQlliRxXPUUb8ePzXYPg0oOj
8siqnqBDKclyJjSYd1xrBSPPTg0QXg9gXtCTeI9l/F0vasouUPYzPlFQYC3LOf60
bIbGh5WWyXuaLgImZv1pHv2ovRdCGC1kJPrpYxOETbwylURDH+V+SvU8e5rS/Rqc
Yzjc9JE1q7ak72Gazk639pY4qp4XibMzi0I8FK25sibt/1/lK4lkoYEStUOpF+A9
Wh17asUl1wyfgjzn4z5Bi6692/Q5OnqjIodExqDQFdzZng0SqphqNT1RBrEHcya8
ioYpinTgtnDt8ykWAwFVJhAPkp/xE7OZSWew1KxVzFfb0AGEINFGDkvh6hnQvI1K
hfawBThgX/RaS3tKjYiJ7JylOplLxp5dOLrwWmQEXlicP6XQOiJEr8f682CLl5Md
zGLpJycHElRcOBiee9QIUyDIP89H/HVeg+kBEizPFEOBD9wzclAF/MhpPuLVDFyy
/wUFOX563BctaO2spRzkIYQd/xc/3NctmG2fJP06Rw+CyNAuN0Bht1DGGUZlsxgF
SnafcpozU6bROaWsZewnKjlIPdsvuVEldtWqjqAGDvEMhdi/PVs7NV5qz/98SJVS
9+uCLAfFnYtYh7eZRxUCUoTnKD4zNMX1kuj3zyO1/BgtuAZUthVcvQxDCNRMi5ba
9Vt4bJIynUeWyu3ssNCjBcI6VzCk66o4hES2viASn4Isb+LO463/HAd8AsTNlTax
8acXgS1YrGmF6djGwCHQ311TcXJQ+bYYB65rzhMhxXrKu8hLmuooUkIssQ0/N6zO
x4wsZV040/8HuKiskDwGlLXWqhWlq9Oh6DO47pEttwHwpY/HMnLSmjVT9HkJkFWA
OWLsxiaLPbqJIzTfCk0AR4NhqF5YEXegDaoB1V6W42d85SHj3U7321cFMXDVWBWV
Ow2PtPYYQtXerpmsAPQHunCAffk4VkCY9u0ccV3V170ZHkroR/S7tBNsiE72Hn1D
zPPa9ttx1gKcsFLiJvwQLa+RRfL5txnhSEuTXFSq5nIofK449BHRibRX5AB2AkNi
dPqyfrZFi/6pHVGwN8gBxVLwwc/G8/IXBYKYIRIGv7AebmFVhLvPoPQRYg5TA/Rb
Equ53jt7MHSeHq6b8wAlmtqwhTiccTzG1a6kf+PALBRs1kvtppH1Yzkm663RTJOo
wW6Q2c8R/JsvAXfUM6ZcYMN/s7kCrjuiV5GVS25zeaWA4CSz4C15+4CRCPuG3CCi
bC8NMXtOMRltMviO3p4wn1XUPa+XpC4QeY7PSSKNtcNO8745jqjmWR13MEcvC2UJ
rxNrdHcISaOKcBD2EU/Pk/HYqHWpztOe18zo+uDkZmUuh6oBDMBo49jM6aOHm85N
3BBxqLcgjVV3sLuAYQ9RAaIHggfjqljwh2HHZe7+RzcY3TWJQRo5XLUSsX+At/UQ
x9TUdKxEP48bCbVNwdrc2FB8+BazMN2oiyxSeb5gXNNX5DYNbQh/X2fGOZg6xYQZ
tEj8d9xMW7RVrP1J4gUi7+gHwLPhSyJLwXoqL1OAE9rKpLUdNuegWHq4ABLq3u6t
fByHPXxVR6ZJ3XgmNGHAEmMACMvri6AGsLJbHaabINJVeFB/1iYHHQEcgO+gZdpg
uh30+e9Nthk8U5CGMhBOHr+8cSroklPc52qvu+h+vg2UIsxDpEo4Tbt4e3ovWFT5
ANxiTRshnTeC0haCop9r8SeXF02H8NlZt2r8GXDMazyk3sVaMZlkfW5rKY+hdDmv
XdGUFFo3P/wacdlkM2Ro9msY3oyjdcFoPRr9udCVyv6dkarYjhpIBhI7YcoqRQ9O
PPgGPvKc4pMD/6PEkkmEHYqeO3TzFr2fCHaNfUSgTMuU4UXYLcwFUsag8IAB6ont
MIfdX66zOfwAzCjFZiLsesFObGeZ6aA7KbgjaSWYwgEULQKgsRxykyze60ldz8jv
MvWMzlKAc+6wQWLjD2M5Z7VZUxmHMg+kGMLFtz5xf/wvD0P1EqRkD8Tj36jjbzoO
2QfIfHdMfDtcATm/80oQ7rvXMHjWRhJ5HxdxwW6a2zViuziO0cLXr/5p4n8eujDz
cNleEROrs+yXl2fny3vqTrOw/Lhd5MVIAUSSnVfPnssY+r6ofRcERyn9BxAQShFP
EagpVRBoATqRzijHDjfxMNMXlnIa1SFwbNzOM+LnS7wYdyHseXEFFu/TT9mQnm/f
ia5Yo/iGdapPI1G9HwcBQ7dwFGuBKxzBp18IxPYSvPn7YkLiFzqfARkNND10/lJ9
w4unUknViWRgt4M7B47Tep9Tlyd/933pMECNji5Ri937qZhqEOJyTcNknZZKXrdt
GPmAcyicd9SbHbL//+x1MMe2sUX/jP4N/NT4QUt2gEEFw06KTbjmeMPjzAkx5a0R
ltmpbYvcKRlnscs0PELI7S7fU9/fOhrq6Y2Lm2xKA4dYkiyuNSeia4yBWCYGZX3m
xySwQmflsq5k6F2EBYGIq1N2gBg7ZkVRG9N76eMPtMrhIMgJ+fxQZWHlpsftwp98
AsSCRSB+C5i26OjyGVMq6H//p1z9+4nFJw7cru++tDP+EltgAUrCCHLLTS2IrWmp
acPJ+dnUQuMsz2PO5aTC2RlEvQhs7hB9q2Cw6wmTl/zIywzAEvUzQdYWG1oU3AMV
s7FQzJcI9xXejRb2uq8DLm0LkBWXZm4FVMhe/FWV8KkgGtX3DKSJdMWMYZV9RPoi
v3dEnmdj1D4d4uAa7X7vrvoD60h8qPLfW0QAXAcovDdecIqNfLjZJ8e3t6KqtoDC
zNOy/Z4M4rWn8NFFYHrjhu/YBxle4qgK24aXVjYkuf2VwEHidh2x378+FmUsGU1P
gtRkrlZi8d/yW95QjODb+kZqYtMcYI/op7jN92XmAfDYylgxqdCsTwe9PfNMUDxw
INuuoeDfXqpFmTuk7nKCuzkH9ZsAjKtnjWCbnW0OWCuGs3iJ1+2Q4xiQwU0omeMM
JJXQ6xmZdpWUrUlGbOQlNsb+xBgd87dvszO2/s4BC+a37LKp2Fgn82d/lIRMCiw/
j4zkW47K7FEkfT9RdfIUonDQr+/4Kgh72izVYEXxgG3pXST6rqQhBmj04WM6ghpS
FpYCktHl7u8yP+kHXvhtBUnQtpnWA6m/Vj5RgH9P2EjXELUpA4Nki4u+CklJhp3s
XT5Q11zvzgQaYCga6wyVx9Ju0A+yeCznTxJSuLpZf0RJ8JFPCQSbr2u5Ni5en0Y4
JE6O0qAEOAfKPqsKPxeraegPqb/kgsZy+SzjCzPGdFgRvJ+vVAXZFeGOmfDfaYC/
iOmiU40nQbSG1/b95oSU7YSGwMd9liK9ZpDRe1ohP9EB25UUBk0G3OPrEOM1fIpS
EqbNmHI4A/cEK/ugMl96oLakMvgKI8l6mtDkKi1HojkFkmJfxRR6TzrSdURAOphF
kNUgsfRFVjsTit4p9F3+SXl0WaMQMdZYNSYX/D2W0sdKjKF2vDlKDUEgpc6VGlQ6
uu8i7SbAvbwHXTaba/a+wEHDzh3u/UZYykULxghQlh5ov2A14MAAwrcr322mR5/R
dr8AtV0ehWXGl8infvDryqgLnhZ+09o1OlASb7rzqqseRepximPvcPC584eB+Gjr
6sBu62cIZBlG5H/DlqQV+f8MdGllnIV9XtkdiQibtDyIvElGv1r9xKjhGwTvsmdk
r/Ght65RoL8IRTGdZLF9MqvTjcH/FNjS5mFvTPpCpx6tP051+pU0j+WrW4E+q0GJ
IyH87rOw3ee/u1a0muBBOKSBYT47OPjgbxPhrFYp9cL84F4fbobdQ7NwhNn6yDDe
m7hZB1DXPuC/SbwHKMQOp2Zrn7Wh/4Y14ExxbiMiploktZ3bZEXvFBwNvvg2U+Un
ktGK11v7D0MC5tukjZi4LMeu1/LlC+OENZczHkUotYqBN4xIpUZ5vSlm8h/BYmJj
Tj7TgU1c1UHMfyIl//vpEHPn+gN83CX/hRBSyDxEDb5c3PuIAIpusGgCzUzu1Kcq
3/nWXufPVa5+E3nmg6Qqt/XNU3yAALW/TIyOR+K/BN9TS51zGrbp/cPtXtQzOfls
Wf+gSYoniEMIn7ATd9e1pKOn8Q773KwI457G4Ymgb/vHUatJsiO6RxnLfFz3Dmfe
xotcU97PUraSLoXL8rygsqoZXf0E/DhCRztwESpNkPDhciv4zflQHum9bO8lbK5l
GM0ji+Qs+YTC+8HVHOwS/USz1P7ihrZaB2dASFeeDExBMi002vATKL7VRgmDZ8H6
7VDzky5XN1Q64Ary2IJn2ttQnXwL1Vk90yD/Drkewt6S/o+1mHL5ffWcoqx0e6gP
sDnWWNA2binbVoQZdHKgUgFadP4leI8IqQHH7ln7VI5ZyKjlZuba7PVeeiUJkSML
/K0WOwf7kGGE3XrqiRfmgRyOGQ8nNlGUsOQlZ+E7mm9vuvnkDt2deCZfeOtCBB1G
0OYnK3Z4VkciOachFchUxxvsywAJ3fYzBfi1a28n6x3/toYXcO5mEJtA8d8iYQ26
wLyNGJr2XSY+a1Uduv4KOOmTZnVzoC5tQjRu9IIh+Uu02l5Mku+vF30eqErf/5ZO
jGLp/M6vS8FvM7LhGdcfgICBXCl/lvW0jkJ7pwR7etcaZQhovMPv2SXFmRekUKer
cw00Bo/WLPG2rNm+ncpJVeenEIUAPhiOrLjedWHSgFbMlzqMGsB/R5FWXzLbNckR
bgoS6AG9UXowu3T7Hs20GmPN348TmJQIoF7fMtHYMOpvyNqb17sr9VTyVGdFJqFz
P1tfBIlW2ukkXv9Irnth9Ld1A6ZZCGyMs+idNJy+0b1h5yDROXYHQRNbLcM1s6QE
Of5O2DOnnikMpXdM4/zwgbZasKu3bNnlcJr9dTyJj+QkBP7XUqfuWrZo0Oa3SaRX
oIzd6CTlN50Y3SzJyPYAgFUdF1x1AIBj0rkfuXQ4dYXatwZTWoz0dm94ABzrdbB6
FwNvAUFcVB0CWqow2zyTsiFPm2MHCcTXTfJaV2tFBLTD+oy4TBpnqgxz7Jkzoc1+
THpW07aBzZrrp5f9hMXoYQaaE1ds6PymSGy5biQoJN8FkCJMYOwA4wCTuy24Srv0
gdEBf04MeN+YThBYUdcZXUhzcLVgHrbWRp8L91QbYijOPrTZLBpfoIxVeQWVQSGE
xVJZLXvYlaoH9TsFO4ROyFG0UJFJ+2lKc3nLIvdLwL99BFJjXEn1yPVq3Hh5etW1
oKXMffSbEafSnUM4eDoMvc3QbB5YGEBJFRn8VpdpbaGvw29xd+hdRY/vrfAspIKD
bNOsi3Iolnuxjhh5OZOpcDAR9bL2WNv9l72/U+uHnnWegopKUdOsiu4UhQLvkl0N
MLRTqeetbxCeAMRz1GYLLiCOfLeVKXJTsXKdVNv9NufNzQPZmVWm+kdmTe/bwt8L
9vaW4Mlmuza+RrEvVWYQgHipMJ246sTSJoC9IZm81VOjGyLlorRPDCx3tNEqY8PV
pSHWt7Bk8z8kJ5U32HNqXyu7TrLQPAVlIpopwBUbaoFsgdxSZQwXEkYk89f/ko6p
Ota0EgV9fIb2GnvQ+oH52yuTyHTX1Nf9dZ+BDBu50OCbtURDKNbfkeGFe7s2H2Cf
ImUrGJ8zYxlVb4dJBHgjog4WBTlXceMCn4aJdu9FCUOedVhWFatw5sIvnTZlt12T
9bTNCYqQQ9fpvKhaKbdOQAlfpteBe/nOh0pa63FZm3VK7TeSDx+YpZQJT0h4MH3j
DS32AbQh9cD0GqtM9V/xpwEB/J53781cb3zZy4VGwyZAQnB3r/Q98oNSQk4sTcOb
EGTxslbBNIejNMXm31Gd/brBiLb9fIfKxwai7KkG8EtqAzUMazVGUItnc8F2nLOl
aIjn2efLglW2cRmecWqUO31Upov/lblw0yd8TcYb7dryjb79M1LN3Z8m5SKQB05h
CTaf+sGoMFBVKjO4t5b7txOHkM41K43vjlMYJ7+uNC7yO1Nlmjk/PD0+cRwyK5Pw
+pVODrURqglsD5KUC9GQ8tbDevdJk8j5s4f8qj9nt4DqOsIk0MU/Nrra5qYWicOK
JoW92yGEex4A1McxjL8LL1fA9BvfTVcWEaY2Sz7qip0Bz2ycDi5EM1OSrljv3wwy
oXBLc+FpXxuxZcRvwzbhuGNXzirOUS3KNH3o4arc5I2NyKgJI0x0GvaZpBjmgfy0
AIzTlSaN7mG3IngtYs0L0GWaQLeXBhp3wycgUGq8hzgVu0kP1X7NHSAKvJDNDN5V
ePUlis4Hb47wR8xiEI274bCCGN9LgZwQqUxb11Ru6o9dmnTRksC+6d/LDyftDJJU
m8+jeD68HIUV2+ccLDEG4XRm9vhtlTa4KhyueSApR9at3K9Ra4lF083N7GQw/pw4
vAZyp7UWqDMBcuy6tWFLbPsCc1yMBD0I/Ur+IP9rP3ScQ1JX/RrVioAZgkzAOivf
EmT9veCriJTwcliTcIPKCubQA+rP9+jmAmemBQ/Ubar7yrQPVNh6HEp2cNjV9sAy
TvKPXEyRJla1hyRy2bxfPOsQxamuhQkMSkYVo4QEK8b+hdZWHXY4p6jC4cXskQHr
MKp9xKtk2bujCxr7cTloEXkXwNO2QRy3kCIKsPshphpEhgT+aeu/+7JkFKDg9ig3
23KQtjEn4piy5dsCSMFaTYqm6Uy+8CtIrbnIM3diRyH7ORPuWle0emCC4+taCaPH
uyaP8KkrhuDSmoBDWFG+NPWJukmw/DxDBF2HbdH+s1zAdTc8cbGFw6ssVaD6cN6U
bUXX+5o2d+9ROi9uuK6/aVxLp10amx0ESCBr3Nzg8tZPV7ta4sG8Rgr4vi7tI1ji
UC7VK6fAXE0R6tOrg9Jp2P55iv35a/vjr99zFqNmw4AEG5MKWQE+EBpznef5eZoS
/cKTwpLbDAvWAAoV3vxJXIL8OLbGBg1EkaY1WlLlACPlcLXUK3rgRN+uLVY+D6ye
m4sd16MGqKUXzsTfvBLW7+Z/yyexQ3yfj2abVMaYbgRYzjrCE2hlovrHnJx8Jfg7
S4ujJYPYVpovPq7mQbu5ChdNpVGUCAUf3XBQC/1Af17zpuLjH+ePrUyJCQMCXb9m
2XdbhDiojuL+U3cMUQIuJEu3JA6IUZC1K1iCmOm9WZXSjJu+anOftj5d1lWvgUO9
YxQ8ovUwDqnbOOp6lqOwEjTgh+J/eVRFxnBGO1DMAXrHM4hJ+lk69EdQsbpAkCBy
XyJr97NND05dXkJATC1n4hYUifQGyYlIJ+ZUGuIG9kRbnzUuT0jGqHCLvfWBSJbm
mM1ILsrlYlvRQg/5Qtvkb7nPMW0LhoBSJfErc07xpNewhHuBKmBbe55kcRbPi19P
J+claDRk5O9f7bEtcKnUvXNp1VqvsZY+kPEXWseyo7AImAsn2e5mdVhkNUF3B2Yi
gfbTTR6Uv8oWBwXNgAA4cpc/WgP/t680EtDlsfa1Qym8UMKyFRCa/tEnISz8CBfH
svzaf4Io/2yZaFeln4ItAu4u5SfFR6LEcH7z5o1seB+LOX10BHb2uq7aQrbwXLYs
H6FaES+Ko3iyC8/7uYGzZpVH9vKxFgpNLoB1Gdlm/wPgZrkZuUbArC44/xq+PQQM
59QSTK+wzucSamhPqYjp/DRazFO8HPZJn+WlKAeGgLb/O+8gRx1QwoWmHBOVAMLU
ZmAR4o06h0n2NwkLTMTgsOLMmKK7F50uOSi69y0T7xmHfz8i/O8nZ6ErC2KCZJPA
thm9+vHfSDi9kOWz41OOH3JdNYWg/GAMhk40DCDmA9068Ac5iwPuzCDm2GtUakVZ
LrCHkVrmHXpS4PK+PFqnv2b2w1zTWuuLvImXlTa8jrTmJHCGVhOz5998t6qRp98j
KAYDLSq44iJppvCLR1ynK8HsX/jeoz3xfNob9evh6rYfh2fyGHoP3b5HXSaawump
7pSv/mrm5EIZYJWcGgkJqcy7pCHlfhDz7vd2DJAeztNglu/EuwVgAPmm5S2t9qGW
UvmwNH8gbbcvq2clgl/PoNtKSG7CkWlhDPnDs6n1+nPJBwqstgLZX7GWCQIYaXPy
ZP/CMfqT15ItXFKdyr1Z0G7bS3XrhofNLWzvVpE/W7vtKZLrcEoHC9Bn8rZgxcQa
eqJ7NznBqMLnNrrudNNXJEZIhZMujrn6zEwHm82WJ3hbKhH0n4KGWvNZ+NNTXvi4
qEGxdqu2m/JmK0EpcIjIEwuLw7Ai9RM4gI6lZyfIK8iLieo9j9TpH1Yllx3bwctu
T33U3qgQNJwVXIrB96puo9IegIaeZP9CP5e1FjMVEDPVZTzsrf8EeyAD0BqSqfMs
ji22feTlHqxz1tP3Qk4Q8UPNJ01zlBy67rWnFFqRTxlTBhCjqEklh/KvPpzvFBrM
w3ove4RAXyrw7btbKZcGVmupMuvkBLmwxp2x3vTRagKX+6TjFpnVaeKVn9/9/25F
Il6mScRL/Dn7qXfMovvaWXUOdLwA4sVz1T9aNgJ/Qvl+ybu9+H2RDqX3A1k3k3NG
PxCazISi/gIDxra62x9UlWH5ODcYOky4L+f6KV6qwU/4fsb60Et/i56a7PvMyxS9
DarOw/WFhq1WjNW0xr3hMAwKOk4rgmuGqoZUoOnKOUtyM3W4sMoliMvRLZpEPQfK
NFGFB/LBO5k3nLSzAy9Rwr9bdS1p2/KSlvfdHkS6BO1pla8gg9BaQLFxfMPTh1UR
TLgh5PoPWviaYX8+5+FSZwnxwNSS0M8Is8gXaxh3sOXMTXVY+J1W5Dsrx3xeozzn
7sPA10xNKzNLviNXZTfuZPCIL7rBYMFo49AQrSY3vUI1bYlTPWFZnAzpV1AUU9ra
XOvqt8j7Jk4wObS/Iwm0ngY3vKgLiBAIJXdQh4c/K0suNhv+GW7PkxT6CLnVB8S5
7ofXo8v4hjU3aVfTfUgnbafEAbKQPwKN4WViodJWt7EYMs1VkmUPwfsbLot5HBXZ
WxmuapgpxJdRo99fhKlDhTH2RjPcv7cz/oQLYygK6I97uOwBgtnxX8fGe7xzfC3x
TPml00O2j3aTm3bQzIYWOKTkCmIbpx++QOUYH29tgt6hn8SUgTG/IgoI/IH7TLno
Ro5lN0bGE0aEjt0SjZBVrgZN37PSe5m6WT43VjX0IPzECRdbIM2sim2CTBwQOGyx
/GVhFFu8/JoWmxBpmho50awMcP30F7knWUUylkFpFV6qIyjoxLd399da2tuIGsY+
9X0OESsvl3AXgoF3PHgV9XEfHFlpSje+IZgpy2G8hWi9d00lr5lgAN45P7p1gkWA
yAnQz7bLmn3ArvlR7KazuM7i2kLiHPUDebqlxB8Eqgk/4t8kjkglZ3BHdG4eAohq
ANkj+M+BYI4bMrtTvP+KU/ORstAXyzQhpSc3VulG3OqGW5AhcdNC8W7bBjMAHcd5
fgHLIUZkVF0Cf8ymX8b3meNJubdWatKK49iMOPYp47IGIED+24rRwcE6qa7c56jw
3X1O4ocjs2qWzZ4bTmAeqtoHSqkMiVslJ5jf84pZrRvYzJsXQCQ1ctbUAy5xf9Po
I0e2WLtzJBLP/CbjjF1UyHFrlBvV9zTnZfBNrj0SMx2wrFwyevp7YVV4hbH3cXc7
9Q7Lqks3KiiUG2tLsJ7FzKvnSUFazwE+2AUYE6sjVRQYO/mmQxxG+OWBi1Rgr+9I
MdmKiqDcRSFLyyuAnhxc2AnCj0QZI8bjJ2+L7x5Z1+yeYAcI6IrYB0fhI+hefGcP
0BTJbzW2FLAX2iHM/gn8VCYOsO+gLy4SJhHgwwPw52DHJhN4PVYPHCgPhTqMULdw
KRzagtF0JoiCxvtEv4Vw+4ZrxT3zhhUO55ZWPBdmFNCeB/aB2pujTOK9oRhjSynZ
uw+9MwUxMAxUqEVzI/5T7qq9rM4s2apZK/uOekMzIW7CgF55Te9xcOWVLB68f4Th
FKw3QagMgCMopdymM/7lcXnm+Jdl5qQe99xBzQ5/ZT3VQr4rnDPOB9do9JqaS9Dg
/Q6aocA3K4hPKJMSMx6HkKw5PtWZSMQhPdmNzbskdgdXbEjvU2cN7LkJTi62sLwl
Ghvo2GF349lnwbN+CvK15Uhz6nhZikEdT4ntLlNqH4egG2MfwXEkmE8Bd9tFH0JJ
txN0jKMMVyrlwLo/ujdQgx0XO8AZv73t5xEAG1+YgKGCzAlwjcSMS+b4OLKB4u1M
M89ljO40zZwW0J1LnP6VKHtKwC+zqQmtzeqQ+9S8PSndbcLIS0F9BvDwnfdEmPXp
L750nmoqYJnhbut3wjhiyY7E/G49GdvxNmJwkb0pV9qBfbtRae6hIHoIRAr5lW4F
usRevSYTZHHhubK/bEvkto360Hx/zI5z4QhjKN1pp3yPu0Q96U169bWWBIykKtLt
TlESfIwQLrnRuftnndyuEu0KZM36T5Wk34wTp4yNlHyF7kJmYUVftO2lETI9l0B3
C3S3/xWGpDeYpLDyxLXgJh1FxMmzA08YvGlk57TfO5GpAUNDnznQbQ4LViol4EoK
VoeofGkPZfV74vIKd0FT2HXr6MEXxWe9j77yZAJje5OehedPB7vOS2tQShKGpJwz
oVl09qPu/Lt90n10ECRBV6B4X0QbHuWJQp4sHNrWVC93wE2yyngOGdksW+j2wQC4
z8Ul2VsghuZfUD3dSbjUkOxtpJSLlR9+mjPcFcNCCHTwrJs5OkdpvUEd5ggTm3AG
/QJ2XvTAkPTkvwofprxjx521x1txjO+rmzN8xEi8CmKc2SKpxkI5rtXm3tCUFjpT
z32FyNo2MQgYfG0nNiwNnccjKo1vOJlgmow6dGr1+ooKTLm5WHYxdm2GdzVzZ4XS
E2C7RdCxQr72y0ZxoTMwQ0fnaRqPg+yzng3tB29735R85HifDq1zeNXotWSrYDEd
f5k4UKTQ47tAGhWUocHPKlFYz7NaoQuCMBkJGBAcy57HeEHIa986kPZPFT1asePl
4i+hsRROekKWCAeDMzTB65UZwjVYKJHZou1H86vDpAwoHHlhnBJ4KwFW1NHBWfRL
yHBaJ9j7uGy96ojyeL4Wxw+E5mkBzPemYNPUX9CSIidf2t18CLj+WlKMHUa1CakI
94oyYoMJ6KlQo31yjlHVFn+45eO2xK1vcoUU4qMdi+hFRySFwVzD5HTqNH75l5qZ
7oiOTYrj0rvKnKx8viTHmk3olQEJyfE+bhTYHqY0FqmJC+Ixdkeqw1XozDPMh0Nq
r2SAB8wVl5kpGlh78ItU0PQ9J45ro9W4NmM4StESgnqGWlreTRHhiEVVxnV1gFl4
rqokLQFVHvCZvpNGCvFiAJj0rS6aUUzlYs6CWh+ymW5qXGWPksbbJ6g/bEU66GzV
G5mJ6k+gi4JR+YDwuMEEPC0xQ264+lw/XgIubTVgpmpygwYFLcruXfqrIeS9evGE
U39pI/2HEE/O2fIyV+UxYhEsQHQKRgDGqZur/s2KJthj0FPCmWfw4Pc7Rzp7ndTA
4TpKtWxu1ujJzxlY2zlzY4EumPHqiAa5oB80gfJChk4SNh4lyRjQtdNMdG1eLtag
NCLJUU0fjgyz+8FBrlCqrryqzVKV5H7gsfnhTch1uErKUsmpfGIyj9fthj7xCyiv
mwVO9LK8G8QtOMEz/XWJowPFzmOeOGvJHcANiVGiyGTk9MstLL+C3Jt/faW8r3hS
yPzf6NKpa+XEPr3DTdk0QDGo4WDAx+ofRbViMLgNzaIUMcLfdXGkL3kyRvrTC7WD
izOmRhgdsBpHiNry9P1o+3llopnKV16wM57Aa3kEknkiNarohe0NqWUD7wIH71V/
aXdtR4kmkFkJ/XwMbPmaBL3PapJsYjMsHVB/VuGxN9QAuGEan+m0kepEHapDh5Kd
YBpttwEfJFo3RmI9h68Jb3WkLzlWsySGZpBrYIPA8RBkwCKPuoL0GdYE2OT46Tpt
h/W/5QfiisticO0vU0OyOPlKrxW5iOyXmL7JreHN2xYEpU+G4LGPW2ydtxst3X+L
mMvSLygkb6hVsoDUWQ66blHbUJlx6q2wfvtBZ1OfwgD96rLpHnceUaHPe6lDbUXM
fBsRjlYNHtzydrj2jVxoE6KHjqSTWX6dnqfgv8IQnHwygX6PAHxVjP2Hr6Vo3lTN
4XRfqMg446PdN3Hfj23dzBfbqEZXSiQy9q7i5puLQ3LMc8q6LUh6Rl7uACS5qaND
m/95ZuvE9W0u2yUf+wgtWTb9UkMM+kJhG1yD+HC2EZ8dRYGOlHw5PB1xExAi2tEb
QXcZgshR6wJuLfJlE6JL949axTFPo0raLCNiLhWIvsnHzopmUQBpwoxtOlaiaa5a
zxzmS/9mEXgWaKe/J7eHKQdNk4seEwM5cWD0TKVU+k1z6ObatL4scipud30IF90C
xfWJB9dV/REjUEe5CJjiFELUSIAw0w6TMc/nAG4+BwAogrpXwWTRWNqj3JPAdi45
l0TkP8g9gHCcy+vFvA0N1U4tKUgbuXvQ+q5e7wcLFL/Vyl4FN+b5gcJIc/PGWEl2
s8hGLQHupJ7rgKHQAStdJlACtc57bMYN+rPYbhq48NpKoSnIYD0kETTAuBo5T58v
kxQkgVY1L+MskRehrtfTrfubCcueqc5N32OuPDBBBjh9m51MCMV0IhNOlRsc7uhG
yFhWRUGohPz2hXXfie1te2mTqH4NT/FTFk1fwag63WtWhGA4G5jUWxxxIKtTV7qT
n66gtbI98u0EEwjfdVGhg59CCZPU/suyTRc231MLb7hNU+01YyGVgRuAzwFe6Zaj
FrYuk6Pn0pnQpfqQnC7XlM6RpotPrFo6gxb2jMc7Qgcd50+729radBVpUymJB8+W
ws5W4JlFYzKQ/Dja/EF3LsmIywAWtMq1sEZ/CjURYiBsK+4FnACIaQVp0V4qc6Ai
3Oz0oJSzCj6App2PQOVjY5+dQmFAuYt/gVIt0x1F7gFOiBlPLPjHsTb0Va+4AHVS
iElefhu/ipwVUQXzvOv7ll6G559c2jrAfm/BdK745nLS9KObti1HqsPfhJoldp3X
rksOc2Z0GnYVs8kkuEP+btu2iAM1HotSFY+vNxLPUnIwydErDBkNY8ty3+Sh8WFC
NHqffwM2U/mUTyQK6dxuUNIZE5N10dQrJjyw/MtQMitvxrSZqdw2N03mVbEVuL8l
1fRqLZG+Ud7doLC28oRnbugKNWuQysTIN0HGkbw1PTT0Hz3skBIJqjGYl72ZfKg6
KcmfDQAfOiE84jOA9xYspzFeVD+QFKq4EWVMzPjKM1kqtPgWEwy1naUde2Yip5qX
UUohEKRUIhpQAd29GyBP7Z6Kfbal2b5AahvybOiVdyG5IgUP1bjyTwnRIJ0aWc46
oEJd4phz0HMMrZIjZDDv3usQBgU5lbEE7DsLmaFA3+ThmkRGe9ZjdOFQ32mWICPz
u7FDpq18H7B08mNtdwOEEA3f04/jELfasKTkfwHaS5BuNLMsmdNUG2/2ozTGwH0e
1oxuJ1+wINmMlU9JFwKT60892Jg4/05+TT/Pvgr29JEpp0A4/hYDpVxh6VLjnkTp
OJcUtMGmQWriQffU/iUInMJe9o9l2Fv5khNbwBwUVGc6c5gJAjqj3ycROtVjz3lT
2WI/eGg3QM9GFgO3xPzJjU/8whT8c7K9hcjDfvkIatgzpb10dx7sWrOWbLMuGEsb
lypdFuBIU/qEdUGS2bCd8okN+2Aju2QgF5NLZ8sbFAyZHBEeFIVjlLBxvpciMcXj
kud6v5GpDjdjlZ9HMybHtkGXGLwtQiExEgmmwEJz2SVaGJ9PZIvDdI5C0bc+co/b
ebcPdcKHukfGtok/dCasKMa/e+dcPho5VzI1+uXC0gEVB/6azfvEijWvmBveUm4t
0Zxy25hGqVOw9+XDdhJxUtm6qFn1+5+lucFjIfK5YD6k81u88D9wlkTQ31PQC9YG
Z9p3Jf0a3TZktiU00o1e1DiiSk5jGvMl3G5jsBQgfMuBriHozIA6R8TqPzopfqV5
n/a/3hvY3QMi5CPplfoA2IrfSRqnmIWmWTt1asM6Gmmy6wZek2ghMFLvR59u79/2
mY/9txQCgcpsC6uDnDXgn6hT3BIj/eycam+PE4fNWiNt+ivguzw0tvKune4DobcR
UJ9sgTEmSHgNmLJEEiP8FKKEza8wEDkDGyPrEey/KbY9XS0lAB7m//Bd6Hy2VHIt
EjdbN3ZMX8Dltit3p+tAV40Zb2GvTxPivBZ+EhoTROcbfQ78PSfGNp3DHJzJtCwK
+ujFw7Qs8vDNu9qcC/Ly5Sdt+CSzBMcjcPPmZbbXyOGywpzp0SuPF3ss4kHvPtdK
C/+KRMzthhkRZXg053xwrIUbdjuu2tyy03tbKn+EJDZnBYc4DGWkiV0WNyyPYr1k
MMoLPyWGi/bsnUgE/g/XETmEqecomx6K6ON9DZYk+gvVn9HcqgymaDorbRHF/dCA
Z7dG9ARKxVbB3AqLyDHgy+WXKBorY9S5DbEfAxQ7UYwJVH2gAAvD3txIVPv6GmJz
3p3cDtwBhitR6Q9NY6zox+n2jGQaHc6deMgKIi2yS4+1xkvXwmODp8SA6IWnSWt1
Yl3lYlF6SjOG+1aq65WnTQARG2lC2dOCtGvwrSy2prsTv2LywymOry6964hPIgY/
3a0snoMQVzftMddI4HsihEq3fPAQHYQ5+YlSTy/AtaSiKC6c/rxRh3DS5iY2Jmhk
EhX8VNDJoT5Gu9vtyvQMEhU8z0hW2kIcrBEh/xvdGOvVia8ZPZuDeNs3R7AquSqu
WuMORhtf1vhPOz+HiseLV3i/dMUDbs1bRb/QOUcsPhGnJ9wugY7HgaCZwCSFBl76
jzlMRlhWTa1L+jK8Bk3081NRINF6AldRt+TBqPIdm0VdwpGAU2hPWfapjNFs9Qtb
n3mB3glnj51WRlsaScEhdq/gVEfrG4eM5bfxyJo2boKvy+tuhuONvNntWxiz3EEn
1r7TDCNRh4bbpnTo2QBF4nRgNqyPRbCclhUy+tSZfuA7SZpH+huUUC3x+rHcc8Jz
9OwooRBf0Y0oGrxL4dmNihX2Y/EXB9SgnARDp+XCqVceVfTB0CVXk6q48iqqk0uS
PFZd3qfVHBKWytPcQfhZ8cBB5pUu/XWnhag/OQ1xPIwWTEzbxYRZHgID3CVPWFav
SmV/81EgDZokSKp/bkLsRru1dYqCTmjP619K5piVY5BmRr9LqQZ0wQlRpDeCiIJf
eU3nyqc6Bs7H51ImRz6k+92GUVU4bn7NW9OaiW8GL9td+EPU8Ul04mQvb2amv8jK
x3N2kkyltskzZlabO7JF+88DB7pN+vtElOe4dWbd1PlWj1kn1EKi+sVapPdUPqsQ
Oa6yM6qr4xgpm3jw9D+m8RsfjMEXXwKGceC/W4Wcdg5TFJn1B7Lu2bRqoct9I9VY
ybhOcwadYim9QcNuUaPjAOVx5mHL7mrYpXU0RXLC3UGvEj0cEBkeMGeaQLOGPrp1
n9phTssMFssTnqIEmsVpsp/NPChb29WvjX7OiecNakYeZxcAj8FyXvoLUeNLhj6q
Yu8SSJJmbnqr6xFcLeyuOb2S9+yqT5c5YHbdr1dg5RbWQNk83BFlvOW/x7PhJmhD
8+T7u/Yix7WI+KJMKuqAEGdj+BufqxMB9ortzMvZZ+eRg+5FprTvvcamTuqF2suH
ZIH/SVAMjvXcoNsfZfobokyWDjznfy+Qghi5RMWz1a90ZT7lACt0kAm5J6Ljg1KE
v3DylG+9UAgrBmmKykBy/LYnjE1VAoy1Ipkbid306P4PkDkwDZEZWmdTBYSt7Xb8
SuGK4UcFHXpifa5KsKso5q5f60xDDTMnld/OCJ9Qq/QHcC4dU9OX3s6ZB8cBTfnk
m+2HX/Xw9erGfn7SZlTyoHK3/Xl3OgmWG78UHi1vi/TIfyvEZJ8nqGkMx7btAqmu
ocm2bVdCI7uMA47fwsyeH8ah/XlRGkEZV0hqCOHh8vKdcm0PS9rL/qds6SgnUSMn
eOPgt+ptlvSWKlJ5Lbrw1IB3CJVMnv6bETutTD7pr3bpi/YFhC2QuPtCYm+l2cRp
D4bWvA6Vn7kuScePGFJCZDUqHSeviPvRTKZy1IWYFL19OaN3/RD6cKra+Mq2dkGH
UaIpyk3s5oE+8YmRY3FRJYMgNsCnbL/JyCaYL5YKvikLR6Sf/yxnevB+4FQTO6Yg
jOzwain6AXMEXcVPnbzOTKLhNA6aTgRGvvoeuHR/UJhGgbK9djK+F8fOFVTH8bIq
E07zRzZkY77ewS9LDqyd+TUjrve2b2GWjk0xKVF2ZgvOaaN8TBb++O+bWsSbpNy1
nQvktlbdB7gUwfP9SMqdV3rswGtyiwjJP+5GDEhU8zRyUlUspuy1OZ3i1vBKo3vN
VPnSc3Q0vUBX8n9a6txw/1vlLCAZTzWr0XtHP+NtjpEc0B18MtY7BAQtBXV0WYut
QZK1c+34iqJoLwpEmEwCD6Uk7rKykveFRwvE7qdYIx7b87Mk6ojCEQGFChT92SdG
B1rvcOTz20g3iYswGZZwHFfmWdUpNHwQmRTXmHM1wKDAr0gWvD/YND2vMUJyQPWn
aEpWMFCVj78gCyZP3/eIKxd3TmSJ+IPFBdg+oGUwttNtGQR8hWQ5udCLQc/Q3rNG
3QkQ6//Alj8fnV0ZtrPb5M36C+sfzbwxnmHKM3KnHxzzM8mhwlXUzyEQjCHu6PNJ
ca6ur2qJk4ejKjysMcdnK1BaynE44yQvvA8S+g37PGGozQpCmXigZOFGoa+Oi3Xr
CaF1Y6CpOXEmHz/9UJGpgiqmbH1//J9hXqmVDCPEQGj2uYAB7ZIe3AfST+PFuUQj
MGCo0OWGWsN8uHkox0qKCjVKtuB8FZdVD6FgeibwIoUDDX4Dl0A/XUKl2oWO8R55
5nh5gvwV8P6p/DD7WOOmv4IsqQB48E1p3n9r29a8IMi7Prv9QTW5ntv2BCiiNXmV
GrdcXwr+Q+vsMuiXYyZBNi/Q5V5psHwxJF4CFo22UVfuxQDkW5YkYX+3kc4qO4dn
nYT4H5XDe/Gdzl2KKMKZoSByUuHCTFv7xSu6TyF/P5Etd6tZSCY/tpWttXT4icx3
PIGp2KYo+Zh7kGUm4ag5BXH7bst5Vhhg4BtjVisyxsOdoGzyNlAmJOGDeb/LY5UX
wuVafazR8HcaQGq3Pbv6rC7EBtTJ8AscNch2OZeQOY/3voXGGHTxTQrJ3vldEb/m
DCRnHFBCZfOovtzxdZ81u1sPueHG29zKxotRLOwz4sZ2Fsfl+QoCZ3Ildrb3t75t
v2yui8vu9Z1sGjnbMPb4VN7M0WYv+iFFzs8+pJ/ZGQ/9EG2IJYecY46J5bwBs7r1
VGtj/RDmJjeuvLajIP9IzEubs6Ksce524kgSp3bJ9H2iJAHl7bzWItPNo3GqrQsV
EGBLp6VQDir0GgqDZ3qskGlJNvk6T0V+SmF1fbLEBcdTa6Queg8ObQ3Crb8JXhYP
PVjBgoIXR2XllrpDM5AiJ4DYWaiQgGnYZVLRrWx8QDDTYHOxFbuwFJQ0hrT38VpB
Iw0enMpu8LndIK/05iXbfavPDcHVghuP9BLZUo0cmU4iugCh7z2pzYMEi4uTQn2e
vbyeNWwCQrijR1YYG5sYHbAUlotB2Fz1D0T+c6y0U2lpNwWlbE8tK+yUkA0mVPPD
yEpzO4IPfq7oOYlekRqqQK7fvwzAC4uvMDM9hbX1yaoMtxRBqwgy1B93Vm1LrdZV
c6DC5yl2KH2gQ5kQBjjNshwWmWrumolRINEzUN7S5YE93xKDWsXZeLsqDQVZbb0C
/zgtFh5RUvLbAjVHZGj6DB/TEgz6d8508/48HEYfWIYbh8gzTLOyuXnxbZKj2OZu
5IlNhESvVd7tKm8o3v+h9ltJ5puEjU3YF2fYfvJd7atwUUcYMKX08XOyAiTySQt3
cEeEIkrZEQK8EHLHQ51zzkVzk6M4FXQj1mYpeadyrEZBdAqudcF9HRiuuyHXQFlL
zchZErwQZSRPrJkNZQAOl2QcpeR7e2jyUkomOB14fH+o96btM1Y/u0ijMkZrIl81
eTiqUyXFz1OvS3eHYvttgfBG4Bytma0qK2yVM8ZZthDz56lQdZhP4ozh2sqkwP+6
ynxVp1hL5QilSbrAcZ6G1c8DpXiPhtJj73OrX+6x34EqbydTuRgKfAkt/CczVkUW
pi2UcG1BxqQo5iZsmtPFZhGhYsPPsYqqJwsMQ2/pdau7EfABfqOONKyl0HCnRpKU
TEpL+iiOWdoyvfIu8UWYIaJSlSH0z6Iu6GQRwj8Ocr6damBxTpfRUyyIQnACoSOR
Oh1rStU+3BiBDHOqQ5dBiSuDUiD7Gb3iXN2X3C58EuCjOz8lNY808XZjVZe5bOxC
Io1k2g9BA6xeYCSWxIyqh7QKJR2CFOb/J6Jm0+WH08uUIets8nfVrn30HTsvget6
TKkoKtT9AqWSmeGA8FeN7k0QZ44dyV5HSoaKj3fm/6HfplL+NCmfAs89uRBDUnkq
rhj8/0HDp9xmoISKrgs1AHEkzkghXPYjdvMeYng77trG8XHX8/33OnVArlsHCLYe
GYDYVNk912n+Ezsn8K44MFh6cofLRhXkfuklIBb0nvRuslKVbTEyYWRQrXAgN+u6
HH2oFz7/B6OgvZwewImYw05xSEzL57MCfYC6/efdNoIatPDU/BJSzu2RRkxxEl2D
NpbVlTgOxfohigthnhdO+AEEw3lVAT5Gn2ntwXcjfSUT8quSEyBch6scZOxaYbyg
8wJPL96rRBCJuHp9oXYXD8JxS2S63sPl0yH9G9A79f2WeJsl6RCrSoOYQwCGlrZ8
BAdU6FiOaxvkfaTVP5FPbb2odSIk7cOSf1LDAC6zdAfXelB+zVs06mcO/IRcGcv2
aksNiJFoucJCiFlcIaYU5GpAAoqB4i4h1NrO1fVmPD2rhq94WrY/D1pwmYVuV63l
n8mkJ8eFfIRcl1szCLNRwKWJ1lrjyxQPix4FlgnZ8nqeOmqKFHkwxj7yG7NSBFRK
uTdZbB8pyaT0tnAYV2A3MKlRHGl2ctZi4Wm/Vv83r5EJQae/zT2aCD+iVHWNMQoE
rv3MaDW3mBRA8ctxGIjMEnuXTMc7S+/mm05WuL4C20fLzKVBnILTP0U6pPStba+8
M6nZG1tX4NzofA6xp4vbd450cXXb6TZ+ifOz31mJ6iwKzBpcJE3opPl6/dhDbTvV
DNQVYXWYOBxSCIGfHa7elID0sAwQDKxyctcXoyixQJbz6/yV4OSSZrsh8Zl/qpJZ
7x9aJMap0AO602gC/EXZkchRBjmAX0kWq1UGiQMfmeUeum+7+Tl3+YTFwuqR3ztL
VgmXd3ZS/0E07HrsXZKOzLzssFEn4622Q7Mpw81uew8sCZQDL6riv+C2MY/6LB//
7ka7Rv29zKLWLoRHn6DZDQOKnDPMPAYaZ/lLcrqARb5GaMdP2DZT5ktrXbPGeysR
Wi9rStAw+E/wJX8ir40+1fr1LwaIsBH+GviTTe6hHELaiXc+jb4xljWhCwBgwSD4
IydVFr7bcjCMnO+8PQ1pOpVOQ4vL9DQwgFHwGMSZW0zTRSd76nM3BHkH58FrwmYa
yXiuRYRm/3X9hXkFOoCiz2VufXJOF3c+yZI4SI6u49pwQQjefEtU9YuUe2wb567o
XWn1GQUAFgL4jNyi3RFmOtKcvjrsx3pF/HfsYel8YmIRdPVq+MWb+oO2Dhi20kPl
6N6O7rPdRAP/iew+uIc8l7oZIiT2I9BwLR//YeNygGgP9pbzSzfRXNC1yB5aurW4
thJbU01/cljAovHrGC0y1Qzv8rajqCwtXiD4IoSsy39koKwAPiXfN7pV0NZdMuVr
Ga8o86vAsoOXpPC5yGqaGTv0fOD5WVmqvECEdsK4q8IoBNhagyNIMkJDKQfHwfnF
HR4ryXPy6nklJdPl/AWc7QrA9p6FNFuF2YGhr8+bynWVEedqWZiYxWbN0hwSRhCT
d78MFw0VYpIE2KkoZGezXlGKF3tsgPjItDcFWMx4W2KwBCW042366VAF92E5KCQd
aSrbRugtnjb8CVdk41nnerXfCRpJTMhs6lJcFM5I5V0/L0dy5z/QB/tcOSelbtWs
8tumZH1rNog54S9TmomMrijApGB5YKxlIgINCCM1rpZRp98q97DLxjXPt6x4O38i
hQk4IWG9ssTo8hIys2dtuzWh+0FXxf11FylogyTkqt0VgnA9H4mDWJdKJfd+uJ2t
AJTUoOhS0u4pU2MCg2HxOE1YgorUcytfu6opKtpdzSCt7CehOURyMnSqEQhkh1Ib
KHu+EIzTxYF/kq071lix7ZND1dYgEri51IzYZLDmKZjjyrgdm/EXH4lGVTgpZsxh
/q3mt7CjqH1/CT0pFaOowoCMQ2wf2YcdjvRYSd+5k51WuSl3KG5acentBrW1AmHg
FfUmchOcq1rqhavG1lLdlDEmlt/EM5x3KCIuMy5iuViTIC9bEn74XhBKCyYNUlE1
lCCwzLhSA1PJ9OJ9/fK0vQllkrNjl0EK0aU0PiHsC8C2c2Vw3GlDmiSuU8dDhJD+
W53a0/+v5ZsEIi9ATScVYiztsWNNAeweYGMypcfjX9mQU5gXUO72lJ82wHBd8Plk
1rfehysWs4iM9oIbr0hgnWoW1dRf2Gs+4P+63RqSA9zJJ/cn3rr9+k620d3AHYMS
kfwaEf0dH02h/KEFMAMsCPG8DsElRFkeut6UVKElR3LmwcZI/ziWQVZ/EBU9LTHh
us1pJIUa5Vs5xGVfWQ1EUOiboV5m7eYNuVQZnoTmQWXdK/eahYmrDXKDwCFfTER2
9FYNQOS0UtuwWfRnOBERBZxCxwxxso5kFj4QItpBaqxjKX2kvsx6TRzJH1qnXO6e
Yn6a4OpZopYJyTgLFEG8AGr7XYe6/14n8TkAWpcj3NSA7PsgCJCgEumouI2EnjzV
0U4Ct2WqlSyByR4Aq6XB4qQoQnE+6IxWtUNPTwqddIK4woQglB+GItPponNBWv9Z
qNnx1bzac4IUQe98JpZwhAR1JD8gHG2NDJ2jA6cVSAg1G5D66Vf0HsgsD7DjXSQ4
LtW6rjsPeD0NrH4PffjFYXRueZnJwARa1/i7WKduNRkgUkxurGAlUeNfjWmf1Dj3
zaiI8eyvzsSLXM44QiPLy3377DczKgV/POH4GVDwJVuxaFUPfOkcasHm5DkMy+jF
GJQrnuUki/PVsUaTk3TuHSqnvJBM2LZzOHvafvfcZ7EdO+nTysfhqViUcCVO6OZo
ctfXVwnai8AQtRLYunk9QqQt2C1WgDRGOxbgjl5y7mdihxWJlqjhHZu+XIL788rS
DybX7PeVrvqkC4BKFw0aKVrMvBOIQ/j4XvBH7mczDc23DfkxrJ7rVZLcXxnDRqAm
7tcigwwTqMzbZ7+1rfCIaYkXTGMwrUQNxyVu4z/onOSPKOFNiUIBbRENWoGePF4f
/HbCsXfpiwzzPVztoZy3oMlv0teSscM5y+Jrkzd5YyIx7uhuUm7ym5SjwGM4MBbU
V3C1Y3CFTqe6GpOu23sM+Nv7JZpgeahtv5WjjRI5HM+oSF0ykDaRb9aSyWjWXIhD
EbMtDl78cgGFiwiPf1aUgZXbnKUpy6CCqBRcVL/3sAZflIGpkTUnynlqK7wgTpQY
fVMIiOgjZ8dHllUWorcCXdkSzrKGx9qWsmZ+BwFK3h4mysOvSIxlyZaRrFtXEHZU
fmQ0HOuthK2Er5iKczTUbpbCABp99l8NyqfYLuXrHDs=
--pragma protect end_data_block
--pragma protect digest_block
YC2mcaa2LGxT7fqJg6z44NctuvU=
--pragma protect end_digest_block
--pragma protect end_protected
