-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
u4yDFqUuh8CtFdxTtax4V9DuFLfyN8EvOWSdZxbAVEGa1RhOrpke6TymeiWt6xFenTTfhr28W8gz
OHeP9vnF5nGqSgt8Ng70fZck439StGEcVzkYP4TFWeeCGq3t/0jFX3KZQCJWYcXwKZAZJ/uPMLft
YRoQXiPULkEdGUYnk84Oqm/JWqwTKWoSRNY3Ph9CSV6Z6F2AjPc//H+79xEPQeHwAXWi9ksof5Y1
2O+V2sGbEPUw+CieJiBQ9tIYV3ioSMKaAw0L+z50ol32rSwpNNN/3tMLvLvAyyD4GtFT2lEAr435
x6Vb+WA+4fxwjA7IRY4XHpwDilRJcKfRrH/0EQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13024)
`protect data_block
S/BTbekQTA1tuq6q/BT7c0235NjRUjfxLf1CsgXG/l1uB3STzZTh2QjAN34qLxjzhcDlIMvOJ3Jw
upfvuvV1cHIpCuJvvGq67ASWA3l33eywEiV2Vm7oZei5SD8uhiFi7mtbsRKNBLnDkIIwbDVTXIAO
kgoNJIKlMA4cGGRecJVV4oq0fGF5aRnceAymi5G64sumVE6L1AHTpLdJ1K7jpKdD1bKg3XqodIKE
Vfp20zPwl4BqwXpRJuwkTVd7/l5kKV0MvJf+bawbLbgtPN0m/bqwMaFpqzO/gWYEwxeYV2KmNiQS
rDUJizfzszNaXDoaZZQh6BeKvDwxy/UrUsH8Y9msIUlg8+PZ/spheLSf0dF807jLYeix8cffzvn1
jUz4hpjqhYF6SNDIaWM0otiaDeisThrx8hnvgKE1XbkISGr7RU4GiqgzHCE08XPA5ZJvqlnZ1mbL
/zUiWpHWuEzxWzUvLWVmALt4xeDwEEPh7b2nlRUbEQLMr3ubVMr+C/ATcbTtFci4AEDDZu1XEStW
wD4Gx4tJY7Hn98l1zicOxbrfaRan2UrPmFF868L2fgw1s5eY1pcX3vdrCOd1XbhSGswM2a7RUFrs
kkNv8BQFdC+qOOqSu8v4bCJc18H4rJTMc/HdgVCEE4sf6hneqpFPW+UHlYGEa+sBekv3w/jihfqt
AxIywacs2KxbTOePWBSJ1zZYI22JdWId6iStN0c5JIex6E7wgrTWTa/Mmo/wk1ZlDloEs88ZwjwB
WGjIYTVvKkZT1eugeCyDnmZYFx5I9xoQmHUauerAm0WMQlCUV2UI2vnE+nKLSGIdNyQOGSHCyelr
FdOMaBlWZnGWsj5I6DJrTi0T3G6HDLrCvQ9riBG1fl7ttu8+02IVDbId/WzHA2dwWxXxyj5nhMFZ
4+imbx1DqAMpspKX28wCnKXxfUBz+IxG8A19kFhk04US3hLt+hJ734bc/oAO1ksv8l0C9+FooPIc
O6ND228xLJY/TYIbGBrXUD+0t4bDrOFCTL2btxdJx3r0Y5i+1ZAONJ3NbpOMbNL3jijjb77jfwoo
IncbCGT+5k9XwL7eBXu7K1rVyjGDZ+Wa+/8G29qKOVxWClNez2Lr98/GQx50/qjPPruQ8/NJuiEs
HbtPrG0x6+miBZUIDlfRQuBYt0u1y7KocmzHySc46DWlbx+4P9fShV387vT8Q07bZNWpw+n//mKe
HGJODLsiuLNe0gHIP/xyf35UCYANGj8DDpgXnxJLr+WKAE1+u2JPrU2YZIEgNWj3OhUrUbKYIHe9
OeK1zSsaUb6wxW3+YsWPNUhMvHXmkHZ4pev+uGCsh6/vbcxfT5Hwz67oBpw+ULeUKrEqxALYhHhe
TGDQ/LHHjMgNpL4RI/epyKxjPVnPF2GOqyxhuvMOhXJqTL69P4dXJNWK1g1DYZUCJC+2EHLTbslb
D37gegEYItjvmpbznWL5XdVyDoGAEEfzN8wRCcXOFkN8a0Y/KZ41CzoYSXo1mvp9MR4mrr3Egw8Z
sRD9Cg7WCPGnHASj2jsMFKw4951wo12uNL9IpUGlHGTuk4kglmto5cLPsdySRJpOjn39mA9xNahY
R9FVihv9T75SGWLGEC2a+3ndM3sUywDbX/m46G42NjgT1DGjRTzX8t0Jr/Tgty84XtnGFtzV6Gcp
U4DWtyU3fQRAI0ZNAcEU1qVBvYg7kf0Sm4zwOvEHMIAfNFrnYzd0PoTO/PPSljpK+8pYybo26GGE
NEWKANl6AMdLuZvQQ46aUj6DEi16YGysxxly8Ne1jOwE7bguRi0o94m4zADJzGPF+XQbNuZxQUGq
LvwSdc77QAcHfIa/ATpOoRyckFPOU2l9Xm9Bs4C9/c5RiUwa2TLR/MRox3wk3e+ZoenUK4g+6I84
1t6SGzbMpPISMZumYIpgJvXYOuXU/M5sx1ICL2Mbe2ZH4spK7ViK6/iDJak0NCA+gV1mXSu/Ams2
JQ4lT+5g05yJ0+ZWsFVkHksT+VdTG58aKzTaqkdGPeLI21oN4Ay3feKH3+IE+yZVWEMEcrlTBChi
ZG617jw7Q8X6MlbbpM10wlgSktz9eyu1zv6GMtlQ3XQTLWOWvr/wCv/1WiDJqrd4maeQEpDO2Lbp
nZhgkSbNrlBZ6GLH2idFgbDKXMPSLiiRP+pDLIpArOK6WmYJAkEPnne/dCk6cRs7BoDV7wEBVz52
VtQaZ3gGi8NYvqH+oNct8hPEmHwuOO5UN4l5waKl0ogKFwYYZRHda1t8U8gs+Ls4TcHRrkrLXqRN
Xp8S0OqBruqZdKGkyPatx/B32gGgbecgTn6FHnruK6LjtUaF+BV86aqlEyJ2mlBOvjP5+ts0WqWG
StQYk74irwc9LSiWt6YPRv19YTIYO6T11XlhUcAyG7TsK31TXqNfssz292S6p/HcfIP0kXsUhAET
SOAkvM8IOZQE0qKz9Efwuj0naJnuRbz+ASPVTg3tVEYSfFYu6+GqMpH2SBltpFhLFA8MEvzE2QES
ctwTjwp5LnTpy07kKXKeXxE9/c58vbZJKFJqMhGT2V+QFK6YA9V8gkb3VtIrTq9hPrFlvQuQ7DEm
Pz/7oDoZhhXXqQLY+8S/BWba0vOeEgX5yYCRGz7qNIZZyT2j2YsfU3JJh14AAOmi4FegUE9+blYu
LJjUDkTw74llLiXMIUkCD3pA6TyCadLJJuYcxW31QM5t1kNqSqQIO2ZEQdSaOZ4eCBPH+IxQltzP
tptt6W7PA2Fn1oqgL10wI6Lm5ktC8AUOZ0bt8Rne2cbh7/geWhhmcBM4M5piNSkKCMamRCfILrNP
17TVQcMVECME26DL6FM7Uw0vGpPjI7kc0AXj04Ckj7XSLWAoHtgqua/9DsV7VwqtFqRBJrko7IJn
M3EakE374rqJpmSGmVHARXh7CuzYY31hP2hcWPHKiGOwIxvXIa5bav5zHrgrd7+0646RfT2aOtGe
ruItezcdwlYkAFMyBM8AwKatZ4XEYgrK7Pa+c01hGLTmGz+egasnhqChRqIx53Xu/BvzxOcrcRSP
R22jaASCNPpbDdHHvny9Z9/8LwsZOgQgUMQ/OejGYCtWupH5lRXn2EBuWZdSRu7NC56rqylvPob3
xF/y9tHAwMYthYg+mBb0G2MlFpy8rJWEZpl9Q8DUCPs6LSHfr5Yhtk5uQlwhgCumvxCCrXiB7epw
QTRXCp/5VP4yrlqtspv06GEhQmq3SBUCMxTveFJoA0vc8jXnQVG+Kol8Qg7JXPZXuOathkQFVIFs
EhOgyjR0lwAFKOPlXzJrmA7Y3ioYbwAPwB0awy/RtEWhon+UvlEm0hSP9881co8iZX4OsmuyaDnF
fcSSYh8qN2XzQM3Zgw+fStJOYn1+kd6Fn/e7WqT2iQWsU6dN14RZToKKCCacjkb3AmfvYgsrq7B4
IpJav5Zt9l4D985EZuH0CuKOnxY1eDTS3Q2Av+jXdC9QfF+Q9F5FqcJRkks//fppFKyrZHVAfJ4j
2vFhN16CbGTCfCueew06k1kM+sGTgmTpmpW/n719P01xFyrKcd2sWrcIs/HeRRUsFvrdTdXQ5MwB
MP20OBgPyYA4O2vksXKjxMdK89/on0mu8SArykmnuZNYR7rF2IqanPfigDHyWmjrShjL++63/y1C
ez1kzX7OjQb/xDWDr5QGM4kVjSli4n0d+mT81hBpM3HtDoLeAx5sw90RvfQ3wDHofiIB81mi9vRv
VFE1bgr60fOxMTOwWCv3LFP6IRThXMNBvAN/eFtEI4eHeTrR9nD/UJHnE658wBt+Q29GoBDPKlb0
ydNl5DuuiEYy/Ue/m5VqIEnZCDudglrh0+MP+vcOA74Rq9H4D4FGKzzEc+5Biq5adxu23kmi2skS
jhKUCyIdrlYhQaXV4hny4U5VvsTYWWYAx6cg4Tayg9oFjb10GK3ybCQk6jlS9k2yX173Vwj8cqmR
n+b7lwd/Z6GIDWJ+HR1nb8Qi/w5JR0/imkGwIGFbxbuNI5Ls9H/Y7vpKrq9mMbyXFDB8+U4gL/Or
ebGrwl9x55fgT8yuxcofMuDzI+zvlToc+a9pE6MJ5G/U0y6WJV0G1kTTeyuz+r9qWF3Kk/G6Y+K/
f1OXciigpGuhw3lt3ZjJYikc6P/jB/JJfQSQd5/qNKPl0Qs652Qi+HMansUl3V720SvTtjBx6Xc6
j7j+6xUyODDF+lwvkNlKZXLQydcxeaIjCp0+3nGBgaBQg/GQl5lrUI2iY/irjnA2vlFed3DqGxBE
ExIZ8nmLqxPnuiqJUIg5sFDM2BbZKvN8r1FCCu9pNOlzebPhEOQxjp+n94pTZEGlOxyHggeC2xzs
JZIz3ASDDed86G9cmJoHf8N2nbtNO1tFe7fkXi6qQmuj+7vz/L4lHWlUKyt2QivzcImeHHUe8vc3
KL0xf1KKySuUx28S5/1n28F3zmP389S2GXVsuiPEYrjiAS1BvnzmbulwaaglOuUjObwMIWpRoZbE
qGFgFVfiqBmDLcHZphBziCDL8fRpWIkdGE6/eGWQTE9IWeP60ZzWB4q9TRcgRSKPJBrQVtySSDRT
snbYy634sWpa/mc8DAAH/asqA9k0/vicBtQhk3OAtzn+Rf06PbXHZzafE5v0a7qr9uvmOLC+4JK5
W8C/6mMtBfNNCOevaMHLyv+DioFsstkI1ICYST8cgaj0zJ2MI4KOwg9Xuh8RxkxMMtpINtOgulRy
aBIhSrcY9RhnGWB8J78yaaZ8K5tGm+W5IYnTTRdmn39zw1GTy0PsmxkJNI9eDysZl8jYtHIlelQB
pnjJtz+gXueONT9rG/x7pFKFzs3/LxKCcDBCdILGk9Ll/hqWrPRowG7yCYCW2Pm/5vtih0b4729o
iB2m1FWG5QnrFT4cCkhjKBIfYr2A2x69aoE2W5seMcPtInCzXN/Zcq9ebnGBE1znRyEmq+plRKoK
lHBici6ztCvXIBGOmJxRATASlEYRJZ6Jr8srRSdALRrbQMvmDlL6fySMzT3UU1/d5w6jS4SQmBXt
+vtqWsJCLpZ7tPdTPSDnrsGuLoOXDaTmD8TKQ1oXIDSZd0wiyzYIeWvrbVqfzRllPTr7c4NwCkfv
zxyOBA0jUFznb15AEnsGvQ9dYZy0sf7hH0bH8hHJxh7mC7A8lUbEDQoscEPDDCyHLx2+ClgNcA8g
/IMTkSzjP4esWuZnxSSN5uO8sVYqWtJ56gVAn1RIjm3VJgwxr6igVUdjsgJ3HIA5CZkyyYBTRhh/
S81g69ABwWsqVU98aAloDEXbyP/tcGBUb617xyUPcArSvi7ZagjhKoAsBlI9xyhyiyBydZ9LrdaV
NWSTg5wzUW7bacdUj7Opqva3cwkGKrOYhkAOgEZWeGVYZc4lYKhIIGzNs28FoRJLb15o+KxPzZAG
eHh/e/18aJYuAzHTmGJX8tF0tCaDTub9FHb0KjEy/brboq/o73qaSg4TPYv1zTpLbTVeek2pfix1
FLeRNrVifEt78zpxGNdCcOqWWJL1bXW73gitpDgJ5KsmHujhb0/UZrHIiL5KOiyurdQKARC5cVcq
nolfQBMzZ6PIuJ/n0n/vJBq+kSsLqDip2ucgtbfsSO6agUtOeb0JgQSHwBMkHzUIEUSAi1U2dabR
dNRv8+dLULqfyrj8F4jdwDQk7pzo1q2yTbz91+t+Dar3hx9y9BSKhrr5cYwPRNAiG9dhMNOh8sxA
OrBrjsyRwcrkAun2Qmh4uqTVHW4OGL2zvpGt+WPXxg+1KAf43hN779Aj6lKOR16D9oi2LW6FbfNs
4iJ/kcjkqeS/jzYyWRftfz3qPFIRdutJyY+Zc4ZZJez6TsHktLok/wcgLVJZnsoR3JA+fVzuK+ZD
oEezyL1vBZzEcfLkTwIDE42JSV7JId1Undyoo4oyJQabGRAfyZP8dhD9AxhMQFwEBTc8fryw0QgP
rXgI+hj5RlMsykGcm8liu8J0LODf/RXtm8byo6RXYS7ZFEzn9KYkc99F17XICEJNLs3pbRGVUtpX
ymlzmFKgITXJlax08pZTgOcBQuVNNccmZjAjw4EyvpKgq2GjhRwj3EyQnlXl0JgrgfWOnx60sFTP
dOgfdtE4ZNOH0sWWw0sAnyHWmlktZbaXyohkvxq/jP8Ts8E/MtAtyFdSIHGhurDgDtDeyaDR2Q9s
LBR6VI5o0d0JNZPyntM/LeMpBm8FGlv7ItgHfUYhS8zEr0StQxuHAvwfElvFkqe9Je3JkrwJPS4v
vc4dX/IRq8cmxaH5qcY+qTJxgzP6m629FebJwjZI8/tT50627t9wAcZ+ldyQJpC4KpxWaDSOBD0L
7l528CWPYpo/amPhOavij0AwXHgM+5ox5Z5xpiASe+qL3xSc0zDOjHNwocomrSTyumxpjylpnDsd
+/f0Yklqq4fPtVAxdTKTyyIuobAN6vHaJuBiYTioVitgbLIBMlq4Q5cheFhkTPnkBu0f3EBfXQ0C
kDpKvS4iCBcolweNUD6Lb8MbVJ6Z/fUGaSvjpQQ2pqVvSMisevWRGIs0ggnMsKRJf+iqH7gQnOiJ
SwA/3XN0jcgPjFPpY7eS9ciquzLnJm8md6E/LYRVK8HliBoi2ceG8CIM+Q87Ouz0MxroqncTD1+4
ZSbXy4pkDMcEkiroFx7H8RYsSMHClsAti42bjfDKyPUbYGX/AU7XtoxGlf2kINoVreu8mALhQcJQ
Za0Ra8PzbINJ5nUFfqLw2fF1ouAudFudegF/yCiSPlJmnwsUyziLxSw6rW1YAEE4oSkgvR0a1dZH
gXQo4vSkY7CW9xhhye85UOApDxUfZZI8mjICBHsvcntwqEbtmMY0oPh0ryMI6eYgYQ6Pxuh7qESK
pzLu1GaH8gYRkh9wasW4THx43QpNqQIknJAPPJoGmsN0EwOLlDyYRhNAOSbZjX1RAEXtMLSZoEbU
9Ol76hsLZVWCPHpuJNGHgEozQNgwwieSu/xi7DVVRpVA0oMesDgnlGp1OC4AxbhTc28HsMlDRjHV
iWu4tkkmS3j4bdJZXGxEma9VopogAH2idNRgDZvvDXTY8+1O2mwJa8n+YFylKOu+0z+B70MAmKKR
qbOXNWesfKA7xujCi/8lANBWTn8ej8B26o3voG6Wa/m2CnAa/BATnJt7PoOkYbWdAFI+1s4jsG+f
RiDjE8SW187y7pFPbP8FLKANi93z8r4R/+IJuSRHCbVJvnaatTjl5/21l0a22qRWpPEQMTF6Peid
0Fa88PTeejUDV47TO0jYJoWqfM8lI7x4J4aab7j7CO+Y2RwdC++gZUxlKYqT5Qrhd4kM/CvDacX9
eW32+pt0nejOnd8I5J7rDsktrKOmen6/fGmw8qzylS4hSLk+ICcVyaAZa33FtNWHyMsYXHpvcpkB
PRY0YDash294jBpebFvblH1VZpCwpDim5wy1TAjsJKggcwAe0S04gkd2oGkWM2NLRpWn9nEiIqUD
q7DRO4hB2WJLdgBSyVDKlIY1PT8k0mB9O+Y4FV1OsRb8Zb0oQddvsZGvTKTp4HN3bBTqBO+UvNKg
0H83DYPqc4QVIJSKGPYuKy2pa15tbOPrA6gj6gSX1kuxeFp00G86IT0C2r7cQIVP5DArvdXnkh9u
uh1+xz7a0/OJE7wuJ8Wzll7Jo16WZGKl6T+MsBCGajON0Gxut+M0kMzKTVwmKvrvuda2O0DEUuL3
RP9aTaFDMM4Caui5J+ljM4DWbyZDfu18pwFBGZO7E1pLA13zpLVEUKp0M4vuhMFLZBRE9MKq+WNX
DrQ+JF6uDgKVW0+5uAN7zxxh4NsqmQ+XbBnPkFBG4o42M+PxLH8UNfi36D6XpBMgqqjqjBc/h1RS
fUEpQk+vDGfz68zC34sctiyUQoEk1RehcO6vv6H4eGhgPqGaaJb1Sv6HCqernpbcsbIKStxNCkjv
Ai7CrgvUhBcXY/EGpvyFEbzaFlfaRrWYdgfA5kcMVy86xk/YABNBU20bQ5iSBv/k1dZKjm67jtrD
B4BGouJfpn8MJfYSUGH0D8uMXR2uouFooS0GVxVmCeSp06jl5/WvJICK+jr0QBM3AoOHllyAkD7J
Tz5IucJpxH9JkG+rXygRXPitC25d8C0U5OAmQ93W5UqXOBEA6zi8o6R66m7ROGsrwDqvyYZ6bzhY
CO6nsD90VvdVKRUa4koWmu/Pwwy59GNE82zCLtrrxeJYIgGhmLmbeI/mc+OgBc+vbnMeolZhFjen
Cd9hZ0bymVa3ISLeF8YDV0qiBuf06THRFEuXEJE7FQhg5ab9SpSUW0cCu/wk/pZAFKN9ckSGeuIK
Y9LH1wdbEV1yL2S0G9ytafxIvclIb196/AL5S1qCl24J9tVkmC0REy4ol3qF0AhcGlBA85AyS+lN
VoRCntM1pDrGYzXiEIqthMD9xpJBPX0ZT+2/DEdXQTvYvZvIxA15oPzYZi86honl3bm+lORgvO8j
mxWF5lsFVZZQ0y8Sdv3kidjNUR2RUfwEY9bCzL0HCDg4ljqqvwkpUJcHJ6W+gE9lJi9WJz1x7gNy
4Rcs8rSNU7dxX3NEjsq+voiffl0IZatE21gHVmuGLDCUaaTXERUdONyWPkwe2pF+FnlUzaaIGV6X
la6IYGn7+s2pdh10GFst2wbcgDQ7MVj2aUYrGDmj+vPmZpnthfUG/i+V2z3sq2VBAMcbP+C3Q+F+
3AlybffPaInzXSkkuCTfkfEnJh7An/z3GNXCW/nun9rzNlR8GvPAKWAq4R62jUUyeQDKo2NpJBCg
yPPySQbADhhg1P0a2JQQT5pBZrhM35GSxuaEAPNcmszomGZ/DZ8ULofj7l6qSvvIhYZRNgT46OkX
c96xASpHb45Yp1rTixDdHYqRdrjOGgd703zGWCS2aP8boLB+OZDyRODM0BpVLW9UHv52WLm3CnkE
zO9eEpYW+6fNy8ub4rSH92Dado3PI67bh+kW7Xc4XLUKCRZ05mW+IjG2ZQQGHvGhI6GYPqybcp+F
FkjXX35OSP7UZMk3N40kKcADjY1BjsiwUy80XoP9u5FCFiOjeNAEOTXeylmSXRk6Sql333i+fplS
G39WyfAb7gHuswJBaE3vRW9ji+QHf2rp52Cp3JRm1WOAlCRL9/DaTJcubqqU2tGaHZFGkLBvKpyk
PzW9ybYoF7CQHnDsYBYGnQuVztgUpcryPBwwMS/Bjc/J+GsrHNwa5cGWkdO112gtn6rEpIMhUCqT
9ypzI/OGN3tBXIkJFiMDTW8WIvck0SiX0Wrubp09niewf0tyZxErjgSOClDa6bT1OEbAC3eTAYgG
YfYtk7lObIkgjkWA1GVhMFS7Aby9/g5tcPBxpVX4aA8+eKdGip2A8Pg+D4KQNRN+IgHNh03uVC0Y
EJ73Zezo04gEAO324HN8tKFb+pfSepO++80tbtCuI158dbmfrTCkTVj+reNY9eOYSbWtEtZlzrVL
o1wNqeSmPbu1h2rXIjB5vNVNYOycZCrm5W1BdcLPa7UdfGqWtLUEMHBk44MnQfOSF1voN1FoSRj/
0qj4+i7eRsaaBM11372ZYoa1oHnTDraM2axPON1fuQ+regToSBAKvduVZ3bW6fN6LFexOh63kTqN
KGH8IpoNVvcHXObPqy5yYiIDFzYC8H7rlgmey0OZDlI3Gkm0HO7SXRWULm1mi/RGAv1Hsjeof8/j
r2gsGP7tXpaWKAnOO0teR/NTay+1nBApfGz7PA3ge1y9wKrixvh8e4tsY6jecV2GFzH3pHmUeEC4
70E/srwvGHxEpAwbKaj47ta2L4moutepisjd+WxxSQM/zJtFVfh7962SQizuUVrY043gkdra8Bmi
PKwv8yqw5a2r7mNAOYa/BLE9LlnuVqhFdNRNdSAzUmK/Yuys9R/QUvMh92wvm+nelywJUAhvl/QJ
0ZdkAGJCt6oqg7rRa8dWI6wYweTwcoCB07n/Ed34eG8Oxu9yoJul1OavdN9Li5nGmkf7Pj1r4TAr
+N//IRY9i4Kbiy1LGiLO4zJ0PqjNa4qj0zSvN3c6pB2iFbee0HValX38CsYfRQmPUCNq6TIUdsK9
4RbF5KMBbj45XuEcEcaW7T/MM9mDspU0jP0ywc0jewjri/TBAlg7XAI189nv0GFQtSJdERULTHvN
JkyX73By+0at4qC8OFUv7I5RzxI1vj/xH2FYG/HQDYx08daWIIkYkV3D4H9FJ98fLkThG/2Sek0W
3wl00d3OcfXB5SEaWSOdxqGnLC9TYVbL8uWaewQ9/ZSFzN/V/jSiIn+MXJJDZcgq9T8+afv5e/MO
D/mN2v8Z/e9Fne7BDnZT3YbrzBnMd0nsqlrqfhvbl5ABjR5mEu+trSuXaWBUxd4NOHV6nOMAwrYa
DhueOAYXRyBA1x7xT34hcjLPdKQ3Wi9MfwVCv1JSI8JdKpsVkTWMYPtfjUGJ/YC6GQe5AbiyQlaG
ml2WgzeU1AAKV7yNCy8RF32VVwx1ls6El9cL5ayh8U4zCPvkXbLH/xd/mtaTqJ/RUqQLD60xO6fW
dQJAPHBP4J2uc/yey0tko7DzTgJ7I8U4Z1ePd1hc8LvWTqmnlmwAAAVBiGWpRNH44bU/FldJtjGb
zahiWof5yF+gfuPyO8flAaNqLyDcEpao0B13D1oz6NkQgU8lkOCZM0HRF7CmCCSIYNyMq1U3gVSj
PetK+nqJ+dyvy8w/3WwcM/3BVcquwbswFNOUh720svOXTHIl75bB45Pke06b/rqkkYb5EtR2blex
IPXPjfgmj1YJYz5rtcdIQflZR7aA8LPVowyhRMlRDaxvSzkpIPat0ZJXd57d6r/9Mdp/ftBTViTa
V6Au2TlLRrGg6FOJonIuymM/5EpNqzps+R+Z4fEpecnsC3gkhRiXs2Z3BqVzkdm52njDHbZZAFeA
qwAH6AGzj4c1X2lTczPrD6Ol3sj0I6yomGPqoPyWpFeNu/Deozc841v+1q2f1tj7E5rTtwu7rQCx
NdxVSrYPEU1n/a6ghEWCXqQ9/N6umt9edFWdvgx0n92lqNNAyVU+BvyLYcJXGrFXWkU8tt4dCr0F
9x4tCgu6JKJLP3qGkBrJI612J/AkmTtRO6SwMLm1A8KjyxWtQgfN5PRwO3u3BGgVUIpGxgMm9BB7
Y+MEPmBInX8VB8RtWUE46OK2G6n6PcVCgPARt+v42x/e3Layk2JSxA64Kt9WhreJu6SDofr13mG/
u9xC4EioPKsma7hn5Ep4X/k/YhSDClV9Q8clihZUnCmUcAr3sezjiCfDSjQSmKe7dNtDNeqb40jk
8kP1fmDkUvPDKDC3dFVYteLsOX4XZ9Cce6cbVSQhQIjsmKrmXusbwcuLUvz37aSvFAas95sOUc9g
ftGWAGQG8MdRhkVjXy2anI6XYELL3bXk2pPst76Uypouga5gdU/Y5FlFyMU6c8S1AZfZJgMbcNug
Xo6ONt3z+zCLq3Rj67qA0jFXJQpuevomYvPmN5XwhkY0lzpB12KCx3QNtMij4MqxUT6ENzd+ylQ/
J6ApwLoOnEAl93qa5QFCoSupxsxmVwTpdJZiNOSFSl6EZZgfrKeBpYMPNvXPjXUMwiANZeqHKN+5
KG22jL9TTFi8BvaS4vxvSEtEI27Ok5pwZWDg1MtpojwUK+4kDvbjA20m0bpPbZ+4B1g8vvyLQunu
kRT5j+finCxp1om9xSFIe8A2pdP1jGOy9aIAfWEomL90mGh/x698yVCL5XBVWzh4s1/5nYHp74Zv
tXo1EB0Hnt2qUSWlt4ByUI/v0hUjQ95bLItmRC/6r3HhZM88EzXLyd9RZjw955OTHQjETMUTBzMG
wX2fx0Hbh93b+1wsED0VXjjNeNtM1XJSGxh+UAmahMJgyD26xlO4rCi/OSaDQuMUlPlCt6HXzgWF
M8GZ0WCMH2sDQNz2qaLRZpN/OH8ZkmkIxXL96foY8dsS13hcZlptCD1ubEvj4nPRq5JaRFXud0Ds
gDKS74uVx+sTw/X9QVxN/qjIZ+XH9zkdsVlsVRrDcxMe++6qaPoXNv3WYp1P02ugb4AK90pu5wrX
236cNB2klet3/hypMUEj5RGtIWmiVV/TQgks8nuTrW6Xe5Wk7T3TI6d3erAL1eOKEQz+hCXiZQ5c
+skm7V2cgDsf3p+HsHKfZwFIaHrFOsp1VcVxza/TU2ukDjj+PAnNk6HMSdijPaLxJUY4x80R1Ncb
gnJ7Yz+Wn8JhkyxS21RBJ5ScP6xwnCBY8zTbztay9pE/QHFSvqzeljOug+cP8YjHfMXJz9ajvn7s
d3YZbXcopuG6SAYOYMAZ7qUm+SVXxYBmBeiB9AUlXM+lVPAaK7i8hNkNEXnUObtm3uKBf35yP3++
VCY/ecqkGx9JGoxpmZB0gvN4io6kg5DX4SsXv0G4WhBH/8Qd1aM4lNt1xOnajdw3zYPMRRNZ0Izm
5Qvu6rEU7SDpRE3c5CecxS4sWFunJCU/Bs0AF26po0UhXpGtnzDQCvcRvDIoXWVFQpMzqXi9ZOpv
H6glAq8NmtGzgYMGgnq+6VMGOa1sbh3KC4/O5pNPyioJMckW8fDb8Z9jAP5ILT2E5oL8y0ecrOXk
FamEcMrjutmIfDWJi+CtAdkb3hB684OMZrkKmHxKEK1glQDikdCVcnCKPHODWsFY4T2gKQ97gq2C
2A/Jf2gMObeRJATML/TW+T03uINXifdt/SlFVqyMYaduuPXBt5jgonK5mA+wdfMF+qHT1vgMVcuK
W5mzLdVTwsVjwT5RtnP/5vbIWh0EpBgbItIS6iVlWP/2l18Qy6+/Bm9uNSRjdDeVzejLswRmJ2OM
RXo+wi4Ob/Y35TMt8poaNjA59ju2otzbQMsrb8kIKNcjJdBCLCjA+iZ/T3VRXRsnEqCLjRs+n9K6
e7IWv3F7IBohnNXIB9LvfJGu9Fgrt5QO5h3Jwj40dcnHUaad4di1yqvu/daZ9WunGXy/SJ+NQ6Ki
uc4aJ9tZHV3b4lAthSSB0rQyC16SQ4tMSsmzA+/e/MXVv3ksZL7UABg37+c/Els4+rc0UeyF2lhE
U0qqvV7r+vjlKmZxlMzsFRSeSaNVrr74nTkElfVxd0C9x5A2/JH0CmWCG6gFGKhGLdnMLSCjq97O
DjedsNtxp9Hzv4WxkJJ10v1q/rJIgKXrVxwJ76h5yvadBbL+Gyg8/uVi26WU6TvvCPVA2nkuP98W
gdZZ8ghExHHteCaKsju2rmezZyJ7EBrFUvoyknhg+6jnAQYShAF5uYVsxcCzoondc+XXuFpz3njK
YQxUct/FMyaWoFFTSrQXlQ4N97XBaTntRtoObqCJ7CS4lvKFPRKzwds6x0JuwXe9IM6oNKERHWyG
D//RG8ObfqS0ZmMEp8sr022nMWL+hOCy2MJm5DzdFvm/qlY0nms40jeLHOubVRwQYJBsQ/NZqjO4
7CLY5uyAC58GeK6G8bbPbc2bohipMh3fY2xIEgaoKEy4t1oRvgwS6VAyCF99b9DU3iIHR3suOzVv
E2/5ixP1IfGTEc682nDcs5HJ3Ow2AsfFB4nxMFstD2kreDsDTd+rHeIOQIiELrS+sFBC4GM/YS+w
hb4gQma4Fo37YQuDs9hRiHd7LP//kWk0phrXElYWKxHXPM6Ltff4o75+uXxhEbPOtV8KteV+lr0U
E3Zbm05EbRL4QQ8u7mM+7eZEZ9eRbH5UpL+XgYsMZXdgvIAvs0ieRtPnC50l61tuPIyAtEUOKyJu
M06E/Qiq9pPrrKmoqpDFQGyxOtY6QQ2yZBRXxpM16fpKp1gjgJkLLFuCiZT5cKxiwehcPrxPqBk9
w6YWjzpCtWoGy+KOO7I3CYpVlwt+fABgeFFa9TxSVrMF1b7p2CcUt0X1NuDeSX1CPITgQUOB0Kpw
yraxGvbE7lsJ3JCuKZXtguR1AnoiGlyf5zwhb0zDBgz2JZd7+jY5xe1X1uXspEtyVFG5y5oTFTIc
5P6a51lHyXIA3sLfaMkzJq8YwPMpuqMHdG9CDyjXJusphhcH1yHFqLiniMKu/HIHdPvnINCemIxr
d7KhhYfo682cNuzuB/P9hclkvi15GFUZwtGBCNxj/F7cRSGjgOceROLSFNckwEzbqf6QgxpwDbdn
d827x2Vp59AvfkoePa1I3cx0KTMafEPvJ56K+x6ayJdiupDvAcPnhtrqaNtpB3RdG9Uf4GQ1iEdD
TgPHmjboOxnFF3HgQRtrC8Phmf0PD/5ri1Lx3EJ6gZ58bJAXbXtlLxB49VnbQWwX1E4izOwLq4gU
8C451oKkVjKgtGjxI3ZccPh71f3Fsr1BdZoVduVvDXcc9sRpt1Iu8llnJLNSj2Xby5sgAioqpaYR
fRSMsDdRXFr7SKUCPDR8H2sI81DSawd/U5m9739qLIFMMhUN4SX71P6DfEuppZwG89HUuSFLdeIl
RaKR1HQ0mQQS6Nv/wptTAYj+xoCCJjVEsAYVnHIYqabhAsixZZsernRBOFGU/OY4HrSnNFw7Opfi
oaqb2n5pZNeH2VjHFjSXPHJC2ew9DCs40PbTFGP06XlkPd4S5BfP29Kzg4BJqOW30iqXTS8JUkfj
+kMvOA+1oAyEH6xJ8nVLFhaxgSdFbngHQZ53VkQUo21NDxG/N7R02/hYOf+3ffChWpccH5Lyqiu8
HKYF6CksmM3/gGviL5MqDztKx7k/7tqk9P+o22uAPG8pkq+2vkTQiTAGw5RGz0+mx/9gQ/T0UMcF
epoq3QWXmILjuvqAwrfLBzzem7XWMdGFUCeUWR2XBLj4y8RTzbZukYYQC75Penn6nGjZyQsjnGpt
iFQjho+XxL2sBOZitBn6O0Cfudw46M+ddyaVT5Zi7Oc4EefXAn2HpLCw9+rHtKMXAqWDTQ4mIw9C
oUNMyHtW8d8KebmHfitDcjHMcRBsxbUeFLjAxw61kpybaI2Jl3hM3OAj7GbveAcBlRC9GIwmSs4O
oSmrlinxdjJ2ISFQ7dzdG5Db5ZHbsyydCcMeosMBxtKloVjsAkh22TR0KpZOibUVZKheHxRUPv8u
GZQ0gj3HAZxe+BlGIBmgSmz0O1PlYzbii7df+c9E8p52jRPYMQ3zziVSa4Sm4bcAsw2sUUw1JRP6
0ucRj8GyI/TMgXiHb+HBwctO0QvUOnnc/7jps53tfhbZvKML5pImlpZ7SI3oTX2vlWkGUlsAUhSs
95wWAT+wVa/3ZrSJh+CthH5VdK84WelbxgBALT4Mp0EuSQ5byvFWpqur79fSjYcqLB6AGqtqxUZg
YcXeN1KbmT/c10ztqPdrEo9fDT55iUb/go2OojD3hcqVQocf8BgPZd0ZlYqGpv7v2fWeeh7QsbKu
jX47g51oKwepgJ+mUXGlRf5Q77jXMGB2MjK1cwPDys3eNxqjEJaUIvC7BMLsHWrp9sQ4SpLPwjou
RKAHDF+bVqUdfyyqu3I0b4MWWqgVqv7qeXPsYd9FkLKG9buQhdZdSE77hC+Uiu0kILPCHPo2OK11
2z2u00vTPSfZRGbPfgKarxho0KzWLolJC60thet7sHfNbV2iIoZSDHlPQbXtjHfizMk2z444wwuT
gTT8RGfBGQmB8qoI1z0F8U/0emwJVdulrnPfWBbmK6QKVpE+hg0OIOEwCfljLnsv5m5Ix9iiBD0J
zVxEPf+yh+LKeOgmEFKDBALv43XWkpl1OLfvyRBNd8jzYSJMvWlWEzfkDd8moj1qqMfM1RycecJq
f7CP/ftasAufGbe6JJ9qIhK+uFY40OEyGkG4DyNmL+VTo7XRTWGj+lHaKlyRjzPxpU+O3gJ0gV0r
ewkYe5B9t7zhocFeGZ1xnQLh7NlK6xfUYW6EEJMQxLvKhccxpX326gMmn9HHQhleTW5THb3PEMvH
pm+Ep9iU3savtKjT08JjOqaXeLgxHEcECGC+mvOrEf+HVR2K+JrNEwy7lKLdyanhj1CCt6i3fWma
lYPAnWxMxmHk+ekOteozPbsNgXpkxweJLPMpmGwFNHRhp1iAX1ANsFWM1d82QH3ePG/ampffF5C0
WOhrMwo3Xl0hCX8LDvphvMR0iD6SS0ROe0B5HCWDjpHo8ATIdeOu3KfeAKGeXjxvYlKOV8mRAcKq
g9VB0lzYkn2AEKUw0MOYxnqKXqVOCRZMYHjOPcXaivQEVvx/jjSt+cbKBMLiZPgOjiy8r5Vuf+TO
+i0+al2L0L64vBthw2+ZCcW8mTtNYPq1MSMebmlyZ9+ftjcF/o7gaUqqzO4ooLgWgb434BVdvt/j
RYm33ND4RaeOMWTvp3h32plFjDx/OoagEiv0Y3Tu1+lCVcoHcs7qSQZYeDmzAKMgxWj5gXkKzWtf
RTXmuSyCZEYTHhMYJU/VWXSeqiL7rE5y1L1tLyCPe+oIODbC4vdb2UXPsu8VJp4fW7ivMt2YeFn3
9JeI+GLqvO1iVxBkqmqwTak6M9kLBXM3et3Aqbad/S/wiPIvIOyvf+Kjqm3K/qJxprWPMi+86i0k
pnzXa2yjsUiusiARZQZh4DddXRoyyoCRO956fVHJh18xMCCdITaAD8qBkbaHmpaQiFHtqT7JnVOO
IajFKy/zekgtMbjBu7ooBrteR2u30cp/snM1R9x9p/H/wCqacIMLVXx+2cjnfHLx1deO/l1sBd1J
e1mj1m5iL7IfIrq5edoVOG8PP6Nu30OJ+D1WoCZJayiK35PjtSAYTw1orCmJisbWLrscah4dp2Ik
Hzu9QvDExBRiViTS9m8S23arQdNOhz4NbvlogHMcWG0HLASgPGxbHQwOcX64/Vn3N3VBJhOmDK2A
jeSZHFcLI+lXb0ubLXzb/aJPSCSmyL3tjXUIVyUguN648VKKed9UQlNeGP6rqD7ZRfwv93nUaThr
9SOZOZp1oCZxpxZ6GF3WtEU6KUo32AaJA6pmT+W8D9689llwxz+9lbhNzimIsConxAP5HBio8c1j
d8Gc8/riOZoMj/awtKVjRwWRPJiKpkLvw979Xd5xVY2mOlHDRlUHjyZSfqLzps2cs9V9xyHUZ7fo
MMawx2QwzcrF6FUL7DOx1n2JWC3BcRnWlyS34ir3VoZx/BEwEPit37Rik1kDASAYRWSu+4fS3yuw
0xNZcOyIDiTU0bwUNFbmN3UQgJCkgG69Fdbwn19Lcho5k1u5Zg1zn8MRJ8Y0mDYEoLJ0TzKB0A+5
ua5iH4TbXpyx0DomtL86gglL5RAolp+x7V9+Q/b2IQA0oik1Cw4mUtshal9M2joCQMRvRDgkfN6U
XfR5SuTkPEOk6e6xKbE1F4SqznOvnHYX6YeZGv/mita7KeNT3NvPhu66ljDR/B/6Zup6Jv0ayOHQ
RyGY+2j22n+1fInot+4gMT3DHVACzVV073uZyYuoL2kaUv3mXyjqSqE/pzqGryrzgNHTHCaWUoAG
hrfmDGpVdZ1o35hQ5IjzlPyteNOQmq41zGdNJw==
`protect end_protected
