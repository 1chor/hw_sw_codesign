-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
L32bUaoX7nFsozRBoKHhqbS7IL4kU8rWcrGNqxmSY8U+ypyKrv6GXUbGusRTg5YI
1HQOkBaXClh8xCuYhS8tk21K2Kf838AICVwQkn216gD+sxsz/xU9Z5WckM2CPQH/
I/8BqzvaKQhfzBqx8AEgNZ1kEp1SOrzBOSKuxWYm6/E=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 79854)

`protect DATA_BLOCK
5t+3kjo/ECajLep9MZhaLEqTbTTEWgHgcCu7YZzOJJ3PtX10fRmdKIJVxxK461uY
R+k3n3x5spDri8+uScW2zZxmoR3XbCyRRZoHqqK8ZjP6m2q29QtruDYBrSRLXq88
3uSLfAlFoGbrWgOOaOdcDoDODubCj2KhfLCOoX2NhOO+upeiM7fKDEdedAEVfq3k
S19Vy/DiTZOJY9eWa5Zi5CdAV8oofZiIHKV48+/fw8RSYJvBrm7drnhT8wwC/+z5
Cp97wwvEA+rFsXedn9KdyjglL64yi8WQqXNlPSPrTqsBVS//B6G8obtX0efRZVpD
TzzuXmPi50ZOK3eO780Yy9SKYb+KJdnHQuDD308mkOgS/MAKvNnb81f1gfVQLGQT
L52kqSbiALSHqtjz33nquFPMO1Cz4MfjsSHMlFsa/VsoIXGvESrvaSKfsw8ejGGO
hKWknafBLOdeSl6K/efMNXQSfL6E8WAI68kZcvG5jZT8EzzhW2Ual+T1oHOGsLGA
RlJY037aVNWqwZs/hLD6DUUMwXGeJPy/oPRmmK5+K2eyyR6+F6EPO9umI7bQDaH4
N4MThxnsZFjVgblcW4H7oQPmaNqC0Ycj068d4ZpeQQuHUoiKNrpQbWmtKWj0gz2P
3omlx6evWLYK17AH2v8NdU1yP7+wsjAiJDiIBzCI98oIXbVPAhnEyMW5dFylC7dl
Zbw3QhFn3MtswU8DUcDm7453jKdE6jBpPbxTvwah8fE7Kc2ohN6XMuFXNKOKP5GQ
uW+okVTOkZkbrjxAv6Zzt9r2CE8NHHwZ8E+Z7Ypv1ArRlXW9uKYJU6/7bvcZlF24
kX8pxF2hSD5rQcWVO3J/F+JNcTGmfLOPUgcsyU6trD6cRbZZfgU3g/Ztu6COIbU1
p17/yh+nvSMR3+54vA8phOCtIaqFGc7rFQr7jfwDY/vJqnH3/hhlpJCUUhSOnB1T
Z3izt8XsHc7ufz86TEh8XvOBPSEyfmkdJZyu3JOC3JJM+ObgiNNc3Wl2+B8K0I1y
LYkrUDtIKqtNAl1vq8FKCN8LFreJ9P7LG9b57XdqwXVoVbpbs0VawRX3ypctpMmy
Uc7mnirpjNImdnEuYZkG3tUQ0jXOa8r//NRmv/FUNGgGb4ZfyTDU5PYNjrKikT8x
tIpTl+dhNFTBTpNrJ2ei86mvPFOOgwjwcTe0DKXWt0j3c7TqeJKWBe0id0piVxlJ
nkd44+ufKQ4Mrp735rfhyLtxWmCp39Xpp5eEJJKoo+UARzTVsq7bhYM9T8KPueK5
lELwUqDwnjPWGA2ANxpf1Mv+sZUbnVDLCUW21b2/KrRHgt7XdNj4LHseIy/NATXy
nXq1q29yM+YWfj5aH4Es9JyGggN8k0Ka2PgQvciENOR6jQ7GBGTzEGmQatP/VkUc
oGFiwmqPG+SIfAjcId7FfpqGVwLHJeKcQAY6hVmXlciKmPSy6qluOeLE+l8yBvWU
9LYWWWb0IJFX7oxudqh7vyeohLbATvCWvsjewifQIfkY8xxe4ph6DVUfvjN7aK/b
kJfT7Dt8QTdzoOem+0xgm/tu8K62Vu+useIg5Xq/xMz27JmadK4P26Ch57iReFDS
uDxScVbMOe0wswYAr/XvuIAj3N1ewjwZBUcbPZrjwTJH1X4YkORnrhi2en0yeo52
vIICSpYmzKLBJL3jGcDvWzENw+rwuHoHj0UqixbsjtG6EycD3HEPKk15ypA2bwRa
jrKJEwNiHtbSTgHSu582JqpKyWCGySeUgglb9qb1SuB8DvZXh6ZxPxoTbozy6M0x
MlvWT2PxACljDFl8W2FESihCXpQNvKwtFAB/dhPkozE9m/2DsEok5b5/kTN8UMjh
r+3gBdJB+b7uVC0KA1cKlkhJ463BqqsFB7zq46fiome0NPP79EeV6SaGrxfzwchH
OkxGAInkBrEwBmc7BGL7EW57unl7umduiH4ki0d33W1GmIG+kMZPXj+/n5URbF5v
RucrsSri/RjZmMz/kHWJO7qXB5hbE7sTZ2+z5OpB7vjBtLBKA9s9KAAYrjaE+OVP
5vsBy8Oj7hNyjyFS4/UJNhiO3zgA8jq/rTYvEyPV4T8uo2D/5ij7RhBvgzPbPUrV
AbhqBCBZSaskuxqoIj+YaGl71z+nO5D/jMiIhOa0TFtnZQBEabpIMM3M3x9RCVXl
iWnUFVWtJgo4YXCbmBCSV3yJZWCLE9JnY3/JXOptTxwyW8X9oTTurdRepQjAHlad
ERGkiPU/amKdRRtr5oMbavT2/yv7/gOT/ftMjDzuBDo90uvbWn8aUb6g20ZYZzlm
c1lo9ddn8g07u1JtDeDnQnyy8WGB2Xp+dFdjQIoaUisvLixoAipW+eqjwHtTaiEM
1Up6uPznYMnWFzrXDs6fnriMcdGGKWOc8NV/oCSiwVQrkKZhZGiGZJDJM1c8lybP
XdIcMyvYuu5h6f+JH+VO4HalI7xiICWRKizbpoFKf6KR1AaA/76zoUjiM81RDegE
KqU1AHPLQGnV/UFuI7KQyFpXoOdqf2No42bnNr0k68oq5s6xzGm6bWOZaWKSFzss
bYs4qgqaLMjiI3/b2CFeFHqqsQVX1y1FQ2U9XI5aLCnowfIYqgDUQUfhNj7Ke4Hv
zvuDPUU6J3IoVjWP0VQ2Lz+7v1DKMCqqfkOMEOdpOffg9G/85nrICldllnDKMklu
U1KTGsVbbejNiP0PjmmY5+vr1JMtRuS69fcstMaAvWLfJgfwFHinKtH2RYBkH2jF
wXIJwHyPMOzwfO/dD7WvY5MU4uZy5D+pIbHFunA3C6rWeLezh8BSpksDZg/hf9jj
Difk8rhu4HN58M+g2R7XTzPeVm8g2Q8Z6YBzmRfSNDCZTMvXwbp+WnSZ23kSTCRS
dLMXD190AkGpAsPMbhOqy1aguUb0j0BTut/PzMvVEDqPHiHoWhZzmgF15iB3Urkw
346gKYOIvn42MhXsR3452IoImZ9G/fa/z/nRinj2D8pEIIPQ0kFq5comwLSW5Hmv
tvu3szyh/k7++uaYzvM6rM1wLOo5a+jicwXCZg55HIZkXe8RovdozU41k6ZU7Xdg
dGL5WPh4iHTPrv0dhAmdjMpIbzx2FKZQAWIBcBbqgt3cGSjPq8c37uCrridwo4w0
Upt5ZnQnVk5T3M2vHVicUenARpYzTrYVzlYtngwTXsBqU3tecpGDrd+DYrZv2qnk
X4qt/ly1WeyuBCdujq9uFFNW0iopFNnEmnBvxcKFmm5x8fFkjMM/R+s0Tl7Fv0ew
rjGodlufVz8l3DEpKhxnj4pTPfHXIBE2K1MIP3AYnBNEvyasQ4zdFloFulmvEoSx
k9Xcp3FUIuaKBDZzU3z0r92ZrmHuJO4Z3OLvzgyrV6hT0T8Evf01cJHC/wy+7Y1t
haQIfO9+OdkSYMmC+cK6g/VXe+cWXbAhRe6e1p5luQzUHq3Hmn2amOVm2AJpyNlW
1T++ERJ1umq7YtGTftQrQ8xnFRp8ZID1HMhrFM0mVpnUq6SXEt8FjxVOPJiU/rPs
em/QLuCMhzU/GaMzHK2jMNkMfI10H5RKwGN1gM+PdPQ/hwr+t+asR1pdh/0XC9oW
8i+SAGHs3Kz5kDalA8PxjSb5J2uWD0sGuqFtnYUnlqfnZZnBKMV4oxI9wgdDBfAc
l0vNkwY2aLdHmFC1vhJeDpATg2bynM4Gq31kcOJjQVC2i9f9itl6F8PybhUgI9a0
cxwS7p5ubs7yiHHVWKf1zAj4Ph33DkWSqjK5XnrkRB0xugyDsjJRA3CeH/DNO3yf
O8Bnb0eTci04ewJHK+u/DuErxpgVpx5u0WagUe5Vy4fJBrCh3gzyFJB38C3ITOzZ
Pl5QfQxk8dkVVZCvA+M44BB0Ca3qSuPiLso5swCI/stS3lTbrnws71GM93DemwlT
5f7z2fcFoiv8sQWjoL1zoUe/BVJov2Pu5GJGTaf6Y5D70loDWVfhjGPjD5NUPhFa
J/ZAPFbiT2nWiq68jjEh8O6mzpO42F8toihgKDTUshKUb8sZEwM68dFIbvx9LCv4
kQaXaBB5nLRFzJV0M/t01nys0a8/sUyxIPZYDJK28vpB+w/6StO0AD4a9njwOdlE
v0pQl6PrO1C1fEtv+HJnpDjQBPfXlOFFLbOSIs97cX8akBXy8EDUDxYKptZzjgLk
915jJ8bCih+uU5K3yJxbOT8RF1urcHAldtuw8it70nijk/qQWce2nlxOCJYLnxy4
31DR/B4o5lAzFiiEJln+uMPcbXIKLIGv1r/J8QRM7Sk3yuJBCxa8In9i/j636oEU
hZUCM4DjffM/iq+havljXabwJMvrCyeVccJUZxYFUemy0quXKjoi3oZGEwvkNz1i
NgCtX/mf4PXYWSoaq/nkKY30vRQR48ABVMFQNI5gpP68HxUbigXgcT83q7O1kDcy
PM3PyYu5vp4xkCCKeXRh/PIrYu0MDIZZxZs6vr5pJ3ASPrI/G0dWDwllbGi9vSiN
EE0AJErTC6CBZeIqjg+RUMns4lBTQAoeI3j8BkxPRljR5uJwZGDm91GRAzyuwTa4
husSs9/dO6bVdTak4mBqmAiJ/4I6imOSpn910KnZeoqdyHHBeppxdbwivJisVU2T
b7ms1QkXxwPoeb2MAe/HHw6QT4QifkbdOcRZ0PPL9H3feS7J7FXEjYdK5aEG9D9I
L852Sph7H57QiI3Ox6cHadJXHFm2ifTINA9UoTwakgEadbF4n54fMCd/RsBoZVrA
toAFocTpyNdquCQiNcjrIVhFnTgoE65KxCGM/q8jq3ZjEQi8X4pX1x+eFFDDEBw5
7JYZfwGu2J8P+UBIyovluqHOCZGP0bKsIFzKeqLUYNXQxa6y9iU0fLqzemtKPKT3
28/CeSJI9Iu33+6rDsdvlP8aaZ9pp+iHl+7cm0ImMCfh3dad/+NMmGilgn569LAK
jaWqJtbxl4MmZwh6GZEFSP/6JQ4aE3ss0oLgXIkd9HBiglOz4nZROiamLiRWyGJm
UmCnfWSnCWQhrnkIq3KKdRflKmp5dONMoCcPSlJSz4GLyWJXQCZsYKN2gMrGf7vR
RYitoR6wlwJKS1fIEN8SLrRCvVyvCL3Ip5fAl7uVb86ZxeVNx9zfhD8POsTltshE
yqcngTlvUnVDQyhTCrDdH/4f43q4WznxmCagMF0dKxiV2YDlPoQavj11FcrJ0i6Z
1sboDnP3WWMNMkdadm1W0iQ515mrhHfX3JgXM14nMNDawwaOsxlmvWf4fH+8FEOy
KTiwZ2qgwa6CfJjZkve+VHpsEozk+WetdKOJ1tOFDR3kDyMJxhGEuqKqYA+NfHlU
gMW0HbVePCp6PCytuY0B44LY86zQ91T3VpDmKWNUgtEwb4dtlDZqhqJP3X0b4pZq
Cdoxegu3cJKg+U8OT3/eIKIlM7MY0R0LXqxZV+MO/oUZSUMPD9NSk0uLOuGcvXDp
OKtaqStKS75gF/ceOG2tscHS7dSKI57B/KcDigJ3LaucqpxNBgWxS+pRoIDhn7tC
+xk22ijmgsigKeuOO/WV21jUEDl8jOqogFPuUoEtjI9+aKBkx8bypzX11jovwoEt
u//1mOAwFm1YFIXDFQ6ONyjFDLFvHmdhVW11UWq3BZ3hsJmiNdc2COHL9eadt33h
A01anma/YnSKYdCtMn8NcIvMwfDZEx9JnPcb3u+95KPrQ/gJsRVruGyARc5SDAco
Q+TFN9R1+nrezZUh7D8q1X8zTc+2YlJJlhc4iQRt41lcRa5/N9ofGeGK6xMX9j+O
b6tK46z0EIXr2G9Eh5Yh1VvFfslExCz03fp8FCUcg0Khnc8nYOsuqiIrTN0iLa0z
nlgGJ5wbbnr3ApJi679Rjcs4I/hqBBKgByimzyT1QjJEoZ4g0/lMTfqJD8yNQCAs
Kwc0KVf6/8CVXDxsqAzhLByMRel9qdwZ4ti2ZBn3W+0ulXQLHrZ07f0WScxvO8AX
VfbX000F+5nrP7krz9N45ax55wOYvEqeBlOPecQc4eSMqioyio2QM4d/IbPfFSZ+
lBy/ykU2DARYdEj+0j4KqHff6l/pzDQmt3lc+fvgFhI0i5E3048yg9pJQhIO29W6
O7VzHqLG4jKALA+7v/KPiWIGW9VEw6Y1tRWCTD/jHjzWg6ssX0MWhg+bpPz+4JO/
1kbUGjrlawUlSbOKc8pTsvBs7Pf/Yr4vwUrS2A6JgRARcj2+BoA/HpKfCNjuP5JK
X/jWSrwYniTt9dpAzogc3YVa+NqehPATk7iV/xzxOxvca6LEvmWvjkaG9ASQVugG
smhwDSZ4iUxMC1VhsXt5jvA89bEIJDBqQvnxsFAlbY9+EoJDTlgiSENYt16nGc9w
8IS2qmwm4re6qkovqjJIDadJfoiDveMkR9GiCkMEnBXDl79B52g/lDg7kkuSFAaX
UbOG3Ih1o7yZOknxlWs1PdT0yhskKGdNA127xO3LpY3E+frbNUQI6fwDk9/DBxaT
lw0pa63F/HHn1rEKX6IFmm4SQg3oyC0zLpgXDdb9Y1UH/DV0PjHNOy4Yl7cWzAy4
DscUTzGOZVK0KS85xlyOjSz7veuKU4JP5Xva65/F3nkOg9I+gJB2h2AYyQ8QmoNt
2Xc1YTvpio1QkHvX4i6ZYaNcYJuwk7cXKtahYe2WU6ry62WC3EnHWBxFWyZfdjU/
FYaf4Ww/qkPSCuUahvAyEt+QoUilNvnMIsWhAG8ZGwuNXVcO8/yOdG+kS4uulkSD
BizPDm0+1aEHT6xrfBDOsglyNvetf+CdVagdsYg33ujHC495c0bz8Kfwqsn4uPxt
rvF2Z9O8JaU4wJQ5GZV6O3nwcb6E8suE2CvMjP36N2wh3HFp8yri714PG3xT6SHY
WkqtLVyNf+kE5iAlYC4MYK5ZUKsBh0PCBZHCj7AAjRlCPPw7RXsnmXssJqdJ5aQ2
Vh5zn+I0Q3IJDYyssQjp+5QPsH93XNuuUy3OgKKX6MrSEQytRbA5TuHBEy/M3f4N
1dcBVEFf9g+jYvxlqA8/phu0VEDWxY4ExEx1B0oLmrx3fZy2YJ5MRY2237ej2HCm
Zb/W7eTweg1JZp8A6U/IQJnm6nTTn3o6kZW5vhsWxNwO/1OqazdLCWaaI/fTISXv
s9w/UcJna5NJmKIyqBc2HhNDzEuxskLcBlbvj/Tqhbp8qB6iOrM9ljrEOv8JVdMX
DS+2frpYjtm1n9dmVVmD87fyIPprEUAIZ/oBsuomQV5UZpSpfJCLOfD0OL7nzE+S
ZlEbEwuYiFISoUMTBYpQu9dDc5bg1sRhDMtn/IwDZtXPpwgGWHb81aDg6+K3RyB/
NawRcPZYx+vWaYguMoPecZ5Sy4dkV2RXC0D/pQRE0IKbI475bb2Grk484ccTmxxR
Gvm7hxmmsxodJMbMMMG9svZi1yESNMErBpzUR9P5JH+W0VenYP6dY9paPeOUV6xt
awEzwoJ++GCMlYUSOcxQAJ53OV2bBdspdJiQlEjkP+eS875vDT9jFXAwBfAzyD1R
sGt+AmKxd4ee5y1RVLgMMh4W3M+rplB5h14MY3nYaJKYfEUHz8M2vQkfhxdSTXVh
wyH1YjLarNb+vH2GYZf97djVPzuehOXcTbdKW0iaYlXErs4a+u6oZ9ottJS+Cn/N
IpspRt9HwG4Zphl/mC62kqGGsDN52GQPIVDp8vHbg3SdxrPqzSj3qG0vchXeMI0l
6XZziYoBwIUIGTyD5JMEaYfO/tC4DqXPzJmYeJgKT2XqxIAtiMHjB5q4/UUsTc/d
/ASEE9zeLJKEkepd/Ia1kb8fmqewqktg3Lj1l/6hg94wywXWLjS4nozPDBHMzD6x
/qJLvnOq+ngrs0mDSIrDBwL57vhiOip/4wwIH1vdJSHEskZHkHJePM1fLOj489+/
Ggq4xoly//T9JJkYqxiVcI1wLeNeCDajTTwrZX25h7/h9YFNJ9C14FFSRhSvnbeC
rB2g0hVVVs0IGo92O7xhDf5E0R8LHJJnMNlz1rt0OaUrqlKZr0kZ1CWwR18Wzy2I
ibE4jOb1CLqwi8ktg9KNDpabDuFnScWATCQUyQERWCKlkKm6c1r8sVeJ9jVKeuZn
MzBllcQgcM1ysjURNPCr3I22lbKZqNH7SBzBeLegOAjMQv4oiQknkJ+7itC4c8jH
uojy2UtRrPC48q45MHPo0fiC1wSHOfQEf3Nmhe6ljp75w7D3FX7MOwd90YFTcoQ0
5RcXmycbccrgzEUVLGku360HNX1CObUchE+jUg17+enc02fmGfdV+v/gN2Vr9F7r
i4kM7WQTtUEKWxj1rIhFLTjgCWg4L8CrEP2WIX/ZRqzn0oieU3R560wEmG9nm7vd
5lDaz2Jt6V9pRYT5tMbu3nx89KlQw0jmkbJ1LE7Ypbe5Euxy6U493EsF+czhi9wg
q9NObLcPnL7ZgF69MZDFo1l8QpoMM7s/p1aNuEu3v4HX6C6J/1un4/JWo/cQfzKp
gWoasStuSn5duC9ruTgQJWpo63PCCZjO2LxzVChSW9JWSH80/19cYzzs0XlwrOOL
v5wni3371OZNjkNeU3LxHciPkW3iSI+A6Cfsp8NeuCut+IwhtyfSwCNMvRegvNoA
QaB6zzH126rqdfM68++tUS+P6OcGKNmFeOvK8Yq5D7JI0Asrtc/jtqXXwFPxtEiM
IpYDISL4VNqhuPE2cMaGmfd4SUfCP9OIO/gl0j8dg+FmXxMN/F/1HV2gxinhAQ/i
KNwEmDINStWWhaM0qho9rT7QhGQIozdhCUBE63O09GHZuhdNGKSfAM7X1iP5C7w8
xqepXTysn3wpYfMqqxD1Kn+7F9A+RzGA4KDwtVM20o++uMSXhkwnyJnp0GSHFD7a
P/e9NaFDsZbu1s2Dkk5lO2jjAX58GUCl2vMzgmAOB36JEeltVaIQ/kV3hcMkgOiY
tF24tRmqxJNHySmOESl3W91chFWPpW8JlfFwxrGzW6v9eTW1OG/9cGU7UfkQlSmy
rNmw+aZIxLGIAcp39D+saUoGWPXDYd5hSuX2VMf7FWw3xW1c5Aw2RPBgKxEA5h31
TCzf5RrsSyHLJbpVV91RY4KSCGsJtVYmZkR3WCxpESVnbjv6LjtcNEHPhCmdGGKM
UdwNaIbcG+5/CmcEph7T+qEaKT7gx9Vk3z0d/O6T+WoiMfRf8Sfmio8XBooTRwhi
YssA7HLlshfAkZ1GOXgmZVmJTSjrgd474wsjMle6WfmgkrBFwLYbck+GGCVyXOwF
L0ijVj+7otcZZdV7eu+Np9yw0maK76S2wqDxxJgl22ODIcbjbqAqnmB5KhBCDi/v
uX0VgQx7JAsxQeznR+xOVEbU1M+WPh2RQ0dm+fgZksCGQhLMATg5FxRoioeCiZTk
H0VBBFIlrSswP1fPZ7T0hNf6Jt3BdMdY9lYkjUhmrxapToFFwxw+TYBdixkZ2P0e
wlGs1xxISsgin+WDdnaAF1oSZ2IuA9Prq7pa5NjfcQFMlZ7jF2PGo3pDlnB6Dqsj
H/bZ/Nsm3RfKq9+HNrc7R7uzblb8Aj9a8qrsIXuZZ0rHxkpVF6hPfCgbvdV5dv6y
s/Tz8zuD2nvpH5dtdgLF92Eu9vZUiSb94bzdA4xg6Ic7Wk611nvFYK7shgX5bxz8
RD9V7MvVE0mTs1ddwpHCYIUI546pvYG+0WVu9X5TXDBRVzDGrZMhaKO02n91cxuz
EZuG1IKJ8eip+NeQkMzFKZXe7mB/4WnXW7rqK+22Fl1wpJa+XBv9Ycvwz5jLuLx8
RqKNjdCxGRljOrZ4Kc09g3uV5oPPQGT15WkinHsFV92S0MgnbCp4eXedZVg9FbjF
TEjNq70Wb33KV3KcjpxdoWdmQ+xBIh53pihQoFmpw04nFB+N/4f1ivKEElFuSX//
LctiHufdfvLYKj1zoxVBCioUYbSEHnpmO9Bfxk3ygxJqPME5X5teNxWVLrHgTVoS
GZ+QH89XV5OPNsBVXrseL68ZJS0mLkCIBIapPxmdn8Ftb9O83EC84ctHNSAnbToc
jCDLHRTnc6qbIbv2AbN2Mu2ud9z3dVNen74EiJC7Gdp9AjdaBqzRp2yiG4tSrMVl
dVEHKq5YyZMcti2i9WeSynZPK/S0RDQy8v3ialkluJU4yDTwvg/i/cEVhk09O8eJ
xThcD8DhmAHF19Qw1axeDaxfAwFzybZSvXC1Qxc+CKddJRMDGSssBQOk+MO/aXHu
5i3BJMn0JCcyTwv7kCUVKlNuHcJtupJABQAqW5LBhpndQysK/OrsZQNgcfYLjOOA
Pj9UBBtcHkOsRSI/64hgbeOrjUnR3I6jPxjwAQUQrzgDQjbHmS53b0rk+l6zXSm8
xLNXPLUlLo2khAjThqj982ztiu5QNg3Y87hCbgaQj7omDZZKEtt3Y0kyd52Tqbe8
aIz7jAiEbCSi4Sb6+9Y/zJXtKROld5zxVkpEGKxKNTqpft84ckGkMzmTgxx12Gf4
MoNbs53JRd6EaCCZkj7NLpEiyF0K0Uhv+Y9KLpBJfxgIhVSGklXuvtEKJ9CBgDRD
B5dp2U5OM8Bzjxy/AOcmn1TwWOWlSG75I6gWOMq9aNNTc3qh/cgQlnSKlHqfIuIT
u/OJuU09zq8f6rK89hoshRKjiFO5I2/pPclx4Co5yeZbdDkCLl7QQSvmVpKZwPPW
TMfb6TB07fi7WGnqkKGhTKkKq11U7iC5cn4tRG30LpmSQKHOJU6Ky5uFwRsxPQR2
UaodnV+BIxpBFjCfa0FFPPVXaXVPx0O6MMsooO+5tZFvohJcleqamFH6WIqK5fD8
R8FZc46s7+q2ggkDTVcUhZ82xaDzRT6T1GNYXhQC1DTst45QDJBgD1EfX7Sqleee
hCyEQY/GpE1Z6N+ixQTzYWBSkbyTXfy65iDmZcpf1IU+N6eZqM1wlv2SnvqOA68l
wy/KUwsWqFURykhcMU1C+BnyYaEVg6vGmhCk1GoSiByreKQcHh8d0gqJCab0ptlU
fbjGIZ+2aykdQMecvcIoE//vqUja87MMKbzBllvpQrP70T+bMp/hPy0p56jyXOVp
lKKN41/7oU14Xcc3ojeELBqw/mTeyT22hQRhAe/hHPbWvB8I3Q3mLEShSU9YzZXz
T0Wl+TJAFy38IGzlEFEgcgBOKqgzMV1TAmeKn/P/liZ/XIAGxG++qw5AWOq9milF
DSTiBJYE2FBPmlhXGEmqUk8E/rJkZ09uAZvZQcaOjoh4Xn1A92ztXlvrk2Gsmz78
SytY+k4vOEh7HIiZTPJz5m5BYAWEu//4KrLp5i2KkXw44YoJeqAJgGQWH3n/6Vz/
BlFMGqyClMl4bPyirrIvojqXrH5yUctKBOz1RV6gFTzTb4L9KaM8TCwiCtw2hsu8
GgRF/62eqKnPZylKE64b68SEd7JQxKn18bT2ICQhUQfWxy964LcQrfFf6NfilneL
j+ANX1qg7baxmoSZ8wyVqD0VsrUQ4jJr3fKJmNb4HYo9HpGpb0EdGor0qGOZJ+Sq
7bScI5oVX5tlinz9Y9fbeYamWcXoHxw5vt8sMJxNVGfFWBq/ug5gc1tZtbYSBxCv
3x0unPeMKCDF3DFiFju3DHl/YvQIAPbT5ddl9kHZiZQTLuXuBOIaD7EBoDYiFRSJ
Gf4a0vyy0LlZX6vIdTzz0ToQpp1qlObgsX9EGgvw+RsZGoVBpodKCIn650sVumjd
r/DwtyE6IO2D0WgsYUAconnkVJSx3KKrtoYMervCAt+b33PCYip4NSZifWICrACF
BVkyfML3zeb1SGa5+ELnj78zx2tGtA7zLWKgoI/+Y/L7h99MmhKimBAiav3OJUa6
pqnYmCA/T4o2CSXYC1EhyQuvJBsl8TFlQFL/iGGv6x53Wx8fCo1fYH7VDKYylvzf
yybCRV7DTS5zJB/Qjs0inM5oJuPR1D35lCwouVCNJoSX6g9BXLBlqtVKCO8yw/QX
eXov3em3VcMNZKN2+2HubEveDjgRCTmOJ0AuhulryIRgnuMZj0ftTkrX+mRUCniE
PZHd2TJgJVWS1u5u7OAoypGHgspgKxM2x6K5gDZPZAZIL8mHbPt74xap8ROuavWg
OJZBLNezkn/scY47Pxk3G3zF7Hoj+d/bLIlLBNaDQmnJEsIcGQbXe9qOpFg3PXKt
5P4NP0JH8IlabSscEmk/eT19BbgjVeGTb1DfW0/fwO/VJZgHOAif6RWipVB7WM9c
EMLBOAKrI4nOjslira9fwi+Apk15yKNOSsP+ES09Yf5ATgQcZ5BUSKvc4auXi8ld
+tKRN0q96uGxd5QJDp/K7I/lQDnzbmQotgX8YdrULKo+KbSeD+2JGsnvVqmGzWD9
35lEHNZP6Ber2rFzkYVoXTAUzO8XPHRIzUSCnOdxz25eEeLyg4dNDFGeqCxT4OJv
1jeVPA6/CI44jzTl/RVVsOi/4u/uq19XDRyDMjiTBgTcHVaEwoc01sl28iy9qYW0
jS9LbtdSt8lx9vOL9PoH6tWqPkDoH5BM8fumfhnKepAaBUU9de6RT9JaiK0DTlbS
Yo+BR18TXtI60dVvie3qxw6aa3KUbYmS+s5nNGyzNFtd+SrlyCucqQ47kYezybPi
js/rB32RiikuUi8Qh7ott8FkXwxHJQymNUIiwHjJJI8Nm+fwi+9yFaI8ZXE4I2qI
3mKes5in66cDo0S3hcADCI3SqREh7m4HDWBSkOxyGwmW67rlUzWGGYsKYArjofm6
MKd5m1htWGnFXwRatUAEyHKdt1vkUC4xdvq6fzjMWDq7ojJQI90nqZqmVACEj0oG
Xxca3qVtwhn037PTqaJUprrdN3RPT+0NfUMb3VncjcF79P7B0yhh8r+EU4qDGxIF
PtGfkSVxo1jcQrcBmUdek5cBhWtz28oHSQHaVDQm0KVdbIKzp0/Bv+9S43lzz2PT
03vfLE/A2h01gOLODgeuU9EaP7Q9xgnKnrotint+X/1GYcrnftXjFQ0IgNB5sz1v
QhwHf8KZmz4qayADlK1ZrbqAtBRaKzvyZl54Zy83R0Yt1QCSfe9IUzhhJgtyA1SQ
lLNWaDNKtX69g4BH400DUYjRPnuBF9S9GNHFtofV9hilP8fH81lVJlJjdcQjryUo
P4zHHh+oHmrvqAJM71TVw2A9Bv0IhOluiURywa+yfVLwxmKZMBHkBlxlVH6neKNa
+AD9RW9MSLNLxH+M8+AC3qfh/JoJMAOPPDHbsA3IoM4XAch8T8cIvdYG70NJdH3b
SdKI2qNJ2s77UFnirZ1ejqY2lZO8LNphBsSNrrPpn5OoP8V+U77Iu3jVHLNAVacI
tQp/RJsXZzYWijTJBCNdH5dJjWYkAenHATCp665g0El+cMmwzxH/HMZMIL8tcLEv
CVUTz52kI8taCcKbGQbVHYA4TGadfXTD1/GLs+Aua+ReEqbpoq0ieWGJXeOvWtxu
G0pCS9eVKlASDfvWafryzx099PiwgdAzsBiWt2uWhLFuyqWcEM2cUy9nVlG14/ag
nxOU0NNGoN6HExmie65yaQnlZUN0oP3Atqh8EADDKdEt6w7UYyDV6ST/ZyDa7otx
X3mThMVUjsaANnP1Rhp4hMzEGguMPOEnkm1hhPnZUgQVKt3Pk2My0w7uxDvLqSeO
1ZQTGcb0GqGn2ZrIRcKDUI5RBfiyVLZ3onBtGu1TFmis95XYs99UiltsA10Aj6H9
BuBG7Di63nMvf5cm07hFVGxqLoKjxFm/AN87XtmxHSumEetYoSOysxrNeIjC8Gs6
57vBDloCc24TIeNOzppsUyoZJzSK548qWieKTS3TP8rF8BoF9IaXRhyIZLSwNIHF
1M+YblRP2Gh0R2nrbSDSryFxPIlWUzP7Soz0MTLeiYMHIw3Vi0vF0mcw455PcCAs
3yzDqCln7SBsu7Mn8iyjbgLFVITldRq5A2u7XpH2fTASTjhNsEOx61uC65cXLFTh
Lf3PxIlaH4lvB/eds5iENupXB+FbLqcD3/2MR0weCO/nfku6MlT+GgArcqZiYJ1n
oiwDSZVO5G9O1ZkIOKZJ3e8ZjVpzTEvuJRc1fV09RV2b5/SzSEva2AVevf5tyz6G
S7jXDEnzh+KDow6GmR9Nhw6v09OTRkJ1ROnziQwmYwmhAW2a9gl2o7xk5RjScWys
UUg22Z9WpJ12v3ebsaBuHENTjJREeti6Ol71kZzhozWLu1ivw9ABYvrWO+EyO9l0
e0ipNHjci54bzJSrr/1nb1IdIjL7MN2TM7LhpWu2BI1tVC9cNvko3NsfTr/UiD+4
7aImnfyDNxUaELBI7WvOJnY/fO77WTMw+FrxjlOfjbuu0DDLvwh1d3rKY0pC5Dzi
+j+5hvhj6NE94InXsQPD2JKUrO9Fs03sHGBNzFvLj9JdoR1+rlkfWPZoFs86TtQU
w4LUVzxN8kLZvDcoUK9RMUJm2saxPSR/31iENW9FiGRUMG+R49fqCDiHZhwJOb+v
PiH4rCuaWRI0cmTaT6Ui3LkSOQjIeE0sdNMxTwaPj4mHfKHcpO2PHGzYkyxZcy6O
dWlqkFB6ulRrEqHKNgNRC7EQzmk9633HxXssqymRzsAjSN+FAKb0sfcbAxHovFfT
M47HCIi9dOWAcPF2idEc0D+jRDcRNVzRAgPK/kltJsuDbytD44kCk4XhToUzzOGi
RdcBJanc/vVeLQd/Pb3RTfI4K/Bjqroyy8/GfRb+fkLOWqU+D0d0GPpNJaefdlB9
YUow+zKxghDIhMIe5dyCbJf8qY1Mt4ZiZVBSbzY2m76Vq8BTpjIIFIpPm8/HwxMl
2dWmaLkrZpAAahqkpU536/4YYsq4C9INKe3Ds0ns//j1D9wRuG10hNosMGXj13rZ
ph8qqfWopD8Lxq/H3nRT3uN/e2sqcHuJFuWydkACSqS9BnScUK68QRdSRtIYO4Dc
w8Nnqj0r0snKvnu6zVp/dEmrkCG0ZeU6oZjFzgAXJATPVQxM2WEoOfwYXgj2XE1z
+n61cAu7qTwRvr0nzbhp/R5ZCleo3ZyVEa+jadoItlJosnNOLXqvDNZdmu7jd9up
Kfpe+awJCvAV68vPhG15dE6ribofrNvrk9ipmYdt15gP29TocovaNR1zDnaxzHCf
tKXQAgpTZOusCgvKejo7gcu/JenZSus4qzMTpF5moEJKf5bR7tDZ6SMpwkNZr47C
rhe7rA7VPXIln1EGHYvZcFDF2LdiMAB6zLjczk9seR4ULrM3b9HvakVQFcLjJGNv
0mpgWcVraFglsk9PGhqZldoNaOMcdzk+OnSOGFMZAcizDrj0P37lsvJda8t4hW2p
1/XoNDc/nFsxAglascOA6i5J6YYqdzAljllyDJ8rPwM9KF5AIHDizZzeYS2qqLIs
uNclqCYsjpJhuxsxnAtaxQDwCWgSovHT9Ycs9tGk74nvQyjj0m4lip788Nx4YqEQ
zyDlWyj/JKbPkP+lu5PxJ/yBwVB9L7RWuCjPG0iUUkv0jUIUfKGUE/dqLtx3B9ch
iBZDa4buEImxbKhhsaSSQlgDZmr823pCtNE9NtGSCrF9LQVztwHXe27MrXbrKogK
2qSo8hXDnhntCKRh5arJ6Y1xvyU1ntVI5ny+Xvg7+jDoY2jaOEdYr0Qf4//8lo+p
OFBFAAkRiCcodoMKgnAq99D2mZnpcoyUUQ6Xm80Z6W7aMLHrJePZpvo3/GO18287
YkAtKYlRl8bmTIfQrSzjsgIJRXuHn2U1Y/GKULgzI23OqhdKwr5G9zKPaQD/rgsp
LJxFzI1AQRCsLtjevrA08g2FU64KyA6QCPHXRqe68NIOmNI2ZR7YwxwxjcvQ13h4
rWedX58rbz2L4BW3YdxARIGF2r2B62xV3AjGrCFCgq8hRILasyQiqEP5hHGoTTqA
Wwwxii0qWXxUGYVA/plhiPf3A2WEvuJXakQTWa20XYvruteh6gt/fqwmVcC0xfPZ
RQjpgM+X5ieKdGFeH0l/5v46ca18MCHgMsOLHL7k7Ou+9vS0Gz1riJl0equAtpSM
PI9zN/Xs8eRKA2Cka49kw/dcd9OcEUmGuR6BSqjafvcQOBaaH7EJanOXe8RyJEto
GJpA2s6lc5Vqpr0C/vOdg9DPD3Jm8uppeyiF+qyVIK4mE7zU4tU/OJANNHQPCVBb
9oD81eJdRSmH28eMueGHdI9+lBq3Ox08lwbnXvzcbivVCTN4skhkwk88oc33CzqP
SqyifHKMjs8UcPrSA6s/TE5Dat8puUHp9oMDAS3rKXbX7LPVvhPk9olRcrvQIIPU
ykfNEDLjQbrDdYkDDuXsmQwC7C5lvDjcDRyggE0LhTFq5Bh4HnKlfP9DTLv2ejjn
pnUDcdm5nhMMNenIOwQ+dBn2rOARpva4XJ3kOcq6XVrNC5+jtU7K9F5SWCjfSjcZ
pmdTXP2+ReJ4gwStwWoZToff0W8/Z4hcK9qNMRT5k5rWUIMDhMFwX7MXfImivI/W
SLY7zzQbOokRfsdi2K+YzlWKsL/DlY98yyn+a/xC2O+uRhNA5oXPX0+F67CvE92o
ghGqkRNaAH8XySfY/6+S7Vt+KrM37QZspdiWggV7cAdrWYA4owpAjnJZV6Kbwg7w
qkMT96wKzQptxB3unp0SaK5toNFz9w6vtdNqF5EMby+/9ZdDo/2YUDjFflRrgpxN
XpLznSniTtZfR9nObZ1NSEfHO9q9lWMZ1y5s26aYeaIgPQwBPmdJRbcX+aphDQvB
/SqQATw7lBv2QdBENmwMCq0rQwG6kaeNoV8UkaCv//Mhh3El+P2LzslGY4CSkT+f
9P0zrJnpRl91ePGUxbwCkHAncs1x79fQbuErdSAe967CjjNjRRt/2ER0135SUICh
82GeCbOhnC6Gttd43eAVztMlHAzZgRQ6X2Qaoh7tO6rfSIttCAmwT7eAaWM70+x7
ih0ndn/SaSAJ3FrE8d+lZj4vsP5GyBjEq+Rf3GSRvuAWsX2VFRN6nC6gqZrsvz/C
ZVWANRdoeu5QqdeyUTE57PZeZlxX0mXObfweD03mdy80Bo1XJcJwJOMDY6XgfE5F
ZaRCIQFve8fRb2X1GXEDigLu/5aXzcT38FPBSvK9sfVVDLDi2LvSWB+zntwHqGjT
KxXYOu0ZB1rsq0VQk9ls9ZttUGpjpOP9zID3NSdXwSVjUqd+Quvki0p/0+2MTren
VrYA1e2SaGmwy/R2aZOn8l6NVeXw1qlDey52Qi852VTGdzzojOhWS28csJFGeEHx
a60EzEKW1UTjEPZXPakdzM4sCkFqyNf2NR1RqNcBUJapqvgZt90kI8vF4Zye7cD3
TfjlWRxQBNIRPb+JDYvDUOkI1JKgvAjCEfdGQIAZ5RdS3wNUhhidkVuW3UF1kBNh
ibBKg5/k2c+j52W5VlkFhWqhorerPPw56DOmCdda1RzbY6HVvJVVWn3Wfk1x7xNb
J9Dhk4QD7WgsVfg9BnFbipVXoxDggxyyo3WIwKh4n2pB1FQO7m8HQGdmZ5w3/95N
cLVOGNxdLZtihzuY3dI2Jd8LQ9VuwEEuWFkRv/nugwz0k77FTUVmHtiJ3af/j5g8
tkTH4WjfzLhQI0cmW7k7222rEzLkHz+QL/jde87xo/eNFOwniOhGjf9PxIS3L0GU
h0KFHw2hZf4f3delUaESVuGz/3NlP3mPUOJOIFtzLUNi6vWrTPmpHQGQyFKliA3t
ty4SNQT8ekNnqB6LVm1RpLwnNYxOJNrK2DgmWJlq9PdUwllXRDcZXkV0DtzIuj3z
59jC+hPcfUiLtbdyDjF3mwfJr39eIuBic7caFCIhdf/kjXcswFQiKzpB40xTgVyu
uR+ChL7LjEMoObYSqPuXcs5qmO2nejgCe/BcFFHrrrxCr7g7KC6jLWHIxt15XMox
wKZyPqOxC3nA/D8XnbbEdhloTizpIBMK0u9PcUh7cTUIdWe5DU2O7KWjAiPm86rh
eOv4SmSTTjcbjOA0j7kV/458nGbFaojZ/kv/318LdKxKQi7KwVATIakVN85cdVrQ
zpTKjcZbMiz5pk7azKK+GUWm6LQHMSFol00GldMbEMmLzUijFDeVQcExx6lJRRK0
zIz88fXCrC8CVbQdtOyLR7GfhC9td+Lb3uc6fpE0CJM8f1af9LLaHyc+VHjemPbE
pM5JPz9H+x3KcXBT0bFrluK2Kez86hOmtIaOi632Brrx5cIY65ZMEiKARlvIeo4x
ydgcnJ1+Aq7oQCgorh7YoEGLe/ryWxjovObaSjezM4LqhX2BA+/SyP+b/JhczPXf
xUun11ilciyHPb4U43qIxw4K+M0QEfU1OC08MxfJJSHzf/Hv2u/9jmst/eapRIlN
H1Ci1jqtxE7EH4xJ7HhNlw/hyhSebtIct9BhjriGV1jGEcUvJlTcSUXapCOdbppZ
2ytOPAgJ3rOvtN5QTfFAdzG3lA5vrWXo32Cdl+dYBL4PGm+pr9Be1JiimK8xx+gB
q7T+jzDGgdd+TzklPHU784emq/BXLuA3fjyLFs7jKZzPbesvjtffiQfKSKnFws27
b/QJOr/6zZrEJXGoyE1eWob9J5B7ih1srBJ4z+RT3WuOYe/iyJCq53fE7ixF0jDT
yPXvqof9x2UPIPiWrBaTcX4dMIY01lXVXdlOxGL4v2LV7/u+JxHpxhAO+fQ8jD8p
EQYnrJEvByyMl4BOCVA3bInDuNwvU6l+pmal8xxqx/AXlO/dW6N6unhiAuSsEg0N
eYWcwEXRW+m6y1lsaa0QhAYhg/ZnBbIpP/yrZhIPpmyG58DS+BW7bVmbiQW04FSG
7UdiLyUJ4AdWXTuEq2CN0RLnGcH5FCJaUiSv+pvQSqu/bTFriGmczfhyK7WndKbM
8FZTBQxj5NSl1ipI5n0GgOuFqHs6WlNjUJDnXTc2DHO9GSzVnsuayVF5O8VR/Kie
bB4CTlTwVcMJuEA4aesloCdcd60VN8t6Zm3iOkhDIRq2CxgOI8URw19Txxwl/61k
fy5uzY9oECR40THoePkUPE3YYIuNFYnbLoAceeYQFQB5LlFdGERC2ip4fFLiKzIM
W+tslUvMRLHF2RTuHHZD1NzESjFs073/Pn+RMOhfmYOJWJo4R1l30FFk/TLAhXaO
Sxz/HYdUaIGjpNu2BP/JapRuXsVcqk7uwWqKp9E3qW1t676DItNEmIjrhC1vDe9f
uLIbAN9NfUcdyCdN4OPNAi/NLEmkaTWH9UYb2q9ATKoYsNoOYvhFrZaQAPlxtMZH
VMiPfl8dl/auEMx+pP1XvhySDNHLWNy4KriZLpdMj6TDr2UbWjF1P3jcyTxAONFa
A7kZDVT21bmrv+jEHjf5LLVuN6dosgF+OdomhcuaNVU5WHvtO5Czl33GXf7QHEkh
5Y2cdpnBQqKzTHRAa0ebTo5ldar7r6ygAzo5qJMaek41+ngAeQLl56MmPNgIKfas
f1K1nCchcII5S5c5nFFWVZ2QKHvzUOJxECUdwACfDatZ5PgcTVtyEBg0iETvu+Gj
oh/xT7U37VhLr7QKt3QoG9orfCtOIuke+4Dti/cJf/UFQ71XtRVsaoJr59+UKiLX
hAdRpQV6S0Qcu3eT3HujuCpgt+spuJ6SFqeoWzC8hLkkGf3miZSbNcJuM7GbUlFY
09YQ/FhOCmuE8nYdfa/EOinfEkGmlPdqvIklFzbn6am8FHf478i07qbykORpZjyu
xgGCNhSjWK2uAxLw7nMxku17ejcH/1pmd1Dfe/OytKXGKfRtDTg+iZ6kMRIdFx9m
q3zosrUEKgvWlCDhy2p0f/RYlzr9nbvy2LejLAPHFGPeio9xCW8YojLFNf+XUqMw
UTOwvQ7AQJ/spmKzei5kCXnlZw9WevP4v1H2NwrHdcI8uZIHcKGLmob5woe803cV
mqSf/+9VnuZLu037zTHjwgHtVzn/K9NtR2EDvgGhuHjZU5GJO4pITsugmOPY1z9X
VFqal6xgKXtzbqqW9xXCGuMucl8xF1Pbf8U9daeh9FSTzmFSXYvCkxVRT++QGmVU
qf09gYGr3sp+E5q4hvLua2DaFCoDglzuBzOC8+ZPtSPIm7eGg91xKF9MBFMrO+5z
fbSvIaUDYpmymbf6tvHy52B0Sob2TZhNT762zEnpFKCTy0wrZixD5Xz76ynbtdjM
DGjlYaVxEZOvsqEJfCqu10VeWWIZ7cSJRL0mJZOcfmeqYKJZJAsYZEJ2Eeo9qX4V
BFIMi09TWx8VxE8B0GLMnoN29M69QyV3gpwV7o9b+YnFuoLpNS84t3sDC/1z8BDM
QfO75LCg2kkI/TdNcYquLnZRDOLp6bwGUmeSIQZB+ikQPmktRinswANrLeq5vWQi
XyotELq6euop3Yu38lniVYXN/P74A4y14nDCXwM6RIjWdDJTf/orOL1i627rXMbX
bBy3pYMRoXFLvKSOizz79yc8IQw5S82sIpSZlJpAj9suO92cV21vBpEbXkLhuF4z
dmm2Du0tRsjUCkL661z05G65aQPiWajqVyhaeqRjcHBb/1mp8JaQ1nT2OoBwyrk5
sk5UXRbz3sK+FvpQr6VPzKr+yEO3Ypy6zeOyTFacmvpxhGoUuXRCcNBet/TQ94Ql
W+S97g3dQJ+OhT1TQZEUI+qSh9HpNEM6Sxcq1cuaL+FyTYGsKkJ0f1WC5gzeBMFl
zNPDgObtAcAKBEbmczswUeD8rDZwJJqF5FfeF1FyWhRUfhHgYRXgKY6WXNb2DEC2
sA6kkD76nId6JF1pkDkwCUQZg8nn1V7MLfjBJMVp9Pc61TK7YDdvNraT1clzVlY4
sb7anxh2iH5/7rkNp/o3rhZOGuQJUJkRBWPB6YE4AMocGFDWIWEM2sKPXhI90RDE
+UHKHT9gcrUW/I9JYu6pj6SoeGBBk2peOHngF8KXcZrkqfS+o77GV9VE6wNxvrw4
aRDSpanAhV7qraI5ASmEoZVcBrtTDieZTzcrdrXHtuOIJa8bJUdI463qF87ppVDt
kckKIIhweJLf8qWHLixG7TjGlQoywL1300t4fpvcUlMsuPP6NSv/TZ/uW05bf5Vt
qI5y5cdMteTBzvNj5974H624Rm7QEbB7hzDochlbyFLJdVFnzjj4ANxsoz8jNKuj
a/HC3jhSP8B2v4BcoGt7NbXRw9M92iqdvENVualCP+ZIjw07KW1xHV+t7N6YmGRJ
Qof2PzwdUAPvcadBofuOp16fxSVkZBllt51A4sWbXvyZHvjca5J5apDTERSSBmHX
Fmz+2MosXK7s7STWI0+Kw1ll5R5hQRF4P48YLyOrEsktxzvf/ga7zn6V5/I3c+JT
IaoBwwHogmFFbklYvu9J1lUUHUplm6oe6ANXL5Ml4svInEA0N+2yYC1BmQY7vIW0
LsjcNOMxWuliB87EOdMKQbU+c54VxK57Ae2k+BU4Gi2ec19cz1SJuAWh8UXhuIOS
ffucq+jH/VaDhFKWYBje8p36CtCLZ2MX14ZkWBIWd5pqtJXXKatk+9VtAiHzaqnO
IKdniR7mhXKhjhg2/+zYTDcaY2IzITXi88O3O4otp1NzrNbTOmrrlsRMZQFY4f0S
3JJ6VnNYyMCtrlQTbaCV3ca7MvOxILevRnVMlP8//wfhDYYIvQG8OrsL0JJnPl3f
z2uzxK+yfQ+aOnrr3mV8xTwIrXxXhGM8On/i5G9rNdqMP2uL7ltmAUuxqQB5o616
JrXcYszhvYRjlAQV1OJ94e+YIt+tACWKEH1NdT0qpse1z5qMytG7xtMAFteb0nVm
C6K8Ss0QxzSW7cIkYN42n/cnMh/Ist5FQV8KIL3bT3ijBiQQQsgWuKMFJ3Lf5mTY
lJs5S21NBTvsSW3py+gnoOlBVLjxtukLPStFHFoflKsQ+n9P3YwL/2q5SaQ2AIdu
CKXqQ9V2YEHvrcTW33EsFrd2luSLqAnzFM0GeU3z85A5x8Ytzn8Mz8oI9ukeLRA1
/5maj5BYTShzfEBXRTaCmAblz3K/+/WQ4bMtA+L89RSXG29CAY1rHjjHm1a88e4U
ddCL0X0AovXMgL3B6qZnqlGdYl9Q3PEXBxRxyf2nPlYw0jHP9o1Vr61ZUHZwZvs/
eBmeYLvJ39IkxtxZK4rZTbylIwh0OZUnR7+vB4LPhD4KFNQOaQYapreK85RhGjSN
nmda51lFcsvxjcgih7XnyPHT174BGZkMqvtWsup5S+y6QUQPxoojHbBdszSI1Br8
tM27mdpeLgDBoP1iCk02P9dUEGZZkzSEF96LP/QH3hVLxdLWw1xNFrSkvw8CYZIM
zJTfJMq0c6ziP1i92Lcsb13nI8Y8UyADTinHESNRXLxR/RhwDArSvylOlkyh3khK
p3zEK0bMgtSZr4Ytt5fvVXfxbtSle39cpXqEfWcawj5UH56QTpZc8NIVHUK7drr+
mG5My4Bt78pj8cEmprh0YRxavtqmgQUwUkeJSVEwnG6NeWaZTulumMMuuOKY2xBy
/CKxgMPidfbyZNyVxMDyNrb+4MfSzSIxAT9U43oXqgeOyoMxbVWWoemGAgsumuIf
hFc3VmCbT8ah2H7gfcwNBIE5U/OM4zIssGwOhwVyIGdaOlEgdxb/wtWq0jla44iZ
Zvl7MUCfnh9e5xy0T6BVn9vA6yEVE6MIP1LIzkcU7Tw9x8NwTpNg1U9PNF2VPauW
9bxDXqJzuBp1sXssQACZ2a91zzstrr+bKfF/7jW+4zJPhuFiJZ51BVPqLsF+FVdO
GZbRgsWn65kdfn3+QptSUhJDgckS9ye55IHvsHf2PcpfFRpdAQqLZtreaT5Dnlyo
LRBvFofeYC+y4VDAd6akoEbilyGKmBKiC6F9zEBMHr1PsNts+OLUchqF+Dq9MkEm
oxpTB9DqLj0BtwisrbfY6KnA1532fkSJuLtTQLQx2DCpn+0XeLkrlV4GFWDc/lqo
cinP2SFFcObPZyZzo4l+kGMuDZZX7pkCgDasa7Q70ipdg2NH7yZEl0utQCKkJG1+
jrUJ79n/44uw1yFjsvdbO3TYzpzX7PW/0CHyH3s8T8UFuxYAkF6NUvjuRPsdHAdq
pQ/z8wxdWTSXKZrkiCVt4PBCEo5E1ClUXHHCEUF3vKcXdrcOl3+ACRjxB+wrijGD
PNwQpyQhgRgUMPJ27/6MpeFWG26d7w8lU8dTL5Da2ISjs/o4i5U3RwXdC+HOh0ub
PCpFwVO7JQTAC8tzUT8x8edizIkRKgKxg3vQEiU//qRO/GjX9iEYZNW9urj8NCKc
3GOTMAgY3EHSoL7cTdvNnz/iVRxKFaQ6MbmiZgQ/BFwjhy/20rvzciJZMixY1wnE
kf/CI2brlRRQ/9T779P+KkjT4Y4FxNzwee96V3a3jktrJRXqKXVJ8UU54oczXfqs
aOZkxNrf06kV4UIx3eyRmz5AHxq6Nw/DZv/D0Nq/7xaBbWOz2hPQPhBL9KjHH5oY
OLb4HDja5tqi6PIjNkHffRmlMDHB+wNCtCtpAK+bYx+oqQdnuB7vyowa7L1xl8ld
fN2g7KU+1wMkawLgYoFgXhfCPKHgPz4w0RYhLl3gI0w20QojqOLSMev/5xqwyGc4
zqx0ZPG/7XcS5w1IkbFkjo78yLyLzge/BR78Hzx3kKS7pogQJHfpKZ3R4h7GVkzT
3fO1sXAg+j/AKSOllH6DLJbWbzrfon374vwbfTu2iAlvmk8npemKGUHqXyB5Ijc+
REiw/6iz9mLmEApyRPNkCsb3RjGWrIZaR2mOnB/VPwH5DNMSn5m9B2zW4fcJIaJs
UZR0TdQH8nM6iNhRzZKX+S76vcQFEtSSFjiPcGSo2i3r4BdTUrTN6EszPFVpDUuC
NIsqcYEhKtXZL5opZpGXb6BEqgkG0EGNZfQyCWtvkxdOs0GlmKxWhX793jQp0Hsy
bQsh/nh1izwQgQMhmyv1UmmbzhhGrJg7hdM7tD8AjMTazEhlkq/wUC6CoBQoXSHc
S9o9ta7rwv6n+WNgUnBA7bnK9D4yFDjQAWfUfiqmQBa9sY264r0Y1dg6xjf+6oIh
n77yji6pJ+xndbNmKF6egZuffcpQckHE1oBZwlOgFYC+azYGenAcqiUtu3yKxbeq
SV0ghptq1PfU5fV0XVltMaxPUhQo3RmN9Vt24OuBFKzbSFtJEYNtWHB1D+RHoq8M
dASd7mM7Er8Y4DjkRTiEgRYnYgWw62yn/0rztEht3xEoMxCAXUx5GE2ivxIH7sAn
FYIDZHX8Q/vRWy8qU994olmXD4JPrdW93hBdJlgDcwHG5QyuekHv1RGRtRkr2qsi
M97GstS4fIMdLx/cQOkruFTOp6H+rmqko155U1lg33vgC4CIhuqzF0Hfi7VfDWwP
pc4/WQtaV6ElHREHbe7MJ4QC7+INtnhnFiZatocZOEogPXmLJ7gKGyuSa7MDRtCq
MHDfQTdHuV9PMFqEmTnNR3sY6gEUwJMmFGLLFOCu7EWrnokOlHziF2TUipGvyi39
n5U+y7etdk9aK4o6D4c5OmJqH0+y5suLyD9ug01KzSjGKS1xTksPBwEuo9rb0Ktj
Hbl22hU4h91DmZXz6W5urqOr0g+7K5jRClIxYxi5mjr95pakTej1EaXBCHlCQOjN
dkM+q8L6lTFPVzcoMC3CHAPgecO/vxP6nB9KGEdPah0Q3H057O9deXyqSMl3zKyZ
3vL4qMvJCUCRCY5mTwVvI59TGpTqo5Q1g1vO7Fv2cBy4TJJuQBl/nf/sBoJNFIf5
hmpbzyi/0ik066V16KcQMp7BlWe5TNHxxOxotv+eqKZtWJLB9d41r92DR6/qomRx
/kpgCbZd48tcez1sS2/Hk3q68A659geCCUuYe7CmzG7WXydO4/v5pWp7SzqZwnJw
O+rVR2CtNtcFRi1cTfmyobDgbvm808KE7Ac0nS3c9eM65Sx7GrmhwLaSWhYf4MIH
QwMiAIpWINZiW+DvvP/SAPsuE6l2bXCNZfFwPCcyOljSipg5KBYhWw3z3GfNu+CE
y8B/EO8Egni9ZCjnghf/2pwomOfPNoGncFuralOd4IIdxC/ve0wfmN9Ev97eREBi
EloCCw+gfH5LwSbCSAZFrxUKlvE2znO5ndmhLcdBJ8EkQEkwEKlwH4PW0s33cJ2t
gaVkeREm+xOMJ6R/Wpg87O/76oEZR9XER0Yp4Ze4EUM3WbjRkp95ZTiJfP4TooiP
8BNhhH4tJR5kKhNvvIGAwymcW+dAqOllkpPhMbu4wth8PmJ9RK/CQ0/pi4YNfRyJ
3idUnwoHXK577AtVYk32T0d451a+K7zPas3n579KwB6i9p8W35F8aUL1NNbZMZyT
t/2Y+iV1p9EkKim0sheJcxwCwwC+LG3OZbg4+FAT9HwZ/TlXhwBM+04zSneS1QHo
wAKikpxigRHRFIzB4OZL6XvtAUMIIAObbYHTZHfWJrQ9vphdCqNWJYS3S6e+lO9C
VSX2G04d7GkGfBadXlGSoffxOlCn0bUY6ASeL/shxMLTigGcJ1yvtOXEGgLv95aq
B5iBOJkVvWXonyZvebTgs9WeSNQe2L04SLbTOGBy2bAt2ZEItbXjQ8eI7nqQrM6W
uPyk/KvrGCr6BW2m3HijgYopTNZlRAN0CXfWnMa4iDTlFvGiNNXS2Q0PzQPbynVg
Y60zVVUJgTzLYkSQqApf91TPoowZbh+e3gl3uKf6iezOBYIZZklaN0SMGVjw7ccU
3Fl3Dw/BBr8YPSiW4+XrC4Qry42ppOTglP4SvsqwxxB5Ua5OaFaJM7A/2NgRimEN
4pXngkv4cmHNrkEZp/WH7yinJmRSoFeq7CkgLuvOe8v/BiLnS+W5wCe+w2Cc/6/6
4YFI72MCqgxo2GDvBxQbclTsTIV6SnCIazxhHvlYIaPMm8Co0BWhLE668Txf/P4F
GI7nOVfU+AY1/Sd8WHKeImJd4JoQiwLiF5XhG9kgTktTA+rYxNKIYPsd6hhlUugR
S7+zZNtD3E3SrAJ1En9EBBf6rSOl0u76kz0BU4Zq4MsQTN4RlG4hhxwXFiUEl0Iz
GatY9oCWeeeh3mQA+APuWohof0PvVzRQmGIpyk9/C/14AiqNNXfWltaQYBh7ZX7M
xbid3aSz6e3AUUvZTgj6Gw4pZ8443zdECqdQG4FR59/nVY79RuEKYn+ap4yR+CvD
sHPFOzHRu9CoJDw0Yz6haNNfUUp+8rgg+Pr7b00upGBh1Y2xLtY6UleyLScu0Qr1
y1iYWndYABPHUxeuiW61xIP5GaWGIaw5tmnpLcOci9jruSEaW16rb6T3WL/u/jep
En45bgjB6+J0gJZnnWwQ+4CL6+udMoVvDv668HjayuWhoaA7wemTwKSlu9eACMTX
0b5QNGG6HcBO3/dwioC6uPkoK/U8GwrAl4b3ppFhQjN3WbWAuTvPhuf04VXVfVY9
qjkcH4ALePfPI/4iQGLgC0EqhY3LbEOyjzy1XzT1H0Nu3tTMCDsOlEq8QmzLNt4L
QUohNQmoP4mMt/6WkxZt8mxdmWeyUMZwt3QueeTP4S5emtwHly8JQ6zS9PkRaoJE
ub+Tub0x1KMUZeOeoEPJhO/L/gxZWLqeTLRWFUQiXxJebujH7CNEQIyUJBP6h8Yr
sLJPvesHySeQ4Am+WNE6Pz+XZQraCb94fkAeWvI/vn9OnS0OVFQAUzFrBFL2oThL
NOVZYi/R+e6bEloR7r2D2aHA1Xm0ZYaQckxUKpDttcr5eMq7FNBGgIYNjuAGJUYZ
y8M6m0MsXCuVPzUs87wQaxLiB7eHZAKO5/bBYuSd7ayfW8KLZVvH13mR2A1jPrPU
kmT5FIihWzcFXbfVN9CwRVMEHndg88snVnrvL79ahsc0ejOhNYyacvyA+cdVrQ+t
Y5aZAFHTjDHN/OzhJa9LlNVJ3pvjr0iy83oMnCRwoJq9X4QxTjVs+QFJgQp2epp+
31BR3FTQDV7y/KLTIpKa7gl3aoXYKT7Xvwb7Y6hvrjAihdOFTMru5mF1g+HUshSq
fMZ2jyatc2cuSIUWN2BcPJT8WXpoJk26oN5GAVf7byTfAxZJo00BYT8x/J5PPAo/
Lsb0O8AI7MGOOHHTqY5MUZTBDGbWX5Rwi3hYBSwHrt6z47qcUZLA/8arqDzVxb9t
pqvDWzlMGsEsMvTnssULvSpeeZqIkJmdUrrGdENY+/rGVwzNnsLuej/AndazymUj
f0F8mDrCTz1TMZD5uVaP5o0NOBcTbdTsnPPMug8eYvec/9si3erACzCNJs+kpGPO
tZfnbDPcxIJ6DbKZ0fkd155S6q/uLuGVt1IfL3l0CMGUp7FoBLDpYLOJhDFg8C1y
8gsu6xPzydNgHBwu5mxaNkWsKrJLriJhh1oZotDHxz7AGycvNfq9BT3AaCy/vHZ+
PvzFgCks6M8QflWt1F1z6OOh8HAnE+ZoWxW9WNU99Vq1rbnC2YrJUvwb5lyky3jH
PffqkaRP2vAdVBMjdcUW6MAscGJ6nllFAz5c88pDSFgegQ/mrcl1Nn8O9s2MwIDU
K8uZUllNZ+ZHQCD3Il3z5nZGHA2U4VOW902v5CKhpPqfAnCORpkjh5eQL+V72873
nn7n43qu9s4Vp7GUa7c+CSIcH0qFpYyKmPzhx7PWUs49GnspPgKkqc49mBp5iEVP
84Hsml+ADGKpbidlMJuzG61+Vgl8A9dhI6lXRKC8036p0io+cwadkGd9cBgvHlwp
haCpIP8THk7nDaGuHbC19mIJ/9gKajomrDCHhxXinU0TmKKAdM3SgpZdpK0ZRn/V
uaLwS+nTvf7HpDfWiFu86hSoJ4FdwF7WqnaO79lMAvu5jTcmRF3Y0/H7A70ZewVM
nAzaGyWht/vbOxOPYELfIs0i8L9Cz+8bWuDR4vWxx1yBddoYSkcDmGXbs5fLoyLL
DWVQC9RhfJiA1YfKUYLB21gaEJMcuR9dgFVVT6lYSsNgohE4ckZlSkBi/+IaMzHB
QTSzqvEdJlvMp6h2EgAgpIZxAraRZohj6es2d5sYGaD8L12vwD4BiPcwVVKHTqfg
MbbAJMmMi61lP5qClcWNKHO7r8i9C1nPQXcGNOWMci23+vTQ1uV03Xwq5/QFe22E
+EmGw4vz2VbpVmaaJ52SlYCDb949JEoFDAF0TbzXE+ae+WlsVhHPftnYjRW8oRqy
reH/UE1HCE74i7UtUxDolodqsL/3KvP1USvQ++Jq2ezqWTVOiiSzLHFyHsCnLsf9
aWrnhOnOUoFLR0xiKIlz/2XHC40sEriapSVOlLmcJlAwcQsssmb4HSu07yDaDeB+
84HzQk8fUKGIpgSjcdVk+Gw2f0s/9Q9XW0mHKPGqzd9di3qlwWeLoJhZ2DnY9fIB
+ytebOEDzfGwNJD4PEz4BVDfYgNllTZZaT8wH0rWUkrX9aiRKSbT1idjXpLbseKJ
2gdo9ykRZZVeMY16D67lNU78YLhOeTPrF56F95Xfa5YHUVm2AXnSNUcHv1v4XcYI
jvyI1qIydeC3uHnsbbEA40YJ2sJabsibDLHtWy6OamRNsATIiGjAeyiME3MyNQNF
4KFRnOj2fMli83Y7EA6pWsoGXlF/d1DidXHDBIfZOUkPLq//jvTFTa69tKZf2O18
o89tph2TkMBj6GSgCzKN7z9ZEm2JvYHtZ3xUH5FDl+Mna5jf27GmB/+aJuT4RD6d
OZC2gASAvaAvPxGK9zVG4JKTu/6ngzi2N3fFzeJllth7zrQBQnwonm2LE/5l7bTV
vdGd5RDBGW5WRQrUUYGaoqGE2BhRkoh1L/58vKqHeUf+A3GemBaMlGYWxg2k2in3
A8FSrAclH0La3vRU8LyGHDRgVK0NAmmLhQenbOE0aeqLxw5eWh3UxgGywIarE4OU
0eAHRJDeB5elDY4BK8cOyz6HlUttMkRKrQ7WQ26KMyFZhR0cOFai7v36d99+ls4e
yO+nhwfnv/k/+rsUMTCa2rBcTjk9ns6p79UQtE53aoDWXfX37KIu5bw0apaRlZHs
kIEdVUVjgNqczak1nW6SGI9DzMH4g4PmXSsf54GdM9KYL+BXkmgfTIGfNeoMd2I1
E0Bzwjudbv0EJQIf26rQ899RiryWJQnhCRdsNKnCbpcz4zTR0CBNF7kykz4tuzHB
jy7MLw/fdMJGPDb35ln9qwYJwk2AjBzDhiezU568iI1Qurq84r6rO0BjQcfsD/Dv
urQHWR0HoQ0D/E7RlxVCMF3XlW2jymcRUwN7xevChmospZEbpV6rF//di/y+5q6U
MCWQU4zbnTRaO2XVU3poWSLn2VMMzLWrusACi5SfeWEslVZKNTTKH+Pa4TWvtVA8
aBQgnC+4MghKGom2hdOzUkG4NU+RCg3WS4463U8rrFR8z8Dus/f1+DlAHmcVLTdd
4PYodAW9tAspRz5S09LwBPkl3hWd8iyjI6K0O0gC7HYLl4Il6xFXks/J3pfKblUB
Y/6bXI9ym0NaPKX6SXQAZOeYabnHMc9sFb13t9fMa808tjUiWpaFUJDL3igM5jUy
rSTGGgpjihJ+UOO/xuZZ85r4oU+50avZoaKLoLX1uz91sIiABYmJqIdbaj8Yz1VV
G4aN0A9oaSFmYxDPVOkmgcV2/S6eXI9q4JT9k3GWqWWtTBia9OMzTJffq560I6/m
PGNfoDXEJgEEMzpuqn/lvYkUrIv9H1hAmMFz208sB65uFWLX27Zbh2G7V4eNnEui
waAdYZFvx1QUMhgxEsdpWkhF8vlGihnlXqIXvhPtziH+RPIYVSpUKBblBSIcENMZ
cLBcGq1olRLSIRKbXLgrhXvxuUNiaiQ6hEh8c9gBi3GggE3DEx0r1pvWjcNQ0OEf
xF/Aznza+4tMOAnvh4B78f6fCfSA/XgP5dmVY5U7ojuaAmBLB+Hm8vA3J38XTN8I
ag+f5n69wAhtfXUa+gCV1PSTOX9DfVfGUbR/MEUpBhh0H2Q5Lq0KFn/beU+gR2ZH
cUzzXCSG/6E0+eXw2PLhA1XGt1ajrXYjQnZUjUMrgTZVly3z2yD3a+SgBIe52gdz
jq4+V1p7DYRT6Jb5uKQTuXAf9H/oZhIxYzUvAlxWfDE8NbCvWLuOtm7RjecNXeIF
hmKjXklb6dYzcJKJqWep7nsRxaOkeaCqyLPDjmqUyoQSOyaOEcXvvjb4XazAkMLN
dysSCQJmZendGFh0Cgzm9s0Sk4zgeI10FaOwvVfQDklouFm7X6YZBJlqy3E6YfUx
NK6IroPORImvoarMoIkr+sAiHLa8HjvHTK58Wa5i0RWus2JHGlprjfkhkk0lThoA
s15p7wWYH9YZbgkPu7PkKRIDtrbaE5yYdnPT3zpaknV+QepZqRyLlXeO3EeZ1edg
4bqwFWZ89gygPQ5PzTpViNj359QtWdJz7O7jxVyZcL19ki+5pcvPUGpx8wUVcQjo
XzykTk7s4SNUK9Vn9bLLpusYYs8RIx+DJpF9NnJlUJDggrWFwpAYWAX+oEqduuaN
Q3oAGb/a+MljWpL5ljgUJrNxNw7XjeNbcNQm3Dq2hG7Y4o8DZiRwkmFrv5nGoqHZ
jX/jvGu7Ds/+qkSOZfiIkfeGT88/AoZ7EvrfVZLMuZMi8swZWqAXjm9WLshY6U3p
UX+KkmKYZt7nIED4VjnMZFSzeF9wYVd9MOfzc8JJ/hQZmSTz0mqPetR0J4EWcdbj
CnG3VIlCVWtvgjq0acTonmggT7TJ00Vuh5ajvY8I/Co01KHyA/Eeywjgo2pqykLq
bdhPIs4zP9wtTp+kfZCD4cu0vKfbrS91+T2JgqePMNsw5yH8+V0S26Y/wu5OtLkm
4GlDKRaGmyu/pIMicmOiXLargglNfOTyuTc1FdSoNyH16KVBf2he1dlUcKWKYJg9
vJXw07beBzUP3UylaFOzby/YdDfsh16Xjhhn/YDDAH5XItKp0LPcTOZRgfSZl09D
qe7q/vo9LBP8y44i+1lahT8pmN5XhIWFutDRmGDoVmUnJ841/eGz9/zh+7QU5/k/
214R3zLbe1YEL8hOlIL66HvE50t3vrriWpwxguyEIEPgPNaTxeYdKg4QACsa8sk7
Cf4Xy77VM5jAf0cF8v623XGQB00P6ezAUB9X/J5EVHpL56kVDkCg2a2u3AFlafZk
E9+pFwU9BZiywS/fxPvLF12pgX2k4JYfmEJw5qtQcj4AYHKCJYUhfDMNQ9JY7SM0
SXQPKSiZClu7waM0Ebbout6hppNB6GelQoil2wpSuw2SYsf4BYASq5hySW/u2wSV
kex+7zHjcvvPLV/prvFr5fR6WRUiPWGQbUvtOuMY1mn0qy74FlYUMLClj9bxTHOW
gVeXQgpsg0rmxiaszcIJUHj05IV6aai7CxU6eLjpMyM6JWc9AGR1VRdcUXPCxidy
xAkAI/YfV9hZo9j48AW9lO9XMwanPxLathSUTJ4KcTpTHGhmnWfGV+NihHeYIEEe
5+bF1amk4LnV/OLF1Wj6IvhSLG6N9Zh38/kIWCvW8gtjDcjp+//K/a1gFZ4i8IeG
3GLu7KlqrkV4eNkV6QqlFNV9gwtWAsv+cgZuHvg33P4YoqTJFfFfJfBlf6d1b9KT
IdKwmOs7ifcdsqD5x1vJn6MqOOFT+l61WbdkZ+ZK1o7CCcPjr/iOHH71VjTXB62Q
y3xosGhIkfSnHIi4Vvu1SjB7S/SLz6E0Je2F2g8i1vqHd6fNYw5TRWHpLL3Pc4MC
zu+eGti3DQU5FkQNtosDkFMigY9gW2jvGPcXzkOWTxvlJM0H6kDnJvrZi5GIJhiA
uEvnZoEhw2o+h/ifx+9mWvbbwFEhZZKxe1OotcRHcpAQkxIJyek06mWlEH2e4krH
QXVYYkh7LsxFb1gLBE+Gqui1Y8B8X37/+lhOw9C19t4R+YKifAwda8eFSQJxWx+z
WDD8PTyDMJxIdnG/0ud4LLw/04+3H9zjWy9Wzii3zSin+FNa3n+ZY/k5gHsNZghT
sMhEdMLAlZVnVb39dWy0xcNsTAZ4Q8GTnknJ6NeiX5A0leV7YkDoR7TK16Brpejv
JqirY7/tBo1t19XzPzjMcj0w4gHIOHQwIlFnYzIlnStntuVKHU6TelmWzEWIvQqH
WO654P6b2mSVpWHhSqh1CZ8mlCAniR0WQtqcSRsYcWo6kbpGcX/6kVLD7gZ6snxP
QeAFmjgWpUB4tEOqeS3yytK5HpWEVsGOcT8koYtFymzr49qu6C6emcvOuFzknG+q
TEQzM+JR1ItEyLBqJX5N4BHtNE796kqKWNeSTDYqRpH4RjOLlaW4PxD7zJ0QAxyD
Sv+JbLBGlbx4Lf0oES+aBbUbUITDJEPqJ65mhoxv1upPJ6DLxt+DwNmMoYCjpCC7
wmh2pr3Ljn5PuBNKrZcBRT+mqOoVe0XAAXO19sske3I/dNj6FoIoN3qpdB1VydqH
sn7LesTrNzdOBLhYQ8/+BussGHnD4jDNtGxP0Ev2LTaT6uvy1FUYGqZ5+gB9JZdV
TENm5cLgh/3TDoK6EWSuFYBc7gZdEG+NZxKXXI7CR+Sp2uWofY2l6owzbk66544P
27hUyfT5MtJ3Ji8UA4/leBQv+dybEJ9XYfe9BmW/CdoypZAOwz88X9P764AzWeal
VmkguOH44JNBr27jaOkKVmeiQ9oJsDggF+iyGuT7et+KwziFQXR4nCORVKOdDzRK
LMTxf7GWoPXXhsLTTOTjtmVHZ6JYY+UuZHzOiQZ42yJvchUlxx2RfDrdpuPm0OLG
yJKy5t5jJ5A9kM/iwUqnivvAvPSY6S+SeziMvgF87XGrsAitt3PVM7Omg4pHilDQ
JqZ0nyP2+r6LVtqqQ6Sd1kSUWT10J+gGmxDhpn2zoI6wKBZhJVIMcBr7H3a7/fW4
CzIZwBAo0nZNir8VG7W7U3QA7Rjv3+IqMRFreHalLqSKv7Hbro1dLjaSN3zO5JV7
Bodoc44FpvkQwhrxjIzqPTHjrcNK0pegiygAIwhlN/SEj29tHBRDG26WCLM07WDx
eWYSx2wo+vSML6/rXgpz4UwKifT5antxDe84ET2u5Rb8N3yaqeCGVbQvTm6QkAl4
aRfS09h1FlXXjXLZNaDMvxI2GKgAi/4P+bz6AtKRl7kvUDLmoBpSgUgH5T4b9m/8
PG3Mx3LuUibI/0asf9DKAmx8RbsPltaGsb+tkSBacP5KvN55BblpwlC/hAcxbVU/
IRYjZbwAFWTDqVL2w1Q8ovp5SNuQ6pFtYVu0hEP2Ut6R3McEQhk6Ey8GGNtJ5fZk
MlexKvhtdcDhbgL+wE0peEaDb4TuIwOhsvq13M82oPLJ36wETn8Ggn0vJ87udm5R
WRkEE270ld47xNr1Dbed8xl/3penfrFzoQLcvvv2PcepEeyOsZfSJ2twenDNPSqm
s5Tzxh+8yupYZFKwYj13LR9XV+XhUf4fcMTkvJow40eVqOm2S7G6UQYnq7n0/7F+
Lpz4Q+JXvtuuaocC1ygLjhSmud4+pypzQF6ez5pMVuKZxNmh0i+d/ZUy+PQR35la
PDEOboM5yaG8XWOgXRgASigFVHCv3Q6RQ1ViYTkX/34XaolndHgcJ8wvcUGo0j1l
NepTYU8NIhGaJQ+GDSotbFmrwneiUiyC1fm7RozbSz4r5mcjliQRHknmeDfPZFVY
MVQxbTTNythv6Gb1qnk6HJo9J+W0S3pPUmxu0sqTcsws9B1RLJ4VWCiIvRsnZyzA
lMTwM64Ti6WCw7+7p5GloY38IIIqx5NRSVJQeyRE98voZP+WlMUvB9RPPGjNLVbv
QzivadRlj+OOpp3KyCvO9hXGfnEy3DVrwKvBJH1lRIRi5cYX34MVl/qC0II0uX3y
bql0Nqnu4WLhO36Kyu3xeA9sGaIF1M/FW93iCe2poO6IeK4GMBa/5mrpioBYZ57m
jr86xBPsZ3TLMx233/q1HB6iefyST44zshKunXgdoZsCOv8ke3lSi2P2brfp+5DE
DGN3novHc+YsrqMd4uLEPGvF6CNIGZ8TSb2nM4eqbMoHtneqJ/e3hIe9Py7OD5pY
BQzd7N2rLQf9/R5UYL11ZH6dDLQzXjoW0BCtmsCuKj7OrE8b5ek8H6EkOVgTfffN
2C9owVA+1efhqdQJRU3M9g0C1WdaLIdhw1/gxBj0CH1K2/ddWKT/Jfk8Aw14wMta
PToz9TF6hAreonmNabbgdgzgK7jqBgIOfW8hCuHA+KfoSsT+X7NLcHXZAwgGNpyj
lRowMJIiQQR6yhN/PWYX/YLTVNd6cvVRBFHuHqzFYuSctQmYnKgN5uatT1CC1CCo
72EmqUf4L+8RRisCGgO50rcYR6gZNd9kD9dNLhHDAcRv1q2Py0p6mlzWfBz8ywwg
gL8pTvVVy2/PSSqFjJBLEHbohJYQzI3N4/GiHaS2SodPlXRrQAKU/9pdpoTcyi/k
brC5/kSj6hTb4njyuct42Yd6HhBaJhIy5gt4yheLUVLEDu2IdK3Db3jkiXGGEUSD
Xzr70OtE0/grV7IK9wcf+9l5oqd7gVPnV7JfscvI9xatlXb6EaujmJYkuFMSA+DJ
HVRTj+IzrBVerA82si//Jdx0+adV0gXM2RDNIbUbLc3oiw40gvxWJizqyYGFVbZj
T2W2Tu9oFd+QLGhmcA7j4vLIcNFu4WgekA/p5BGe8QYUqoTNzLmTYVssPYKVKxRA
JW2TdIj9ukaOEc7YUWArbl+nscHZIMQogF7VxJ279uW6qYaWB62IkESb4BXkObSB
J099qrQy87GORqqTwhPdohlHzZMmTqFGUBZHYzy95rQyCAlY/UOAWEWRJz464zJ3
hlhowSZK7EQBa/B9/LmAmJ6p1a21tPkEjYgO4+SKIjXdTLosDGqHGJZ25KCDNDWB
p4FbTTJ7CiqxKtaDUNpJB0kCEPR3O1imGdcvqflgfonfrotqBw+74LoxSeBn1vuz
PtjO2La3e1/rnQiNsdHpYx/uacPpBSZXFrg9eEVi2uo/9QcA0AzEXp+RpD5Y5YML
AuDK+PLiG/HNyB345jhKP96N0JFBFLuDt7ngES/IYBtKTHakIter0J7Phi5iFjG7
CWYYl0oEgdHfMm6T2QD81TOBVGBi+hyjZ5/5oAB5GxOa0NgFPRAWsPL5YOp+pSsV
zFdJe6qz1vTRVU48BiePVxWilSOMKrIXB5/dCF/zv+j1BMJX0V41iF1UJOkzqozv
3WlwkhgJaca4zGIny3kXm1eb5x4LciKzUGlYylmsM3aTYloHP8ffFVaDjo/fjrFh
YmCXzQlTVe09v/RzDpITFe/wGWuKNvplhVssWu7ujGcXSh7evAXZ4IAZtGWgUH8B
n5a99DElSkaQqKK/wRfp8Bk8/wXvs6CiCq9pUvLPGY8L0D0DhXfDqpV8LukG/s74
QcrvxcZw/VqRaX5XkM8AZqKlVBhbYQq7kk93Zu93rOosxDniGNY50kGZ4+uhdxqZ
mH4PJZ808pRXrLnHAaOGUqOmiMUsU12z3OPfg6lPCvGmP904Bg4M/5KDxCDQMIJj
gEa0u3j16HPk47dYQkpmAjNfQ4q7J52doxqh8L5iZVavJzCG5b0w4a4ZS99ofXde
Xjuw9CLBnjh33NdLglaWJsEeRBURMVowiAS+eQbdNrtG5QsVABlKqeTJ7ALwuSEY
2rZ9wGNL641EnFYm+UygXVAQCQu6FQZ0Jlr8eLuUykGHoPaWqc6Yy+KbRee1ie7P
NL8dgpLJnHV7XvfEmqwFM67Y6hq7WfDL0anHRPBuk+bmoGvQ8ShsBWSf9YeKz5OY
/mKIX8c89rhYhF2gnq96ct7eVRzCTBJgkd72io7XlXw6R5nW1Eg8pu0P4xp0huIj
HlhcbjA3ous+DrwkrGSNqlm9XvvgDzosaoHwjbRSFK3Oi8gXw+adtLjV7e0WSA54
Kex8BAhtvwYhm7fvjQ7ALprKI4TJkizsuIhR+l5+aWktwh9ECTQ4UbA9C41wHBxp
riYEyN4rC2WRIMcAT/DrTFvCWF59SFWMm7otaJzhDqyQGy0eCtr8ANsWhI422BDK
jo2Pcq9I/3ozKRfHyDQkpFkVuTjeyybeT2zs2/LXA8R50Dk5AtNSr11MQG1tjktu
b7jB07HzKFxE15aaPLprlO3BXfRwg4vweN8WwkXTcdYee9ulq7jf9dXroc/kKwvP
8N8ep1VzVMPDoOfd7TcwzDbOFNqmQKOUXIgBEP6oZmWl00jYpWJm1PZUBOsx/G3R
M27cGsLGYjp2LDV4D6NFuUTfiVreUjEUSSMdYVbJCYWu6EIoN+Oq9mzcQirUPvct
ee1CjGFc41mCuF0FYav7x5MMCTHoT71jbj8jLXJJVh2LuWRnhWt4HvIFhAND/OC3
h5mmNBd6nl520TRkxn1XhoRjVfdJFNYZFCFPHBYlkP4fjy83mxHOLuw1ljQ4sWFl
RPtvsDvz/xtjWL5zQc8EdabN8c2R1G2T+YHL6TTserVOmDSZbSvlXo37HM1ScX5w
9SCy/qOBgJR9WNCBVw6zUL7Nizkna38FWVpMLFn13BZdXEIZjJiEbVGpoGODxI6i
i9UgJvvoH7UbVzmRuqzY7Gc3fPgHBUoWf3OVkh+egbKEa2hrdrto25In+EJyLrNA
LVmqPYRlD9jFt4Vsk+KaBoYG5ahvmI9GsURa1ydAv8E9GbO5/9NOhRRHopiaCcrD
euoRpnhiiMT/AqKFCGJiQM8m6t+3qcyHiVEEVlV7Ujs0E4B6Aqb0wl4yr+WuPwWY
BJrbgwKWb7SmEgZhTPq89nBhpnNsYNT9NgyiGCwpf51ugrUos42vEDuJwoHwITtD
CemhcugN+tTlY8gUdxYmjmo05q7U14ZEKczWFIss7q7TPqskbc3/+hjC7XoNjZjF
ERR8jNsbdXemxer6zjsAmvhK7mUzMsGwSVO00JwiT367ioBMSJ+YrrLl1nARvnb7
xgwmy3MBlmCXnC4kuMANOP1ZAmMDBEHybtzSf/VVvu6myQ6SRwTWJMNmfcPQWnNG
DSP/gs6j8V5Dp9eR/upb0DDQ7JEIhU0rdsgamUdVncQ8Lw6jUOfkarntW45bRviu
RPzFWzsOkrL66OEjNUK2GegWRmScM0X7MyBGyBNDb6OygLvHa5sWSXZLBIk4vuVo
Aa43SifHdnt0wThKjeK2W+AWK/t2pgYK7k2OUSos3dwi69R6ThvtQXdYSW0of7jm
ISgDQVEpTEzgJB+uA1aXJdvUtLEzIBN5oTKM7i/KoVezYKNS7S+UojNxaxLO6epX
Wc+9xJQXLMYAnzn0/vw5ZZ/QWhMhhTFU72x29JWX/DZJ0FXcKRi0VIcIwKLro5DN
PkJap4nCiENIsG2MQI1Y6gf1faUL7izTpr+jy0onrp7IJGkU3s8RXzoC2pQLcYQD
AKmKDhKq5dXg7nneAmXQU/5t7OrL3/7mVDoeKWTU+rwXFI3ZwVg2jKj9rhFfLy0r
eWTiFLslpHZP2KfFKvXnToDXVF7CSp3PEahHGs3Fb8FrFjYcaHY88qEbkJcqV2GP
5PyvjIIh73haR/+tV75kSZFLd2FEwe71SzccDNOHlj9SiS3F7mgReCgrxnOpJ7r6
jlNHHh392ctwwJfSkolVmZFm7TuE7/SKfkuEi+8pz/CLHwDMWH0QltopNHV4IMW+
PPeR5ijsdrqoP3xYagifM5+ccDketIcP+QAq7UFe4uBM5VdYFXEOdnpqU7xPEr5D
LlGGnV5su/fisZWXynrDbqW9Z73CepbwcZWnGQRu5zuZoTIXjhahVxzCRVmVbaAf
tAT0SFvoOjwK0iNwm5Y4MCRjXYyBTp2Dqh6lc5daROY9LRCU+pKRlZMFo1hUkfBs
ekbp9a7EneRcOx16xDkmrQFzJAiJwD6teRIgWrgfn+ucSQON6B4hkzAP8WbryNEI
NPJMQEIpBkjGhOx62t7rTnIAPYc8Gf0nRRLIQM7XCRbnZgwr9i1QhGuZmOb6u+6S
5uS3ghxYr4aLMCLdXnugWQlla/3afuXTmsPyledUVLp8PLd1iGYqIX0thkbqB9Cs
7zn4ifrm9GOWou/dos3TUTO+va/DMuKLfdx1ZUp+/jAgVGnDm1qhW5EImzIykUsV
YA/kxUnPEdcoCM5r7h1Ytd0PglM4ctKXKq/3jBHpK4IKqJba27XkNff2s47kqAUd
xfDnx5cZQDD5eU5kTbrsYhaQ0QAWzRac0yS+Hd3Qcst7rwA1pQ8JOGTyAnvrJXhS
G7qopBg1Z8UHDlVVst/MPGlt0zmOlp8NVi8uL2wE+NK8xMjpzRCBhjT4Z/6D4BcI
rxqcljWVNSO+/lVTLcAMm1m9JSHp2wEd5V80YF9QcFH1hZCwc1baU3vzpWwYv/BC
/UJDa0Q9tsn+gn2rVKFAoQd5qCEg5jPj7nCjtCEP6pE0cckVsnRNhmMD/twG2Fpq
61snO/kUMk/NIFUQZL6JE0Ud5IGtWAxcknuNMAqcqunf2whWsCy5KsqyothvC+cA
oRMR8qjvcV9MbTY7FhsbTTN8dv489lh43roSaTakFCSwwv/Cdm5XSEpo4BUdvd2M
nCwQSPLZliWB/4h2lDcNPcS6Bk8DLaGsDT4FqCFiDPy54DVXyvnlsDbghw3epNcV
oq8+K2eB/PtbD9/KUoVdinFMVrHDTGkY8NNjn2JvpoyDMC5ILHWH27Mhv8YVJpI4
LvpvuMKO2JqPGEcnj+HfMziKliWdx6dfZ06Iu9rDyfpQ1nuaBhC17FTLRiyOjPBH
4lCDaMFJC4fi5IwPySYUd1sr0g7fuv/39i94igvgOaanlSnPhztRoHiRKbgIo81J
x1wn5xt0enZY3PQ0Tgr4Sfr8aFPmBmF9MZ462fmm+SPq56wV+J0F2/CEDfQN8/ub
4kVb8VI4vSO7CR/7KEi80w2F2MEi3SocXWdpdKUtqf7mSRSem+KOVZ8kNo3S1vDT
MOimMQB8fm0PBMqZiIT+/Q4q4S8K4uXXwVPfp+DhSsPIkWRkfP4myujo3bdGFKHc
m3a8tMrMt5aemz5i2qxQxG1phSJtUYjctP4y40Ag+8kmQYIsK/qXZm3WuKEq8eFs
FI2DGCNCWGtddybIPlhQUWmEwqBOLb5ohYjNuPBqj7smrjygYZJslfkUzfmFBU5N
O1rQ1TJ2OG/oqFCIZHO0c3AnCfNfUoTeF//GpWIbtkbiK1hBhrku7+P+HXrRH+8L
GVTRbD0hH6qErjaYD2hXf09RmKmTKSQFtUAx438uvxfOJ1EjVJQHkPvlslvMZwzi
0/C1PqFzKN6N3/TZuNKEvhQI8qKMNI8XQ7tVPca4jfaIRLhNEXXEm6AikFZ6oasU
UQW5OwczT7NVfdubztI1Df9IeKh6aXzjn7GEWEJZCLvBGfpE1N+LP1IhASuBL1QI
0iakpR74IaTBLKhHw14w3YO6HBKJV93ISn/7+Fih0K3kbFuLGmMpAdt9ESl9ntuB
qJzCfkhrmfcalR271B16hIDXKHtVLdsol0INZCMPBX9/Zd5cnNtoKDy0KtXUkToK
+ub2eT9WVYp2FzGg1Ggpq7lu0RImfu1iy5Y604zA4HpMt9DjUSaTkM9kBCyhdZ2Z
frgzU0wci8+p76OsZSSASkXXPu9JtubWumLHJAQqxYoHzlJMpwtVTTlAUPO8Rpl2
sWtDw5QK2lW9WpHNoJ9wQkH04Trf1gWt+9+qz7lnemf5ZhaLrP0mCIrPZWfZkniC
BfgEGuOc7Nz/Jj6BzrvRST3yPhh4xUW1yVkfMMkP8j2FkCONMePiaq25omgvT9Bt
yarFpq5EsVuuZ15msCWazkPJkLs+Bbye+BxdMB4EZU8TfDirlPpkHsdVgpK0pMYK
amfl7LU3fqEmLfsrLA5zwdfNJJ0jq8KAQR1i+73So2COGfkBvp6kTa+DadRtZ7DX
esCWlV2W0aX2aTAigVZWieTbivUckCz5Bo+Gtuoui2UTW9TZu2i/3+2k0xFvq83x
ZCZ3VTj7+SnMWlKqOfuRk+YDYtD2s4maqZN8mpPRBJ+o+nTJn5XGTNLDdl9mO6nc
8kaigVKB2m+Pu6CbWXVyGBibCuN6dzTelzc2sJZyDTWsFcWIjMNmR3bG58jDLdKz
hB5wOXk2bSd1IfknnYRxh3U+qbvjCUSdaYHHvjstkP2opdMCgyi7jntMmJuwsBJD
Deq0fIwyiJ1O2WeiApruorIIg0HOq5lwd6LNzBcFQRhqWH3I2KFFxYNmwQGDcvWB
8ZykU4P5iONLYo7wwOmHmekYVsVKVecWv6Uflq9dup7gmKiSM40yyViyR1NKW6It
HycOUYAou6RegHy+apZ8oju3AyfsdwExj00yIuzWVwsa4WpSiChSLY6Bb20yWyky
JZhdPpaMKXJtnCpisdz43pMKpZOurHDUIYrTAAPEqsr5cQTmEpeYk2PYxJIUpVed
/S7ik0S5ZLvPuNfXbvzfCqvzJZVYv8rw+xpD53E2C6co3V2FOhSAVFQcWnSPbsBb
YcvsOHlOEZ6DBmh3kIZz2HzkizF+x+AK4eeUNW7B3XkLx9lpTdTTsQXz2FlaBQJc
HLQ6oEMAibd+sa7gW5hA+pF73WJyZg+RhaGXuiLKzSQyniTkamMPTgCNsI/KzrCe
BXD3b9yo9f/UMSTvqFI919dLBIDbDMl0jzGe8UC7eKz9mtC6Zmoi9kdXZeKs6hdF
E/3rHf99RZuO97RyBnepoZgCls7sCxd7uz9lSYHGJ+dK15YxPIvRHQSuYSY5RoXB
Lxp6TQO4DSrbEuqBXnA+ubrK1hvOzZsvfwWmyLhAWQMyey8siIFGrg9sQuVPdr7y
nojlXuANDR3z3JEpAd+gGsNQebgkaTlPhPkpvS3hKdxOSOJMrKbBRqrvuxRWdJvN
itVNJgQzr3/QTjs6XJXuCkGQHWJ0Yr9mM2exh9zh+qMZCc5EN1ZUZRo349r1YqCc
gm0tZefeI1iFvrOVc8iwQtGDJgI1FioCpphAE5Iij31Wxj87qugcmdbOqFwM8kp5
WhP8RzfOIzoiH5DCVg6l5uX6iOdVys4mKsAoGeVTsazVY2zqF4T2cb/d5EpqNPqn
2jp03QDpYjbfF1A8t0ZeZ1Avq3XFBuKJJHPIr1/dzWkcC+dtaZN0XO5vTdcjdXVQ
t6fUs/RiProkb0zFxPvyC0IVFSKnKEdrcrpvewsB9N7l2KlmZejbghEHIpZA3tp0
j4VpcdsEIPXGe5UymYEXZhzssw/srFVFf1GBzfOT0gGRE26JUnXxP5kDwhT9rZq1
/Dtb1miNPwg2+JL36CTEdKyopJt2I4vBnI01hpPfq0r7mVR19uIXg2lx4Mf9Hvot
WueAawaTyQEKqlrMlx5tjDEn30UsBurRyxQihK0KI6obEeUQwCaVtFxQtA9uiQd8
+2Q8EHmpp//R2kIihcuhobu9/zbJS2lIrn41tfh3irzO9bmbYxoRc0fuWo4pxPHQ
dLXd4B/PPxGnprJXVhi1/0VH1N91gINs1JkxOt9Vy67gUi1AdevDhBMz6hszsDMG
4qbAp9wsZoe2+WovHqSBdtsfG7hqRykLZXXSM8tznaiEYSGlkqveugQg8FBu2BK4
XBPE+Bx9uy2aLc9aaecRLtxOQsVRCpMD8YdbR386+zcQagMaTQcv5AAkKlNnUHTw
VRzoXNoY1+uUaz6SuqHR5dklIOqe4ELG896TeXQRLgow79mhA/nWhMS14X19Jal4
OzVr3ONBF03utisRSNSgrKwVVveo5O/GAHk2JROShZkcCGmBE7Df5zTf/1WIDCCU
fIMbQkG/ouCXubxAn/DJTF9Yltv6UL+TZviR34siDpgvCMJ1FLRMFjTgWXoN4dca
nZukNeSsPEMO+DdiI2WMPb3vW+pivWrp1pMYtC6FnGZiWIQnknUt2bgNH560HkzW
oUzeR/vd8x2WoBva3jDqdv2PEucpOFeSjSZNH5P8Kb+/xE51cbgVGZzoF+TgCLFk
vOl5zRwP9J4BXHtqua3Pw+wxQYqB4R+sSkdfc0zSrKb8lSSYz0ak8Eoxr54ko5Jy
3kl8Qjd03VqXmPP6ZqjjadVymNo9jOxjQTpQQBkxCynIiQUD30kY9ev2IfegQSZA
x59H971IG6/3o/hDSJBv1Aj468iijLASMfYupYS3CnWQDIGHSR+06iPUwYEbx65z
YfPjaQmomRCp6NgNAuJ7EgwY1nOWNg9a2D4d0gO53ebQ68ia8OGtvU9qe/EHJz88
GiWuBdaN7S3q9au1u4QybfxoVgY2uOQaeDhTVFqiCI+Kg7OXDFTfoX8ACOJRnH7G
DnZbosi8RWxXpivzajwA3tThLUfNMgFn/lsaatbMi9lasPW50MZVm0nGnLq7Hxt2
yZ1WdO6Fi6X/NsCXyM1wZAx/EKvRubcDAG0wxrOQFOVGMbDvVb3Lokj4voII0S1a
GAqJEkknzRcltWyYPU//V9VX3dk/2JcDMw8Jbs6KZ+shDAEjnpuhnf1bVsQ7E//o
GL0IIs68gBivrCM5jSyREuPV3CckXk67PliiJal5t8oL2PVRum6fyNG9M1jxWouZ
Fu+PaW1qLFbdMnto3pDfMeaSbcdb6coQHFGPypf/q3grmcoP28Dxf1h/I7KLErDW
Q3AAHK6CSL90akpxEnMrX8vfQxFKzqk9C7se07owp6EeUpVVgfp5ovlBYQECz3jZ
XMqxlOLzXU8MeaGerALu0x0aDMdAvIL/P6dr+o0kqKTEoP9cWDWOKZFaGATBGFGO
uIrSpHLzUSrJlOakLbH8hRflEm+XeePhnWnn+/XQlMzkzBB2fuXrI8EU17jPmzbf
8olkHqXxzMTUlxrsNXiafr9pi6lfuo5/YHxrruUMs80Ol7MT8vgP6hfIYoHISKcb
QyrHBBBCVETdG7hGW2Co0iPqkfcng3ImLCMhmCukTX3MJG4dY0fA3V8jm6Xfk9pY
JVsl5rjqip43EIcZ3/bmLZ5+FKKNreSMu4JkfwgDcgusFV4tx7ei3twJVew8J13K
ouiFS87Hmjb0KZpNlONyCWMEv32S0b90laBEdnisLit8htZbFEjtxlIZg1Ofn2TD
df2bxkyAi0RaCcdvmYysOMrXrZGav1R3tdNdOyIZSJyDjFR8RVXUPGYznscGU66e
SZOah0BnIpyK3XS1qN8GJXPyFCAH60M0zKAi7DMCh1EzEqRqc1vR1u5DXKrrlffS
VHq6dR+yiD6mgFWuKqde1SXq+4t1SWHwVJKX8Y+habYTjVbEdnXI1U5YCN4FMUwQ
k0+U4WpsztkMigDsbFq2loazpuzg5B5wCRneZLU+eTzlVJRJtSbPQ/duSwiou/Lh
ORfhb6ri54+EcLyAF0n20IP9GfPflWOqBGdrBjdlDnmOHJ8MZuxBW7kRkSBdBHWM
BJ+SS1ozaT/KyfAVl3D1OGEhbpBqmVms4zfGzAsenQk0JhuJAkrcOSGYBuJ0LOSR
oDbFDKohGmhKAKxrsu78wprRxDBrEQKl7lmlASZ9p/FAYg5ieS3IVXHEFDSTMDtl
uY/k91isTDhtKrAo4kxXEanjO7CJdiuaPiFlcUARHU9Qm3xkk38DIAx3FNGAezB1
cB5quJgq/4A/SNCb2fG39EzPscLXxhkW3BvZMF+R8EXLQYziHRm89FJtZ4j3s8Rq
xpdn2Cx0ni4YrjQqww+T95QMyYGh1IrvI7P9l5dJcArF4tvIYgy4fwuolsto5UGV
VFMojiG2X3coubayXh8EXRywmVJ9aT4g6ICKWZ/PZgrLigoTXYYiKWZ0GUufq+Mk
MClB0oXORptVLP6RvCHrCnjk1JUALZGmmxjqXHKU+Py2WM4tvlCiTSit20UueToL
/Ar+qdYDn7rmYf6yTniOwEzSNNUzyMBneO1sYyOr0X6rSAAdoWmP/UHKYGrKp0/U
JXa/AoBwOP62V2inKiERKt6jRif9L5Kf0+MY199Ia8vMIMdTEsRyN8719QEUYO8d
4UjWObYmAtDQjComnPL1RcKldJVtU4pGJHkFGd4c5MZFSqbYWA06+W/QmFO2RlVk
c89SlgUMNMo7bNne+x4O/aCObwYskC0HgihxzLr0/N1G/nNCM3MiKM3cJgDCQUr5
cnDVd+q1Q+lsuh92bdxvW5sjSe6f8497Na1M3Y8mfqyqDdnS5KlXhTX4Zgnyb6Fc
Mi5oJwoGkZIO79jUGm4cDXaUT1lnExgnE5DN8UrsbbEEWyMqShGwnTwU8wDwk6KD
+k178kmraI+BfhgRa2kNh8x+zxqa0mq7uWf3aA0PSu5bBtAxYX4pGoFje0ogbwbf
LnMvnTiSF9VadCxAfoMpvLJb1i9qB7viiUqEahwrYJBHrazf+/KeIT2JXfD6WYQI
/e53dfEDVlUIIwBjASufY/tjCOCCdCW2z/xOe56OW3FPHomM7qaBZbX9syUsX/mr
QbjjTtuRHsaybfoV7iYGDkLdy+xSTmit7n1eGiZ8DHnILn1eICadW7uB7Jpb+Q8s
ky2zGPAwCl/g0I3tzgZhnZFHKTJTdO8ZA/xzGUfZuI/xUHbdNGl9CkfK/e+6O0RN
pxraRZNvTJfwUGMzM68WFDB5TglnilTwkZnZH9KiGpoDXYvuHC0JVfvp9cvzk4zx
THGXPzUw3keYblThVDbnZDz4wgtGqWPo1q1SmhiaazRe14xDayVJNZ5+IrImSzW5
D2FNQSqqnWXaFkhbb6+8oMQRaxaIY8RqDtT7QZqOMA7uoEqsJXvdmKI6HUEu775z
D8htWE9W19zu1S56uDv3MM2egGocLLAsFPrpbRyPLDoNVnUGqSao6gO3LEMEcsaL
qhGZBgqCH5LFRzlbDwxIBnYpm1NAxQ375lU2DQ2ctDHAZi4CNdOqaS3u7OH+z3az
RCQ1beodRQrMD0RVGxp6B6LXaeIMzdcoMABk7vUZ0xE/GF850iNcGnsDPUG24ega
rc/MeVNiY/bsx4ujHh9o2ydRdMfzBKghkSr9lM61IjBjTQbA2BzGEVUCXeluoG3I
O/ZgNjz6JBPXUDtCd9M+4eAXQgu3jPNqmDNlBGK1B+ZcCrA0OLcK6J6PqrbrWJTX
yTVQTKy48ys0iwVPA0XMeu8I4wY6wn59Ccgvny/XM/VtnD1NKoOfTfIql3HgRarQ
bFtsxF06+5Ciub2L+tAArszaoQZFwZNadhuFeGEG8eETN5RN1Z6mjqhWRvYVYaYH
0qt9U5O930BS6M+Jn+emYXiYfaGY8V4EYpUGOrStUQQm2Fo37IgyDRAhg7nVi8ht
A7ZCIFUCLSBTL36xgWaHHENKrySLVBeOpP3xeLl+IPM3wawpvt7ZI8KYmzyc/+8F
tnT1xapqUl+znsh7NPZb+Dv5djaoOFf+Q4fFHpP8CYvxOpNaz+4bjTdY8dBkAj0r
560miLK7G6zdHaWhFSIY4OswGDm7WsL4b24oWz6UOUdj0Cm6nQdNX3KQCOYHXQlS
4VUbU+hsW78vOg9qJ3LU9iSaPBwDC/hSiuTBw8p1/d5wBSvnAkME3M627tAqCwLZ
jb94GIl+CxqQriW3hRJR6EkQgPDrTgeE8ljS84FFysJNs3++G7vhINbuph+L7Grb
TitpWZ8jBr/7g+rDwXg7OlwPlld4LbhYjdqJnfNcYyWJFSzp/pWny5zrcjq4kneP
N9VMWioqjBUIkVYkJJ7VDBNrYMx18f1upDWupoYmbV3V1Dxkch+MFfupRmyVmBAJ
NSs3WxcROaTzHbW0YoPeyNZ2QEhvKDEWchv4/zUjUWQSxUh7iF/FYx4WKwjAC2Ln
VB9yPYCp3hS7y9ZjiDeRiygul2BUnXmWo7UDI0532DOGZaQr8rhszMzUcDV+BW6X
ZLl3yWPMeiHn4f5HNroNvzTV1baIqs9a2xecWoC2S4zcI3VFznZNyJpkrCtCxIfH
xmQES6ZUmKjBK0MrLDZBYedvaQTZogzCDkOGEz2e7u1cf3IG7PtRrvykvXe0BIIA
8JFzCNvThbcYEG/211fUsepLuCKg/jKVKdil02eqXcOfc/k2UrZb5nNHOqlwyyCV
2AqYWjRjehFPBaVGAHhpHBBiX0Eprw9mHsO2ioneV+CTrpdtCgf5HyEhXYVRzi1J
QxT3UC6CEu1V3UAjo2j78j5BOs80SChBr8Ql92VHGTTDFeW7skciH1d7DrfL2qHb
rt7QKQ/mDMjTjgif+mTJr6A+q82j570uD6qMoVxkAHjcscpOE0e2Zq3ITfQFOf0F
kzhtMO+h91CtVd+PhD6Tyo8yEbQEOws5JlfTHpss5CvTBCbLGJrPwRO7xSCpVgq1
OahyrXXtSYHe7m4sU7akmHzvugxRXOXqqadkpHSyG22QkUdcH3F+VI8fPEIMSP49
3AhWX+Y1XP4CTcEVVA47SpJLrzZU5i/sMEA9CdM1gFOBEQulE4R1uYW9v8jQPyL4
sEdlDl9xzGt7zlhOy88SNdPJYkh1eHrmY/62sxn+drVEftKfsU6mKB5HZtblaCw6
uBi7VQbr1DGrJuAAGrUMYghiEP9+XKR3j/QwpiBh2Da/9ACUU7TTnyXQGzvKSaaM
XfwDJsnpT0F5AIkKQYhc7R97IB5nzDl//xjyUomQs0gtR8evhXKzWS3/Q8gZAtzv
T2Uc41I/yZ0qQkrKsIwmV6aofeeFG2TB+ggZhSWz0YKE9L00N851tQ9/3IofYHPL
PTZh0/f6geCWEbwPODJdCTcBmc/7XhqBTe1yAspP9cd3eRcvj6fja4O9zabM2DVX
fzg2XO0NJrkOHIisRaVDameYWvwGZ9Qz2KDEijDF3JWKDjMD+/hmMzQcaqiPsIkd
MsjC0byBFw9PTTHfvj4L3yDeIMJbTZ3OxZGk/UpKhfaJSAFA7cO5naWnprupehKb
ahAvV1nblvvLmXdWmM5O778uFl9OT4uzaHsj51nheEVOy757zF1dyEHLVQHwctwe
IF4GM7QCXJ46QLmHv9hRCDalub8wzRW0EPj0aHNyPUAvGNqIGelFzR64oJt698GT
LGcLlf5h2JLjuQ4AyukQ+WW9vOeCec/CaBrjzXYLHit6MbiOYNOgKWN80Yg3BgPF
XwIfJopJW3P8gYOz1Tmdn1KaO9of6hHE7knpNTPBPbRyX49swDhIV8u7jSdIfE3H
X2NsyCf4JaEWwwY+jniweI6oKNwPHoP9i1R6G4KPOO8xGHHxtsNIGhUj/gbxzxex
6lsy3HjHAMGIT2bJtVgKFnJPg0LU0sBkOdanJja2SbNu3fipsi57k2gjDJ3O3xmr
VcwPF9CBc/Ax5eKwEYT2Ce2omuqRMJfOahubtw801xG59I4Zi//ea9+W82IpEj2w
4YDYIzRhCmnD+yv8V8+uXtXXyjEbVl2CJZdU80OqAksEFYosYVlFXQ/O2Nt3bXAM
sMQhItG5wwUbAsfgtX0UdDGv519kDb99NZ94Tt93ZBEbCbFbm27jyAndlNFPcEw0
U7DLKmMK0cnrTpcW+/PbhRiDi+rOduC1tAaPaNR/3RHeTOndO+kT6zQGw46h7ail
3ecqLyRa34WRJ5MBHkrfr4DdgZMQSuNNOI3+pL6AhMxuSYni5dgTahhrOuD7Fj/i
25+jQId1/oimBnWqQeYG8pUqTBysMleM+9+8BplLMStJpPCQOaD3dL2cm1C9yd71
XfCqIHXg3eqA7GNsXGOaW45Ccx6qKFHOuRkltczoS2WqVBHQB4K/uvGm0VAs5fdT
utNVT78xDNMsV0NfMPQ4bZwGk57H09uM6Ykaj/vPSe4VzVoVDMULnGl9YOoIBZXR
BMqHZKq0nD9vpwQSQ5q94canjhuAVKNii8asX5+1HqNEp+fd1kWcR1plc05nYdTk
XCpVah/F4EEoXlpmvJvCoZ2eIyKMB4sX+cpLmV14EJ3HYF3Q664H3S6ptHa9ztHf
DAm827mop6Ngbq3LM11Y7Z7YJ7hpZdPGaODEeVROIxzceeCU5zvRItnKhf4HgUbd
xdXaN1xv5mEyymLm2VcVWzKB2x8HukculYBsbogqgprIIqMUvFBJos3KmYiYWL2j
9GuHC9PReee+mMc7vQRAOPSg+jJ5/d6jpesTu9NQl3MIO83QYWyJxQzbFSlHV+2O
xortrh9COBbVktqQqCdITjmkMg7u3OH8JWt8kHTwYI93U3ePVsd2qEy9WYkVQ2ST
MkOV80//zN+350mxtDzIjQpXPF6xVtBJQ8SkTkodOfeU7a8W4Mszt7gq/cuMNQoS
uyM0gphFbbcQ+Z1lRGb2G5PNpOVVYUMZsC9vljLP/g9p9CJ8rBk3vaSZZY4/k7Rl
OP994pgZo8E3lVZjeyFRomLf07mOZGdT5h1DkYOGeJOvW+tB1BzGfJ13Aj93gIot
SqdcIJa++sBY650uhEAm0p7puSEM+m/33QFY7mQPSYO64Nhh602Y1ZqVzOpgzzP7
r4pCPqFOAEerJmPxcrPi3v/qTUtfEeoNJIOOaWmVekRrXB4yX3JTWS83r61Okwyk
OSMPlZ+h3z9rG9pbhMhO+4MhwpaPOVhagHaAGSEgq2odIv27/LSv8qbzY80KvY/Q
2XZ85+IJ50a8GB1Ku6HdU6JJEiw7EO1fNvXZSQ+IBEN7EuTu+curXBh5H3FrT79O
dhfxLplENODZNiroKsZMmsRUzB9Lf65i2BdkL+gFDa5oYhNJ/URXNJ5fIz0RVDiQ
A9dsf6MTgAiV/3W+mDwxnkDpnkj0oVYNiEUyVSiFGgFB0wmXzKrAsShC1ZpLVNKT
81A9Jp3MrWuTTOJCGXX7Q0fTRCLBmTpMA3r8DDP1N5UlIcR4nMFETwoMonKYYLTu
+Nx92BF1WB5U5Bj8DiB5j2/IMmbFUkwoOmJxYeZnWUrmGM4B7Xlznt+amz0sLPVW
Q+ziXVSqv+Hp2O7EB9kVuyPG4mzCSfiFSXYGzEHd5HZEgYEysgDEUeSBDe+9ANUt
qsqjee+pL98TdjVUi4mMqu8+zDNc6uinGc5GohyD3j9uZydSBln02XpE5n4h2w02
FVTSlg1ZEYVVQnqf+tlrXtlMDrsJvUMeOxV0r+z92mPfQu8balqvfKKSUaBKv2HE
npg3xLiag2+xmuxdF2PGzu8RAeVJTVqAItOhu7YDCdXHhPtHTqajxWWMxY/4H6ck
Owrq0ITbS/cuaIJNx8gFVdgy7U3PHi72Njlsjcl/PJBTqIV+lF2qwhVljhVt4xF5
JI8zeNPFTQ/UG92gGjVttZmN1dZlYJnZL07Hxzb3GbLfqyfcJPLlfCXqopXBw5Oi
xHJQVrLtFIdWJ+bOuw9pbLmyp2LKD09Qz6bJnbOlrOvRKYKdwT7Oo7piLSwE2w2L
nhKtQtCShvo1mWtJ4uEJJjfhH7RCKLxw4ub/23i3Ht6I/oJExor06iiFFIGadzAR
eTqauENq9JFpexjgT19fjIUGWltFHMNnIH6rmApFBk7etUitiYQOpmEbZgxMRRiu
UXBmFNobEZsp48kg2KIKyRQhps5hwiM5bbiv8XvAIiAQ55pUNHcB3v2iTjjj+fog
VBIzs+kTeKa9yW9r+ok3vHuVYc5L9FRwSFzvI+KVe131JsBYEOGy70Gm6Wph+8cT
YVLeltoJfCyvb2OGvsAw7nStIuhi2lsmKf2CHYzL4blDJCf404BH7rx45aW69WKz
rNlV0+5WzGYLWU5pHOabEHZSsVkGNpr3wKYOeIvEJor08eettgMhL5GwbLDT7TBB
yzbaVycCVdvZ/YpqQbJ9tT20Jq5jjCwIh0u7X9xuQG7LfagBJYUmFbXFOwmasUCZ
giSMuYU39CepoyPlhwostDajhUmPebsXtkMTkM8HJnskUQBwhJ4KWILkYb6nKjRV
EcbU5QplGS8eWB3VJrtDUPZEUXHtoMiH1tUDOeu3v82pimnX/xo4QXAHLCr2HVOI
+03KMMIuTRD1yZPf9MOkWckBR9Kebs+FmNCbMgcZ1gUpA0kqzq4PFijH74VUKoI8
oNnzsPWsSsS2FemZXEuTJOkxrGMXcgcPQoRCVNipwuVuz/ORagjS0S2lFwFgfzCe
XVVGf8hC56TvRni3R0LteB98s/sKharHiv/3cxWvlO6p9sgoaZ8TVtQ3mFWPrGCU
oaGTdo21NFTsx9J51X3VhgPEznMQChKSludvzoruVpCtd03/bWEaUgpmMeXlt39X
u+FVZTSM/7GJAT7I6x6+Rarn2ArLagtfUCz3CTvqAIdRfQtjr46j/+jeDJITO4m4
Uf+AW8NNKDvrozMMI4YJGlWUPCXNCh6yGG09ojKeGRPiSYFvzCYU8BOC+9pQugCF
P3nryWU8OuOpslS423fGTCBypizUyiORL5J7Rg69T8VtEpjVIlxRJq+y1F1huJmo
zU7FLq/rQLw9fuKkKogyONs1qB10leIqF0SrR4rU/54zdafJ5OLezsTC4fb25sH+
owwHha0sjfpcFiDARn/dm24y1kBpmZNkBtVRvRYyo9um/bj2vYuUqobyFwgmwZNv
m8zlANyncGi87yDA+n58OBGLyzhm04ESsrSBEprpzLVo0/irHvhSXbxxf+qgBhRe
jwb8FVQvCekHJD5CpqHSDTyBYLyGyinj2JvvloYsvYSb+U0PP/QcQbOO6d9Y/Nkr
/o/bLuAOhc4Y+Gks4VXhOtTWOFnRPK2EnV+CVLw+MvcXyIocAshDlRIdSKMqt054
kpJKdW4snZ1Tg//KnQiKAiScmM6viNW0RunCWDhfyYMlQlAi004b8g93uOO16IQ1
pVWakQ27V2wVRgzSWCyBLjF++TxfI+UwdKevOCApJ3UGL2qpJNCerWZFIPtpFA0f
WSRkQNS4pwuzbgGq7eiBZcVbrdJccz9ErJJ876bLAT4rjYn0HE39ZXS+lLytP+tH
I95s/CEo7xTIxKOJ2Tfcrx1OCEcEIpYo7kstlm2kKqQwYeIMs0K9+V4oXTl2uzfG
4ekZgR9sFaRjSJ4O5/L0pDR+kK+1PpcBmWXNjxy5UGLUcgmRAemuamAbnE/aecx2
opCNCwpwpjJNXfZorhNkAuwoW7Q4QUKuc1jUlrNqLqh1D852UjkBYX7TO//nuKwh
ESoKSbRxjmSZvC7aeaMHFHbkaqSc+Tcyy3uaAP1eLpdkXI0iJE3XOcMIcHm8XyiW
eCQdC9L7nYMmlwYfBjSwhAMmD85miH11YGbqkchaf8BuWp/8vJuwfVlsrhqFrAr/
10n/x1WLO5l933akJu0jkLx5PPoknyCSMp7bzNcaZj87fezgeQ6ci7Xn94XUA8ce
1jfizCT8ApZ3dVUiBSZ5uCbj0geCRFOxyX78BmyH8apQ5P98M1h+Q0ciAUNSqeQN
xeOJvxjTxYCVmlvHuU2kx6bLmlKYBIrErZYx3cK/FnXLigDwPZq+Y/l/9Wn4NQuO
FXValJmNux/6WcX/6OJ+HWBD4cKdUwBw23Bp1ZmzICKENxlj/kwV+azXtmcK9JUm
r2oqK0h2uhY3SucRRTuCzJvLVcrQ7/lQLBODzxjxgckjS60LvevrRz61NZXIYh2H
7e9vaYa3O1kGTRKz+iwWOsxlKDHBrjYfqv/8phdH9GgNSqr48fLaghkhPb75W0QV
YRJj1elUL2WxuQ5l05pwnjn3M9PyFaySl1GzgnYDCWQeJ+pzEm8xFlVI3d3GjrtQ
SXuzVDZYqrQP43upGzS17eKM9qFhjDEql47lduG6+BXFNV2c/BYtA8F0jKMuct1D
kzAJp6A7lnDIw7OrBZqWYf/PQojlnqsPcyujC5fsneMlx9nclIxwPaeIzYLGjzap
9pDPSri9yjJ2DQTZh+DosMMTRaarqnSbzIAGSU9tt979xwoi27+EBpKDN/RgU2Hd
tPquIx9ejEvKxj9RTkzYnj899GpMJjVuZ9V03H+do7MUH4t5UNSy3XSDQ3CX4e/m
hMKgR0lEm6k3f6WW2ipzkljFM+x35X6MJ5BGWqMkxBvObpfIGTG/c0tLZRW0QZxU
dyXjbXX4IF/pJ9gA/o6S5eb8dxM7hyB0UGCHvbZIzoqenBYagm2OzEmK0528i4Hc
I+dGWn+qfQO18qNKxpp905twtcJNj/FNvKfGfrvn/t9r6AZGpHwm11R++qGFEIT4
7Ka5meAu9bui0ZLpjOloema6JbDP4gCSeqi5piPK9KQTAHs7DbdsfKe/VQWZRFXY
N1KlDNQdJPGWv4OLh4mrMe6UX/97RhrOtRnBMYXUzN4D0j/mNbUp8k7ik5y8yAm/
7pQTKbjeSqvlTWKagVnu4MNKzFeZHNRRs5k8vHbvh+hFCnyBdyiVCd7j12VQ7/IW
mLZWcXLxAZHozGG/MbRjShfuPKyeBwGk8UrCd+nh0Jbjjn/wqIjx6peB3NWRFnsG
W+WHQpukvKuI/VW2SHEZpe8rs50ZzmZCRg6Zuj9lpC9XMw05toxOnu9Pw1oEjv8u
CAAQvsuwzoQG7TNJrCHbFR8WXaS4oaN9xBHgBQDncGwStsOQfWYxN57NOy1If3fq
jfmxtm9l/pb+dhfplBywnJHt/rllcPE9ZNSLPSHgVWje/7GDAobP3B3dXudKWz/j
S8761+5NqTKKE6jIQHTangOnOmqnYwL7V0dSeeg3WdOVvKzydoLcBqElTWXK3UIR
XJQU7l3buyq+6P0cNjhtXmEkzKnAKZu9z8vl+l3GLH55vlLKTDvyNOfE7MXAbXp6
wcTDsY/1YOUBEbACJx3QsToijtCc6dbZ4mh5vqCTMhQwFckHQxTCT6xsSK77laub
aX/JPa+KSWujDZSNuVIQci+3N3zWZ0sxqinCapXeWMEyhHYIhRJ9DHuGPQLQjzYz
s4zes71RQZXVk15coVHoFWk1BLYuJLT8m0A7tvJzENib9FBNVVbr6cRMWdbYn27z
4OTNSbmgJ5YMLMrK7MhkzobJB2ETZDg4jduNylREkb2dLH35C2iqE4TvC4NwhZF/
pXucOUB2/OCPoFLkONFprRl/BRDAHL5iXGOIEiGgunCIJ3Gjt+YVx51hkgAjFTJt
K/fopHO6VJwcmfwLT8ANo06lt/yJLmTN4CFDBLt2MsoZgMZH36xLmbXnRFRPdGR7
JMV7e2TDMmgoR6V1yMaCnMomk+IvEHifiK0sx3An9ESfn05DwTI3NYDKqfXAq4Z9
aTcQcQgxyg9KDucIH/Zmff6++suEFJiXJFIbEKu4OfgMEf4yqROtEVrazTaYCVpP
dx88EhyZ2L83eY72cKad37r2PxDyjF05/CUwsjpKHgIivWhAxqjk+GWsi6gATkm7
DVNTRIkR8UqfDJ7NkiPFujL/t4XJAFwXOY6t4dMgHq+0huuh+FyJwvGcX+NqAooy
oFwldcIYnejJ1wiYf5t8KnME+4d2/TzTF4y058LQZtrthcQBVHE6p/mAZdSRkflI
vjC/zKDuHmrKgpCx1FjwSO8RaExOD9mL8S5dT0qDqxqQpmGpPewq69/eAxUzjTh8
PyJ741lHGb2gADOXC4EkassasEa70GSWnaMPp1TTfX944kyphlbXIngLOid7ZVa/
8dlf6h2tu0NXvesFTiMiXDt//6HaDifXj4RW+nPtSk2Oc5khArmcd/6/ON2Vabdf
LB8i757/obf2IhJll7QL8CGBIiPMNN5vZ8+k8ptzRGOjlF8mIwSt6kTKEJOUuBca
NC6ktzWcCe+L1Iet84LMpfU1ITBgKVa/bPnfi++2E5+A3w0PCa6+hhhVud0ic36q
/mQiM1bDdeszceck9GTREJ48PaD+31AHrxPTh1g82qdX6DZPfgHBEa4oDDZc6ibb
eYT3MJ7dFuW87m9QdIWP8FuDSdFvg/UvceQoTHSTKO7+LGXlCg+2uFfUJhwUg7f5
0iBCcoDGKq/pgNeNSaH7OcjXLCz2HarA76onl1mOTyiDmMkLpgHcEL/NmBhDc2+M
L2EOyElagG6J4x5PQo2w1lu+hzXFVE3/gfg3ygHNomE/WVS+Id8ZwsFgpOuWrZ9V
BBovBxRwfoHrawAXRLbddM0XSvrrar9OMV4roaPJxOnP946Yj1O1+5PwJ8sxl89i
d2VjOqgRBcbBua3W1eahNKZxxAv7H+m9WuL9+duavJ5kYyU2uoKBR7vw0jiK9YW7
da4e8Fm3DZbdq8lW6WlfvguOfctSRIE+VfGd5SUqOw5ktbz6cv8SJQnKs1ksdElh
NAp3aWpI6ZnSCSNQBVBv0wt2Jxlw59CTzq12XYf1W5JOCaPZvvDrbRGAywNeoHXN
E3lv8oKFvj5XEDSAi3fZiRn15eaHYFE1MgKuUs+wUyOvubTfEU1Sm2w2ULXnBI6h
VBtCt67PaTcL0CEYHVvyWS6qLTVyfMr+3YrAXQl2iaQzWe8VX5vrEKUk6jMkfm0P
n1MtpcHP+L2UkdNMqGINcfPDKacdKP9OWQ0fbpB9giVQaHqEqyJzWo+KC1LCJeHl
ozxooR4f2xJB+ubutwW4jDCUCcEn5x1oBWJUfG4tbacT6D0BagVS6vRaY0EMcW0k
t7Twg2TjfUV4of84sf5PyDQZJ/u7aPe5/P2CnWdzuXxoV49rtaHePQBqu/HBt5+g
L4kLnNTTP9KaPHa/c0JuNkO0ftlh6x/ri77ShKgiFh/e9rNx12HjdswQkaCSWEI2
BsrsHfKnfixW8VNDXfo3INuZKZLG9edxKMrvExG6VZvb6PxvJH/c9ZJ6HyjlK8xn
hqYeHlaVZ2f7LT7udpPHFdSdpd8Ml8H6FNXecnh6474hrUot6W6KoFg9y+FWcL6Z
wmuy0RLf8tWmAurCcVres9OAvfnxIQELZTv33WiD0soZk6hQcAT1rU/WPvqMw+X1
GwqzkI8+zOi25KEibtpY16v+/1dVgXawBxBKje5LlOCRLz9ZAvYFLo9egossdPjO
0Lnkc4ed88hSgQjOZphGit4HfU8PBjU8VScshDktctBiAVTf21lbjKw9wwDW5wAh
s8O+iiapPeR/j6lFM6ThBRDkAHpb9JOUBx/xpSJMB//sG+8vx27n2s68ikz36wG9
WZn8cftmMngd8ZbU5+/nCdqyhpt8j155SiuZZOwcO50jxNswJ1qS9iu3mhFJA5/c
xPL73Nn06mSnZGassdMiR2cYm/PTFmpCJEyGgy/q/SaWDPgjRR3WJlrU+Id9MTnU
1E81hnOyuS/UiQDjT/muF04Ycbk8TuRqxL7NWqaE8oY1uBezGf63R79TBsQS7owi
hyg3uKhjWTrdw4HTHuICbodkGRZoUsu3Szx5ZPHtQagAg4PhhJeMY19z2gzg0B8K
QnHNIk+ytLHfCkpbxOBoIkiWs3w7/zRU69gua9jbjka6Hws6vowqHNsxCPNrzwoM
i/uBObahIHDdmdimXVJ7/XFBnZAAViVoSom740kQLBQ+L4B6CAxhxPo+PT3lUx1u
6vW14K/dRj4BGGA2wOdLc3NVdvJestlEpbUFmF6kyNU73Bz5P+7DnmY16pbX3p3O
LQuEUIuPO7+WrFTjvgNoB/MtG3WBh/CXCJsyOCQu9BBvY3T4BTp8pqK4YMvRaQbG
INhODehSc8rRdilunycbZDTH6LUauxIZlP758g/BcUhZXgBg2Y7SJjBeLuVeajKi
nYYMVDiA+q88q6I6oXOUxM1/QmkJvnEKYVW5KuOKf5CePyccM6YeuIPG6q39g2eq
aey4Ui+mjFtg2Oe1JZ4Fj1KpAhXGJx5otTTITWr6eTo8hzfwM43aTrrhoHguDmcm
weJ6+yzwoNKFeycvrVdAXFDs5m/QkRo0t2Hogy6SDUKnoy+0UsG6kT8NAOhpZQEw
HVC1VqIHK4szsNxa0iCJZudr5of5bw9llgsog6MgG46uX5cx+9/SYSmNsuBZJivT
382MfwrFzEvqlvTqcYHf/2b8ujqPwwdrh/07nu3+ZmoItdBq6O1PTYr5iGmoRSXl
SLjBDZi/DBe7mssQTm4/gE6V5X81aaTb40Jme5zwWZ7Btf/VfuSFWbFjTas12vpg
eaWwfQGwgHad1dHpx5cJpfuOaR/VpllVmF6xJ+RYPJiNjf9WC/NQ/dnz+44R0L5c
4ZizxU4YvaroTxiEPqoDGY83df1SCzyxVuS+gUok0GxROhpMgKwirJtxfBLDFkak
FYZUbWmzzIAkr6H38MR0wznJaOAwdUnv89vOMGtIwHlR7dREAZdsXqkSdCs7X+ZD
LR5Q36raVODTIwq5oLU+bPHJmPHaWkNAhqVYO/a/UWb/OMm7owoHmv72xf0bZMrp
D5Ju8ukqiWsVApGNpk91NT0NEa31z+irl8UYw1/QBNWoOU4nx8Amfa+f796ijhPM
EgIE8CFV/+BqKArcEGuKXWQCgxqipw5ItwP9AB6cYlaKtVyr10s4XFBN8YmdHIKN
jhRfv3RVgSUA9cFywaXy6e4+DgarL39gIUNWwlBaw6fBhsM7r7OW5EeF7xkNKzYA
zi6A7sptC8S3RK2ov4epFa5yb8ICMslpAuEAkKg4WXZXTJhugNkt/F5Mr1E12PZ+
6A2EAc4ilsPI0F6WDaBJXP2NoNqpfvsn6XLceqwvmLD37u88Ja1o9uppTKpuREHL
kNj2MJlY5qY7/N+LoqEA6ctHRS0X1RpjL33OqL+reMluhsIQkJ2fgtZ6R52B9XRs
zqL1e/DhqA3I6setF2dtW94SM7hVyKC1G4akRapl+D0B7v0MgyyqE/5Tfud/D2k3
RSpLMTF8tQhQe18G66k61UUeCC7NS+3UrC+QsxG4pn+32orBoQy10iBXAy75fm3O
QSVdbJbIhDzFEugB/J4OxjYsAq8l0jpDXxoaCzSkC7tQ9302cimL7lmqlwFcRCw7
6BNoOQE7zbaPLsDUbsuykDu1ZI7XJYld3M93wYX3t8e5BWRfjSJGZhWQ4Wgmu6U7
aXrQ5qfkwPA+XHVhsDNmkfrB0k1zws6gPxUXZ/+aLA/1DW03jmGGLvYzhh5noslN
Gk8ZZ9pObkLnCz/F5Ja46C48guHaDMS68BhnnHOqvReDDCyY+Lgsxm0le5TjuLK/
b2lTb45Xlnkj8UaudB0M+lH5Kvipwl0HZudT5dB++0/Mud0D9MfhDB5UCKmpkPjT
P3SQSNjVfyR2aoUxl7XzKDw65LrETVOah3SkRP64+yCfCAE0emo65I8Q3HZZXWPG
l9fh/KDDLIHCBP7tjuXJRJS82EvAj6QYFdP87xgvDypFZAsw12T79loKqXF1u5iQ
7s+wpLyvXC7JB6OdQEAg0bZtD/gdnMpNtPNaJGLGFK6ge3bi8cIvx6g4OqvdPYFt
q94dcw6eSSis2gQQzgsftSZvi/icHU7pRO2w8tN4q05UZNreziubHRDDZ/m5X7LX
4WfTFczZZEHGp8KCsQK8qD/lzid8P5bXtA5mXBir3BoD9XSCDDW4DAZv4KXwA17Z
uekbucpTaHqrGD7NghmWxoDTtx6FF/bfUP9RtW91SZyxmQafD4RtyzhzPpkapakY
UOCBfAzIYX8URcVUS6L6NBzX+x6f+JucLpmH37VbiG53v9UI1mrkWZbTlv6+rsGZ
GOw+8uxEsfWjgeQGJuOPLY+nxUzb0JRSy+2IAGS1Lb9z0CfgwmbgZbrGrXwXvws3
uxIgaLpPIv9o2D4QUK0FNi3ZFciz5vpy2JOoCHsoyG/9pbsZJsai5+g3txCDrx6I
us1ZhBoEb+BpAfLrm/7fNMp96ZQBjOA/cw74CivNu6P472Xx9vR+N6bikKuGyQbA
ZLudFDFOTDB0rxqpf012VjWUZ19heJ/PLXGjnD1zVCkvdgvt37oIitMob7J3iUe9
3mG5B4VRVTxz8xxJivfceXFFKX/ikyfoNTCEC2WyGKbTbcR3CfZs/bHijaHPdz62
f4YAEvNaqituK5+g2trUdZhogy56G7i8S7JWJHk4Am2cYcpHsMYDzSedOUOaLlij
k6Rvvs5iiDkWDzOCl7EpSHG65fZBZoQSYHXDkKKqqau1cEXkDPWxHh+UaXziRz8R
J6ZI4In/Ezwb9zgBU/3xqV+qtCc7Ohdzl9tjgLtLIYXT2VPS7eZbZ9WYFGvP9Vyh
ONjUF2pulhDWf6lijpGpvUtgBE0q8nfjp9dvIa40PHB2j82wSGr9UL10QAB8I8LS
Hr7XigqbnGG6nIIX/s/2r5whST+XfG5Zhdv8pMQMbPmdCJxGjlPxeNu1kORJDmNe
zjPPKfhNM+jQki0mCHfnEVXcmxmSR+cNwhB3sKk3DtgaiM+C6BB5CIWT8r1SeNa2
UBXmRbxKq/y4eaAl6ljUyY4sk51BiU/DpNAWDsS1QIh7Tc91BcHlcIBc2n5fANZj
UZoLYLYXl7AQplJ6QsIcxlLG1Ei0/ZRUFbtmvGgwsserrsIbOwkdwQsSbnIoNOhZ
6cAcpfh0LqsxIL2OeG8gtuxt0yf0NBhsj4Q+AT4SB9bZhlNVNfuFgLSeEvm5pg8c
29ZfVTibHkrXoSPZ5MacjSfzSXaP8a65blUfs97YUBU3IElmEaMd6FL4sFqIcfUG
WfUaW4K+XTKNpeC7Sfo3ZM1y3LOljMNg1yg3puJfTeFmJ0kr94yDSP6ps5dA369S
/srmiMEr0ehJH35wNCGJfLPLV0HWAHkfAW3fcZYwbjQj+gGOoV2n7N2mF+a+e/0T
xVLixsrwVUrZnn6euY1oarxZqbBFRyNtsOfIRYhpXZMef2kt8v+gMZiwJNE6WO80
NG33EpAYR9/6JNrKi63Wes+mWHnn3Xn5gdtVUbFfoAj9OBaljYk0s77cRwTAnvcY
WLFvtUZ5EKhhZ3SJER5Gh8lTtpEZDdxKSv2XB36O39g4hTlRS2JjUafff3jYn+HW
4tclt+2SIe+Ly1eK+nuQHt76blstGqjeVWiD2/uA7p/v4UibbOC0b+M8oKhU3ZdA
E8uUBbOhZAY4rlCeKbctPR3d6usmcNK2ttpgNLsrMsca89MrR3G8OnySKUdmu2KG
wunO9aTRTfmBGoIpqJjceX75xqkGsUo7N9Pjs/k+IFXfCYAvTp7qQL57VbqC+frJ
oOIDGnJQhE1lp8VhGQOluOmu2NtvB6e/GPmHDL6WgfSvoGddQL48WhOJvnJfcmLE
SxrJMeZCqegyuZ4dKx7nYn5yv9P/7TbCfgQ47+qk1pSCNutyR5qHPyWFWHlv4aeX
tCujWTNNns5sMSDj3yLJMHJT6FPBdeKFvu5D9YhP6nI76xHoYKZI0mC0wZ2oRdLF
wJb/HIa6l2Dpce35C4Q/hWiGyWHFXpRh2IHGE/AWadgKjCw8LyoQlUrZuVdH0SYf
pszHt5DSh15hK6w04IYfXcTJgEWadH75K8tOOVDGmCgMOInHBCDVsJ0TTo5XENre
odUMAMefHwnyE6xpbOwPk55svLaA0tenpqOiamv/I4fIKNUJ6/eix5zR4TarOEpr
ZO4Bkj5VgtayOfOrWrQCFVh+WY+KlC/Cz6guYZ6gJIOYj5aqgUEqN/DmLOjMyJuH
1Y5uEUo1FaO1YLqkWhukp6KkQKR8Q+UHwCkshSft8TGxIQTDs0YXv6qKmFEFw9I5
ZdCPhOaW1Ti1GlS0/2CoCehem86pwE0CnOpHLgDYwWQsFbj/198leVRTIdLAn2tE
H59Swxa3+AC6cDE2wqbTW1VOOamOQV0vnqwQifiMjJz2D0merJ5fXpBklU+bydOy
FOxFyRz/sTsY28P2uW8YDyZ7X+yJe6RGkzYL/wQjLA1+WNcz/JIPzaZ9JikEmnP5
LvnT5TpVSQdGslPv0W5yW+QeR4H/Yv0oNhzRfCh/UvgpjnYURxcWdyX2EuuoZKe9
v7Aq3A9Yab9GYt9CSbjUSFSxlnvHqr9Hi/B8KNqS1BnoZ9MFjyFlUGhf4sEpRg5u
GBWgePsbL7cTGBDOv5ixt+HOhI4OvaujE69aokFf156FcjNcWD8pmB1NaEEe6JfW
6KjypxvsKx8h4pazD7kmfQTDyjqN0asbPh9uyNSkYlanh8bZIqtv5qJZqoBjjQsS
Ms6zlieTljDpHSl0O2QjKnSpSceJtwSXD5Zpg8uQUGm/ouWYmIVJYghqS6y4etaa
rAcvRrH4jaf+R6IwAes0wbuiFvLFg85vTOd5HYaxoOxvzoKjVep9sMI8gLw4VnZK
1CBilLz2FsMvn1sYmEQ1B/AtTpPrBhT7hCLht6b8jtpPwiLfS/t2Zmt/SNjJJO4S
/z38J35353S50LsZkHW2D8O/eqAJNANMcDFfDvuPoCLVSCqbCA8qbIMChkGOEaVA
pUlPjvMXYvhl1apuKAE17T15lRey4izQILnIKQB0r6nSwqJGZ5RZzzc2AmxG9Qfk
diDd1Qxf+syspMk7jGM/npaJ5Y46r8rIG6LCQep1/Q8fvYtP1HbRcj+NhQbOfGMj
OCD7qtUh0+C0aiNrEaZxAn5KzHFoIgc6DJvXQKChCuJ45TcLU7aM4zBoWJBkYAWW
Wp2CAOMEQ/JSSeU1Haa0t9+4NTe1T2Y7RZ6KrRGHDjaHHTHEJ2Ltue/+svLZ5BDp
LrItlQ7enHGcZD0SvrbAUfa6/xuKJ/zB3WkZkWyhz2nwOWL31AGxTeJUJlAhAPEm
BGp0wgh7UGzEjEL7FtvYhVZN770keVulFhzOc3Uj8UaGBdkjX0E9H6bwfj1dW8DZ
Py6OE3shvOHegVFevFQvcq3asjIgC22w+AgODnylxgEY18D+j9r3ecPby16GxoXX
YMgUlEXItj2mmpRFZ9mxa/+HuLLimoLujkBPYVDfe+c3j34FoY1b1ZLvXuzZno4g
PaNq1qHbLHid55OpIdLJt9XwcYV8TpW7Eq4KZfKbHYPBPNv9SmlJE/mfWPLdldW7
X69I42yE7BPdKCwjozT/l3Dl8qSAFqbiOck8SdS6xPexgXnieF0Wk634OhYIxDFW
VSxtFKI2sWgrg7SaDziJSqn2K96aSk3o3N22+mHEPynYib3/Lou3PB0RncRc018W
j/UnDyPye/26kE2OBhjSC+toKrFoyegdI6hvpN1ki3p801DLiTN6Q+7leJUpDbm4
iPYEqSxCZ9qdvovxY6CHWqmRVMx1rbtrV2eFgcXOZiHuqIszFl5X/5JB/GGWCYy4
VOryBjaJGVf7sXwj4emPwXML1tCiB9eBeJkusMTnNfAmDQLNFqv8aVPDmB4LBk4d
d8g763IutYvMKGWtD9ojAA+rlhBiAc7OJAFwv/u4mMBBUMfjOoKo0ecUp3K3U5XP
j+fYJvc63Urqihw8Kk0qu/vigysh268IbA5y8UkpLjfOjve5P9u6vVeU40tWrGP7
Co+uy/+hbuD9YJhRVZy8m1rgtY6Bbchm0upEy6v42RJYe5SthLg5jIKGjZdAd7Zp
5TIkQ5IXzz4SvzdWYFb2tHHBpEHiYrrhC63ltsKs1jZ/C0rTHEKlI7hRNJUuF2pU
7nQzQYp74O9IpoTyZQ0upB3DHfB7I4qeYOGLAeuYLrrBmPFQE/qbc3yvbIjuVtCR
Ng8HcouClUGGfJxLTYQ+U/wlwLwmk1augnPyjkpdHx0Q8tHNHLH5FoRzDVEtKenP
iKBc3reO/ua3j9KlRvEgI6yTyUbKkixIxsAAadaVV8W/wqlG4TFq1cDKUz6t+B6o
vzqSAGNdSuou5/uwaX/U3UOD0ZXGgkMCT6lyvFGRf6vUKvMvG7I/ICRk8mtEa3X5
ZsTRvfZt9vjHDK/RZaVddz7gBrsR+piYnJh4KI9x+lwf+3DzSMw0FSOCiV1KNP2z
9Z32aPmTkRKu7S7qEZaVBrSW0ZA0oL4SIjcDRD/ou//FFp1dJAiUjrmwQTHgdpE6
87xyearUiK1b92zUm++9VIcHW8YSALkhWu/UJ+EA6zaWHD3kXB8BhmdyrmZu6dMJ
XU+Ey5twEzG0v/N2NJVP056aV9gOp2knyAFO1aZCykf91IV6Kv3JDHOXYRiFVP/j
1Y5ZgFoBnW6d10MQ4+eAUe7IMQ5kBQw02KJwy1MgqePIn5ANY0U1bvNYzBdmQrtG
XmUNkHAg9mCrm/x0+4vKU+u1K8tct+ja/aFRrriDR+GWyed/ts1cqkynuzGYbTLL
Y/qcLbav1+z5H/pYm59fQl/+7o4QOxlgNmkVYOA2T/y4dV5VqEZ4SXLvM3O6EtaK
C/woum8Fhs5gn9osot2kA9Ij93WzerQLvdF75dD1SezXpeOF7qJbH2JWNl+7PzC+
yMEiT8m+iQ+bNn9Wm/ABKV4qLxT6papsQ4q084nFoRrpM+KzsFRZtQa8EyAokLOQ
8yoER0rhuZ+UEV7VhH4pOGRl8K271NPa8N4z1hHq90jE1nnuP7xiH0G8TtqwSywF
lduXoQ3HU+1KuBh0LPDmKKkdze3TlgmfPXPV1G/PBzBSE9FxlTs+zoxdRwN8CUnU
qVhnXc6ZfffJWf0T2MQVOpIFHdIfnxtmIzW0W8epVDPu7vfAUt2Al156biJRBe5h
f0OjMe/MPQPjIPQRRZ0iy/W4mnDTcM8QzC6Yeopy2i2T3r50zFkphTEdt3mASI88
3aKD2v636D5u1HSfBl1NNuzP634aTdmX17XesLOdTupmCifwKy6QyRl9eMgnySSi
vHZpVrQGNFrD7uQ3YhlB1GuRcuq1RFDe2xUV/5cPqdFlFvy49aMAqQ0zGjOulcED
FlfQ4PoiFKhCQHJR1RUmZ0YzpQb/fW0jW/oi4xREIl+v5EJ2RBE56R+dPK9m+ObE
fkQ05bC/tD+hjdJyTNYx275xEH7aOx+roU0O76z+ru9KbFTtCRr7BGh7vr5Hgn5I
a0/rwGPyW3CBzLbAg4GfEcqh1krkV7rmdSqUpDZEcdU/lh5vhnNbFetf2gndv7vd
58GtB3BvxHQWGnDv5Mjk8z6E60TZKfHsM38F7EOFi26+4BWKF9W7son9AOb08AL6
Z3pgf+zm6hNx3Lf7js5WStvQfIhqbLQfJE1kACBjWj6RMbrr3epvTuAsvxP6Htok
p9J5EbfkkWDyycGnV9afoABdB4pdcH5CMSfjxPHJotHTEuU+C5C1SAiA/XoMuHNj
AwGdOuJ+cDvVf0OSRvjm6JXV8e+Gi3F+w7NTdBnRgr+nzit5yRtuCZRcneMpJaq1
29oqrBwJ+0beu6NjIUZDbhbL+S9AvYkbRk/97CpPu7AqH4qnZ6a1dr4qPLts1Kl7
v/SdFwE6R+6xiY84lnwWmxHmoT2IA727g2U7+lA+dEG1kIZfUj+wCOqH3zks0AMF
fItQobUzgFtWCO+r2+fObcC3VX1+GZz0wNEkhzgbfdzJroaQAfxGosvkVCd+9DlN
hB+ptlzGpcFOKcYWp7vL+Pn8vi6zCvqZrF25bEusef9f/uraj7ff64tUQm1yc51U
bro2AdKH5bBq52gWN4Sje9+kwKd3/UqI5y9VD94vr4aKsGRjpTi3Xw8mN57GZyuy
s6Rwb1tfMhzJOCrmCq5Lhv5gOVQwK3oeEljV/Mf5jvujq5DD6ReHCz9NezvHFdgN
ZmxnUrg980kY7zM4mlhjEjUGoyK6fbUgaUMMWEZalLlVjMOZQfsEfRObpptnRDMC
0RK+ejkBiToJ3UvWLgHgEe7WjD/ii7qMlZADqlWR0BTDiNSIcWRiNubIkOPdxoIY
jWseVH38H2/EUkrWcZxAdmfDNPw5VWXceL6uUD/mfF+17lpPEKt37Jz0BHGY2mqZ
uFaJ+UosPecb6F6rNpngBXGn2NIIuBivFmzNzHFaCZ4amEl2Iy4HS2Q6Pp71K94u
Vv1BirQ3irRUdKqpvvqOpvGRCu8sEQExMnnB66dAQ0o2sgtWeXvggpvmauza+EdG
jTat6MUV/qs9Uzo5NcztHfPineXK9LHLB2pdojfpNEG+OOZEBi7M7B57xZmqlyVh
MSol02vYIbEt86CtYPiox3Zog31sj9WUEZ16uhWOsLKPV1rA3Qb6l9BphEfihmUX
ViacePviLlHHqh4tjcy5WDQDVuVz+1FGUj9Wq46rPl3Iq2Ll5U5RZG1rBUuRLcyI
DhcvhaiVEilzn+zh8ctkjeLlzPMePw6GIkVWR8yacvIWkZdyUvOEXzYdE/rqHuoA
+jgM9EhY6sJ7AxOL3ywP90XJVZ40krxKtTT0bBGsYB3KV0D5F7mHVaqPAFtl/YE9
3UK5Oec6PlIO0iB4Ks498pEUaxeY+7sUYr52J3JkwHkbQAU/BlvREQeJ7bxQhaWP
X10PuPeIQ71GczCe2k991rIuE7yItZchaVSQcUs6n/QrfI2gNgOWtOwVdTqx/J+Q
i8TiPl285hUHTgv+q2c6iU2T4xv7JTkjLCXv4VfScWjzOolJrz4wNPIhLYPN86wV
tJH1sxyLpHw93AGIQEzbBzKHFqPWW8pUv2rpNAj0Uwj2SuvWC/JVc4mHQkDUZLcO
Gem0R58/9+QqxfnrivaCTqzc1/37UzGhLi+7K9oHfMa40EHHkj58D1BGk3UvABnE
Xm/8xsp4DH1S/Tpq2aj6G+XO8LXj0KCe6+ZXDImZNsgt6pITmycJ5R1x8dlu/bM3
StBXrQcZag6jFshAEe2vzNLkhYTxb9lbIZsQAM4vDjoBMTNQwWSgxc7UVQGV+TEk
ZmADIXZOn0SphIvzYmksfuG32o656iZwF/urbAfrxXcWWgbGFXZvhS/dbNJMdQvf
u8uFSJtAREzKPTZerxS/LOXhaKW3KZjssoPOpZ83Y06xyK/HAKp/DaOS40XI123S
PV7KP7NHcF3qcLaXLV4KlJGd9AFRR75vhClxWi8dh2DSsK+wDP1s1i+8bNtADViB
eJbsG07HJohVocgWwRd6Ip5uqETU2Tm07TuuZgJ21SzBvSc8A8YMIK6UrbTyif/s
D7ilGLP5vvTjU6etos6tF6pRKlsa2HGLIWf8azn8dbX2E3e3Pn72T+LyGJvlBCXV
fNazUSaxM49qmuOanh6LgFKkIPI15fIV2aJw54C/ExBnmO3/yeSBRIJrPndCcukl
b6/Ec8ioA3U1S7gT9g6nW9mtfXuvF6Sb5euvgYS9e7Vm64UVwWqRWn5WNkUSxqzf
KRFiZZRg8Q+Zd5Jen+9rpHQMzQ1vU2gHIAEbXwVW+9AIRJO5tniAdFOvtOPyXomM
UyAlaowIm8e3NoinHh76Dgbk4CBfL6OxOLNqE3w+nIySDRbA2oggBc12E3JmLcRu
XotvQEx3TDP1J9ql6IpkIk8lTaa+JrKShvt2lMMXdhT9K7Ux1Csz1upQFM+ecp5o
QQymmx6PprPkXwOkfGKt9DeUsetywXL3aFf1s7TR42fOJvcuPIrc1Xl/ZW8D12yd
jRVzM60drrvMQPq90N2BtrQZ9AGhzAkVGFNWAXWYS8W8HKTK8ucUDADccr/MvDrd
ndbVHqKlofJUzVcF6BQPk3wZa7RjiKM11Tjhozi/VDhJ/Zi4oey6ZOWe74YeiQLx
91wYJMc40SGXAEJqC3B/kMBo3Ik2Q5GMVfPXPZDKvFqq+/zLuTxm8uSqEnisiCpM
8Tt6TEkN9RvDGUwGn/X4xTM13nsTSppwrv671TseKiYL3VKT1akNIVtb/jWHOXoc
Ri/Lag0ftwAbO/gJLbGg2j1GHmZY2SWFeC+YkY5cC2TsfKwQbK60q2/u8Y9hasBK
0aVRzelGxsza3Dyc+Uh7QpVC55aB1iLzh1H4UuCMauvdwKDwrCVvOl7lky8bKCdT
pPrYWse1ZSUg4MzQ/0Hmb/pLCEuvOWbfamHiBN6zwedHAM7EpvGaFd6sxFkJoQUa
6FaniDGTyB5Mvt+/q8eK5NQBNQ5AahjE2cIi62feENA5s/K3PhO1pDbt3zmFvxAc
3OqdWKJOd/GXGyHgHNmcp/yHUMWLQZfEn8vcC94SpyNWhTJlS4d3x1HQrTILj8Nx
wrsExued8iWZkOzHcz17p01RX+IdDd8pO29GkND+2nyUOzHtpoekJgcwt/evi67N
CAxtzUGMfb6qvQGMUH098DhZNJ/ae9zTyWTJmXwYNoTnakJF5kNohDSfVjf2x6XV
V66nc839Kf/y3QmTspTZ9qZU257cdyIW/13uInOfW7Zz7kV04GGV5WHJjv3SBOkA
Pjh6gziThbe7GGRAHOMOC84pU/EVMlpHCYnbg+8prELpAMdah7KPg9LENH3nDIoP
Bj6zb0Mb0naSsENL1iNEmd17gjaw/8p2OwxfqV6wXgecRViO6QvTm1Qpa/nIPW1x
bcrtHv5lj4m50uIwqhEpnTSkY/9i4s2xn6ePiQZzbyJwxWuzD035yQJf5bcnGhoC
hHPsJeovdYC+Xqw8MeVd2vaW7JdzgGRA6oua+O0J8Os3ZTHCN0yC4VLR/dTUq2D0
MVPQcSvPhAqhu9c8xKUxTq/arBt1bY/Bu4/ZmOJexHMI/Qt2E2RHdw3UPkI5s+mC
eACy8V+QnuKec+NpXhtuwsZXbNzdaG5Qtxn3kiRMcTb0KuIpMPXulP0/dsKlCYM7
HHfONYuU5nSSrLrH/1iDL4jm++z50At14g2UYMo9vo3NliqhvkTIJC56PT/MqFMZ
NuwuQz4OSBc+ZRyPO2OMOlcKBar/vdEczH6lhlJIL3Z0mznXDzALpMeL820VlIq2
z8WG/rN3GFhIkZD7Hff2ClzGvg1WnEtg251DaeSNNX7fzAhafta5InYmqAZzItZH
6yLSfCSGHdiOMB0g889IsFyBc0+ObXdR9vKbt95ioiAtFPJ+o6WBWZgGDyjpkjAO
/f91hEdBc8YKNY1GJgNJYcUCP2G4ciHT9W07s4ACc6PFzA9uoSZcHJiyFtrVfOQ7
/MJBUvPf+ELBtfU+OsY6EHrP6noMwpJKdZeHIjyktW2mWX/Dpw93KESJSzUewmHq
QdtRAHBxcJyfPCnE9HrWmDAr0KU+LisQ0smsgydTBeiLLu2xhHJBsZQQrMQAruGY
iZ3Os1n884PQjTfA8oelIzwm3NX3qKMkA2merEVDqX8NAojK8cVeY9Iq4FHcr14e
z6bmuCPKgrVLqN5FDPVNeM2bNXyvN0r8ASbZH6WnZb3FLZTifXNWOv+9UvHkJylt
EyIvWxJzrnmJcIux5Yx/xAgbnXUbJ9N4ErD297P2t/6evKMVQrXvrSWEA+tc5a79
c0Q+73t2SpvFEgWVikR4GaiTyl3gyjR0qmJTIWlYpTrxBTCs90/Jj8dZmF96ifW1
iE7tNGYrihjJ6rBFDC6Lw/cK1JLZ9x15bRug9+zyCrHfvEvcS4iifVi3CbJvMMbN
BoAyRTbx2rMU8NgzrGX8YUtJw4vOtmLAxo0dYoP8D1HO+ZQ/46iB2NCTaUe8Mw+9
uMxCQCQ5YZ10LYXGzp4x9RgwKFnb138f6ji/PxmKV/qi/baAVarjHGL9xIkQDyPZ
0QKEiGYeqHa0S9aUCqFLCImzEcLMCEcR4kmaw01aDlN6wkhYbdWxAQaGuYv2Jr5j
1UPVH1DbwRhm/mJSHEPJ+MkyRMdH3w8F5C9eCJ+j/U6s5Gs1y1poXIOA06/E9QV6
LKvHcl4GYgsKejiUNfyBBJArNrHwMOtOmB7863PzZEJ3ki+1TItQtgThwxnxHwEp
7DKzHqTiFhwz4hTFli2Xqkekdz4RwEWuUwW3tweWE5lSPJjAS6KxFrHU39S21Bt4
gnxA+FrHhJ0h98rVnA1/9zZodyolG6Y4Hny2Ta3zH2bLTUdQgukRfIjYXeg1VwnX
l8dI6Qx/Bw25kXmprUNVYghwHoryS2zL9/JR3QZbotsY9l5adQcCQEfcRzKLH0YK
0RG664sxjH+d5mZEVb9sW6fcv/eBOWZkO5ly24lJTECuhfCIqEjOiInXQcIjYUb3
gw8BEH9j833vQC7CDjKb4+W2RT+VrclXShY2iFouiOmI5cw66SgX/zLBUWbyD6ZX
D9NnwCcM4zw+NWts+Dw9hBmx5KEE1+rxxsa4c7CBo6EW82XA6zXyHAv30VPFOvV0
cQFLLPBGEXk2N7+WuT2UEKZOoEXOjHu0WDh0+N4dJyx1jr60J6AsxYdS6T+jsica
HfAIvbVX4NJz0iQ/XlMMB0+2qJkPLD1G/ZW5mIOgKurtYmb5e1iiTMjOsOIMBnKE
84rjXIAs5eRprIHZMYFd2+hT0spz2sIf4A3ECLRLT4GG+s/mPfp1YjLuMfiAwZa1
Py2sv8vIiyinWp+GcVM3TCiBKa/nHH0fV8waJw/8HcuOA2VN9oYKyL+nRjCQCvot
byWq9ucbZG4d0dLSzazQ6UosqLC35qRdPgiDRqbBMrI7LDlCv96YlrM0SEFvmWpM
gXUbtgbPLw1AcfeUxVpUrsN+zWBKhuOb8byzR6lgYRe9b8NoYNKjZWlyZqShmybH
ZOcaz8d561MqHcII8kUEMh7gO5kFs6A7VJSt6XnY9Q+vSNjecE7bVXboJ4ief5kJ
9B7Da/MhxZh0hlDFP7YQjArt+QhrzjJkbil5TLW1prw4ZKkrhmOluueT78OKypTz
x2Pu9qGJVEdvs1NRyFaeK8pAwQg+ebv6qksTzTEWySJUb/xRtzQmGb+GwI+SWjBE
7pi6R8X11mQBuu7nThdpykBe1ho/8f8/4cubUTfUS2Vkl8L/JycFAdVsOLi9X8ek
NFpYANl6KOHy9CJem9Qglhyaw4SX3sHpGjSPMopQp+4ddQwPIHjHshLVKioc33Fx
mSd1GhM5MNf88w+kNiuqYjhMV8gEtXT+dhw19JCQlkSZXGQpuWBx91turf/y9oeZ
rA8J3luUxX+rGs/nBuzIla8aZ0kh08tBhPfXF5Ym6NvcT8bTVaECl4yAZOZXdFr5
VEOOyrCfkt0thmcsu8vRNd1RcGAIJMkTCPNdvShw/x4WCUj7scZf7F8X7p+/29Iv
Du8pcqQqz4RiCH/tCChFP7B5RACh6kikY1imovRoUQC6pKjxjLDp/WPl87rxKC3k
0NojCr2gx57hLQS5hhHmZ/FWgPjP8q2Xszks+84Twv4cOA6Jo1tAmBLZZ/Zn29Jb
X/W+cEMGpffjnzn9X21Pe0yvt69IvYWdPaFETa4oFhwwRaMrcDhuy9yf6dIsK79u
x277qhvxgBToQuvREuHXnmuT6qkH8aigSar4TMicA90R6QMYoCQW3aLCSWRy3hYe
of9kH62n2v2r71Pxl7838qeZOYKhQ//SPdX5K2dCuCmmXAG2geQ0eAwcO3LXk6aE
FvAh9yvAL6nXdUq+Eijlnpv3wPF40m1MHkbkHuziXUVbQgvcHprh0cpFb9b1iV8b
j5pTReU1KOp2kS78/A1jrVsbrWeju92PHie9P28J8c3M+qpKfK3QxGAqg3aofWKF
dyF1b26rJ8KfcZC7e0amE4RkoXrwkWbOswMspfpblGCELGvzdAMEPUnX1nQk5y3f
Wf4O3PBZpjAAVvKaDayhwo8LsUvnmLtcOZV+gb8MJ3zXSn6iKJe5Yo8hgYZId2SH
FEcGxMTj/qw7oyFhBL+Ay0aWIuZ1Z6cDEZ/hx2XLkynQxKx/Lmb9mP1OnTHvuneS
2VBP1G+kNpsi5JNx9o17RkWbWdrM1UqnRq7H3A2gejUS46plzoSlbrggAY8W3Fd6
iDB16b+CXGUIwkf5Fn9E6xluoR0aX536FZA8Rg/Q3aWHaJTntgLWk24g4U+bdDwr
AMboR3pUN5WgD7VHT4gJ4ZaKwb3AB1ebrC7btJFzCEoKUcJtpxi2puSWaWRVScjY
XnH0g2Bvj5/tlp89vZ+eOG/6QzvmzfpSGkgBCYyt5IZ8+CBATta1DO+pJbVMEPRd
c5uXoqdTBLToMZ+dhoPKR2FWHPy3LaXhw98Rb0BT+OXlsxgiplrlVvzJsRdwEJDs
lujxX/BONRv5LPIK0FloWbhFY+nZf0qGoKK9CmRUnchRxBVOaP2iA3wM+aaO2/hp
l9wxypnGL3tIfK9gosv/5RhCFBVXy5oER1ah5oxqax/HG2MgBFN7mMvwoxLCpXSC
iwqvKhEym9HWgjF4A2BRpNfW973PTMKy/Hs1TYncyesiBDAQuTTzsOipVMpJboTR
+VLvpRAeGnfYN9RYI8BlgmV79SSNg3f/3s8cmulftLMkV8I0yxxEXMJQRueTskXo
E5bIVKxEJxJvKUAH6URFmWaoeJGrlN1yOI3UA7B/GVXb8ZBTPksKUquKSBdJf3Y2
idzrrCffAnOLy/vPKR8bttPwAIStkOZeUHWvglc5hfk//w0G6IbqptGjiiY/cW7P
ynUxzQNhxwVboAQ5F/7cCpLAc0E62CJsxYE0oci9CnzLZcKfx8a4iiA5JIyJSqFc
eldKOha9xFDfwFdH8zs2Ui1N7+VY23rAg+Xj1a+42K3Qea1FF9S2ZmoRbOWqpqwy
cEPVKdLhSeL1NBKrrkWfAjFHPlpHF7IEORXID8D/yyH645n/fSIQ5biXToDiimXe
SoYv1I6SER6dTgrxpH3Sr4vzqbzqK4QJq9+vRG6myRs0KzUfMqMtFG+r6bLi3RJl
NJucUvCNtdOl1yMpTEooY/tFnrr61SbNDjkralym14h62zj6HePTwIfSJg+O2f5L
/YG2xro2gsTLZPCyButYNzG9iyc7sAVBXqAdUc5uHts96nw/JQzO0vRgesJor9bV
25H1Vz1SkKUxcpM6qtyDvh9sBjaOrUqmypTahE2l/gKPZorTCb+LC8eNCz4TC2ft
eJ1K5MaYhtwkqyVNGPxCgKX77A396m4sHR39QEb8W1UT3ZmesfT8wfko8szGi6Co
6rNCOOJEDEIbcx1N6W84kWG0ry23cl3cs49a4SniNilT47ZEYlXn4oJwl4fNkjNi
R2gInaJLrmhFVQ11mOl6dQF/O1qRJWEPyXATR6S/YqJKkJUdUs6m3aWUanCmSOL7
us7pXZqQg/r/lVla6gFTNmWS0/v3YTrHFhKyQZGBnCqBUlKdFMlIqwzryluFUC1T
I9sA2LRy1SWUYxDqA51kBuhBRrG6NiCW1Hc57hfVOeT7t6LxtIv0xF8jfSp12zEP
1oYvgbhe9a9pX0yUvyQMZNOQczazGU1HK7Wi4594f24wYWPgF5QwrDDBgJt6B0y6
s3jvvqYAZQvnGAwEo9JR++5cS5k5Ml9ssuvHR+pKqhOUz4QU9v5oMf87XmvRhERq
NmjCmJ+uWTfMwNLbKZpCPmH4YYtIUgSg0IbFbCwpOGxzgsomHf4wSX2NypMmhU19
O/+f9x85mTn8PvlpIMKAyZIOCN4blBdi805AgWeogY7IuQ38YxcomWX6xZJmvWbq
uULW+aDJNipwhEubXFz8jVOhjrMU2nsppw7b5mcUzSwYITlk85B4IOAt+7paadj8
LK8fhYkm4IOE7zXgX2wFZQrwpanoEp2dbblCjrFJ1eO7FckZwecK6y8FPUbSDjXE
YaUh54SxvqjTLV+rmSauQ3JqN4tQv+P3OQYH1E8x2C7rtBTcRXKnm6hkweh8p+2L
Zf1ILY9XK+Z+ohiQcnV3RxRzc1MsRJeP8GAlDa089j3bySeazIWAdLof+ckzvnj/
k89I/6yh/68Q+v9J5X2D03fnrbNMCzWkYXGSCaZIwicbPFatZZkBxAZEjyUbA9+/
fvvku0e2AxoECZjo0b45JIDNpIZfSpQ4ABzV5Mwoox/rTKyukTehmYmQc9T6/eJO
Ky5nISnQ8HaPih3xOTCI3GN2CX7zYei0qpkPEz+UNMPG8KGr888nl48/utLjJcLx
YQVtJ9+ejJqInBKeAGCN3xkCnIRzCh0T4D/iiYGS22dmGwQl3i66GU4Xs3RGvGwk
B8+7U22K0IP0+lCgg3D1U8Oh6yVvkLVJ4cPN//vClo/3TPlNjh4KfH+VVow8xeNm
v8Qwd/80nZy09JhUkJSmel+OhFHK2ydXog1tz6Cwfe/BXMPNCHJX1aZOrgvWXWEe
18MQXIdPS4uq2C8At1J+BPzt4SmHtPVmeSoKcHen2t1VFnIp3NibbXwjFP4C73Gl
VUQBwR6wqssSATwZWjV9T7bsLlv7Mq9Ypj98wK4otQ7S70ppgyAIQwBR9fejBP51
zi0SDNR6SfQXC52K+Dr5f8rB76AOBHQlk8KdVprM9r9sIn7JmU/6EdyEPy15MbIt
ZtCRR0yWeZRWi1mJdqdimJG/suQgGOaaA90AxeKWWtIW3abpull7NpcoznIQqmGm
/T+hiri3ds8d/hZkRKd1cY/UhELp8w2mEvpIescqWHJTVdAKKramLP0pbJ6lepFo
lWk05r7zsapEHcCeqN7xX0rAx64wHag/0U1FSUCAfz2p+SjdSEnobVXCYe/qTjjy
mKNXt7EslzRzrwrjYso3irvsRdXxSRhZaCc9NkBqBR5D9Dj3P4lW1F/p8O82+hK8
oGTbH8Wp4CnvIdRGTdH+iQkGUcwSoILfV+YgL2mM/WF2lFrNjiW5zf4lGu1+3Izk
XV0ibFlKionw1G+sKY+DFAyNU5sjrh8HDVTYbtle5XMlwY5RfnP8LjFW3P5jh5PX
AJ/Gw6XOz6kRl+jn05RGDlrnHGpWy8FVSN2HbD1qHYyRHfsTPdYY1C5ZfeV/XqHr
TWJTVL7h7D1syPfLu1pFbA+4u8tLEsd0MGp2qyOo7bhtk5IqgcHu+o6fMxx7TEao
8UA73qJa99mqtVA7fKtfX80VbafGpBp3DHX3YFO3jmEs7YJq42fL3LkmDCobKBiP
jq571e/H9q5If/wVGvA1QJb/sUfp59crnhV2Gl0NVlJVoE+IjqPqki4u9LPwlAzp
vF9lGf8P+6hhnk3TI3ZS5THE2kssfyCkukw7a0b+vNWNerka3zgkoIRJzPC3QL4s
yQ5pkTnnaqV2Gn3LLyrqHexII9pKRW6vB/LZl47XaHz+LBKY28RwWxIE2JWzqI02
bdmNEmnUxwO/8kZXhMRlKJc1/l+3bO9uuRiP1lrTtq8il69CadkXWQqJR4s2Y3Xm
rdiDKBnDDHR9ulAmQ37+2cNlfa2kyu8lOGxHVXwDlDpdXvsFuRj3Xp1nX9zPM4lq
Cb2jS5jPEyp47yQcp8U8w3qxBon1ZXKsGFDUZd7X7qdkDuaCnlvTgA75Uo8Qi2OZ
cDOAho45LfNS7o2OUPq3WG6GD7Wop9IBIciZgZ7e8sHggaRlbFS70NKd3N4ggH+f
rPevGZDDy/nc7q0OiENbo3eVWIhizsgyr8iFAAxgYfgqX5HS3pdXJlQYtAw7WfrR
L0WN2V6qlFyhLy7cG4q/n6MP6dE4Zi38lkCJGU8zE5RTAktWOmudeDBfm/ixoB/Q
o/C0LFskFh9G7BYnQng+/+GixdJac478R1Sd56qCFSzxFr1RoK39UluNwNkE0kza
9jO9tvux8ZriOaX4F0hH/kGbb6HoHdBOklqzY/kG5oT6qQjx8gk96GmrWWZoajRc
ZglOC1XUoZt71uTCfFqsK3PUMJwTEMGP/20Czeq/F11Rl2sUiljCkTi4/Uk2DbxJ
3vzAMc4Y/YB0tY884lkIPxjbX79glYj+Rpnwjkdja6hzQ7O9lFOPySHDFZ8vFFjD
Bckwj2IXEDG3MuM8hJV6BXnTs02VmdUPO9EaH8P3etu0kN9h5Qsafn+bozQMWi2p
0CQgzsk7W2lCXmAszf0HONFK7qdF+ftn80k+7o2k5XaGczu7v+/233GjIcomoUGO
qjtebLInfT/V2e2gTVI/vFQclLz7myc3Q/iMW7TCivpIymVfi73+0jj1bJh7Ew4u
75oQesdtZrtD/Kmb+U96lDkVCTm3nfDS1NF4s0APd0WnEr2FF/7in8keXy+VRcmb
n3bxbW/HVkwZO/+ylvSZNZMtJkV7RWnV8AHyg2eBQJg0h+VXGbORmi2oBkLbQMTF
eBvI7/vneU8Z64UN9lAs0Ovl7s2M31YmVByiEKCzkAOkya7N49BofL4cs/Lxl4aN
s0fntvEKXTFbQ3W8OXhctn0H1poIfnDqwXnaZM/EwW8vCKlDzG2pnEyc+eXAmYcP
uDw4vk1/ayaqtMmqWrMiPnWDxozUDXONLlqead/gqrapxrwdG2SfMZrKmm7TWlz8
/mBtm+nNvr9fE75vIk6ns3hPdt6yd+o8ICx2tIMhgR+XOKh0VFHjHfDDmYNQKu++
REj8tqtRZMCYOpA/JtamG4cqsEJAyCnFWYo6S9EoQ/WYhamYQ5ynkttoWJhWo3vG
UlTmubP7fH2efFpmEgRk6S2Uf3YGXgfiiROUW4aVF4XLVue0HGPATqRNkkVUfMdk
qSZ4wawaGdT8t8D3TsVIETESOxXANa38lRERJVRgOqJccA1kQUFHasWzBCohw9/N
MpMrIwf7yrAL4kblKWfcEfMguX5pZCNua4tJzU/0qdWmkAgGG0f4Yyica6HUYfG4
166tFpzaMCwzZoF4R9X3nvzdogPNT8GJdTzakfQajlLQTueJLjtnYfasVS+lUHgk
+XDH4HIykLZRZEDhjWYARyTNoHx3wfXVldA4qm9Agod7m6PhY5q4dVzri4JEWuT2
akXaG5TjGvojTbuDj6fec4yEGAT49Z6eyqI28hKcErlF/BUUJgK3UPWkSIP1Niwg
W1y6Gd/euTAw9GnIEnuOol17smjNm4Ijcci4fYDPOy6ElvJHTB73pfAw1hucQ1lE
ztYcNLdSs1RO+cVKzmiLPmHx79zrtttCiqXEeGbfhIyGuRG+DnfLT6VtG3pil0sE
FQhisTNEjZvgHUNDyyfgvo5ncWoEYwdwc4lSaAU9DT8zNqAwGkeOE7QRIPOXkE3d
oI/0ejRAqYoUGaBVOc9zLH0CttGAKhlDtLe88OTMorZCkN+oRH8jw7MJDuaPdAxC
LGmKZIOsL8azG32vQmAVCzrT1nk+SAIXCecfxOkzQRpzUtrGyCzj8D27iNhJrHjj
oQs4YzNxywSMb+Iy4e6juwhLw4mSU4oCscKwu/JKyK+vgo5ernVHxL6waRXwYwgU
oTt2oJ4/8Bzl2QuprsO0ceLngevCniWEm8t3dn2f9SekOB4X6e3nVOYgAuFhWQOm
Bb/R3e0mrAXjzhM0dLs97Fgf2hmIu2q0RU8cEa3Uwfv83203IOC7votrmMMxbt4c
SVwXds2CD2XWzO6c/Vb8TePTT9jVmK2SWNC1OtqZ4mUeWFpby7bppAsfGF3TfB68
DDm4EJ+Yv/0pYoVHDloY7uj2nb5bEanL5wykLTrXQKp96s6GkqOW3N8rI3+REjCs
Wpn1cce/nQ4tzOkHAsLKXTzhISMj2YsV8rd3pWrUtAx1k80AUCjtm34QbvYGzwB1
xTaX9N82E8xz4ooVHXNOmjyM3MQtm2NYLnccSpmP9Wd7+MVeFmeQBmPLLt/FRbHi
2DqQK/smeFLHnrpMRZSuZXflBhtut4dmrVZedZdUgSCNsAG1C0C1JUyfwecf617Q
D0vFh/TSv4LYPgcqQPVl20Kf/PVU8AcdL08yAxU9ZGF3V/cm8z4Rwf9vyAHob32Y
F6kCLqBpc8gsQF/AFlAmwcNIo7dJYfKYe5JzDaytDKvmCT/PjtmVgcp9eAWXG2Dq
SzEZlfvkgfr3DYAOKCfsTM022iBLJeFyjjmVb0ZSoOyDj0oBdJCy5yjH/VO1ehDZ
CkH8gPC/5k4c2/QIe2Jj4/7ifSSOjx+XEqKb1Tp3nNIs2TG8ev5q5kuMIToSTAXT
AuVRf8195EK0H4GN1uf3LNPr5oLW2M8ZRRTE9TJETWdhxpCwOOoCAmqABkW8WOrD
CYRkJ3mpEqbD84CEPLR7whmJNebmH/O3KB89iTASn0KxhPaWx/XpRPJ00WZb6XXs
4pk11iLQqFpUwpucAwH93zR97HUGciY6fb7pd+RM9h6NqOr3E7VDhyfp4jO2inOd
gMzc5Ug0oeGxPkkHm/GSFRd5VMCBgoAy6oa/2I+M6jLpWO5By01M19fGdhQWkx9b
xq99h5y+Ml9WYG0JG0+fTR8+AaCEwq5CaNel9Yq/eDJX5HCij+onjCIM9u+l4yW6
cliflZUN8Zoj+0oxeaEV0doUzNy3WIsPn9DlAnIVG5FoOg4o0H4zIFNMwu4V4E3B
RVTruAt62iFnHuQJY7wDN72Zb01gSzAziM5tVfKVxc7vJolAOBTEeVJkwyF8Lvar
QYhtQQrQc+APz4ley6GpMElUN4o5jKcilgnlJ7mP4Nnu+PM5BEyrWGEKG41SEBBl
DGfabsc9tmRJ6vmqYUI8sQ4610XGwNwnbTKBazdr9Cu8RT9FFnLW8RLOzuOFauZY
Am9Rgg3WQfL+wbC37HeBfzwrq7LWOJ0lesPGjRYqHKrJ7ITnMczxIXYA55QBwkKR
L8gUDP7soh7hKRWxD4dYcmaepXdKlprUtfCy0n6VpY1yjFe69l09rmyDFXeQyoHR
iSwuOQCQrOzX6uz2mMBv9+e5eXxyFCxRRJqCA77Xd7grpAtHK91abtHHXZxuXhtV
JtzbCS6ScXeQ/96ZrXFfYcG7Q9vewXt5JSSr3O3hvu4NhpP1dwOYkPt0W0qH/Sq3
P8z8rOj0neyuoObF24ckIhELGH6nQuzZ/H8p3M/hO0aN5D9hlr6UVOUe4Yh24foM
L1MZE9WBHgsKMpvsDYVujOOLZddXmDzeDC6cg5EVjtU8/fLss/YDA0iXMBVW3j8M
Z1L2VJsO3xpNHpGtmm2pCMV/5Frxv22B5hVf6I2SKx4Oh627mrTo/fZT7IGa2aWS
e3rJLZVD6oQymXmwYj0SNSBi8nyzSEsgdOAIoIB164Z7bbqMrwMU8dsq2A1IJ1sr
7MoVHSKHxYNGMbgmz54fjk5joVAtrUNTuNnmJQKGiw9mAJY0lFZsFgS8Z/HoI+7x
WIO0H3O7SuJnxMDj6s+l8gKSpl1Zrer1BL6vmAgslxuTVjBXqtmRaBW3dHw/ohr7
sTjejLrOU2Yz3en4xEtO+S3igyBoCRqF+Umj6YHZRLctfg8DoQORFJis1XezDUoK
YUSPOJkZ3LFDPy8vrAT8mC12+n6BoTIVkjZvFKee01eg6QBfwyhpApwbuthCHFGz
ZK7SjmFG/L5HbeAXTKnk9xzyqFrk/DfNgEXB2gPfrr+zZk+O9r1/t/1f4pbOURK3
uNMx4NaPh/dia4yMuUu5tML4+uc1bkrLUFDzIRlWSD5m3s33iCYHxb0lpdJKP+pN
BLcnyRIVpkKs6QyX7tWAX4CuoyVOv1NH+BkpzKofQW/FBv4EgpXYvuDc17EGG7WE
7Lq58ojm34ftuAGFwg/XNxIWdipYVoTXxK6yolNqCQeW4EzYBWOeDbZOoLBjF916
9bxkkOlfnMTtofUvDqw11A4LQbSYusFwALnnaAdMpYYGL/2z0u8ysf39Ein/y+I9
DKQawO2w7uNj+093stBT0XOh1iWH1H3PDiwg+jgHftbqGMyVT398hfmO33q0B4OW
ZVXl8LMNhkQPYiNwlARkyp2jFmEtiLCDEw2YtjptAeYoxCsW08EMImIkPzgW2foD
N4WGEZKKuvXm7G6/jFPVkD6qtn2tj0bS+gFIyRaqUwkXBaDuv18aZpbuZJGqwJmi
bDLAPe6XTqObBip/4AAetO50d+o6mTx1G6/mpeCk5hkWo4zwQt5IHiaGhuO/gw9G
1JtLcG957CvvfMiipjviLeH1rg2HxXAq4sXbt3jqVjCdCrJ2AjkINsRmNzUFyZZG
gY4qzW2PYnEcdY8RnI6zA11yyZKriIxYxFrcqxVfrHvQeCWyiSlVoQ8Lgyd5ZzJP
7K4RZ0BJWcrJT7FlxhERIjfEQzSNj7BMYCDh/Z/VTKLJun5+7dsd+tNCP0b2ofQW
n0EPyROTRuUl9+a1IAEsVEzlFPcV0V7PnouU2/flgm6UKoVPMrX288B7Wpw36dXK
VV04vVHu2mdXkTwpqMhaVFTUvmVpfYBLVt0HKI+9pLPunffHHs+SkknHtB6w6Wch
+CzSbg45moqFJn6F0IiEbHi34dGYXWERpJe55OkzeCS6OFs9/jI3dg5X+SVNYBj8
knRw53JcpGTwbfLaYy71hBMqgW4ZDAbam03bcPVhImt89LJXG4xJNQE9ihnDTvqk
DcTY4p8BTGB4arTaOd04XQ8FnTTox5YjFaoFM4431B48+hRiQXufE1L6WYSZ16Dd
e/sXe7E2V4cqyXhE0QFiVH9CqATpeLfybbJmTrTEPQeahp1v5d+Pbojss7y/YCNV
hcOC0MP/z1cmNBUCI+ZH2BaTV93Vi1GLUkpgEL1H00hv+0NNRdA/Bw4We7GsA+IC
Xw9LwnY/QeNOayeW3qs/bbzMHRbMRcsw6+6VToUvO8lzmnc3/aGzEbPSIfSZijQ3
E/BfDG8GkbVEmkyaJFQJXvEVLIVem9m589//ZpxlcZN9K6lXVNzPxhgTcRj0zC8s
pbz7EYmq9sR78JgeLnWfbAMqfvEong5xuE72PE9BJLlUy9c1QuMKNUVOhIvqfe/u
NinhC85b0gT7kNDXYFpq9BJQNXxXFrHNbO9Mhn6kwU8b6yTntoa5DflSMxQ6kN76
wYVCThTww7lJSWFmLXLTzCa20+peSXqrJn4cLDDh/j2nDSZMXoxHJjiY1xUrMvsR
+Q+ZFAGL/o9Zq0EkbN9CDqrl6ahZG8kR6zz3nBhtxcbpizvVTxblRVRUiFBJYRgb
jTywX8MS1O1N6mz6C5A8ImceDRiS9QLl2UzLnixc74S6FKAzJIYZQRXzBI6spZq7
WBH35CtyWubnNQtaYovujTsDb+kcWHQDiY49j7/nP/mROgSBb/YlpoRGbNwNhfwK
yPu5c82cgrY8YXwaNmXzmK+l6XCopO5pJ+8nKeR1ktI+chS+xfjlNJxDzsMEbMwm
gvmkHbKVXCfPDvwrTngop+K6UE/kQNwDALmNBK4CcXGuB5tlT7KouZusjOvpYlTV
2inpXxtEWaqkOdy7fbcxogJbHwCDdnqwnn+8jC17GQsW+Th/8F6a9DYj91EjZDID
D5DYCQwTeAJShJYscfqBXC6o6OjrkSl6qJsgSrjRj3jYQz/mZmpzMRkpJfKGw1AF
hydn69G5Kzd/Jo9RvThI/GZpjim1dF4oE/q955t27WqHXrFLCVAGOpiVImhhKLYw
aNi7R4fA+6MxvNIp0gMmtgaI7gwJIx3Toir+LVpvc11yKnL0RWGzOs97yVCyWAU4
XXIRlaDauFAEHAqi5qWs3I3sEIcfC3ys0mrwR7y23j6yN3mGqftPCgHt3SnsFmR9
polMUPS6LreCou7/YaB5IOVM6RuQvg/bAob/GPqW8AIcH1pV6NuHq0icqd8036m7
B1Pw/eQs/b+FvwNiVU1djeOO/9vep5gLlqYc574kAa4XseED16rMJP3U0TBhBD86
OH5Yk/7S8RFjfAHg+HSFqrPwrvTncGi1vEfERdOn7pZT2uOHizQH3jGcSedjkwuw
ScDLDWLjFt5oH4joZ5cuXGMOqTE7meXwnA0zo2lUrkVheLcfGcHbBSkitEoJxiqd
IcwcLSWzkHc9Pm/Za2EQRqQ+d0Ys/0uOqtn8A+ifGyiro8MnsamjfQbg5rF3m4/A
Ik0xB35uuIl0DlYBqHKtyDrQpDBNDnj2rcsFohA/OKD5YIGuoa/Y3awOr/CKDCCT
nxZe9Qeze8uWewQ8s/wn/loD0QyffFyuW+LSR6MyP+QCon6sdIqw4p9FceC2IjYq
y1fnKQlqFWED9kxaOgZgQwL920aoGT0KPilTVaMFqYUcGWzGex+NiDloNL7POfrE
b65U4o028hH5GUt+aVgHfP/PIFR/K+aVzmVjVUVEX9ALa5LAvLDm1+Bt3aBB4guf
fo4m2BDkb4sqnFpmAxredoA/BvrpiMT7tWUc4D9k5kjY1evf8wKoTSv5jhh31ErF
MI6eZUZzXhwdMwIDTi9IkrgAvtvqDR2uZXeBRsVkXEx9QK8bJ/YXfSo/vAC9d6d6
2S3e/3c8Y4CJBmyyCyBxyvESweFIyqSRrX7nh8fU9vyLgXfERNZFpoPvTsPMNxx1
5p41YPexv65ijnznQ36Y2EcyRfKN+/J2dL7VaU70Ygg3MlL0Aa9rlV5EpZJxoLQs
hxJhUGHK8QVz6vmjzMwmCIbsptfN/davn88DKbiPpokAUZLnnAiKPPKgllYE7z0H
IRskYu9s3oTpePT1CofQI39nwJ8yRAzJGd24xGql65hHOkVLzNFvvQw5sutlvkH5
ujal+CRH5P5MS8rwC7sLhWiD3+x23EV1VMcfE6Vq7sg2pREKx8lCm+Mm+ByZjv9R
cPbkT8k089cG1DlJUrbLRQjLsbO9NmE9rdwDeDdDAqv9wKgRKMiTnTBHTKjjUT5V
H2e4GPIe/korej8FKktOQQzcqlrfcexXQqG0wT5N4sgegq17E+0OZhGuMfYriKoe
FlEihRGZUPkX9zXZDd8wPLF17Z4bL7b4dfdb7M1HKNERWtTu2pxzdyrouB3oZKwT
RlgfAMu4c9VMZi/yotmqGk7171BnplEXGQijOrRfOAE8ItXrJDPisOdDtWfMYoVw
ww5vuoxsJiJIfVLs2XOSZxzOUEN0X89RWLjZOHGkvRNi10QhjWj7mpSwFsPzS1Ix
H62JTanGmvY3J+45CMmCMmmzDxKR//NM74SQttnM444PIdi+zlp+oo1BepodAaEP
aqhzzYCUjH36tWFRR3IEkTRmnhNK0S2KNHkaC1gwnGIrDaFLdiajxwyDcMrLyebe
R1JFJBGG4kmTN/U/3AaM0URW4g29dof36BzvGPylZieHIEL377cU4HfmleicJDh2
4SZbGjkgqyLO4jqNo17fV62ykfQE/zck8av/Kpdv3cwFFBmj4DWlFflpFB8q24Ph
KArQZ9/3iE1FXeV+UurdZgCSUi4NF/o3YrA1tqNV5F6cY/I2VDeUpeec9CuEPAGD
efppGS+eg7QiYoH4qUkNaCAWQYHs7DbaVverOjCMDvfwVbLe4GINVWDsS1wuMbXv
cpWJzyGYunNcowHUf9w2Qw0cOKxVzAqTzqvRObTg9OAzrLyxnpYl1Otw/H3zjGHo
KDlScBDPSnFoTYiPndUn+O3FWlcW3Z1k0r/CyKUhBgnCQ8G9mbF+b96XobdQk2Tg
3CT8rMucVikY8QRPBDl606huL3EgCiHzp841Ym4i5me+WKggbXWlKF0mqj5dYWBq
FRA0iyuSAT5w4HfCFv4bhZe/5fxkBR6o7Ty5/dzAAeGUVA/sV3omQrt3ROeGwIrl
yz9q+h1XHuuS1N0Ua48lpQoNMZVuHFt3doaMIx/hnfywE3rjOfskgmnY2NQ0W+Fe
kU1aCiQ4qBtAQQ69rj3wUQIJTVxqJt5jMOMqRyVmNCQzqNCmW60jXgMHopUvXINg
J0zVNsdAHIkFcFa1MlehfajWa1ZUyTGQuqbOphqKlb/OIoWvfuA8Xw+AFHMJNWaU
tp6jbUYVKiyjFpY36kaid2oE/F9diKxYz4dQcpDMlEbkisOzXQ5aM2QBgyu4imAR
msuwzkHUDC1W7HP0NYIQ/MhsGirR8sshdJSs0JKYdA3ypx7UK99AD6AsK1bUSXC4
ZH7STmyJj24WUyOUle6CXOjaQi/VUiQq4XVJkb6yftKzXxazrJldanlLUfKvJnx2
xD1bX/3Uf5X/3IigRWgyNfTS8NmXvCtSvdEHhn/jQ4oF+yHMbqn3wWFVoW94yctP
U0lGADztrd1E4CZrqdiASA3jRReWRV54eCpVVQvAQuZEU2yDLzjzmMUqRkaCIPA7
Y+P5nMw0qudHg3NvQD0xeqEBoRwb/NQTC7uhBCMREkcCxyIlTrWc61S3n6RgxcWy
fnR0DwRD3AKTaYf4QmzRIZlZOLHvJNXQ+eZ5JS0/XrFnyzuJY/3wcSErTbyGvBcE
knQIKYe94tgXVzSEszb60MojjHQKuEs5bKpqtq2JRCs6SX9gsfp1a7PFJgYUovhM
LwSk25P6LvcU83UmhCNTfgSHzVwB+jsO3XtXwn3crc0IAY23HcgAIewihddC7Qvs
NAiE4LkE9yGuGk5mXU5v/EyZRYjUq4L4zwiXb/fczhuozJbgu7kzWJi1iZjIFtES
v1MHgHxTFwsOtEbnSnJunDht5g6rMiT5f4OdGdliP0qi5fpZPy+OAcM0Wo7ON+BN
OGmwEJdtcuH1J4kcokFebm0MICy2UJ7FEhb4TsrLP6Tlbg0Ugq9htyl9060kH2rf
FM4l+Zhe+sR5+PaUz3yfO8G22uUm0EehEfFdIVuqsepiJQwSSeD3h+tGxmzKL8IY
2BR7h93QfxBry4oT0kREW1SaGt6JHIWFnRnoaTpmfbQJpPat9dp8VR00R3WOXmuQ
na3Y2V35owVO5ejkE6m5+TpySqjSTLqPQMNaGsUydd+phGIgsMPS/yhwCl3rH8Xy
BeBklziwPS6vCMxwP+ww7AIIHsh6pTxfnbsgsBAtaPi2p4yYBuNf3qGa98LuKINW
TPxv/2BXZh2I+ZyRvSnj04rqT4y4pi8iFikcozYNqvKL5DMUDIln2kWvmyWlyPBP
QZKu9H1/Ccb6S30Koak0YW1KVhBpg/4nrkjWA74VCDACGjRw8MaQZmmcm/G0ELMg
RnzKXuW6IwOjD7H0iXMBHWSRsjnH9Yz6FZ3KfcqWmHeqCvEukCT4a079LZAmQns5
46DkZsxp0H6r9mzmhG3aeaZlnvO9ovAyXf02Ov/cCO4qu7rAD03Z9DdP/lAEFhyh
GaVGPc2XWVYnULVGGDA6mXG29RkjLofWrr1QoaexespDVju7Qt+oRKlb6u5+36Yi
qfjrFQ5+jd0RfQaKPkN/PZb2tDKyDZrkhwZiTnXCfPmkYidYOsm4ExxYs0GLQz0l
X4W9QIb3MqwB8QDx5i413EEcwiKqWYrGATN5TB8WYlU/M3wbE3YrAzbaupfcCxnI
Tel27JjXFs450YgWCU5wUNutz6Vac3dkHZJKrljmqVp9ffidxdDlkFfDH5u+ihQ1
PDmb+lBeww0IATBi0p5/s4WRn1moYdgmgy7l5iDGjVizGc4cWmgFAmaJ//19FcvD
9a32g6kGeTGfFkhzxGXzRFXdgHf3GWsftDA8Vz3PfDIGwpcVwR6CUtepGaChWkys
1N68y9QJa3uwx3EIPXfXq0zSsQd34dbha58x7Cd+ZiHeuH748b3je4+SAWoYB7n+
gKpiAW2uq2SqcBgUPIbQanqX5U0D76J7dTThWkbL7yZcowV2dfkwtNxYbK53ohpl
Kzl3nz+M2woEsw5nbIcE8ulIiiOeoz0ti7RV2vcZcEs883PXyHtbBtnCSBchvNJj
q4nm+a/tfScwytCUh8M1QksGt1cumKOIcF2kmuv+D0ms0Db3JOu8uWqOhef25zNJ
Op9O4a7B/LKUu9Y40N8qkPdLOL8/5zQglnqJtaaDyV6BfV5gBxX1ZYy2NuD7ktQr
Tcoi6GMbDl4r/BR8YYPcCFK3xrPqPbPSllBb5fK4YvrEvbhvHonsWIPj+EyBiWro
jTd0VOaNZ5V2l8OR46kZZNDtA4Twuo5RgtdRb+25jFVh5IMESvnhVwEVht18Vh5n
3avjeDxEezCnWcfroTKytkPIBlcTvQw/c1G2vKNejlJB9IItepWR0QWiVgcjaX3H
4PvUALWEWpwWmDHuNsd4lbTV6ORSYXYy2HWfEOv4hSMrLLRji5U8c+6PYD/yeqTe
NI832HSPPCiPBpEKI3Ky+/bFjE6stE5yQmiPicpJDUtSrwjJStDTJdFjVtfOE1GR
CUPvmxat0hbDM4vAbIkNmo3nXGqjAcyFgs4+Q9ozqnkG1THguTzqhVZGdRHsQCIU
S+Y8Wn/0xgHZX0zdQkhUjiid0+fIugGqTrbnrHveL44q88GKHgq1qeXgJ2kXChtv
+vDYSHdliWeDLsXY0Cme3s0IH8mKvdVR/WAJfOf77l7TdT2Fps/n7z04HfRyh1pg
8ovGjzvFPps/KVF7NePkwcPo6t5+VvnYI7UeJo3Jf4BiDmfXYx8j57ypyRqOgttb
/fResIRHuoZHJ+7QfxXw7tneGQaZe1q69xpX78wkg1yaexXyYuc4gnMZutY8EXgy
WcibXSLKx3ebGfkT+uKjX8cQmb2YVLfdttwMCyxvh5HHslDFVcxYjplnpt0w4BE7
qj+ANspR9q5dytxZpytfCNd/pavfE3kUZMvg+Gx6nrZxca/pnuj3D+4jIVzxZPFy
uuuWZPFqrJUOGvTtFFKC/Q0LcXLTgm8+tJnJ8h4qHrYy7KKfbuzyjc+QOnkn0EZ+
6hj9W/swqZkJsdOkmA038FGAFmntCyXJm2ZEg2I+OQetidn9geDOU0HagQRniTNZ
+5uxPeXlXePxRT1+ZW1UotC/vxPHWjrtTuEGDY0rMSCqab0G73QNrX96p1G6z8uq
Nl+A+fgXE4ToqVroqN6IRaQtR6yfnpprBwr6187GIZu5pjjivbqBbjFBp7uwE9iO
g8PQaeJigX+rs9LSl16wTjTqvtZb8w3ZbYNIRQoAh7//veMJR+5rhjUJT0YVDcZ6
guntb8yhNRjoZ52VB6sehDcdQdPYFhHXxGww4sUYTQqm8b/e/ehSC5Tev2kg/IEF
z8bX+H4AtJ+BiUj9lNlGGXV3uB/w7DaCLYarmdiA/rCWxOa/59OWrPcNcIUwj4+c
oCkzFIv1mc/TUfwnlgVnLyJQAEH82YTfrMVcu/suX0GkW2X8hy9E6As1F1AZsKN3
pGthTGlmHMOM5rdjUOceABzSOFPxx1lEBv9nSEEZ2SLJTLVImskamP2GzRVKvW+7
pQBFtSNfJXpDDu/4QiU6e1vgCM1L8fY5SWoDC9OX7Re5AHzwrrSb9desUpAKDWK4
lN7DKtj6m1w/1qmlf0hCXyRckVudLzqPHiueoF7IsjU8B5r0XsCb6CX33OxzEWYW
08O5dhkbq+QBLu7iXPmsuI33SwtXTEPYKi+Dj6eydUqsz312c7kSiw/R99i7VTgd
NmZTigP8Cf44+V3sOf0QJ1xoncr4tgmRkI7pvadGgRXlfSiXBNTNkPW1IwsLZNfu
f3TCjv2RutzHEGGLpFRVha8b/LOKEq8pbJON7hWPSYNqWJxjvDXBm3DKfIA5LCUq
R0KdUGYaAMXnTnKm7LNnt3rn6u6Qn3phYTTYvCYfwm+vG4edqksHD19GG942bCqA
dxVIZW7KbpA7pM7w1jTJIcIW6S5B5GHdGiG0QkkShKDD5gylGhdwTq6UIRUu8+IT
koUSUOuy0BSRwwPMAyF9tdOddYO22SfPAddJeINRkiudqehAAiEautuMw1wXSasQ
0G+0Ya9juWmDn8eSTh10hZtpYb6CVzRoXeHBHMvXnzRXLdruYH64VJFXDY9qDI+8
DspHETscJt1Ok2gOFX11oVOV+ld3aTKWptlSb2lXJg1IjjuF/ZxabCNDR3JOniL5
tTPOhoDxbdYbqI1eH/2txQePGBJ0WFZXdMVIp1/cQUjBvOLjtIwuyBxNSQiAI2jk
OMa6P27C26HFmEQHxFowsdJ91gKPPEGyRwq1Mx6l5OWA5kGp0YFaVC8I/PEamRJ8
W4KyKkgxUIv4BHfmkVNBCJ7ytyhVpeU+O47PXgOaLeOI3Alec260L3Uy+lIsmkQy
QfV57Q6J2G+umXNwAulAceVSMQGm86/1VSk3IZaypt+Nz0ViychpGtAZaWJ9dOWk
3K6k+2myoHeXmk5jNVwNg98LSjTlnjXME+6JNbE1TyFFkVwrklVsPd8NC+pyC3Ic
JH5YWA2Q0c5YlBsSmMBw55Xyxwwyl+aHQ8yyrWcj/+WAR7/7XENHE/qq7hBIPqqE
eWJAys9NXnlG9vxGJN0N1nqJ284JqA51+6zunLQq9JIEanm7Y9bYV6+yj79rkeb5
wpovnmkNbVH0pl0vFstxJPGs4F2bY712rN4ihBOk40HUH62UOSm3/iFSEq01bUOM
TMVjBNiGndXpo7QGzeKTwWq/SknET+mKLNJrYhMO4S+RwufuYcvgAiz6msT5S69E
h9aRrUN+oBgZPE84Kxyh4iSISy467kT8/kMYxrBFmezwerX/nAZkqYSTdEI9flMj
bA+ZPiaSJJ5H5OF0J3Ba9f/5OllyCkhqo4i1cODddlqekK/kLeKuxYJxOT/GgtBp
tgpMd682Csf3R6sZ5onJ0xOz4GQlCuNIu/3Ql8ft2kGFwrGz9/u0NV+4OI+zvFEF
SMIL61JJjD0RxLLdGH+fBCPWNpSvy3DGRDqDU8UG1T5DBXdx3A5HEiSNk3J21sHp
/v1nGX3Nbp6u5dAuQl0c5VJiJDnFg2itG3EZrkqZaXYwnxcIvh8K+4l++uXT6q5c
wDheABvXEOBeGTXDgvyPfY0LcopixYxQ5ld8VXPdqLB68A5Qm+Rap6KFbucfW0zN
GF/SLVOXpeiCY41OpEFIK9AHKHZYhKSUFLRiU6NPPqQPuUgDHIrrWQU8PN3qLakh
uO0YQoptLgHf7d5JBnRG3IdlUlGNvMi1tPV/iGP028MJM8+Y+6nP0e/LnPyM94JA
v4nZ+Fqw6VYvBjVfvKdbJL8aFHvlwdOxMNUrWUxRKPUcp2zr9ev0+50hw52a74iY
R5z97Rs51Z/rVxhwncX4erm1rnD5Tfmfq5aArmgGDahUIVs53wjYibyfL8VuPQgK
MDr7ZGom3fuownG3pmfGmFS9yiXyF++HFlUsjJFaFbcrDeqLG8h0lWHTBBF3vGrp
kHGvQMZAsWJm5B1QE9S9ERkOe3kpI64oTybXdDuVUcw9X1HFJBUwNr5QlKfMKhFY
HNRMgvcCmuGd1OKOht0d1/nCdj0ZHvfrBYBXKiCxDoHlVr44HzmOw+K8ydS5fmNw
2eQgEJvUFfv/K3pVN7gSMgzPuMH6rXhxzDLM16Y3acUdNIO1lRqtCR1CcpuPfRT4
qKafLiZFo17EworaEy8TKt0zq65csGw8KpB3T2dg2Zh6+BrCpju/T1NCeAsXFgMd
zTtzOxIl/WHdyHeNA03QJ2p4/Mlt8ItT+LfkSHVDy3VFwdmy2beZ8C1eIeb3dhPA
hYs0KwJneQha4ZHBdfj/zWHnfJL3Hh0VU8rqceUU0+90gzcbWB6mE2rC9b+W3ft9
9UiEGiTMad8D5eiZAEmo7IwmmIIgSZi45Xz6kZcT2jNBYstH5V39PtM4vYCgPFWu
nVxpicj9taemObOWdfj9v6/aQrUV9HKoADy/iGUPbF07FRxhDcD+bvY1qwo6QR+z
U7V73ZPPDWFVO5DwM9HJooxhjnQVebVHthaTGidBP8L9mH5WWhnuUrU4M6IPtDI7
0i2WnQxnN1Te2tEPrHLkpv4fom3BlyQmy7zHCnzzVsrsGmYy/EtqcLQb56629u3L
Tu0+yIHdPKA9AMxaljux+tB7FTPmN2JL4F8AUVWeTGymoqnmmb49KzJvo/goK22u
xS40WFenFheukzmXew0vueGuQ095GjSIyGmS73hDr1Qimw+tB5MtQsr7zb5ZyVf8
tYQ0I0gGuYiv6sd39ZNdn0uh1bn6Yvgh5jn97Sh5VRwfapSyOuP31YwD8o85sFIt
PDQkHeE23vN5kjb3hFizuGX6mSNku+GSivNGDXYHW/pQMVccXKck1RM42WFb6E+x
hlYswGaI2/uVmhhvuVIXEUttiQhv6x3d4ucIcyJp81t4aywcb10xyZ49LfptS+Vc
Oi55wdNPsctL3rV/yV0Ia+CZ6bufMakuCbJzESuKQgUNH4zYV9CJC++G5vYlDVfH
/A2Chxt+msGarp6ehuWx5Xg+wmT6JnEtUN8rPJon420Y9reinnIpT2z0z7Eyd5Qg
uf+ZE284MlS85orTfcttlhiSfHNP65qMJx44YnHOjXEqrk5FNAQAaofpMZNFGcd7
GMa4o/te4LKydTtci28WMbQwMUeDPXY7LVvdi3wrPDQ4w6OCgk27sDFHzcQPje8s
IgjIJd0PMFK0N1HMbqwUQus4uoJLi0oKtKm8NIvALfscs0Ant/JVQu7IlKkxAXi0
316s62csI3djQhTs8roT0HTSq5LcwLXhRJuBRiSiMwYVffi1fY0SVAJCk8Y5OGY6
bnriTFsw41hxt2ETHIMp/hLEpTsRdakAr5z9TOxYyRk/qODBuRYSdrW6D3UNoX6K
f/ZCu0uoP8y9BWPWk9p9gHJo05h2XypVamZoo8LKUXBnRdRB11nVXFcCht18TqME
YoBzUI+vs9mMMhP/bJoX3TVMwQ+58s5/dli5mqrVG747XwjjVIn7vb7OhKuG6Z+8
TlCTozx+gHCLU+4DuMch0bu/cSPyvB8kzg+wSeQ+xYNo/n6QupskI1UIjC6NVfkH
lnyCzcCdSpUYFv+tG3NKoZFfpvAbEQQ+sUHo7l7IWK0qU36gCxZ4PkNewFDNSFqW
z6TvA9FZ5wggjnFRy21+E/fb148szQDGcqzNBUp29VbIH4ARb0ubk1I3f9UtJDd+
cW8g7Ifv2Ztp85Jdj4CmZIY4pVhNRKsppr+H1ZDDVn5Q70QQdx6EHB3Z+PlwiyOk
fK832BG1/2NME33nTgyrWD6kX2CL0+yWTHec8KzdRc3wPm87zLrRVkM04Yqvr4qZ
8LGkbJekCeWtWZnAE7jguGqogmF7irHW5rnuyAv2ngTEJv7QzsM2gG6djb88wvTT
l1o77B54lH4pARqi7PiKGzlupFIZSWEwqlhdUna89vX1o8rObQ8L12+0YpzyiVpG
MzTYvrURWZvieg76SxhRn7XE0LRkFyu8G4HcPkKjMEV3XDrLABFDDx/Ob7/62e8K
CNRR+Y26uhSnjlUhV13QaNd0lKP92JK2TiQGAHAf7ReaGnXE4nWKUs4EMzqD6TJr
YTbJ2ZO93JPBsJDvIa8cHQlbBntI6RXQFgMDX8qPZb16kDOykthv7qC/7V6xhJeL
qpUgRQ8UWHeYybn6ktYZpcTuNKlIQ09XRctbr5Z2rJsDsaoYofL2oq9EkLMabvM7
7yC7ern3lhZi/qaKpxBJzb6fYsxZgg0mX1HDN0ldqG42CHsO/z67t4p8O6XW/ihp
CtwYOCEvfFbAGe+Z2jAI2nHM5UQQuDJk6gN0U/sTvQ4Y08MjACYPqoTuUwamm+/l
yyznwK2PfpYN9tNOrbSg67IoYH/ctyhYZ+g2PjGCRWtnS89RBo8DrjLZoLcEZuD/
sGVCYyQrGk6sZ5WMJsNIqA1uLCYsr6roO+mgGSui0a0xQIiMbkmP4BYI35cafGtn
pHVU5LeeKrvVDMn/+WwsbfLCBBNvKvNgwj+2EOlBW0O7dYvWwGTS6sCVg8y09V4X
eGNvKYHIORAEAXWPmSmnCZeeIj2KcvcMliNIdoh1gSOnmaVjK+D4Mz+gm8HB3YFJ
IGOBNVLfE2igtIjNp+dkeebZEryhAn9nEvgwb0s3DItVtIjJSWpWSdwVDCKQSg5d
MZAZMezrUM5RrKuFH6Hjqd4lbjCemsVoYh794w2T76BpOAp9yApINuEdNORNdZw8
mmhsfGydfYHLLC67fgN9OQpt219ygB3By5yzPQyYA7YbKmpqDVBFVYgKJ8bx7F6A
dmxMuVJd/XyRzfyr/3RquWdINdNWxlpT+n3VTzxhV6X/lTxPeZJ3Xxt/br26hCyT
wxpVTM0KGOdKWVPj1bzLe1d8HSzylszXtPwG/LWo4EmGCZ26WqGCWYVdRf7xOPZl
hlTWYUD8pycnvbzI1WwEaarzuOG6yzQvfWOey8rnPUKGHa5KHhMXgaRz9XGVuzIh
rjwN/VLFFSG2EOy9qbPo9XlxZQi2Jv3cLdQQwryLsaCg4mPTFtGr63U4b+VDlHuw
Tx2D2HzdekIf290j/K9toeZE+/3G/gnpS/53XaLn+V3LkDufMsV+r2yqOjE5mLhg
tLYDWx9zc6mNirBbXpUQbS9mTG11MTr2gjTnSJpnH/40wIPUpgiGE7bA8i9J8gIm
lS1xOdc8bcroxHd6Nzd1fm7qngBqiKGXtL1z03HlLkXwS1mQuojbVcAsCqTcwJeG
2KtaQv20RcHnzP5nsjLgMVLtbfy0Zox+aM/YQc9UaOMedbVkdiL8osaaMdxQIRv6
GV5+jWotUhheHKboY2Y/Bsd5IW/jwDA3eYOllimwPrNX9IcPWXp6p55uv6OI0n/P
/cT+W2ar1o1rf/flfkkKKFF/AvLQ9ww07SVSfXVlfr7kEH2ujZ7oI1MomkU4rJtt
10XIGw+PEaRwGasCqrNQ1DjdEK+VmhB3aeIw8mvE+mL9RInLe3Cf82oTW5yEU2Ev
uPaa2KOV+ml8l9cyyTTmtm3L8RSnRe4xcX1HHN6UAstplHB5gkCeWGu69P07eJW9
tEqbSPozvqT3DGBn6pTQA25agOJLTuCTXom2mUuy2h1RGsymJtBgMKah29j+SGpe
DJfiqUvEYDPiAobcKuyyg8JCGAGKTShCNx+oTGRpYImilgiv3KoqbxAc4ihlZ0hP
HDdUL0M3wwjgr84c70G5/CgPba5m5oS+4eNybqBXDmcbg6GTW2CpDljvABWhRNQR
Oe49rrj9YRQVeCmr235hL/WPeCnm6iE8/ZBy3Ch84NpkPqYM2a2LRjvbFU5r2cNC
9V09f/hicJmwZCqyEYbg6gFPurt9lVtJrq2wKxHRrBqeBG4aNpLb3wWA6mpewh7/
wfiziX3bsqT6weQ5ligeMbCRKxwOvmqEACAtbCaz/m9XW3ACo21cssA/WcnBKX0M
LX3TRWylTp3gQicZmZ8mKagPZpPIqaHkBSEcRgLn2eF3JA6MCUsDb3WapP8tm0AU
hB0EEFd/QUjxtVmwo/CalVCz8bedEOLL8s+BjYecqiIX7XbbmGwsJEXrw2bTxZ9s
5jdsgvKIZcGMsJvGOS/rpxDfnVwPoT3luIxGfU+6i4DV5Y4jbvudz5+Iv21ettBf
6ddAEISpHRmTQCpmzQKiZHg6LQTJonVO14jumKjcfEPuYi+YZabooYV/ATCM4pAi
f0+UZJgINDNWvEs8apWWqf7+5FOcQ2HaRUKOquE4SQAu210GD+gClPq/CVaC8W0V
SKCYXlbcuKtXJOqpbkMWw2/IEGint3PyEqvGidBf9T747tzpNzOZ4zfdBpain824
YOdWvgQ0okT5R1jkKqwUIo83HLBX6vFV8z/MLw25WAFOjsuwxqs4azpWIXvBmhpG
4Nv52tNCzz3BEsybJYUQtytTK/tL11rK0oLHZf0nhp5Ruqz+x1/3FDC88wMBwTRW
hSxxksKDrD8BTKZY3ohHlmmvYy2KTMzY9xjNU/kv+x6tebfHfd1td9UuiXcdXP/m
GivYNcVjAptld9Z3us2f4H7j/y5Mnj6/LXlseRvt1vhGYiLy1VXweHzgND+l/MaR
owsEd1CHkJY3WsLbCSbFfBzXfG4pWBm1MWw25fA8QWnM+C2fhPWTHhAcNvgMovvG
TeWy4ITwp/EZIXu/+r6HxsyZfJPNeVB5+2DTf+fYschrY7d7MAwPpMULvdFnUYLj
ow8JuZ39OQde6wBACx/uH9GXkfk9plxbJus9MUlYkIDAsxBd2EMnQA0s9SH+F6aE
bPM+9HBOMo+O2ZPjl6IK4bguqRwSm4rIByHpJsSi5Ldfl++qtUc7j5GsAuGUdnvZ
KizzuNxC3HX5MMvfGqm+Juph1V+obTWp8VxhIAzGGxpqpFqF4EKlJtNRJ5iPUe7V
MpJiHt++Ro+DJGo0BU4fStp/5zPJKRkkvRk0fytLcG95sodb8LJwptBHXhVqHPbm
mejhLKFxy/Ee1R98JLSUJs3ZFTy/rb61wC395G6R5CI1pVNBF0pf9x0MpZlDc6i3
vgFdYda10sNTOkkAv4VJzMS9PUFYTWK5g5yWXmDSUwNokXXGYoHQ1iSAquBSbJU9
Tw46tT0zM6HmOb02tImdvNaXY9X/YJUleLLzWOjshecCXVGf+XdqnHKIJMKztPwV
ijplNHV7kAqsx40WVt0jQlC4XwF0RfQ8zMDzLF9hTf1zl7NAUdQSf8SqjNUkhvVz
l9YVS3SEw5qxLXONYHqf57GuWNHETQA+8tEK3RAFnTAo8aCsSoMFPskB2kBxuo8G
KuTMIHzrZWy4IxMYns1qITkUEWCUw56/rpqbO7wJbB7R4wR6TboxykEsTJzzGk/M
FCVzN6dptYmXW+434IowpmaWQLFMlT308K8a4PSs2VftmOa26LxR093x7JT5vkco
wOHE6edYquBNHuufyr5aXkLnrGH3C8d6MvMfxAGVLGS1fsjub1oPm81hIfoGt+DS
AybjOMKVncYGSoiw9WsR7bs1Uiyrfr3Kvu6UmHZWWTCpfs/STYoeRTpyR6Q05BMu
pQtBpEDpYJFQ1gvtx4yUSrWDu7SuAXupte19MiBHESGEr1QJdin9oYPf3E1z/hOD
IWfdx4GOei0fWB6AlQhj5/BbXuBhtrRVTQIhrgaOzUBBP+sqsqiN3CsJOWZlqLp3
fxI/VgVuu6I4K9DU4pd58UySF2kv5y7sAb5UBrocaf+nqZ1DEp/1Dq/ZcaolwDR3
3MopEJ+pn9cQkOkZqhqEd1V7fZrrtR3izV//jG30nLzanK6RXOS05s9LO9qFOEcb
JFOvIjmMYlt4uFYaFWm2jSpFgaDX+4rXcl4ehHkFf7fMRRgKLHcBJLv5LhBgvpG9
C4wvzidzgSugegnt5dkIciGvoZVQzWZPy70GW0UWH1afcKtD0lBHzEXc8v8aECN0
s7E4nxkg8e3P1V4QL4Gkf0NuDLmShoqV5+w5N9z3uFTOTuLT1updGEZAt85uqWYt
AmZkh8lCb8cu5mjMdbibu4Gj5wXwat1EfM+umULM/1UqGCuxkKV4s22v1AQLZikm
Wd4NEz2Su83EagFPnZ1Fj4MRqCtTqh/TWEeWHv/qsoiD47+8kkPe5s1B/oXTyApg
pWX0T+ykGv1wAilLrmZeq7MWtmx88BdVu44AOExHov7vOFTbjuwfujGSRRylOzrA
fn22+bqLmsjPsRD6Bbfnr8kPEDOUNG19JMfeu560Ou2S5pY5zXcGAH/PDKsvRB5G
XRiJrZ2RGSFIbAUbTE9CjNZns4Z9H/8FDOhpi30AdIxHaeQlNGELcEY/rSUpoUrJ
x2reTDQV93oWk99+b+bL5HqdoDCNEzKfeeNVsUiozbgCmawNjQbRsobOsrlq2q03
z/Rfh1EsO5f3roZPyLomTqI7WoJ3sOxqbPA81VOv9L7ZbAxPnukj6parNthqRmRS
C1qfCtG2/B4zfIDjR6CC1JRpBY842YtMk1d0gvtipoSfO2UCePi2TvunBm5B/vzS
NIDK7/vxDC6ltfE9+jZhvXkaKucCogpKs04vrqKTrobW+rQSms6pBy5WV3/dIrHA
TirLrXlW/l7HkBI+4C0yBp+1yd20RRkiS5a0srWin4JVnS6KRFUIuYZxZwDhXRkr
f/phcpdby11o2gqfXMfZ8SqsR5EX54KqsrxUae5tufPOEUFQZvr9WQ/TkvUkyV1B
PqGTmfDiuh5TJmXEvMyiNLxmZwSwNYkOaI+xCHJqmDjmpEeOpEfaZF7PBQHGhBDD
yyjdBFmszsL/z4JV9ck4e0x2KGHiXwVqoMQlYFusDuvJAKxbUDppJ+n1/y2bIqxj
KXOkS6WgGATYMJcl2SYmQLuuGqxQsYqobPJMWB7ylmXQnwBqPp5tnQPJUac168+W
IZOxtsXrnt438DiVdAscxvLXnwDC0M1uzbf+xXBoBxwQ9TBSlPYC4NeWyV3FFW50
cjfPi9qPz4zv85o8eyG2kQEQgTm3d/M9dna8SEZmCMecA4cq/4aXWwRqQyOS6Wex
3esOmCR3XjbBfUISsUSXihP9LCPr2EbpUkt6UJmpfxoCDrXIbMGCn6OhJp7WXalY
NpZcmz2g+JYhfROnGtZiV+C5inVpmNa4jB3hNl/3Pcf0/HJvj0ksXCzhjlZTiO7I
L/E8KFU9l8cKJYrHVu7twG/AfgB+I6+kODzERJUDTvzn+vw99DBxYh9U0L9wIl6R
0DeO983Hmem/qOTRRj4xC8qtbGZBn1xnleCWMKWIG1KPdhrGaac1JGvnNz8aJ246
+uKoEfrw1mjwGe1xxh8lcIGDIsHRbaTW3Lqk+WxD0D3oAGAFvQ7dhJTcJSVzj/em
1Y1e/l04Qc50UwHidlbeaafiUTSCRRLdJ11SzrJK073s5DPRMEKwz+MFcuN646bL
5fPZVdGOS8EZ4FukAPx8qrYz+YNI2eLR0szEz6gFlFQGFkN1gS6iTfrcZNpc6IiS
Q99av0FR3L9aPnTocY5oJPTMRfCVmUfuh4y1mVlqLXy+oupKrAg3kISqNE5R1uig
/M89uXDnfXf8PTL5Nu5FG/p8LPaeqEzgtA+ncryjXO01luRmNtdus0IzzieIRBTv
XvZRj1EYIHnDsRF5QSCBAbaPQogvhE58yiVpwfLLFun6tQEykDvyJ4zZU91xWyVp
KxVSyIdCOSOn4/1HH663wg/bC3qk7TnvCW31SdNYKyM4LesQGdq7DayNkeiLXr4n
hOYk6XTKBsTFrh2nK35hzASoAfDPvtJkLG4pgVrVCRAe5/y/JZSLS+b6sJ7hTQPT
/SldFdaaOeHkdaJaL2FL+z51Gu7JJiJDHeZNwKh6gpE2x3zeLtzHlB8BgaLRSVga
APsHgpBMJ8TbnM04OMF0wVDVzItRZjecx3tBnRTjKet/oJHvPPGwe2AOM9F9A6Wb
hTUfgdB+OqW4p/yvxPjSIrFt1OaWdOepa7pPAcvR74wjpOLENI7zozhs6j50rcZS
VzImEN/IkFonAucI54XUO7QmzmVWJgmDttYzVs4K5lyZUsvRjJKpBZLBwbCqABg+
q3jAnmJX+lXJqCd3qbg+bG4871lsiMlStOLhmh3KzmwcaBo2KxUvNbS3opCEX06D
XqhUoVPySZaMQgvsEqZEIUsKcXFk+WXIz9hL1TVxYsGg5rf/ikZwBELoFBvNdwx8
jNEqh6OeND4vEQoqsUciBj6AVjBBKgpqzgD5p19lnkcDU3Xv7y37gwNxw7C4DqiR
taLWbURfAB/HwlrIK9DGBcJqIB8br4sTTzT6N1YWteos1HukP3iHFtkuRE556Sam
LYRW3bsbcTAmldkWpVaLpn/RcDvEEN3vwb5IrzoCciTuBvemlTGdeK9r4SKRBHVB
pdsS+JZ+nhpsDYuiGiTalHXVcfOXbAtqPFQnnUf/u1ys8vg8hZL5lHDfk9cvWJuL
+QgWVFStch5u1GR5sVVS0WVuV1Qe+3VKW20+/QQnCbuJMt4q1m4iISr/rZO8CNgF
fteZeSPrXO+pO+8p+qEypYij6XQqVMB8jCEydI0xSSNyy1ITMMq8R7Dw0Krw2vEn
dgLSDWvllokHtJ+x+puAA7Y04CcWZdz9I17NJ8RHiG8mIljbZgqYHvtp959o1GUF
sK3HTEUwd+tw6SHw1SQFp0P74efWTppulbN8h0UkyHI3dNfV0uQVPWsETgJUQNuc
V8cY8tH1pylH6FzdJL9RLOyTas1uvcjJGiFY0QyDDX9eqKzQ5cnE/CD00yxan+F/
fv6Rk+ic9TZj1zPwpejuuqL1ZDK65fbwDz5t0D2bP/990nCmFXnFi1q13Vr3LnAz
Z6NXGneux/zOWfab25dOqZMKsmbmb8ufhf2oe5dC9QPJCu+4/XB04VMSYTkoZTeR
kZ4x3LcG/vlW4NY94TH1VFfpYHWJs5AoQrNjQvBpY2rvVeW/Nsk6auIWNMUylOq/
BRSedkfq8BTJPG3jw/WMScFrJdmE6j4ajzbtMfoc0CjTAmOXXuZDreVuOjKQtyW8
aJpG9a5aNh1Xa3x0cKBQ0acSeQk/9Uxg16GWOYGpv1gcb3mF09uVVagycjbU9IJu
XYIbWeDQK9SjF2yiR8nnfqiHlywMSFwdmEDsSs0rJmxAO7aF02fRTXN8nFQRbjsF
9ZYDNb964+79dtiWfo65UFdjkQ74bvn92AO4KUWYxkOkp5FkYAWEYZdLjgmJ8Dap
ePUpVmTdvZ/YXThJsk1EiX7U/vB8kJY2jPsXBY6cl++B8/2sTOLjQCZE8AZgK8HM
pxPluZBtL4TR0cV3nimJ4YMr+LOw8lttfDDndIoD/WLiTi8zpb0lWXr+mI1Adonj
GEK7ajZ+pCZqI1W+8Z66FdPOZysNiu7GANzeR1U0c86j/P7kXTlOR62yzMB4+l0c
f5WJubNqs6pNdU6wbXRnsNJ6SU+0+VJa3rIQi+Wum4+NWpskyR1ylxzsbXjHuNZ2
Ahb09fZ4dt7YsJLGQX4qqlHObGlHZdrhAJujl7yGN6VrHeyl80L2VgafdcrGZzxk
5BGWL5RmvYiNns43Ssahevk+tLWiZ9gFgPP5D3BfNDwlz7vpTrzmp6gwQn65lrFg
oR+17xHiXPjaaT57hPJOKQszmVwSsEsHuAYcBuhSVcNjR5Hx2yr194okV/QnumAO
kDi9mgo0dXwlDU6968BgX2g0dYrA4jGbD3VrTABQjjE2nS8z/S1LnwI00b6iElde
hYLn4fseDw/CrWan2DHc3GB8TgzVK7OmtnA/Zt8PQHQju5yG3cwTpJS2NWixmyja
JBFjp4lLONC8NKqbS4UKo/rvReWmEZ3f7Vlg4CoLRcVChH0pDx1UMMR6dkAUzpIe
vj09qB1NNi5tv6PU3MnLNevWbadSS3vErc80/SUnpPIF3bTC1lBDAkAgfK9hOfEM
1bOJvxJQQmLLNKb67lSXdhn/ktr3ZW2BlEy90D6j/r6/8zK+lwq/odLkIR1aUAQC
QQAtsKzbOWTK5g69T2qmeLLZ3CY0DZKE2EzogffOnmjMb03LeaQBnvjbhZtXVKnQ
6HvEpD+PttSFUCBW8G4OwvJr+iqYWovJMLKppKfIR/EKzM+yWUIY7RKv01Jcqzs5
sUjDBm0b3XFTCZx40THVAaegLyEOy5So0T8Y86ZzDoWRsMZT8vWQud2KxlpFPqc3
ARLRoLOIpU+I0W7tO3BODqVNXYvFsElQT/Ig1UXkrIGQ5i+iDCv8a+M4rsyWjykx
4ncmKtL5wjTiBiX4RER1j/rNqDdFovIdqgu8li1+m8gCDMrSVY1nTEJe9KGAkC9p
II6xqdbIRMG/Es0ANAm9q+snJNtz3LQa9a1givfOuJgvddpolMSqq25VMA7RqVYv
2HT8UsbYF7QfngvB6sU8jfv/L2imy2kbdFoidtOBhjG5O7rsF6BiI64LhnbIztdm
6P6mwosD5HKFF0ea7j1jvcxx5LlUmRoVjD8zLKXHYSxiPeS/UPlHaJ+DbvCyMmpQ
n/Q8q3g0p3g70Bix8DfphFuNLBxTFXp4cenuL70zmk3XZZ7qbguWoxynqv7UjaNC
/178gZSN7OTn3tK6RU31mjz7c21wkdcvPUSTJR2j05E8joP1UfyMeG+TF3DuH3fJ
mJyy+mUTxBBvKBOzqvAmZR4TEf2G9rBG/VOtCXmJl4yaLq9RBfTVwVplBEdBN7h+
3i9a4dn44VvgGlSFiEhIu/rJ6JIOKamxcwm+DpxwpvZwjHSqvjOddKUMlHqi7WZx
JMl/DCIv+4zB59NHXje+1yCbAketo4JvECZ0Iu6DX7HQ7XkjN0VS2gtnT591WRUC
NihI6E+0+jZBEBQDxVNIJBg2ErwABBuvmLIBgszroyhwo8cqw5AcvHxdvXfvQDev
9HpLMdrg1V+gV4oNc0IYZFlz8AH3la9wfuyV2j2vQv9e3gNrAvRFO0ox3qunRsEh
URJxikAiw9coQE0tX2up7qm4j96P60b1iQvn7KJ+p1uTw0DhUnmD58DVVodhFaX7
LGD/VM91xkCW3Qrx3iG+uZabkJi7HYk5vhQKZ+2/xVBpU/9kcZa5PfEmRqdFxBaX
pBk8AhMmAq3Ue2cWU1sBvk0ZsK6SuAyHc9uV7tMxplphM5+yORXsw6IzRuA264J5
rpBL6u6sMTrxKYviT6n3qnZ5rrdqKDdLnvkq7irSAVJVEXrHJqLhYODCNqOLXPgO
66Dk4/uArStVhUWN6tn18La2gDUwsSfEQdFWGDlFPISW7FlG8UcJWBNI3AlNev+/
yQ1FsTZMSWjaUM4VRK4M9wl2DfTW1xSau4x+Yv1nqM3jPNVF/aq7BIWF10kQcHMN
DCQ8iapT3UeXLmPdGd6EDsL0eNbfsgnVIiyv7pk5YObihG7WoPVUZxbo13sAYV6W
Jb4mBcJdY9xvNc/CYqgScIlvzVmbo2H/zZLHR9Sq6vMV66BZ++jUVO9XZf8OCUm+
qtlh4ltnlv5z5vDpUw5HzWoW7ukekumwRU6i+M+wR4M7tFLepK3KdYHZu2yFzB0f
50avQg4tP1JFR1C8vERNfkAVTrvJCM+9fzWqnWQJrlDMcnsjYrVFcqLmn05Y5jbs
9BXVdGW4H9a+ah62iHnCQVQA92YeKNu9g61N8yGI9r6v9lPQsZQG4/O4y5vmoqRc
5fw4fMC4cgkzgLj057HsWqk/q3YMpq0EYA7KfO5t3KILZ2jseMFjawf1EvPKctai
9lW7qyUMyk5GkHKNGm8LXaoBOXqwgGSNquCMHXjrYj7Hsb99uVDBaW5u+liKrmrT
3kRkb96IrKT8cxkso1rdIvtxLZRUmTy3ymICp4vJsA5DtL8HH7T6qKN5zA76MGiR
fwinHCZ5CLTy/5ACNnTzleuCwaY3BEtpXeDU752AStwo18/I24TMpNxi8GXB/puW
YbC6Y5rjFwjfRH1DO0JJG7u4zXLcylkP358KLKxLQBghl3GOLyOS0yGZUZokip2b
jEHb1bXGrzyQOwp2o/kIcgaFS9iT1zqDyrLF19NmPg9zt9UJqD5G3KuQQYM6Colx
/kOGswMBBToF1lOz7coY76j7Zglw4K+TRCgFcAwWOQAvBrh7dY393cNC7V77hUZb
NWz1Y3LyaHZ0c34nB/fKRVs+jxOrUX0Qyj7IiRLhqfSlSIL0kPgl1882YTHq4ZIW
2c++6uYOn2zf3Hn0tj+5zQME7fC7sp87bWYZU4qrm6MndmSxmwapGfY3eqVD+90Z
IdC65a1yJqQNmraYj2DD7rmOzcvpAJKox7aoDZvEtgTMAiMtiMTDOKC37S57iAhr
UxHu7BEy7wtwMnONvtummMJWBOD6MCjjR7Q32Cg8xbteBiYuWZQ+TcvDnHUF6rEz
utGDytKVuYRhs1iYuc/XHbZOvvsbZR4A4Pe0V15G7TM+uKntWl5ByUQo3RLq/ijh
P3wTm5K4/atIi81Fiq691S5nG/PqGuOczIBvZ0aSjpEGbWNdYg0+mRLpoRClfj+7
COIbnWvWRnKuCAdYdLHDVi7vODofofctpWtiUbublgSr5a2cTHKFaPIT61J+adW9
dPWh65infok2RmGX87TCCqSmn2ahOYeJRqGPRRjeZUAqWFXNFlrQLhx6ctfKmNYm
HSGxT1CcyrIiO5GjkDIWb0cJ0OmdY99vnXYfwpm/kg+iHbi3YNz6S5XRay6u+Q45
qGjKnAEnuJHgYU7SkjyqE3vEdfPSWsS1FT6ectvb7A7kU2bx2ih/1OkrNg+beGWV
M8Xkj9yU5tQ2qmbyLNMLqwVR/oQP1v1Sf9Eg//IxkL7laGXpyJOj6LXxDZFpiXah
Y5NKHInm6j2ofs2x7cfk0jOCFND4iV+LboFnFz9l6NVL1gNcyDpGIiw7v0HPRP06
2+CqgSH96n5UT8uIQgwBnWeHUZ4xDcDAbwNxB52SfbBQmT38taILM1dKCvQdMhDO
7F9Fm2vOriQToGW7iEt6V+Tv2rwrAzHk2LNGycXlvbP4qbxzF9+7dPk5c3E8MJre
uXu8woBYWKyZQ/gnwq8jkRKHLBpOp2Qj5BDBwjAw2DwwrSOiDC6Esvyurx6Vmxzq
GLv3Z+6BSLFbNisdxxL+lc1egCsMH+EushtduLeTTrfjpzV2QrZvf4tLBrM4m1tv
8RRObL6periofi1oQ21QnUzomT50Nknd+ks41J98oLl++M4XKayGTPD0wTdkYJwk
rqFkexLwS6aDOYK7rg3hMyOZMS4HBQhdqUVJ7vt8bebLdXCly5o0DK1Os5XoTD5F
/+vk1adFuN7lbhVNOhyvpHyJ/IEcytDp2r/MDo+YyWI9okuU9g4aGUckKPo+q/K1
tLcLHEcPzjOohzGbEI1sFgBCJma1JxZD3gsWQ6EBFqHlT3m7wmMhLbc3dmfUi7I7
+c+MEdi/LvEcFKa+MfKO1XSIraefBf7sLX3+qaJkxvxemowlAcoQRCOePjNcn0qP
DxjE6FnxYYBQWhS82tWE+qYb0kvJBVeVyQpnkmZqvLReEM3uOmAHvtzAkwvch6fs
mrZ0AwE6mWbe1u97GOpmaWY6KFrBaAo/CgCZ/Vec1OcGH7T9KBNFCIHx7sYL46C3
CPv60ZEL2AwmVaF0+N4IIFW7nP3vzInx94do3nR0YM+S79h7+5ymSqM7b9UKGsid
x/w3bxqHhvsXUY6OcYsGET2wJMlpc8JUtlCcrlI4vJdCVlQkAOifwj1ilo8enN8n
Yye1dx0JyWyePdSqBwhXYz4XGaOspUfFmF7hEHUX1IBL4uDXDr94OxBOa5WLOnVg
h19uqiDMsGfHBzyeDXNf2nBZHmcZTCfI/ck15UmmI+fCir+pZI+33BSJ6NVvxk+l
V/JCAMAJbtpr+LD3g7zmR9UonuPhW09COrrviV3mz72lFKOzUAjyAiL3mNJg/VBj
zmlD2tKXJE8ZGQhOwSvQ26pmaFdnOLAR118agfHRh5HrtVVrIOoGSo7Vatex1AT8
opTqhIsySTuhmeh3WP1rbKyfbbK6+/TBNgRERX5S2iBdZv6cvtEfaUoUx7XUoyYE
dzg+Na6NRF7gBHKQ0XpHWHHhAfsUPAaeJ1OY51Id0Pf2/mE/JQsHGYotnx0dt2+w
Ffr+JLwqIuJpQwCRTN7XgMqTSJ8G0PbETTc59zpzL8R2qoCHT92IjN6dsIAgEDJ9
qOnk/GOYnuhtHj7uh7JZ+fJD4uf6tz9GuY5hLdlT2PkfOoB6KQOq8DaeGSDLkHBU
sUCZWs276N3GIXHyEc3e42UBQFaGPb3OYraD7yhthXQD7tIgxPSFfmrOBjVx4ZQJ
ayp1VOBNXemWy2OTERFgwphOfKZZQq/l7MBoCBLx2LmDF3J8OJ72cpIKl6bBmJ/+
r0hYV6RawVITqHC0BrSa3SXBH2dMjq2LdGF46mrixywd5pYV/onvZLXyd2I+KwhX
XX4GXCcDfpPDqPZmA1R4nCFUiKHJ2K2tguBkuF/FD7xPmhvTw+zWkOwF+i354Xdx
Z567BqBTJb07FmxB+4F8vMOVhlBCUoAQR6kkumejMKtO0bPUNqsBOHKccwPdeXbU
s+8E3xNNOKn5oo7GX7nT7iJTfIIPMG+hpO4wG9Lb+xqCg5g29phOWDMvnYSRKMIu
sROgwhGsvD7j/fwSHaZjGPB43t02qPbH1xGc4JIRs38emKpSoWjv3x26lL2ZShwQ
zhZ1r4SjTqjrAaZiFlL/TihscYGLjCSg9Ptqf5PWJhBqiay8x+ileAl6Q/WFE7hn
2g7rH1/k4yOwlX3v8mJ6SZdWJc8LNDhRhqD/X0uGf7ZRCa7um0+owmPVRThf59N6
9uCfCOgh/p2je9CDCttwYFa7xvItMa847mt7hYTiX0gXd+ZoBmmR/pp5+2NGOZ4i
2yptsgtdVSj+Cjvmo70lGvyA3XwBo4suIRubO9YPjzNqE91WxwpdZg2FtXUQiUGw
xDZFGuaKw5q1Xlkh7hdceBprG68T2cxTkkj69YPKX9GQcyGNUil1PlPlNl4gL9R3
QtLugJB8Kw9gfA9TrNDJKiWZPC+hel04NSm0mdw/PwharqedPATV1Tm40SOZSpyM
dWZ3dqe3zSCLxkQvocZjejYMlpjG5KrBibWYjDaBU/6wnXZNgy3cS81187c988sw
+VDYtvkSJUmgdKn45N+dmD8r+TcGUfCJFN/Wecc+r4eVd3dyKiDv6FQ9UjzEIxm5
A+aI6RiwnxvpKMj6zRcOryzZFZoTe+sizc0HovXPA6RhdGfQ5rvkDie61hlY3pZ3
zW4/IpHSb2dbSrn31kLq+3zabbfpz7lG3/CzB6TmUHTrKSCY7LlNsnFBmhC/KSuW
uNU6pw53xf04XKqgm+d3WZ+zUKAWAEfdQuTsgcosodm1w9o1+rXchUaXjiAmxXR4
XLCnh70M1riADeKkuPFc7dEJ3Lx8NVyHintOY94y75qTtKiYaBAuFEexw6FJWwuT
J+/ict5woRzjDk+NXrnK9r3z5I67d0hlxywrGwdVJM76Br+Xo0w6+tm9RLMRNImE
RnCN2Q+C4h3CQvphGWgh3cEV5j27CnAYKBxPMQbMlqUgnXw/Ss7YGbq+cInNClc9
r1ZDr+e6WMAFjMAPK+p64J5qB4FvOKxU6013HuE8VQrAtmTE+hRsRiYiYUf4Axwv
fmceZ9XhM8T2LPxXyRo1/uId699bRzYeQ8wjaY2EmtxvG8cqyfZGGHYKIru6P8yv
FO3/8EfvRuRVMnjFhGEgW/OsnKIrJ/SUu6zhT/pBbct9nUbomJ9+4ttJTS/3vNu6
VerItcCaN9rn4ccnF13UVIt72e2/W+TAclpWkXAdcnwBB5akmdPAZoMIw/vB1isU
eUffS2V7QGOuFeG9XhH1F0Yj4oDpCpcsxYmks5E2zBXsVkX0CrBDHdr5mlc39sdo
AKS/V2NManBC0OMSrAHjgN80tVZ/B4fveazQVe3fprU1DkhsylcJxNQIeRxRxxRw
R3wyn0Cs0ZCWqqj4Zt+RmDpG0QC581tzE28IN77gaUqDJJW06Hq0Lxj/NSNG5FKw
9RP9CpqR168yd2z3zWV6Hi2t6vBW4MnL+/5i+0gScW297HR+SNUxGiMLUSncKzTm
90nvyY/8QgY5iJRQdxja7d0cXhZZnU70X78QC6AU6gJ6rgx2xCLkTkSyYPrO8Ihm
hbO8RYcM5PqiBaFmwCMoe5b3HJzLoTk92IfJaSEV2jkvd1LZSLrY9IDE0pmcYyf7
tBwN8vN0s0rzea0326qFHk3kz5ItvwrGDOsLdXDeFVi+1VvjN4YLrz2wQVhFizXz
xDAlyxzo/R3AZWuCMd3vX9wu3i38uHTWeqVXcOy+vEkO8RAXHS8EE/JEC9tyVM3r
JQ7vMwubZdcflDwoIRzMB9AlXbhl1r3FV8o+C+hoRu4bA/li9WO1gkchaxk7ke/q
cc0KEkrpTrrWpJH/dyokbljPws4dXw2ggJX5ITwcYG8axDsY3T+BBCGL9gYEGiDW
ve5q/JFP+CSyqKwAobhfozYvtkaepTb7U5XJNphZ1Gwhm0MUgiKMzz3SLe/0zg0u
z5Qw9UIOkfZQzLar4ffrKU1xHsW7zgghHZtWUqy5f3N5xN8IXGleUM6SVuumOyXK
LxTj6MhfA9raVSjZRIvBu65mWXx5ztyV0TcbkMak8dd3MRhgUupMdPU+hDcvhKIN
+O7ZNqsF/Zwguzchvc+9nh3y6O5A86/FC96N+QxalWguYS/nW6kzoexdYIw45UPJ
hJiIwhrr/jIaewl6iWIpQ+/4CiYERH5An+m4OgXcDfRolXQm8GmbmfPoQS3/MVr/
NxTZ0RACsNy8Q62ZsnH6CUfiLefuKdbTxleKEptkYNTNEIIA9/QLMu8k7+QgHDIh
/BkEpGtRsPjuKzJE9/HCgGM3iUemAv7qWvrU7dMqaGM1ruGuH8Wlqxq5wkTOkLw2
5/AffBGJ17lCUlYoJGlM2nrWtqUk+DqRTi4IrLqe/LN1ishd6rtifhETQ+8dxmj7
g7JcE9l+X9vxIuxIEUYDUpvV/KnP27pnClvuGx9Qfzy9G93ND+QRZRopNWMKOyBA
wiXkekql7IvM5/z/+8nuOOaWxdfYRKeW8vzAwmzJcNqfsIYc8YeR90p3z1qktaMA
VA2X/CAqCrMxda0Okx/SxnoDfatdKp5TqtaYR8PhCXOQj7QIDeH3bACnpWnLr1sx
I2rHVLYag/swuS442by/MRjGRPjgn23JCvDC/CFfWBBg60MahShv1OUeBSpP4AFN
d88aLzJdax1H4v+t6IxsNy+EpmxyqVsEt+85KtS7KVKXBpdF6AwlBHj40ghBDcqF
82nE1rWyqK7sEQhq6AYmzbl5M8ct0jOzmt/3pVd16G4dVWIHOk5XGv+9yiaNzHnc
Wknmy8Dl1Rwc2l8WU0nY49inQYE8RmpOTdtYXqe1Zbfid/OE5zOSdDW/+/CWyjl7
4AJxR1gRybzFu7aBm/yZLveUKTWjHn8AdEQHZ5GlpgtoQIE7DreDVaNYyydfoxcj
c9rjcNcHdnLDLulDo21tM+fMqPKa2U1fVsE3QjndAfFLiBp14e+DAa3ZuTSxZwu3
8YnTrlQ5nqq+deN8HslsvUBKvipMX6O0CuG79SiUTVKRg2EdwmRTiUM/jDj5njor
pLRwCvkB+1devhCcMuR8ZaJ81yQOlefIa5HjkgE/IOmIUNZt7yo4I2BPmgm2eRZ9
PHm4rxHQzh9Jl1+YctO5+UkF0MRL6YJxJYUn7dMvuhO7Izfa/OZ0pXfz5vYI2TxX
0/4g2LkPAk/yVY+BA18ioEBllyybPKgLYGwPHbfqS5I3NmblpONanWt1yWmx7Pv9
zuWCSFFUn6Hw1NItg1YlBXYN1HVXCbNgO00IRAcrxZS4axDvcgtsstVTulxfHpIs
SVYqgT9cRPQ7/0D6Wk8EGmRGH+D3g5BySzr5iWLi06mseJKOolKhNr7RZjU9qtX0
uo87DvHGv7DFjZMbDMjgUxP472ED9u6A1RBfY7Ub9da7O7q5sAxWvgyDJMt+yJZL
eYbl/P3eTBwZu2fkbSA3i2w1xDO+OHmpoAagZwkvb6dVVtGNZdTZy2JG0VnAFfpM
oxaJOu90WesWcVy3kdWoV4UJdW1YHI/e3PSf9dKgzSGI/e+0VJf1BDtXY7OGjK8X
VfsRN4MVv29GmL2gTRBt+Qm4alCJF7chyiXdoTMZHxr3FEgW8LZo/StWR6Bo51uo
+Cu57Y29CDFt5JP1CqpuvaxRdqoW//kUMx8PS+mvca59jP2Zo9OF0Jy65zwdZejk
yeVn47/np3ANDpNh+wNOxWh9UuOOXvgT+6sRdzoQqgy7pz0Spb+C5zCiNmhepi5V
/POkRt1H1DIU91Zs/bLeI1XW2Cslm7CWdqmoXL4D7xZFwmPPbPbb9QC5BKTHBIOy
f/NU2rpwnWdqVYGQQE/H84irzm/TwzO7shwnM9VCfo8iQNnUnUl0eHI2QimsUidl
U9gwHk4jNfOIrkTEhfRiqiFzWDtTIp2Lg+YXXyW4ygIYkCHKaWAvcXLL2h1ViPvK
ROIOhH7WLJK+Il/79Jyp+r205kLbUT9vbjmFaZhY8zmwlRzv72OK38AXE2B2ygIi
4LjacfKKEy47GWVWYPGUe+rXgPc7APeKDaN5rqILFO8DNOjMqSIn+3Dq72q6vQl9
tJ8jdKWCZtlXu3f3VMGY27X9DXWcxhwREl3QI4ERz25xeL+4PKzD2XRvxNovghI1
qAG111GIzlDTsyWHPyzmo/h65clNtfQPpzyNW08KyBID4K/12He779vz5Ke8vLOC
bRH4GPcZzivJuVYrrjd9QnEy6uSResEh3Xxiv97iLLjX/NVG+SCQ4wJOwHQ5JthX
XHYYLTVSzi28j7ifvdHv0G0yIz/0811EcoouXfl2cBhnxF+/D9RS+ae5U7d5NKoW
bXWRJMBwdegBCFTye/a/DC+7Cb2OiNv87v4YjLVFb6K0h/Jjqyrh/uOe9QCFL/bK
gLlnDV313qye3UcIiPwAXATKYcHfKy2FZnRlZcdU1VYxbEgIadiBYnL5FlA6Eq9P
B3SKD0zzrVS2Q+/EZfDuNRUzeshoMeafzVeFL+GJniar1dd6zFb8nV5i3NZYr/Yw
oPUucaqPX7Sm/Q6QWDy6vzN+ujT8zkUJKnNry0CNfH3EtId36XqLhadtgOmvI8fT
TSYu5BA48z/w1BDgg7pS9ktq1+FRW94pYUxUlc35Is+fNXTzPEk8vZnk/yoraxMN
ius/Xgpd7jeGl++1t1QuNObUx4tDtvqzLQDD8a6r0RF4f9xJBzvOym5TqTSmNzPL
nztzk7jluSJv696oQigV7BAqVTzTpOeDMW2KVSirTim4z5LBIE7mTINNtd277ZRs
mkoHtFe8j4C8BHO2de+g7LQM9N6iwlVAunYMm6FuVBMXaqusniLB6jMwvafg05lh
eZg6d4jmoMHpRYAHUu7jAtkOHL/GC/b16Cv26RByuY1wpu6f3mDnl3sdegEjMP8n
PdPpmRWu4Pd2PirvtQmRzSByRo9W2aC6JNGxxm9Auez+D+a2XJnJvWU9mA3qUPag
dhBJORDfWGrnMOMPuXJr6MY2n+Z+oEIfhO6NDkeKSFLrdJz+xKCPxg9iWzTQ6N1a
KYosiJWLJx0BAo9LB+fy72ID4Lb2BhyVX0sFo0jt9P0elHf2QveM728Mm4lV5PJy
t3F59IDR/CeulzK206Z8bvLSdCLr+p2Inl920AochZa2dPaspnp9YuV4SzJfBRjK
HFWZ8ol2Rvyp5ApHyWxNwrqdun2T6zMPC72spFmjIV+iP5ZXJZy6r2kPD1jPtQMb
kQcUrZl6HrlEMeHboqq/ljlNWG0emzpe7RKTRSpE0wCXjmpkmEvpGW490SpnwsWO
ZI2jpVnMfrns540IJ7r2pBqi/V6VlS8pypEzgTCD/ApVcxx9VcYJAGtObUxMKy+X
pO9buYLxHjBBcYCvoD8d1NpZJhiUdaglcX2LT8RnozDdH2Mkk4FZ1pXmwsS7gp91
pPSFdh5xg+FqsSiMmpTtG+3jXxlR1QWWuOlrV61syI3cJ8WzkY2UnO6vdGsvnbxH
aUkPEF1pEw36+4WOedaK37azHd2nfCVnmSi4hBwW7AhMo6fkadKjadAP5u9Nhtkx
//SzXvupFiXaadNt88RCJcwgkJprEElE0T/OMM0AqvB4kwMpezm/4D2vq0dhlWdr
HctyBCM2AqYqT/3cydf3B7e+hpVD5X3S8fQT2gkOl285qA8l1J1eiGQMm4AHnoGj
17sKhyTjPg6MsJLuWlboC/NuHXWqnOwa4ABCWOLSo2ezlllyu272e64iyAdM3WqY
rRXo2s1qjc0IWy3tAVxINDkqhBX5cAnhfiUjk9XRDM8qG5CDAD0PXWcylwH/fYQ/
tLh17dzRl4LDqQ/EoF0jV+xDhmBX5I4bNZCaB7umawcOLBtROZKWxjnGjVf7Y5HS
9mDwiqMzbczMhPi4JlEX99TM2AaIJdCuAN+kQnnqqzeWMvan/l7fFH3GkdefZdPC
1ljt4sk3S+VaFtJZlsj54xygGqdxBGvJNC9qOLCQsOLyR9ZtF8UpWMpeMe5QXo22
`protect END_PROTECTED