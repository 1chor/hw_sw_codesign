-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
iJOzlpm6Rlj6TsZ9d2lbvTU1jfE4vRtKOxPJsStQGrxL51FWduLbTxWK/v4p14hx
rMqVRL9qXP26/E2EwQcQ+iFAJNSDy98JjSkoRHR0vWkx20hyhhLTXT10ae8WHPoL
2WjlS5SKk24kX9VscbqkAKYx3V+HK4nlOK0mQIYhJN0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10313)

`protect DATA_BLOCK
6W1va3aBVQzl8/+IbZjejnb5sxlZUxOQse0R/wJaTCJqgvXDDQIdMfpPZ4C5k9I6
E38ZrS0c4jvJiBpKAP9jRD5xp7mfU600qSPycS6KODJooAIpkmX2CBfA138gInIw
Bktv/VESRBUlOetinBJT6fHEv7r9uxSE/XJ2kXyEe5StKPQBFFq7vt+AA5FLndrh
W0vwrfwkM5mjvwIGisSp2PvntBgXyXzngpbCy7fjmlU8wZi9l2LPt1QPn12NtnT8
agBueFoNOcoaLWu7QeJKpAqvq62qdAKCvOYHVIGylycaxOF+IfIkjTHicj+oA/j8
tbtSeQk4C0DXlsfyOUOrpUxcUtKnJUQj8046spjA1bMfbEwPKltOgmod4OrtfAS8
XBi/7dBRnTJeP8VWglZWKnIzODSh3Cv2L3rjTiHE3ytAikPKU9oSYK8M+goSy+vJ
wxOO1RDrwvU+t51otjqG3Nc7D4hXEC3PIa3ICoCYJbcb5FNnJn7ivSdMKIDwQshJ
26qhQHwGNJDcyr1Nl/yjwTnpZ6KeprgYQLuJCEc3R8EUvGbS9waUtbKik4la3ARO
ddrjuKa8o3Y8BvwVXlg39U1FOohUzdPGpVEnL5dVfNRaZx5q9ci2jW9Tus+0X4FE
Pm4Nv64kg/hBIfnFHuNzOETyeqDpwaylB5IbH83isiRj+dQL+MvMjXKJgySZQaSd
bYSUqtBdsYh6anvmHXEGJevnKpfkz9j6yoZMzJ5ccg4gdihw0f5sdtn8e2dek2km
im0Kr9Wp4vTJSwRy2dW0kNpe03SQUF9fF2WvQVBXBwRNBPFzKcJMyqkDmHTjK/ER
qHky9mW7oeHvCiCvVH3/R1SCqprFxQ3GzirxFafQXm2szSYmFQSjbCbeq4wqm0Fw
kwpn0xZUKIrdcwqCi6J62Vy4O3UyLkkhPMTmrJVcOSPtFkaFvCjFzbzPEMB7R72H
1Yql2bX821QnjdCKE1nP9U/4iW3Hb5LtuFbuKyamzx5k+PYZrFeyL3W8F3N24RrO
aAzPUiL+9ratP/QrBV8nfxtbYsGuM3gWcGHspUuabJP6vIUChWwK4ZDUY951tmqm
Kg1NdwU2IXO9GmWFvS8NAI6JZatwd01s7zdGu55dGeOgpWG2QYIHTT3UBqBc0xk7
akNh7SkUDzpcY/Ok7YeVi8oj8g82/VgfYDzyeTmxgMCeucNXXKlCvq3skSs6KTqd
sCKMt3VGmKhCR9zwjI8bneaLvBr4tnl3n2yPlLR3tbSa9eNabDTOE4uJ8r5cKJ2x
lER3+0i05QqibgzlfYouKIwiKHZ30RGFAKHzyA18Gkj4tdEW+gUJ8e9T9cqkXhLJ
FprWHaRMfq61tG2J9IjewQaW8bKctwdLMfJxTFPn7+eEtVULukP20GF/P3UpX6PU
vcgINDYIKyHU+Zb8ZWlvzBhMq4hTV6U/9GPYSgHpDRK9gHur5c7TL/pSHXGC4ZBx
hWDt9hPzS9JVZXzBxciDHpDxpINLnBugeBDVK+Hc3amHnj28+fymukmqabretSie
rmSLBd6ArqYg2sxEzCz1oIXJnSR6kJLXDLS9pc6qrXBXV2qCQbuLp9v47ao91jRA
TVfvppbgpuco6yg4l3qUO5dPQEsKI5eiFJFznEikkQEnqb3u54VNUTKxgRAjV3Xt
0jg7ebNGHi/sxoWQKQBdkUKKBACFHS4R7cFg64xlqXmI3tcwEMSo9BxQ1hlZhG0F
QzlrKtsKwrwxmHW8Yr+gmOxRAAmpqHZOiIseICWbNTQT7rIi6gZ7i6qmF3IDiuvB
hSe2m3X4zXYmE6/ywIO5BXzPwZHIoorNLwBUCWtOkr6uhGq0HiSMEu9rY2+Q1jZS
0TvGw31yUTBcE4BXxZiXDYA/anvthMZlLLDnOp79Moko+8jwqSDgNME6tR7DYqZ3
LZ8R30TgAW+nUzQ8L6JeTkhxmB/S3KL8zHz18uJF/VS8P5EXYDZNNnuRQ6yHnFgy
CMsRJN+lkJjwIoEY0AMb4n0WY3Ro/RlfxGrxtkpa3r1vJt++38FAnoWFdOX5ZDrG
zHhSzwPC1WXDYFbBQvnth8Nixl41MrmS2+dnpsE3SzK/RL/2PFxf1hm2mPqH/76i
SbXefr/W0L4Yr9Mw6IPhM1TPkox1MC8Y/zv7L3DA/XazBHL0U66AQnIqooOxUqJo
ul6FWXZ6wnNsfU5SL/OIv9D93hDp8zI/WUvs0pwj7/6u0o4dsOOq5tamXgTT26Yz
i3gOZ0IzACnvTetg5B/AiQSaYQtFqAr2zUeW/lRT7WVrZKbHrRdp0J0lX0RqChgf
hy/bMc2UPftuycIxdBdGmNmSazH8Ghzawf8oiLxeoTYzm2lsVG++AmV4eje4nUVy
4uBb21SJtN0rzTeYTilvfCiditH+7UO62OMC3phIKOOoaN9pAxGZZXe91ftjw9E6
dx5VVouMVyxQ75LdgSDWSWtZajpBAnaLuhB443Nx9uDiVmpVcIKyUOIZ4wbbi8IL
SnJMBlFLRnfK8tBRXX8ipjs9YPt5wr+duHl0cZoA12reRYLtQsoe4vHdNur6EVHm
QPGc/4B2huffUdkNl/mFMhGTgw31Ogc0jcfW8BnCp74kPLJtjz3WUvp2naFnPa2o
1Tb9rwUPIflucvAj0FwJwbKnZBINTvK8227rTvlRnnlqMuRbPc44a/ZVA7a7qqVz
dPwiNrZoNMfZr73m1Tys98OzY1CGdF+MaTm7dO+2jFRfghkUFFr5VvqhMYo7+sWh
xUsijd0pDYRgg1VVGfj6hK45WBXz3Ojy7O49c1f9y/wCfueSMMFu0OA7RqzaHGXJ
9FYjKMCnXvw5gZefjE2zQCHQ7CLRoFdE9zhKcN5Ts9EGuOuvI07elennu4WClOIT
ard2NO31Hlm9SqbBo2WfpbcJ5/sKl/P/8rO3EA+yKBX6U7JX/LfHl1b9h3Ee8LUS
o89ydOeDSO5CVbEgF1g1A4F2WNmquYBEEtQrRMM3VLFcROkAw2nf3MZWr3W6l3qO
ZeqGHeDTXNTGYT1UCkaFpWCd82PJ7r93theRjMxfBP7fkZrmSJ+KixFIuXhFdI2X
q6BAOFR+KiLPah0XoEcyLF72wsjrzhoSvY0XjtHNKt8KbfztmCKSh/A5D0FB0b2d
yy85/w0k7LV9DyVztaQ3pVAQ1bK5e2Id6wWRCHzwqq++ep/0bPke754NxQTyhvvt
o4/XSC3X4g11KaI12SF6oTRWYYGfyp7hKav6NUwBZV8pwNFGdtm8YIUVHID7cYjJ
94GNoH/02vY3R6h2LHce9e+4QIOI3we8PiAYwAhBhzmxrA+yQYiy1R1s+H1HWimx
8id75eR/nnXsbySHoYtyejPp+nkcJcN+mdUcGaBYNuihcYaR8e+bU0zWOB9pcjiX
vyLyWuIogLPN9KzRsOUExju53+2p4uowbBvl6SIIuWoj4cCOSEL/WKIKpsURdQq2
fMPt4n9OgeETs9DimZpyIjuSJvPYpHkmdQ/NeeLapzQm2iLc2ZmGt4OCa2OrbZQK
9Khd1fomDbiw62b2r7l42UcHAPNWVBj5BphtI5pncMy5cgjm4Gd2APNZArJmkOwi
/yZGkzQdCG6sPGGj9VOXMbidgLFwUeJGafeQKhfPfsLmOEMUqEdwDhmcTi63ol2U
ojKrqFF0Weccx3NpFRbU/RHSDwExFfwytGizMY+IHUfgrN0IJzn1D5ivSSIqmebb
7dvA85tx5ZeubenjNN9nx9j9ov9SLnYetGdX3BKRcA0WWEbZxEZui8v0a37NScxy
QGlux/GOrEzLlECacpK8zMM8QIbb6eK772ECHQUFOppXwB+1Slr/nWjzAT+glfrG
wTWxyh+zGzPSQjL/IkkfHu+zWfC9kmXrkC4CFWDknrI42YwOAS32bP4LXYE0cv0V
LYBEmmZ6XzoC/UHreeVwK4QAknB0xnRBrv89YRFlOetr8/RCY7+qYkuTfdEjuwOR
OoAG61WTgmM8w9WHhGuONlCSSdVhJDPy7XsIfdBXtrc+gpF3eAk2mIdIzcqXea0E
SpVK9kaUIa+Mp+SWfYbUjACk7eLe6b+1M3dHL985/eODm+7UkDmqh0QNSJTkR+xL
wQ7ROlxWuyS8BJCa2WWVdxnCNgdvPWPkK3Ylry2pHTRL13ROC+uYeZV/cLZBxZDO
wUxqkoNycBlONnZ/HoH031EsFp6Q4T71rnIffIdN3UV05ML/L35dWOVG+zvwaINl
KoR+3+Q56q/1ADKdRevebADmGrTakJUBpl2rW9jTbVQ5NpnYfRRKYDEJV35FMUeb
lZe6lfSbyWqvEZ81cvVdfdyRCeMMH6gw2YWuPGfcih45zGvu7543aMQ1l72IhPWr
vwM0k4ff9uhSmMaBovPgN64F2QQn9zNVsNX9FhX4zOcbeiROErwoylHfGeWfsGYZ
wPEkK3cszfspQb8Vs2NaNrCyVLGPXrXJGRXvCG9d5Ebp0fxoDZP+UPQQE7HUbCko
rVhyj06SqqTrmg5CUdE2VeqZZJAdyKGFuxDtX4PYK+YoD7xO4CGzcZu/hdSgvlhm
tisyeMrbA7bmqXJfcijYSTjBYMtO911Vs8U/Rkf7k4wAhWfOl8AcrBHY1RrrhnyJ
Ai1uRkm4PXrK4qwvyZoR5B4twtYq+oAQ0CUvG7UFYb4nOntae+0sVved+Xv2gUaH
1JkLC8i8aGFipJj+4Vn33rZeR5eE73Y83USRJ31WG9skPL9pCTEt4h6mMeWrBkjE
24UGKKM2cxXuEzUIThfgZmbSbta1TTmjOFb/dfzDP87lZMJHMJPDF81mVvWETCm9
VYCIGU1vKmEWwpn1553G22YWYroY1PoyVXnDjKVPSFsjZYu/9ntgWVuqI52bLWU7
GwgrTBeCPXnPsV62kaQhqtjWyJ2rifJ+Xa3ohNRaFxhtmmedwOjzQUSQ4HNkmIV0
+3t0iFLSBxM+5g95U5tHcON7DF0d66AErJGaIBT4sxTlawN1QMmJX2VsnTgFdC0r
31Fb9776oWwtu4oJjnUNHqhPG+b0/SOkn5TmIekHVAwNUrDQNPFUurDHLrbvonrw
KM9tyE7qKQDG6h1wogTpW4tCVgIvvUJTJ1vFoUOPHkd9BTzys74mBKOhDBruFPFU
LtaITtra/toqwURudVcY0xDcsWhv7T2YbQvPgYBeHtLMRvx42JJPjEgbitSnRe9M
XcKnExgHlqB5DpOC4zmQST0hYDc+ZErfDGkFGxUG4paRJgndAvvWfpec+/5RRo9m
5CBOuU+nAQy83JehpfGhu0psIX1ZDhypB05WX50/p99o9J6n+yOqvHUumvb6vt0m
KUGhTKqWpAzt+MXyVS0Rl4Tpc1dO/4TnGyVeX+xzKslVo8+901w6vjoMQAwS+OWW
1P+xoJ6DUTFwKSBbIWKkRJvYIUVfNo5vn4P6iE+BFVgPx/2BVkTdqkK4GoPtUHkg
y1AYJfrYMSuRkTWu62RYIPU2u7AWSbj1BTkaOSs3bRhWfyw3zCF7V6RdzLUfEl4j
lfp7ILIu5kGd6vjkh17Yn5YxyHGJ0YogV7eBVJYnDCr3Zn9ef9ab/aedhnI41aO2
BbWkHxY+YNVcr6Ywx4PppB1LV2z+c52Z02jy9seYPlGeP70ZJ7ljBGMYUhPoCnaF
4FrSImRgye9tVJi9y3UrdlBykOtVAUcGeos+xU5ovbHB/C3Xz0bJbWWxlFhU+Eie
RFf+r+Z6Yqyz/uEds/SUFnHLpev4FZynDaB5uQ854xfKtsfmfEeHf8T7RXRg0LcO
qQ1Wt6zNvxvKlcRBLab4XSjI/EfM5O4Xq7vNt61yjWr4cH2NlNJy5oMhUhbpwMPF
cHh/jzJVX+5HkJy26/8D1XMu4FYbpmfHBgS4/66fpio2UPfs7RXmu3czQDVBcoLZ
47tJ4EJFBJ+5ACi0L/NivsNqc8s+mUlsRJaFMSv4Kjh4KQXckaMRl2VlPX0Vbv2W
jWP0MiB2wL67Yf5b1HoBHFeCbYm8E19QKFO+JNLixX2/nc39OLl6Dausnb4EV4Xs
53mkF0Wc1OtUdB3G4ZI9utE6OOkImQ0oli1IZk8FhgMcFSzBeu1bZUGoDc/K3pWh
E2AJn1law4QNFFPacqNDz7/0ucXw9oNNFhp4+ozJE6r62C+IluRH6SYZk+Uq6L0w
qXbpRslgaCNk3PZlIpzs23hUmO5CRGLtNPSI9mOtX0+suvJuW5JPZexSfqDuO3ZU
mJjyBU4kmpeSvCd/DnlWF4RhL1867wKnJLwlf2tmHv0OZW5NRkOXdGwrnxjyuuhq
cCncs35vjo0I0jVaptWFI4uc7ST5Nu+RiAoqGN9yoezWDAKOw0CyATe12eFxmns5
h5Cj1x5JcISbePRmS/WFFb72CkB5x/5Q53YCLyO9A9Q7YOX1OGmgf5HDDt1RnZm7
zv7D4PxIfXdd7KRLaesofLaUKQ5Ix1Y+nPCiZcTdXh4D0rl/qr1IIZJ0VOtQAeTD
irJlpQ2LFEWpbXd1CArWDsYKXnwYVXsVmj+C/WmBrAUGUlGE/akRxW9e8N8dAp77
NK5jIOjk4ZL3txMBW880NaCIYRBzJbO7xmKQ7faarDTyrC9Onjvl5VztRPmGuFhH
rqrv8dM6kC1Zw+oDhQmkqCs+lquz0prvOx6c1J71+YO91W8w/uNoBlYzSpKxMlKt
EFVpCUu+RokgH1q2mUGVf/Hjr8k53rCpWMKsn0JdBzC6tjLGAlWNQQHgByfAE7jC
vWFSYF2my32WzmmLn2rUF2yEeEqHBLJQkEaP6DO3dvt6XAZlAVgm9U15slqNX1a7
YzvW762z4CgVQDCIfMHknH7USTep71ArrvDM4Av9uNC0H7mcYgQUnE/BGzMFU0ui
afMC72J2gaIX5vuowblaUnONfwn1iFKDLnepZRPOVGGBAir6Oi1jogHyZdnvQFnQ
TVlSmBFZeQcS5cLI1w15vUc/R2TKIhmUp34B8WsWCcF0jHDRjUX335ajX1ZypHbx
jITwPwK48lTQEBAQC1nwivOLv/gMzYEUfsINU8XVkAq6+1rHGT0oMQBoikzPmoEG
0KJT9rrlUt5cQD2N4HT3huks1fXMneYhYLX/0tELOtlWpUaMuLMP63gx1ro5/PiU
6k6zeNVtaaKSTX+CNGhrKSx9AAZlPpbZgX4JV4NF7thL268O0f4kHGh5Eh7ktHSJ
NZ6M8OcbblmXyGcS88oKNM0eVHq3h3l8+cdG9qTljrScwIPKdi8yKD52TBv3XNau
fbnzGI0fOoIToRJEz8C0/bXu34NQXWtY+k4dSv0Eu7OCAw3KzXV7qksEsA1z077i
C9R3iE9jBPQ5JC03PLYvuNfjX94+SPIrVcQlFsZaYJxGxtNJxSw+Y30F2LNCV61V
ShG7aeqz8qotvY56bIozRFMI5XQ5Kqyv9PZGHEl1AYOc8LZJNWR4DDhUGvsohnH1
EdJRDGVv2ejH3dEg6l9VGhTD4MUwm+XXsPNqxlx/G1U1E9pJ67k8t1Vv81gwTO7Y
P8js3GhRt8dVog35wzxIeVAj4sc34Uv5yzIEePwcDAaM2XghZo+P300oOvik+EB7
eBGPHkDA0nKlNHVjQA+uFQVW99aPcr/YOpo72N8JEqW768DqlZJcX+91oP1alo8w
nAWeQudNWd8vAPn7CbEH9c2fkL5hOju7Y9TUluszCp/1pDN75Rlp5bfVhkH/hIXx
r31mny1IqlUPbagqNa5vMQCHHLgf4567Mm820tzd4Uk4rTJ0zMC8ihQR3RfOt72t
2z5rDzc6E+rVZp2OW6H0t2glKOL8nGKzzVAltY1z9BqFH5OcggXW/bVdnPfSiPKq
F/S37WrjQSN7/wX1XTIVVhVm7jlduQUXJpx7gpcTuHDb3ia+CunFWulpzcCgkSKo
foWDZh1Vnl2OtRKKssUFjifNYzVBGKg9ENfP6UW0VKpNzHInxDvN0nSz2nMoUFuf
GEFAFok+/Cib65zXSIP44o3gBTj9DvO35qc5C2JqEr8rodWMdEj0jIgaK9K/p3gb
8qLWyly1U9Sy3nDkPMJa2YSII62uMXV4HLj0aUI2l1zf4UgV8RWcM3Zr7TV4iVsx
dkiy4dnxVIulKquMPNB6KGh+LbYgeU17eq8mvvPDzwV5/Fueo4mpo0004vdP+M+Q
P3WLCx61ZDHmpd1et0nlJQmCwRtJjjRnB6b/jeQdnJx3cWtKtnOSV9LOCKEnECBb
TR+zU8fWen0RZuxt8AOmB5bSvCdiUME+FSCB7f6fQm+hzPuz0pQID1RGuAvacb/X
sx265Af42ncyahFuW5GyCDOfxWkavGhL5wfC9jg3DQjs4mlXFeFQZ96cgaPa0KpN
S9ryyhzLkd0GOqWjyybj266OkXmyiM4VQv/uNG9Hn7I5t4+Frdfro7UhAqVdLnhD
ANKDzpHUb97cz6NKOKPr98gTO8vNNTT9MdFz8U5M7Z1Bz4n+c29zEueBUyAeQNlT
ADZo2VE0LTVtiO6j3tbLsfZFctpob/ufhJrkwe6yVthQBembhyZD68T/GAm+yPYo
fXEh+D9bieCuMmpij2sOrhyasRJQ/O/jBByZrf1pO0/I9mtTxnWztlOisgqptTIG
1yYAEalkXTmvTr5WjE7qlyd3J4nW+Gwupx9VlbIwcVXqtjqEiaWOF4LtU7Zp00Ht
d356LREGDV2zi/yiKOS8iHNeOUwy9K8StquKe5L7hQH1aBpha1kCopdK55stSaFb
RbjbNbStH2K07kJFFREm4p+vdIVd6iIluipSiE/SApQB7CMnxGVSWwMiy6ftq6Gz
VXm23bm+CHuqPfMWkseeE6qUDiuBXFbtmD/6g+L5I2fQWP3YVWg3IZuNXLYZLzDx
kPRy71KThoTCJRG0QcHo9ljMMnakzF4+PkSWPDlYexhaZKdlfZB4zZMGSaow0jdE
tbZnhyaYx6xnNKDM4oL1JDVgTvLP+4kviIPJTYJJPb0ke6dhPJNh5t53QjoOZQKZ
zII+BxVasYA92DcEkwRvCnVTAzakr/Um/Yqp8BMOCauheTqYBnK0nHROYIc5EKS9
/VZbciyOkzvHRlul02QZMOseQHxytADs2Yn3bT+y4taIOX5WVJ1SXqpogEmJUaha
CnXChvKsKYi2fzU2ythRkYq3C6XuvMMc6/x3WLC6nOK7a8u66uZ9w9DKrvCeAm+v
Hwy+oOI4a6pymQAStc4CLnjeEn8wFD01YI6AEZ//u1rOHasLQKLy8WTKSYY/dhOg
CkssSNyIV+ZPwnPb71rrAoCSsrTVUK/T1/ari8CNxrqRtK3SNH4AdWP6Ut4CyhWw
ONBgrJGNBA928zB5RGTltd8W6VXfpcZ7nIfdEp5usSLMl8BBxj0HVwxGcv2NXqSZ
9b1G7Jwdih5r67cQnIQM5QOkP/hJETYxdn6LcBdrLBrxxpayIlaYAAgsPjjVhcVf
n/EXvXazwgFldoLkYXduc6AArnlvAcR6p+KT5A9tTpg6Zl1dGaW5YNMfoR9I9kLc
kV18gHBzAv4z3btnlcvy6UmP7ZlJKIxN6LB/d5NWjpsxjHqdhVwByxeMBKyvYxPy
Ti8CRC5W5pRFjLduCeTs/UciJyrbh7kLkl5c+fI1VBZO1tejFgPd34DKa51F+wLN
Ix96yMWErOM3P2V84oQ2QdpEBHM77EjAaW2tazP1+zp6GONC9XF447ZJWTvu84cd
H51Z8mOkU9m+mJoC81jjA20NvLzvG3w6G2iLQ2+QomnqCLZVI+s1oK+fT1bzXPyp
qtFl1N/5+wG1CKgtCT5DB3+dWHP+oEu1Aye0ZxJ/SACvdB4DEqkaZwbrHKtB30Zz
3sAr+25bWrfIs9tE06xfbDf8rEeJOd05CtE78PZQET7dniu92ltbA9/YQRlXlzHq
12OfYVt0yIiqq+o93UK0o3qjAW5BzTkOn+WwkhgkVBgAlfQkGzHPgn8dk6u3AeAl
Np+RjsdAr7hMd7/OhovzPMVtmCYIimOu7r5c2UdKhUsgh8xpdzbmXVN9DqSLPk3+
990xm8/X4kDOCg09487I6QNkzpx2ljtHutF4bq2Kh3V9yCcJ+KK3krL5lVtu5WcB
EWT6lP9vROm80jOSQp990EkcOmjSQsDEjvsBUCuq3uDuwbUf9suBGvaWg476oXFp
8Plju/e0r1HxGSo0bHiBhBd4ggpD2xqdi4A5Bur7xwmEzfYBGa4b/aRp2CI40u4y
zrq1Vq/cFQF0zQK1zPb9Fh3yBvsvadTVCaCB8fcuJ6nfkuGTvHrSNaYHypBRwern
JrhTMGwWVQtuYs1VisjZWCcb2T/XvsPgBK7g7pl3gdEPFpXgIgfw900JGFWrB2kp
7NjJP7vjaLCP5MzEIOIpsm+YXGvzQjWPk0J86Gq9xxCNG4tUcAobTD5El5RRHr35
TdDIMh0bIn+BhWiAvazb1o+i/hQs0dzmkbzlEER8/x4EArBfkSVGXQkkVO/6Hswg
D/qmbNgjXLxGcJPVhJ+Tgha7bwUF5eG0AvknET/8FLxyrz4tXu3ejf5XCcOmBlF1
1ju3XGJo70+aqoGnl7H00LMl7bv7hQbqXDwo1B7iQESzuA3MwPc4ifrXF2mf8EpC
MosmuQzdC5sZiARHhFEqUayHtwk1OkkeJCin+dr3591/RnhnTL42nvb4fJaNHHNV
d3l5bwdCB/VR3CpTfIc7IHoh6mODqxtThzOAD4UJaJuF9v9Emfwd8cNmWJP8JEfC
2vablxwVah4pOcT5o1H3zI0OIXgE+1jsLcvXsJeNQuTuQRM4ADCpzDE9uIG9KAYK
4e71e5RjHca8MW+rrYFptLREh9PgG1BjNSbfgqyLs/bJfF7EYYGezY30GOIC+qWR
P9wNYq7rOqQPFPePmEbnzl24IhVcK1OFFJFFXgwkeyfy55mo4aLo98ufdl2cykBW
rlGpZVDPzmCSJcrDDLTuNw6EHMJatPNv0gP2+HLfOJPomofhTov6yc29XMQZ6omt
aqKZf5VtlTCkneUzuKXzHp5H3uxHQEyC2oA+y3ELZrrM3TJ4BN59V9e/qJO+wSpD
0gS0XKlf5vkwP2BuxWB8/+jqB18YCBlPttvqA+299zLVzkiZDMwcz88qAMCWBKSJ
Q/Y85xWOPTB8qMufvo/YNrYMmC2/IV9pqyAMO/eOe6l2BfQXAHgvxBvokKPgO3GN
htMEHmdGVlqlG741RZf3hnfISOO5AA1BrHvoeubcNwwSNlEutuYhx8/4lRBLYTiC
D96H3es8ln2jVstbnaoxyRybTCkDmZ4DjYoC+2Xh6uB6wsjgxxKPCsbJ4wKCdc5g
lp73cqgQPAM+RVHuz2+GMKxIhIssOXm6BsOJDMjzNePoRUgPt4xuj66yIoJtNSc3
nhJGakBRdupflokTUkqUso+yRYd/q14BvGhtnKt9P91vApTwseIpSOuJu1Z/eVsd
jVVN5iIgY/a3564hjMc9Z7vu3hC65YWeHTEftlViHFv4zQodb32ExUiRVQg1tlc0
ye6hmQmm1KefK/0y8HFC6ZQ/qZktpT5ZBluwLsiJIj3nHCgBt3L9BWRrgySXx5mD
rsV0VBkVCsCMAFxigsIUcTVHJIwXc+5uYg1cMHSooS73VJQU8NO5KTkr22WVUK6H
Q0SkThayqUDCtDfyJIl5B9+ufSzUaNwYTeP084svBu5OWUvjM1IrwYJJhH9FvN+u
bsX0GLroTsk2ffD4QpxYWKdrpfdPSxbpwHeQZTVExUfYcIpNzDvfPsr/xE/QsZIB
6oXsNk7j3avRXn4Y3q61oIJO0A/GvUqrzrpxD7WJuR8TG71m2Av/lZ/0nmqB2vrO
OVridcCjD4Q/yVdDaaf5sXGTPGHWzjxFGB5K0T6+Z1EqOMDvIr+9M9tMBOYiKUBG
SzxPqcSUz44AAm1DmG15zFnAWgQwfteQpJQIaHS+3DEnorBGlKoWmf0uTtOrlb2h
fWjSSqeVlFVnJEHsHD9GVejHscIe5JduURCcJffyA8fvb5tG9YvXOGd0Wvb2QIp+
VUvjY2D/iM6yLbVqUXuBkWUsFAbkJq62r9k1BJCz9yzS/mmhATD/aZp1f2H1Y8C4
Vor4pH/U5d7sh3/Mp6iZFKvR/a2nUwk8ae9yFIUodUdhz0/zg99t+0ZU2+YqI5sf
WKZPo7aIthErbweBLeAXU0VKSnIDKmF4nLkVm6zKxQdlnWOm40FyETxEB+M79Us+
RVVlLehdhIpduoIffkYVebqHAND4NTfTHbsGbKzieHsce6GKM/fulj7Itx8Dj7XY
ZvWpFkPsUMV8QnNVI2Qe3zzoafsgVB8CopKzmCSpLy1SklMJf/OJfoKNVboBxHfC
4GWrMQnFMZD6gbu12xUbFUmqdRQWCDAfcxbXRrUywIFhaD7n1N7T2bD2qOYNu6h9
kguzV6vZuis+V2k9H27kCqD+WDAF58Em6CyA6SgYqHDtb2HH4q0YUZuI6Vj6Ad47
8lPVrlOPj2+D6ZEbaZ7ZHF9HwO5y7QMRs0T5EDI/2Ais3OXuR0EkdR86Kr5gs25U
LsxktiIu6fVEpygvZFoDBUSun7EztaRarYY0UJ9twSvjYgw1dZcTSYsdk6jv1Xcm
+Emz6U7+Vd/T3beK74ao0n/hUIKfok+hjVS0+g1uUPeBTdB3NrCuLyMStkxWmbMh
kigsfsWb8MEkYQoPAUOkbvKxVPB70djjKvHeF545iRmklUCSAoSBen28jyoqzvYR
WU9SBo22x+MjZCv+pt09JIc3Us2tGrjtgCA8ka8LCfqNwiAsgOKDVYA8GTS4uX5F
4MF0y8cjAVYYObdz/rMQ377VzLah6aQ27Q+rLno7yHDM0sA8VUGF/kqnF0Dv8wUK
Obl1jBxlXDF9Q+NgRMl8wnatF+XAoie6owPKcCe65aUqWCCtx20IJW64oqd55RJZ
Vj0lnNk+kIOUCFhD1x1/g1/4Ii3OfIhp2UAcSH1+/W/eIqJ43vN0EWIACj1CGbu8
Jux+kV1Nw90W7NMIPWY4A++Dlq2W85vtwK9N5+Y+VaYvKRhStSnAyZJnspJGpbFL
6srr9le1PKNaVhukLyVvSvWySNRQKmsP2IbdGbztkaAWUWMTuuHe45iSQD3hbbzH
dhphwCvHvj7i5CqQSfC2wfkCMkNOt/w5islnPqUN8kiGaea88g1ZNrQce7J2IhTF
XJHf4ztbgUDgHbHZuelV371Rfso5AcOUfQiFR1xpGtoHDvyMcfz7mfX6AeRlaLgX
XlKxaPDWDDL1JQaOHfTLdRdso0T7of/jiHIPWRvSE/h5fPdNGalmGlpkGq8F3xm9
e/Ksh6VF/zhV5OdExoA1dKNmmy1ZxDqJXjSnUERx5ulPV52gOIMWF/VnpB93xj5I
DoN0vYjT6x8VnQ7eA6oIbiWwa9ReKtEsKM2D+u8mAn0nYcMTzNXb5wrL/Zraj5wl
397cr67r9k/Mrtk43sMuABLN9wTIAymTWQa/5Xs7chTBq9X01XbFnwo1YPoPTnMv
6pSkQU+Kt9ebiRTzDNCTSaZg0E1oMOFbSZAm3DW+lK8cfSlLlKdlq0scTGDxCtfO
LrRV1CEsp3sxa1iMDdFSWTqt0K0tiACl6MDHIcdEPcKt35srgoWLnk8pVysZNaWz
ctpy1CHEVB6fbCYcwzj/QgMT7WV/t9Nce76VtXP2vOH4G/txN0ZW84JPCetzY9t5
CdvILgL1iiGBXrhmRBM3M+gxdZub0THIGJrTVGip1wmiKbYPoITLI+UpUAEXRK0/
jUveG5hmcy3wWT/lmJJ2/c36ObtGMAAjZFAzKm8Cae3zyNcguHcE6WDNUXXJENp1
Y0niMtd1FrbAnovRNQPHzw==
`protect END_PROTECTED