-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
u1bPCVYgSU7O5UkHfFzFEWR4eNRhDyJBuVFP5r+gzavnPZSf07x8UrZTpD2nFvl9lj2sI/68RcT3
RfD14L6Wph28xqnSe1Fxiz7OZDjkkzs/r1k86u4vDPrGqZP+UkV1kkqARrrOgnPBWPbbfQrU/5Cj
t4vEaoZt0vHq468M5Drzbq+TNky/uEpFyVyLb7ZDFVM/o2WgmSthfn2vEUxLmGTXCpYgz3vDNAcI
Yumne1JBrCufJGrU33yRJRxUcSrujMSiaw4qqpoBBYzzwKW1X+rb4A7MPOpa1NaxDs3LIjFBo3Hp
atOrMXCG4NYIgo3wDsW2S/lKh7/YtaEXrQpHkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12496)
`protect data_block
QHL5xEjZY5/Q0FLwLaRnNrf5fNTwtMHT7EM0mhDcrCs29hvwEXp4UUGB85XcoFP2nQN4UMt+xqfu
78YI0z3xHpYmOuyIXMtqZ/TRk0otE6Rob8hXYc+67akuDZvk7qQfz4OBTXWV1607FIVJZApYakJ0
2TuDlcQ0HyxCzwOJcyheorNKTudwzfm4T0t3InpsiWkdwLc9SqHwWwpb662XewsglGpO+vZPee+v
/7AtXVHp1/3EyB9Rklaznew3nVvLVCgoKMblLqEasfC09Xx+N/Tuim6At4F1nicmgPlvIRvTV16B
RG4RSTaHM4J4vRl7l2hxP4PyltB4iFfiXlVyuF+xPRt6kGMbSa0z+7Y7/ACXyFupQeJDetaEXF84
tgwcxQYy1BRLUOIcSbpw3/Ddv/eM57WdYwF0wsUmFCLKHlED6H6q4XFz5pjMF70e0fsFq6Y/gItW
yDEChis0orICJWKv0LSTdOe1OCwr5dhymfFLdldj1VxF13NsXCDe9D5xozG8RAEMG+aLEK563dHv
mp7wVgkNHAADUc0+YCzE+rRXDI035eYbs61eUWEUH3ATkgVwYZaLEQn/xRGzjpK0ABfjSdm+bFOx
gj6sKy4gK7uJUzCP757vQs4aLQBEIQ9Vi105OkAP+kkrj5sqEFW44LuMvcvUq52oNjoFmq6jSBNT
CXZVYX8S2hR7LI5PUoNQifY1U7wiye7vk8iZXgoTs6GTVs4sv/uSk9BvHU9fT72/h481TWaTL2d4
UEMzZCnnBtsWXklrDPWJBLKrOcgu3v0qIyipuMHEWyWJvZ7PhD5YiNy81TKdAjhpQw53//fXlBbK
GipZdAD1p42ySTo3A3sNkGPb159NxbmamkJKDU4Ajp8l7TYK2aGWKS/kUMclm2A9XB1yx/faBsv2
gSD04X8tCSdqixd44jyPgqZlUjZ47s7gCQUUhvGLcXHdvqZUHKWhBLp4snQV1CtMl82YGoA07095
/5OIpRMXNJ+dMkhNu8uLUj92rCF1p2qpCvRnxGcclh3rUS+LjMgxutjmyNgRK744oaNmWCcMapnp
i+UibVRhcc8RUXktIGGOWUyXd3ROwDOyUkk16oEwBL6ZBuG17b/6nPJirLdFFTl5dBX4HrSL52bn
5T2/WGAuI/tS7QtfqHQbYcRJ76PUdF/UziQCcpF6bfB9q0ZeXD2S6XjZVhJ3WHJ6HH25hDWC0PP/
/DeeI28IaQYm77vgAdlfqhyji4CezsePbC8HGSXo4Gr69lnOlSFcTANc77lKbjUDBCZZj7TDjxAe
34MrQrwMWvHJA3q1kib90+jkzrvdHVwA9lH3wXW0wmEx1PkZTk6SvwCguH+9FzN4/WuG902pgvDG
/T5eG6jmRUJNNec+hDUWBSnNg3QaqosZ0qUyCCjUAN3aAneq5loOeHIc4K4C/R9+DMzLB5mHh5gy
h6dV+5XQfHwL8fMhV1pKpwhwcAVVwGHxwWQFFx9vPXnpVJoHd9hkhllhTuUNz3iiQTG2oQJgbSmP
uKUEMxt2AegtgJBTSeWELJu4aZ7gQ3vwBuRGh8y1MJbBxXvz0OhW+qCc7GkZ4hONpiynygH+FJp4
nyorxCfq66Hygpvgl3v3LgMO51qnlMMTTvf+3apcdEZLzY/qhd4UNuE8/A+GTh8PC3cdLgq4EtKg
BAy1xLorqHSa9KVEqKuvDw1ROAn4SOZ4uvNc3xOLC26VUBURYqqO6NY2FM7d9tz1REFZY1gi7sVZ
Ln9HPY0jv3jHT0AJq81qIot5iMKPfG4fb0wIyHkfFoRx86+WUN/5NJV5AhlBV26qOks4voXkduaS
4lEMjlD/FZBtxLWLx9Q44c1dPni4HJs1YBJ079ckdsyXmhswfPTcDN2jbt3Cm0Yy/Gy+gXwGK383
Bz6TYZ51ggS1u/l+1VROwJ7fg8BkORUFxFtgkBn7xSV6KKC2LhG2wZ+rzvckfSbRWhKTUpBTz4Zz
eu2U/TOIwxxLcb2gyjCIrl6GxfhPuDj6lUGUd3idJfiwDlKN1R7ZBp3MHgTlCKnObd87lcxwNNdw
BEAMSt+C0AgoXV0HJ4xNvnJQdQQSs+g8vDV1G36KoquwyKtD8CO8AuwifaPhaWMABWoTe3HBhxsL
etDZIacARCprEht+bshKshr4TmvfSe7T+OKLrhbj/KmwNvTOycgg3fBtSVM51+jGKdzoywJZqKLy
NAUMFZcImh06aDFtfC4OHooxEuT84IFmXpiL0SDDCNrTYAmRMavgoXYve4Zb/5rz7w9NYFYvPDlv
YuF1e7s1wVHDhzQY7wuDfhwy3KHavcS4ohqlHHhhjVL++euHAq3pmAGpAFO5Q5hP7GLCdTcpc8Wn
S3wqY03+hW/UgggCLg2N937xrzpVI11wgrH+WR8je7/qTIRFQddW9VNekSME+/S9cvpY9R7SLZn7
kRZs0f0+7yxn260jDgQfqYGZro/ds3deGnJUhLK6NGvLPpVSXySXI2DeGnglLAtqIrr6SHAvFu23
sEni/xlSL83q1hfMQeFNP2ICe92hQoqmdYy/hYEqguMbacLtM/vr+J539ZiyQ/DJ8gs8SaNRuQu6
AK/AVYiK7KjDK9RAdNxBLXVv2DNgHpP5fK9c2kVdw2ZkB+C6gs4rrvFguerYZkqncNSm+1kebjUX
G6Z5RmrgnpYYvY3WYkax8OFp2e6QQX1T+MiEpA/QCWTYajx0FgyEFD0lbldUYiOZy7PCt0mHu5cH
Z2pMKcBnPjE0IHLlBriUW5Tnx9O7ndlqF2BaRxV2QpePgoF8YOhM5dEpxl4xbgc/rtX9Gts+EJg1
xridja4HOQcyp0wqG2AeEcLAWmxSNQKETe9IvIolk+YmkTJ5H2mIpBRYiFchXaXlK8tNBNQJInwq
d7aeNDpQD59C/X6MMzuQJ2WmXDSDa2r9xS7hVlOQlq2vTqCt08nrkZFhwzJPq9h6i8eY6ISNXDql
Hq5F5J4LGJeJ/y4U5P1V1l8wt4QWdhrcJSA69WbYQXbClkPiFn3eY+fqB0E92sPCwwiCqu0mzzx6
VKXxjzsrEEHrKysCPuLh7Txb2aSYGvQ8+HwXgh/mWcrIc8SWSfUPen9/He9KyIMOpkyheKY49tjo
JxYkEYibqky6O2B/nuZyruUy6TFLVjeesSrlXxrrmcbMqFVkJQIk5VNj+koofSddE3DlXoPy2NXa
3KTdctwNvVYfA59NxyinYA0xplizhRSJmewzjgr65YcuAkvt3sy9GpCpfDiaD/T7uiRvLgK/JTFE
Fpr8eWCHtQk6UAERWh8AAhP4KBW0dS4ra3VVsztdylz40a8qGEQXZGHcCd9t8z7/D9wS1/r9q2Rl
92r4mkvb7nJsPuPdRkw8nNQL+XjUOceekGaQLHNswfaV9PSYT/RLq3HTW5H/HGJepiWvEZgB5CLF
Ou1hjeZKaeJbYQFUfe5TF15NZieGapYbobxYC0EjSDTKJl+fM4c2V9wBeprZ/Roiudm/jh0v0bYP
3gttjUu0kWZ54c4Yffiv6XFsLIn3iSS2wugRkGZ/QPFzAuZhyaoOvX/mjFrfrbA3hyUrWwyJngHV
Fqi/NQcmqust6XCXsB5s/0oIfQ8FGadiQM1VXZSeJiBeyM3XtvatX3Q1gNdI7RpMQCcvUJ2z3YYG
LhTurqhIlI7DvDCRloAMyiqpzhJOaqe+KYIDDw+Mrg/LRerbxIP/Gg+hlfiBqVmq2Rs0nU9/4c0n
oGWLwlETnNSCKZ5ZC9JeRMnYK48t4RRGhvI7Hxm/y1X579jJmdBfP2dlNihj35a8MPwX7shl2zQQ
3Onw98/IW/crzPWc2+e/GpqslkmeTuh/VvpH+ZG9ZhLRShbtFcN2++ro4JJZwuOJFbtqn9C5zuDY
PpHYtAi8iARGwOhaOQx64HDRbsDtE4B4Qca+ale/KKDrSIxC5iVL1WG2bRcKptvPoPona6GmvPd4
ynkIpkOs+VE3RYylJu8KyByByvFEbT61G4N2mtFp5T6iMLhMAPVPNzJ3Vahr47NDz09zCP+RFePl
76J9/cyDCjpuO1D+IXKCbyL/7MNSqjDwBPK1gKiXTDbVCNgz37c/lEbuKcpzp1hMTULtPPKkwo4u
HzDwSUflLbWPjq6kJyLETQm3iCmmZ/O0UCpG/WijmV1bX3oST6axYt0J+YxazN78/O8tC3LPxylj
sbc4hjBBu8uWat09tUkfih4DNVeYN/dj4ebjdqMgNoEka3bEWDS5J6sF2Gq+yElWmbb6gST+Ec9/
2eMC7EWl1UxMD7jtCqd42z1xBAGX+5l9hx14sfcvu8DguO5YeVgW1xfK8hKqBRVrnyRLPiUZJCCp
NBp5V+lAUDyjM7rBdFxmPrRxKo1NqNCjRSzvhGkFN7sal93hHTUozO76CQvmDYZlpV7ZaGkuKvcQ
Gly/tnIa017MnqjgBPE3glYtAZvMXk00ANCYqokjH0LJjlgekg1WeQVcqOjThXrm5tUEFKl2FnZj
kx+D4dLVXatmWwiGyxPlNmunghVOGJ0QKb68Iz2AvmPDnNxNJGutJq2quCoFm5rLExOuxb6px1N2
ZhOLIw/sBqtv+R6601I20B2EW+G1ZEfTckMQdV0hYBo3EoxkdtswrOuvuO1f8exlsTpq1KYtBObz
s0vurOhWq3a4P8UYGGRgBJ5GUQPWJh0pbEhwlGN39qkRDXDKoZwI2K8V16h0SLtG4LmUXAPdvRPF
xv9EzeigeLl0ZSVeDlUW89FYJlYgFGml+R7v+pddroydmFza6ayHNywiIqRPJNpeM4b3mO8gw+2m
MsVQIKmMa4nywWJv8GywkkbCbJHZDnUwsIri3dFHCzlJxwmjbpdMgFXwBVTnZNnnbF+vC9KVrEeU
O/+E3pWyNaTh5c7iM/BibmRVGVuWV2BP+gmdHTmMvmxzPIchoVQWJCtZIbcL8BD8utEdT7AO8Zjx
vr2Kx1D0rji5c28Z2rBZKjJ1G2MFKTpmWE1RXH+j1HMsuR1nloSa5lGpHKJAOAMpYqH66K/4iX2t
ygZLex+0I8Wh7XoJNz3LROtDfF0fGGSgNnWAOci63nUCyEiKo3VVGx5JWv82juuh6mdAiYD4/pdp
xZmldGeuzZpafvBXHAk0fAFqOVjIGy1k66WCRfKkr7v+Sd6A9gpS/Kov/CdlDELLva+PO6WKs8Eb
1EjIgz1qpXQlghcZ5lIYypB8payxl70qB8lwc6T7XiV/W4SCH87+euVSbof5mjwrco4XjyHZCje1
py10AktBb5Sd1CQ4bXP+sdm2iTslJxXuv0QMM0Bxce/rnwhRtX6JDYpeEv8W3WzpjBNaNS4v+lEO
H9/FByiYo4abXsalBh82IzBWus0XTqjMdCf9ker5AjkviDLPBsAa7PF2IbJCtErqzlgWrSMIKsGC
AOVwwYu4Z6MrVI0yWEBAN3lf7dxhR1MgGYOPlN5rurtLfOD5WuReN6r2PV5tp5ic07t2ZotRpY/n
C1yE3InL+UkN7otU2k+FmRRQ+NxcHF1NkfdQst1c+Mbkg6rYJ3V3uuevU8oFiiHalomYaehCJ3bn
Unirru0SgHcqLuHWDxko7otnaz8W0/nnHWqYfl8zwOnG6a+00FKM2YDve4ub2338dnJFek4a060T
g2bdw1ZMoO3onMnY6DjXK2e8qYsPDjR/ac7HZc16060IC8ZVcAwqPjMCpNcsBGZ/xa6cK2UXOANi
JxvrqCE6TX+5Wo+McE4MUAc4gv1BeTQ+JijaWVlxFwAarWPTSrCXzrXOa3R2WyplcTkQ2G+ncbV1
HKLEGTOh1bnSObutXtJ2LEm+oDKmwLCs3rgSDvjIaqxIzy0QFahbodpGdpi6JFUHWGWJTPgdXOvT
N9WLomcSiBaRx0QclBSiSOdNb0538QWgb2kSIJ+UbueNBYQ5R4uytSJXceiBlPkjxc3AOm1yglV7
x+TR+T66wMv75ZlMghX231NGoJCDoSmbjM2FMQ/LOvIlqY/qtW9J/EYh61Sd5rIg5WfY83ie4VKD
QYrV2bUX2PgUV8ksuwA2cUnyAiUcNKP9Zgu/lpJPep1L8Los9/O62Jl3PvwN9zF+fr1v7boERNar
+LdwBKpRUFiUNtQG7YmluSgg6MFqRJ0JYK6+VdB2Pz369o1imIvIDi/cQ3tGGj6P0kPEXqDZqSfZ
gCjgKo7GRwtEJi50ZnRDJnpZrlQxPi/svOvaob5P55hGUt1m6jC8zlFqshACRnf3T4uTVqgNTU/z
wizQSdJjRhZfTGYke4/JUCW9F4rKrFcQtxhblAWOEIiioSjiRLzoZTvVGSZ6Q5nOd0F8iGPcd44Y
ZGNdwR+CM4KJwAMVTuo4OHMUODZE6mgCRp3AI9VFKSeIN/4lqjb6hxrTTpJMT4ZJCiUUfR0KXD1u
A6gFZ/yR1EhKAEwljhFZ7+73R8vRahGkT8YYpg/E0LRIMjA06KpSnYzwp/BCmM5rNFbqjfZUv5YB
r4pwQIIcUVYjvJ4ZO6k2MRqigZ/IbiBgK/HOPtikMkH8jBoER4zZkqWAuXvuzApOPSHdS3P+vLzd
PoBvMO7m/yM8m/fE7F6lPXSihH/v+oIbv5VOiuA7VlkOTt/38PldOGD/P8i8lbUR8qLB/+OD7TS6
d0n2pXvZ8nIfswVOEOunUB1YLy+ZpJ3zG1mSLtznv1du2noxUCmGeSofcbkCRqDMr2tboDykcmDp
VQrhF3PRuVRgeA2cPolCzx/SLNlzgFL2HmpwLfiDN3uAurcYqtKJdF+txUZo4rvM1H0AnPQyWrBU
qdp+eQRwSFSZxLDYvZ+wZcYLt6m2ZEEO4XL8j7POonPPXYaxWHWdMflyEb84+zN3q80O5iGCzL1y
bcsYPObYLTXQX1rSnhF7g0X8514KPyGwW8DLF31rR0yNYL4rrXvdVAtjo5EiHVJMLqkObWFrbAX+
GEjv3IoJxCHSxr1fpjvftponx/c/Y+FY8SxI5+hyk3prOJm7JUSS0l6WACdC3p185kHqoBFwB843
xMjhvORUr/Dwb3iGzGXTgVyuMDTw+hBT+2NyE/x4Ds+wt+reqCwfptnxTD4O5WL2wtTsdhknbfMB
OkEu16JaTaEtpfWkIM6ifL+3Ke9kTf1/5zm9LemAaJ0/fkc8KetPxDtArbtEWB15wN0DKfzBSCbi
2hIvwNgkBHg8RrHHVb6gm/86zcrlepN0WqEGe84q+zGG5trG8aesRlYJCzF/SkP+VU/ACShbpKUc
dgWPRwj3dt63D35rflVEOKEH0RUfr+3nfiItAlO8KTo0IdddaykYy2KaXNagEMe18zRuOYAqGkl7
rBoAsmg3p2m+c8g8kxvOpqfqkMnnX8zqBecZlM4Up3gB5UQswkgf1Ew+cdYez/8cUipmLshvSBz6
+2zl+8+kDOVRFjTWIJ8Msxooc83MsWcnIxH2F+YoDPMg2JokiBqbnVCZLVZqPy78t25PmIvGE/G/
nI2h0s9XSFn0gbF+9I9HVbWO/f8OnUP6T5R67xQZCAh3XBCab6QIQcs1XeVufdmzTJVafa2LwFTC
RbxWZjk7a6pO6RNVisPGag1vwCzwQNkvND0irB7KokfonmD91cnZ4mUAPHkWYl7fW5EOz6Zdzpg/
ni2Ln6w5vw0WFNU5Hitag4Je+pzWj72Gyih/aen9taqUDogQ1JRKVFUx1QiJSLgpjb3ylYTk4Wa1
DsiA/+llWNodvFdgQawKgizirlMtSTFCfokkCCwF2vDwRHac7pZG1RQexCbdtHsi2oLPZ+D9pb70
P6hS/sN3FJyJBvKeSPWgv9ZUAXB43Hmeq4BGt9abZp9lyuVJ1Jba4vTCHN7R8sYweXPnqljCEsyp
evQ4oTePgffRm/XeaAHXoBf04FVpL0Z5on0PaOAwsHco+fWihOBnojgYpdwiRHmf3i8Qe3SOePMq
TV8NQIDE6iYtlb+Pc5rxMvmY4ZjPAds6J9Fx1lTAshj5Zrx564RJOzA2uPyYparahNn8KS05FAo1
HlUYRmF6aBraWxcBejracsqA8CoGRpmcGvc57sTfgv+oiL5HuIzB7tNPnKEL4iYCkaA9LirQW7fD
hhhlNXB404b3xzWTfIcDZ7pIiCO4G+NvxKvHGQDX6rHZ/YTmn3T0T9oYp5UcwAF1jFDN+Bx+EkQW
9L/HvvF6Hw4T4JqidZr+Y4EgfjTA7EBDt8Mo4nBr5ziYBL0Qrwr0Dx6hLM92gQUbj7zu9yEsuz+l
cPCGsHBDGBcc5vvajNkQB2qSWkVwj6iO9fp5c4KfGXkdzhY0sV+ZTZshxW/hYDVVMQoGdna779+G
O+gSLUvhXMTLbMbesfrJJlt536n+mhVXaX8n3kkT7phoeoihfaOtJvGhnP0JJ4TuO/eLI1G5hMiT
3feoEpeSYmS2uK6OoJmhGwMhglZDhuGbFRT9rrDFC6YC/J2FIHl36IAYizdlBsLBoV2QrY9VlvBo
qRWmWHnK4BQU/CY/x4y7je81GXySKZnFm7qkh+0ippRGqlnEFaqJ/4VZ3c16RmJ4bjaEdbSEEwG0
dUZt/7niIfLFqep2vUxPZ6kIZxkZ2aJB+wbWNPS778k07GHrj39tqdia1L4Qx9DDlzVRRusyt1I3
ArIDICdpL/l3vUd2iTW6WPSzdEguogxoQmw3RFJqTFDacGnGJIYXTi/v3Zx/PDC9hAVPCG1N6qOg
5xomH4uaID5bPa6UOmH82OaNxZqgYUydR34+buXm1PLHEJ5toJT6qXGfKsstd8wcjel7zr8FVH9F
Le/ZmQiPLbX6Pg3qrOLFXt3ixDOcFx1mxU1oENT4RkzE4PUApTv9haSfStUXI5ESgIUU6Ktdzycw
NDUvyccv3kKkgDqy1r/kbP+E84D8RM6CW0vWYvzqFeRzGbWQJ11LJYaQF6wiv7998p8lIHDHwlpU
I1O0Vjlh+NorJZDKdx1HtSWbfRFOypZcDMqwNL1tCP1n3fEAy5ResOT7x7rHKZw4kraJ2vMLIFxs
XVXfz5PTzJ96cuuNnKx+Cd9h2x2O/mNHDle/k1JH8YO/ZhminYBazPg1oS5vTmMQm0lvdYbt8BGw
7mVUVJzXsFb/xZULOhSRS01soLXQQYnaIwuvjiWEdSsJ+G5mKATWe9OtZ172BBk8raBN+LmJJBUa
TwC0RRZEOogwFc3BputJ2+cAeUigUWpw4j+ATALRD2SaQwzqnoWbQ5sIjNfWqlAFoUOQwGuXXc8P
VmXkgM0FL06Hi8zy4ULJlJicIkMNQLeRfo0/YtSH7pf9RYqB1zjzaildcHuvO88QoHnT12OaANFN
oidXtI434XEh4oPuXn5vAuz3/tH8faWZwzNX8CPKRZlAOsYCXpoxKX+nVAYcDnoc25YQEOBY2V4p
aZ4WrMLMKPp1fw+KjiIuTy7BAaZcB+B1Dzg6c9k5ffSfPliiQJiLQDgmTs2wI/0Q0QNPvacsYO63
3iRfHf58ls6CyC9JVXkBnCCGjy8pvnwv8NOOlYzW21wPB9AARcJDu8nxOy/hp76dENDDpXiDI9G3
SmyMSjTHUeDzVkFYCE5+RKXLNVgSAlLky0HErGJgxvf36Y2MOG3MXC3rGw4cSuqZ5f0K1MluYvil
NoMC16dHkmwCSoxJxV8wSRLo+iOXtPCZhHjaHFddxWfR/ZBDL2aoNh3546cOSv4lAzI+79NC37+r
6nNRv0NcvBHDnFz/uVJnNizt0kDBd9VXAra5fukrYViGFckfDRNCAX2EdfTTlCTr7pNb6VJbW1LJ
UvoNrUoE2+FdUsV0stXwsGPmfYk5uHcHmXuqO9lAanzz9v2L7P4Y0PvGtYfjxYaG+o6tMBeT8RvA
f26tFV3Byw+bOjoVolyMh6BhvBU6H2JLMIt2UwM2mviNrR1rzEc5k9Yb3dRUG4ACjF1cnhT1mimF
T839HxGIvCaLKFZKO4C0f0Ch90hNvGHy7p9saWNUWnxCX9H3aentU8nNXVLgQiT1XUO+WB4qR8Uz
Mv6pPxURCTobL5hyAqlUzLGichieeLUd86JB0cVry7PA1s+Hg4BeHiz2WEcGlukuvmZRJEzYtrRt
farY0eIJfT8Uyfsl0M3iPvHNcprewvqSXKz9eDW7CcftYpiCeagwO8qroL7XqQTgx2WdgJ1poTuf
Bw9KCmBGGtBgcLCg6aMWuv9pWY1xqvWHe+pFLamHMvoz/sJ88//ZjWyqq1d8aLSXJIiXJhNkeJ+l
mW3pfC3uqRlyOlIbjpopmwx89cyR4eQ+5pf7Ng0Q1bx/junsIkUNu2kaTlgG+fSI1VzF9ltSHJSu
3RG+mR9Ip1u1OSZU3oMaLewE1IZ8QKnt9kvHxPJOVGhuh8ugbcxHuAYOadjDmnTcJKRRtH8pUY1P
nXrwZcSWNQiVGlZFiPdfWbyC+X66kyFqLQQeLSjEZgjiLOYB0fp/Ni7T004KH/FloGwerAeocfpB
cvolno2fBTGQVwOcfg8EDb+qX7Nm4pW8Llt91JmM4mb5E5bGMBYZImRz79egBOuOLQDNpGDkFNBq
iMQIimaFOG/2mx9VDaDZZ6LSCfi4jeV9t5dculhOonAQO0q09QwTjrXukbaspnoDX3KLoxYHeilG
kTMxPFFoTZgsnmD6zX0Xov7ryvzfG3KT9sMXlOswx4lRU41CqI6paRzIXFmLyxQIxdhKxUNiPVG8
fGeo0hKFhKOCIi50F+i2ejo5FcRhG6tvYAR47bT3laeCEkJR/de1ZFGoa/yGvPaqEI1/nx6y3Bxt
gRMUHs9qs5xEZIuh9dMfdQavyIiCRC2txICG8XZmoz1YwjDxN1QNVbOc8bxrQhYeXI2iuS725BQx
1NDryjmpsks9pVhRpfLfI7II29YoCnA5T3GIcf8Jsrybx0pQYEBmgohgT/QibedY5shOsnd3l6/N
nKpMp/xs0deUJ7jxSsj95+b/ghq3j85XUmkY+1NaEvSOlgb3tNBl20hZlkyshG6tb44EEiOx5rvE
TO+IaSDeAkXnNvqSXo9/czdCdqQXPkr8MJqc1ABobBraV1f8BQe2LxZQ/JmSzAHYzInqeLmaBWWe
0WQZjfKx+opdZ7vshmCxEoOF1ONi+gUJxzpypr0eIIMexRLsXzWo/f4o8nHMoRFw6QmDPLKAI0lg
bwIxcarlKxE9VTm2G1UDCbSlrcn7QsNoq5Z7z0hMXi801RsLBLwgvnJu+3gOwfUx6hTXGOHwolgk
nB63VI+7gIZaGbUeu353gBzq5DyV5hXYHMbMlpQiH307F4sKinhzNXnG+1HZtcrpaFlGO1duD9H9
OpVgIZwwvrLwkTIfdDRJwrGJGbTkvWS1nRw7BJNFeHsrSXemOFPxtFZe043IxGx4D43yAhlea32+
oGYl9vyR22k+qh0mSdMvItwvi7JghX3QYmwVGcReGJSUoE3g9k2SVW1/ayH/2IxURZExf5bcPeGH
PW2nmRnkt7DgJmAB3NnnhcQi+JiROEvqNDnYKwWppbvVmDfiFtRt9kcXSlNHbhmFUjnSyY+sAqgc
fayPf75UO/fHuKRhcY6z4e67Fqwvl26svqmbiG356ohMAzXLcbm53oGMlIHCv6NDpbfv7uy8SVdo
0Fa+Tr9rzCo+lVh7PCrkrXQbouSd7J14GPBEjN8V3aXYtAhK+afbIXvrzJyyBpkRZjXPgr7lwazP
99azUpB4UKwCJd2X75Qf4SNTm9afSlJ6zPEbBkUIfk4qme3QqSRjuQk0g6V32zH+Hue7wkP1TcTt
K9yButtfanYcDgYfR6bXTp4SHH2YLk1RKLpLUqvEHoKaYNOFrqxgFP6TfD1wlCIcSQjYLW1/Tb+k
jVNUbGam7p16s9DKsdZ9YOxt0507Zn3rP5uIabyBhHhi6KZj5g6CJw6qBtWFZjPg3BAszP1Ly8bx
m46svGM1WL0hMezZqblAXi6SahJz+bRmpEWaVX1EMjzL+kldHsq9s3t83WowVsdZhJnRKn6CsTxn
LWxdgtLfyo0h9Qt2oPI3P72hdp4B8Ge8Xu5RPHrwCuqb17HqAaJ75y1Ew81EtwgNV/IG0AIuv1bY
65OqqU+4/pGR93I9GxkRBFJb44JifDCGUKz7n9448iAtnrCFQHZzfxg8bbLKjrQVkDRFvgLzb4TF
Y3L16JU6sP7aRsXHDEbB/4SHuaFhcHTtAknZNLmecxyCWrghldycxs8zd+PNzRRkfw2qPB4xPzfn
n8e/fHdTKAouFD6+VV9Jir6ET5AG1rg5PQf9mH4BYJTTBt1TSLES+1q7pHPn0g2fr5DrvHPaIiHB
OUZSbKq94bSk0gj+L1RP4LiDaox6P2RDRuAfNXLbMkDbnMqRBM7XrrbJa3QxtdYwP7tbDtrUcK8W
esSRso2GVOp95WH0r0YrFIrlC4/BFXYf7jUFDPIpJjj66C+vI4d9oodvrG6aBX5igVQI7PWK/pn8
w0pn51Kq1lYic40nGTO4bCNzYmOdz7n35PX8iX4dn7k2cfppXWr2B3oC6oGyiFQrjQJwYU20lkS8
nZ8Vcmozu5S+sIB0PnQ88mvYuumnpkC0sDoTokQYghNiz9ZZ67lCyA7cgZYuu1T3Uhz4vujgN8fO
xyLp2YTcdXffmTizWx+3gUQVfMWcp9UmdBkAXKJ6XalATnrlfjjqta6GmDcqguBN9uATISwxqSIQ
Pap9KGPirP1q5CpUaHSHyyA6Jbcd1yCaBBUp875JS1JTupBaHaK5c6LgnrhOP8/nu3n4mOFlvJY9
jruWaAiKB+LXaClU7rF/1A3nejw38lGeXIfdv301QSWyg+Wl486sysOua9rFjI+a64FeraO28UV/
rg5ROBtlW9YDk1qH0MKipkpUA3aIGBtcVowNAQY5hMVkTL5Ex9CJ7YmzLhWy0lUXNRyKqZQNCqMQ
b5ASQFxq9nc5j2Z5AMwr7DKEa3Fw86XmWpLVbru2lt7MGu1GUC4y/BuIsmTOggodf2TYXeFsgw3n
UnrcHMg9L31q1xNZHa0IEYZmp5xrlKMx4iP58viHKIx0cssJgU9cXtFLHWJwXDyMw4A63mdPSMWm
ssRejocaPQsSiqVl57s21YsZVNWQK+5yX2r/oKrBxqC57MECXUtvvLjgkY87QkqIOadEvddok6Jv
3hzx5oJVcRM4DvSZgwMw41/ZXt2fyKZu0IxxWHIADKSyWmtz4othxa3ENPrLPbDRvlbDoA9sED2I
/izrMQ9cUxG3acTRGT6ukoxsJubnBz54RDDOmLx4P5Vqwmt82X0OsPMy7s7LxnFVT0T3kztK5cI+
ifPEWqRKNQPzFYXyOC8cPPVd8H3vghXCKLFM7RxazpMMSep2Asf9KF8logJe95zaHJQhhEwdrMwG
93fY8ANV3R/pKJGNiPe/qZcpzF1VkM8kAOP1Km2haZdRP7mvnkOgOyK8AgeAEEhrkk29yS57i+PC
KDxqG8oMVuIntDhjoPLwwWB3czRf5ZhEhzOp1/no3y38CGA9M6cSE9zZh5dMPHP9xkdxX122klEy
2xIiR+jyyDXP1EtJzY5pf5ELIdSfiJaSiJG859IsrU9lKz8VMzk3BiTAec0SlemhuFhZsCE32jaY
aPxfJ1h92r913A71efr/P3t/SlX08+/cZVIYsBtbiuSN3c2ZTCRpEPy5JEFvEUd+eGJnLgm+AJop
YVFb7JUKF8S0h/TRy6EkJeEhqWxZZ+VutLFaXuPPP94CjM4KVpa1Rf8JMbGPleo2PheMGps4L439
KMTdudGoDJuyhfcUOPai4bo2fHo3fymBP1zQp36bmmYiqvjXVzcEOhYKOnDpoe45RooGhiJC1QQl
Q5beBvC+rq69Q8XQ+77tkj93NLOBmdAihTVjQ4yKabfqUJL7Td+xokxx2NF3j+M2mOFILzvrXswS
8Wur8Q4ZD88EpK5Z0Z4CVvlCL74u+J02Yw8MReREDfiumTTVEY58N7VeJYaYUSO+AX27+Ll7HV3U
jSUKxuxaneuJGi897q8PGTFR0xbS1e767prXejpRJjrVt/UijICkO8U8/l7kdYwqWJoDulkxvR7C
EBqi+VtuVDH+1r722Rtoxv/IHTwt2SU3jhBtJ+4xluCYZX30ZvpuOOdKJdcIp3UB/1fp/UjedUJY
p35G3ta7PMokAmfiT8Od0m0RRj52wRhUer+NTCPM/KmfEN+UAdbd/6ElNmTP830Kcn0ArjfkIIAa
6tZQeBTTmIoD1p6rAqWUkDOUVOeWyJWBY3594tIObcMuGsX8W83NrcxXiPRPLfdAiB1CUX7a0lLi
yR8CevDR7rMxDf3/BhStsdqOkhPh1EfQ3t6DqRzpgQ734SBvLM4PYSXDCQRBVvM7duXqaMbSyf1g
MbQVYtvP4ypCnEmlQvhji3vUtzocmBlfnwkiMbKdBPkjt25BcuDb1ZqMZez3PX1uL9rRZGMgpEGs
Oet8jWNLXsA2xN/rdOnWYQjK8NdUPzdIfYUK2zhTTpfslLdYqAKz4u6LhbrrUZ34Q9sIU2WnCpqh
Kf3Rq8sk6HpfNngaNDv83TcGvowa77v7/qg6isqiYA9bFVKLHZjU1py+xAwMXBAXR/CyL4KjoDx0
59gHvGtzAL06ksB9KtfQihjLuLkjxrMKQg4AvrNgTkKOLczgcbxz768J6oqSU+0hvg5nkzYbW1DE
CR85mFok24F89X8vxyQRWv8PuCOUVz188yeczsdMh0h0TSLDC3EheJx2coYKL9QUyHZvB6zywJvK
gqoU4kuzxwP7cnA/fbM7pNZlbT5V+wdCTwY0S5z7hSwQ7Drr4rAHnl5uFL8ZjAbEr8Vwla79rvrP
WwwrBiHstlJwZin8imRPeFDbVWbyZXa3XChNUL75/h8439eo0Y2beTUTZuq2WHF0vWPfSkOiXyuc
P+NFpA7PO/WwFPwESBBTaV44sPeUInXLcHURAFxLsvfG6v5VzqmCoL2TdMTmm5YyMgMY905h9PjT
jJp8h+Ww9qOwHDmyyrP8JubR2Ss3HEr9zbubUCz+suIMqqYWMHAJPwLJqgGsLOP9/6jdkSSzQIuI
/SnugBficBtSUmPzN9Y2Iygajz5M5Gc1XL7zs4U0PdaZjNuafPV1JeKnVPtd2659yY4lKttobAQV
Ym3mjNbX7WySCVpdUUmcPuWaXB3PryMyV2Ufo5tChVwBmG66krfG6Pb0aruFWN8zQ4sPSX8pzQoe
HUvB+ybU0qc+X19Od5FcWxo+XSLu4o5kJhJMbzrXOaPG+EoAGgIAfFc2mYJLwxU6x1EiLtj3/vfS
QQ6AxV69keu+B04qU9PUKRiq55/A0Sf+vv2MZ0adihpqMBrol3PPQqHQdofOJMRSFQtiXfaaNs8m
GogOaose/kJ2AXDWJA1m8es+Gj5blVNBakYpHGaEk3QwccTpNiinogGy3ozOZ5i8c5R1n/aZdInb
i5VihNtdeO2DAvhYwBLeuKvcip8oMx2bMhaUqPPDQwYRzlQrfkjJJ248tJRrN8n2yIPJL5I9ajjd
zt1kL5iGtKiJRHQN+n3XqmYZ+iofzYmAAX7bd09Df4Ur5DaUBOk0QkEON8llCIcplFayfwOmYU4P
o3pvmSyKBOUEsXxkB7raRyRF1wc1ilUkReZXrjDBdbMW830UQkyAbM1hXnM8bwq3U917rNTUqzDx
tsgA8BkIiPdk3wtHhksjOeJMpwCpADWrS8g3KXmQP+RBY1/ZJQmI0fJUlMuXDcX7yE+q+qEGTk6Q
m11TeK7zxwsMPp2mn0GrMMylTuY5TKJBSWW+m0UBgkPRAUD9BVV9TnYNWOxP+OzNJQcf/MEGguy4
l0WP/wmmaSgwegNAuUQRB0yBBAHEwxChHnyquiHI1ICLEN47nKehzuMjMLq1BYXzFMvvOpl1RVSe
AduG5jshMPsWWOMotY7EQ/A7Odg+TjbkveCVJ7qb0saekNO4rBVblz9GkUcGpsMDxJNawV0nfUZM
P+R28RNnFKtiVeSQQ3IAu0aHtcHZkVBVRXRUhEoUW467QB4rFoThXT/3CUYh397f2BKVDjfWRH5m
9cAAJv2M0pkwisnE5KiiKWmwgx5T0iM5kIDS8bVT+dYJVy5eaEGJ7+dii6VLr06xJw+Gbw5bt4t9
hkkKR3RCxm9ZWZwfFvsWanEf65LEGm2kUdWhGmaQ3KDoX2oTKko5hnMfcs4y0df3DfWTZHZ84eAo
uk7u1tJ2ISn7BWS9c5RGApErdj0I3bI79c02HO1XzYKo05Iabw4M3rOKMncG3V/+6hClXxUpHGfc
I8APivpM/GGXFrX8hYTlOpErTfVz01k/OaBpDwf4P+ti/WuFcAEqDoNCD4oWvlWoRyWkO6Mv7Brf
c4Vhxebkfa6nC//xB972wSgBSwRWoLag4X8u9oEW/eiLJ+sw6xI+/EH0M+bF31AxuuuEWs3naDiK
eyqDuRC99XlYzmh1XvNAzDjE4P0fJKE+yhYPbEXU6J+WuIJ7RPAj7PDVS21z0tEkusgpUprRtGce
2tY3v8GR751H+fq+mgBMV5RXygq3HARAMRJU6ybSgHh6GtLkF6rRlcsadUycLhutgtjxFPc9Cfdp
8qnNzBWyJyvv/J7TP6lcZJeWWxngzCfyJ6BwATITbuxaueg9AyIGWYIEcOmV1x7w8njG5A3hphWz
czfCfE+sylD37Wfz2YchWblqdM2oIsD9N26uMrkjVO52w07Cu7QA2Uyq6h6rfBXTEXiM9nuxhrQE
6RkrwgkCwHmNNmIu7A==
`protect end_protected
