-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IN0REBcUVlc7h2wslB2HkIkKFceKkvQeVuAszQXTwErG7j5MLDc1XaTSqWUYPR9/FzNsxc847OSL
sjt03GkVtl0gjWrdhX7rAMuniq9RqWqz0m7093osI03AH9QQv7Sk2UH7u+glgDXYAurJW3cxEZAQ
f86O1MARdW8heZtVqjETutpepMliSD2nEAYbYervXMWJ67ZC401Sx7m8cbroohXzjiLBg6FxagJe
ciz1F3/DKhcMriy/ecwTsj5+R5faix0xUoNPxT+suMNSdvFzBd2keUQSQ1vxgILnPzRHhQFxwukH
Gg86dt/zyUDaKuwnnmqbSAOoxmaFN9XYNKLqzQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
9kszrfWCdn/Q5Gg4KXh7cSCvv9mAysSTNBf1Il9ITzDsnmnsyDON9+PMtQKYaT44k7lKRpaE5zUp
y9gPgPdg52GsgPOavQzXqEqH16C2S8bska8oOz3iWsW9jrdKk/Qz17qI8G5sYCF7F/LauD1QJ1hP
QBmGtp3FeXZ01Lc/I1RR6ZFGOd/ZMMvacu6eKMFPbfLtf3WHtpz9LlYrZ7OdfQ9j4GeRy4So1H0p
S4seCPL8sUSFB0oLUFQ7JKbsbDMrqfBxZt56ekzt60ZtItyzy/Kr8jyRLLdm/CVhtjs70Y3ilKpr
Y3kRi/w8z1QEkRhF0hbSqbTPEJgOcgLVEdP0tu3A2CXqZI9MjmJY7wUnJxoOOjBdgNeLmq2V2wk0
FBwVZOygpp3uj7lQv0BllI+IVRjXM92YwYK2lF76uE+LFWvOWLiJpHRToRf59wCje7DJZNIAzipC
RPkTFHtHi+eoZ9oYkKx5i/17eBNaGe+H3DEwLCasV3IiyuIv4mIN5xEibvuG0nRhx3WAAKDXPbsB
mfqmYuC76C479EBx5veyGi6RHpI9h+Ek61cjehYnMaRlgaKsNGzzWNEDRlJl3hnDELHCqF3lA3rW
PQ5I8BqucQjNQv7+nif1Dr3jomDZtaNdkvKqC69mKyIsHaGtlFCKiy/XfqZEH51D1nxSUy1y3idc
WaqqPbrF55xBcKa9EFopi148Jjc05oRxn94PJVA8L/+4E0RSU0KsBxHZhQhJ/NmvnXvILoejQAlf
TIsK77oHsLrfHxpLyFlTrWYLhtn7yJWUF0/F2qrdjhNnc+/V3UXKNz/vPplOq0fh2b5LZDyQ/rWy
KvPp52d14PozJX+EwOKvlDlTrqvtKYOeyAKsLsSDniLJ3M39WKcO58kLGPU9RJACUtAd7j+V+0s+
WgbujxaaBcMzoXDSOgsR/wWXnLJZLgoRtANUJjs50VSC2o+t0alsRlpeFYrssmKGJH0RiI7rnLUc
o3dZehi5QmByG7LV2r0z/UIzqnBAZ1fMCS4agSrKzD4LRn2zI64Xr3mJ1ZuKBNgcsuye4KgOIBUG
pWyz5xjObSiDZNCv3D/5aH1aV0JFtefBv/DS0RLZ1vreHFVBshfBeCUjCcNMxyY20Gy1jdpse6OX
ckILYKngoHLJVURbN2XJvGSbFJJDZSl5IK3TWBzvums1DKCrSu03M+S6KlLTeiVz9lpTx3M5keXu
KqpExvkGPAmn4QOpdj+93TQF1LiEQ4tSmxNUy2+yYwn0CJFLusXBwUQTP+jGs8sGolyVPYtTVVn9
Qztj452zqFktalnIFd8qP+pWe3f8pU3t2ewkIry8wfCK8oeRFVVDnNSkARNWTZthqkL7/eVyMXOa
WK4e++XDCBag+EB6ggaSuqXr5AFggFzlB43pxitADdwDnQsed0DI9yCQejULr3eC2aT7e0CBPcy4
ga7cW0Qbpnbnzg48Qzt2OUp4NKGpJRMtbDC4LmNj9e9ClmCY2ww8Xd8MdjWjRQ6wWwGxBpRWKfSa
F8tL5Ex+MqOByULQPqHqM0mEQAwCRSFSvjpEK4Gnl0vwNBYvpMjRBvPIoRJcAejuO1TSml22Jgip
GYomtTtEP8Ne3cqrch5vE2B3KxEo/HnOviabRznjnk0zyC81qRn/P7BZSe7wt7asRivVYaYWrLH7
BhajHFiTkKIsCv4OvE0koKnhVHmNzLTTZU/y/4niain28KowZKQFGCgaGePp5QiYL4tqAfsgcn5b
2caEeOrHLuEhLtX5waEcbLR8t2Aq5v+2pwAPUOA64yX0vj6pBO/QUawfvRPceeqB9VkIWaIgmx+k
I4fwonOYmhJLavmJ1Yh6j2rqxE4d1MzLGSXzuAQre7IV8nBEdvoHQuY0wtX7WlDO1bFPFZq5/H5p
626N+FKuHeARXOfGb2K52WdUNXYnWko/92iplw6dF644L8eAhfaCmFdctEaGWbqd+tmqijUZrPYA
kz+OgWxvfdLFef46N1QtnnerKu8lnXbcbjwWdlMIKA12u5QwHPNrqzmDglTC33oyZOuXENXrPMsP
vfTL1XD1/Dy/VMoQjuhi3j8QvvaFgq18YQtjaEAREt4ALMeQmlchr5122hMtwvIOzRaBjYuA+Vkf
ymvjCb+21oM1lF4K1caO25eeVxQ9R5njCrrcycum34dOklwoC2P3OFDQblX3qu3eeYja/Zx/oSxh
v9IZTPSj5fw15p/Jx+G056eUX2P6/vrNgOJGQUfdOyNjjO359ZrYWv9aryFgfaC3Oc/xRTcBnlJG
Bp8PeChg3lG2YmbHTdFXQiN5GwDQJYWt8bWPhKcINqrqgzJIpW+HrjMNVVdVvZZAPAI/o1biaErN
VsRSX8Y83kVEq877pHfnP3KPePIp1br1wKApDA2+7iKu30HdLLcGaf/i0tr5ib193ppzAbriY0hm
mfSh2mwQaqzaeB821LknsvCZvmg6J1KrSsGFPs9+fzx6a3oZqWYCUEfAJZaXtJ5uf59Ry3SyEUBI
oCr0N9oHJeZPyA6o2dyRBmylMxvoRkSuShm5OCET8gHiahDEpv/ooQDRkZGwonMrIXL5OnJIKlOO
c7/UowKrUstDrkhXZJ0E7Uytbq3AHE6ZwPNx63w7ua2lI/3s0PBZvDiae4Po9B3k9ESHFtbIj0YF
MuN7w15Llkbbta1II1W8vccKsNZnFZBIx8dreKWGYyxhCoriNIaz7hNPyMCIfJoJXDQoAlBYkM4A
mWNLYvZqNF5T8mgM0SnSUylq/MZqOCedpEQEYZCHugIBeZphxDRiPW3mMiQtnJtqinLITzKdtu8M
SHqSiY3nXQnskO7d2a5s/sSlYSrw605N/Vi72/v85N8YlrmpNNHklnPHQOsnb5Op9ZveOBwGA0cH
TjIHpCZlXYmptFnUqTdw7lzx/o5SZxEqPuYRJGxyNv9+4KAukinhCrDxS9TwrL/JnZfaCqx1RHla
ytp8FhPLXymjZcu44biXvXgPuEpWgAlkzO+l4a5hKtwz6cfG11wjQMbVmFURQh9TaIMI3QyVnze/
9iTYnpKVjs+MUd3TdhX4TWweatxT9p/yICklh2xRSy/gUdv/OJYrqH9y5eP0c00D3xU+HS1xOSY3
0fqZcznFRyqooKtRdzlfDc8g5Hsk0vAlm/q3qPZMNmwXgaMbduUCcbOa3wyUlANbCZ7R2pb81el1
yIsA4dk3RTRkSSu8bb8iNzl2Kl7GEM+mWUftCZteIcEo55EXkvfyoKBo5J8z4v5GX7SIq7eFFrqF
MYT3rFDVVufSOYgAVz4Ki+dxWOXZHj/ZxDJnK4mk58BQcthV3VYi9JdvHSeFJEFAJanhFgKSYDZw
b2yuTLgJgGcV1SO1HJl52Zc9p/Gs+Q5FteJ224fg6GKarC9h6oGGd1q170G6UT85bLo98Gd1Dolb
UmOS2JJ24Qeq6yyu4x5Dc2tY2aRU+XAkes1RZtx9wKhhrSlqaLiL8Fvgv6J7pAtN9hMgkIpxlh4k
iMbrsLPbdl9gILMXe1Lf0SpdmMXn41XrS0+SBSKzAtls2AeRiR/zvmwv7vesrhXOblePLB7OYLWg
j3N1IVGmDGR8BM1ieqC9Lkun2e/TduZjss7ow8FYHDm7IehDYreiuhFVa8cXixBEGHUbSIITgITS
XV8Sf3LxpAToDHlK2oHKtJsBDrg0AXeMuVhyErinhtnIMBp8CLLx5rlMgGL9CVygCAI8RWUi9X7i
Nvk/ZDubqUSwnM1VQtXJa3aObLYCTDU+5MbSW6ccLs5PoJ7FXJmacSE0HbZyJ0X1fEUcUS2ayrT3
aZw8OEUNXbeTotH407vwZHdfYv1lckF5UK53M0TtrZSc4kHmc1okhKukZnJRoXl1V9ZVp+m1AcIk
+LtdvOqn9RCxHfuWOS9lOavQHwbHuwR0J0LkKZFjdGuHzG2fN3RLOvVt0kqDUBZ9kFC+cFqLhdAH
5zQEeOGdTA1vg+/jQ1A6dln7Vk2BZy/WGtR25t506p7vPBo5EXQHR258a/xkuAAq+GfnbqIzPdru
PcruYsNBhGRtKngNV8hJNUm4vrUS1Fv9dXOKlABI7luzwtA+GQXf/1CDSkvFxP9DSUioN5h1naNe
6zIGADPHFrEhlXeMwjcLAASc0XERmipax7sUQJG7QdQ1T6CpF4AyEvno2ooGi006RNhlSQ6sBzeG
EYGQGjAjv2UWV+FHqYIJVduJMMcSRPGm7motFG268fS76erloD4+5aeIT1EsEVK8bDksjBgsDIDD
ianwh7+OdRflABY/XYdN13wJLk3913sQsx+mo59lGS6+xDomzB6/c5QtAQet3012uZ+1axKdEAmM
1XhQFHTZytpDl4TbEDpa66gstZT0DP8sFGpU79O82GHbcNSXffyY+/d62sSG2R40g4JTXXGfc8W/
XAn1bsru6E3rPmHevonTYVDMvlhSAqrVY6INaf2o6cD3orPZ3a3M4xMleuGIBsrA/UZwzb4pCx/S
trNkfbraRIThRkacoyh9z6BR599k7/JigjDbaabrTJCP8C7HaddLFkLr5+Ix+EqujHuBMORhp8U5
FaJkG4Z8ZDnkXl5WqnU9FlVxKQJuiLFc4v5rlBSLcXrLzMGwI6ap5Nrx6YnwyIl9uopWmnU1aU0H
lRfZmmKxp3sWUDVBu9oTCp2xsnP9I9IIu/Jc+XvngReJgMpPoXMKZKis5tt2Tur5deEJznfH6cQj
7EWFNOsJXldmrwFcYQ/6UYnfWJ2aOshwFDj82jnE6lHIbEW08hC1YKXmX3tDiIYKJ4c+TsJh0DRt
AN8WDz3fXCTdMuvXzKZzgxuXPKShxjif1cIt54P2O9jFAKUzvGqjYezYDT9reFBLIlifu7yQ8A6v
o4h0pumBcYfT/Aeur9MaAO8xASnM0Ae6BTGH9GJNfR/IsMigNnRKznRSskVUJLWS3ffye4YpCK0S
ds/Sn75CfugEOaWKCzMmDi/mwkgm3DfPmc7TGYP2yp3R8LPy7rJmYur+pKhNS+EVrhcR7cymFRmO
3sG4X0qKK7oSulMdhboMEBwZqskJ6EeJKqT/t33XdaReiieT7nQhg618dNobRNv69DqzltBt0lSL
TvKO1qYnyOyJ8TeiaULgWJJOm721YjQU4lrQH3npEb/POV+Sb6I0oHF0Zbqk64qSFpdgp5eMFU9p
0HnR/dpUpZyZ/x0+sMeuIm2Dya13stjoyEB+LahoY2COOITdK0mVKjia2xzzZ+UgD3r5Zz8lYaiB
mMXqlhXsbQgH/Al35lhrDr4QKi5rYNAhe7hQSXzkmM/JX/6OycvTJn+qFmKvNKH+PjYolBcIok5U
byz2lccROtrLl42ct2Tqm+YBhjDIl0RSa1iWZK0m/jDi8HUxG87TrpgEs92z2rMvqErM2UE4j6KL
Dso6q6bTo0FFi6cwRsfgXMsQa+7V2cCFXbfpoOvZCo9kLxR6x+w2aE3HcHvVkqh6BNT3FUgeZMo/
P8JyEMQouoP7pEeay8+n5Pxx7sgp/c3D2PZyxioiHlgi2d3yjIZx3KVQqrZnrCaN9MEXKM/FpFaO
skr2aXl8o7sPRm/2P0gzENdFHrQv3HfV1QsX5aEV2tN1paQSqCg4C0yUJIi50tWrVg1lYpxooXse
HwMR0XtiDgJa5WlM95xs26eO/ps8FsrdlBNauxnA3mdq/piA7osqZ0b8Z8etXcE43nyet1Y7RMVF
PCWmpuEZ3+UkJgDkDwNFa0Bie5igAx0mwBPxQdDdVnTgj+fcvX1YDlVDb2aBuKMstYMCZl7ltoTx
X0nkslk3yywtYqu82g4ZKY0xWnexsUchjOuAk2NKnBLzr+pmvsd+VjafWcPYWyis9kFtuYBZ6blt
EInC98MdtDI3lXO10fIsvU0FkZKomaiD28R7nEa/17TZGQR7wuQJ9S02uLqdASR9gIm4al2+Yvz6
lxM5UcvyvQsiM8sSeDIPkFjc4glmMKhg5bcLEIh+KDoCo4eFDXeY41RVkc+02t6FGx9+G6bZPZwj
LphD6XcveCyqRqgkVKvdtOb7mVXzgs+b5krYgG2Q35F//9CJ5sKPhEoF3bOD6lZOyIXfPmh3kc6I
KLs5rqyuABb7NzESDQ1FwYViaDHx47qwDlQ6Hjc6sMJCWdgT6o6Yvetv+I7C1bgy9Um8c3o2lzg+
TU3Z8un5SI+TPDuLEm3WsBMrwr+ORjXd2BOSrHCEFx2191h9PDaM6+DRBcdwZYPSmWd90PuDZOKR
XUayRXrvQC+dPpy5YFcgvL3/YDiukmWhAGyBOkBWlFX7OF0RaldV4aQ4aHrtGhryzRrtAxfhrJ4F
Q+SZQaVvsEHPDDa1BiqyGQ6jWGxoicJI/OaTFrhZhNmvakn5jkD1U2YOTkAQcb9g+NBKu8TzOxJM
DM9EkOZ7RIsjkqizdIyM/UjyPbvLEGemaD7VZBhulLqglcCbE+OcoJ947Qg6RzU4vOVg2LgLf2p5
cMWTpSvZlbc5kyhbWt7+Z8CUuLh5PKiQat2Q+9Z8VL0C7DeILB6B9tTH0H9KJNFmBtQov+AI+xme
dPJHn71uK1E8SIeJiVHaTafsjXVmUbK2PD+Kfl9v1fLsfiU5MMJrbiPJdzasg2+o35IcFVVghNMX
9vVKC8wsipTMyDnE9CzCCKDsQph2WGsPR3uIgQf+eiHLGPmoN1uBIgOIZh4LljYo5cujf4walOLO
cQz2St6R8Tvbr4AVBZ9vjh18irHHrTpUDNAFteLsT0nrWJbv5IcrHoA8Y1ebWiaPh5/xTV4wL26Z
f7KVmw8tgXHrxCfFd3l/VaSOzfS7I1utCt4SRU8u75DBR+dRadwQjbwVyWYogpV2v5+pHNIiiaII
I3GrwfSEQATzwnqJXwMXJ1tBmIgvRyBUKXrpNxEZKwSzl36GQM8iR+HnKMzYMoApw7XDRUWuDojb
KyOhmBaf7Uzrx5F4VE645v5fpHjaid6Rbb6vzyi+NNr2lnut52ACCVZaH6C+KWSr72ajKIuXCXT5
6pb/GNV7ghFLwv7CytCcjKD5EdH7djKrF7Z49ujcK+w7pjyhW05V8o2GOyDR0wSlFdU3dNhEcIkM
o8C+cJRNHV+pL8mWoFikwmWq0LZV5w6v5dC2C65Z6y/0Ioh9ytU/5Si7L0mu908bxq6WV8c/FYSF
FBTLyIuD3Bduall46YontVwG8IBRVebot4cnQODgfG6mkyxWOMsQkO9uOMLSkbJnO9dbEK0rfe+a
jTDk5I+PXzCb3DJrIFy8qdWThwofj8jscdCoOb22DpV07hTd5GNSF5J2imjmvfE1nRSkX56k8vva
PSKbiSmgGZK+7GGNHpmiEvEDYw0c63yIMml07UfHMCeqwU2a1/dUhOgFXLsKAegr3LHCWDGDwxEZ
w98jE88lMQM6xIM0shmdrgzFMgG+VShSHEVNVp1EUYu6nvJAHVnlJutOQ+IF2zmQXl5hyOMDQn//
wcvX1JUKuypS22i/q29oy3314D7tbfAdBQ417f2wGakidPhFO0CuvN5iopZOEmgaps4FgAvMqIQD
TVCYYjhJGTSDPWA6jFc9iLvcZ0KrkFqVoYyRbt5AZPPh82uirInkx/ORDV9IlnQDIoi5HembZ0uk
/NY3WBL69dri816IRtBR0FhewR5lk0P2u8cDmP/vnJRWROTwP7iazu1WtypCh6UrxLaHNakJjlRa
IwJoVCk5TgxjTXtH7YJfpHZEFDBbYZV9bKwv59Fq3/xH/5unTopw5LDV2LvyeoI9qeIXS0cU4URW
LTufyADcOf/W8kBDte+f3HSb0D1mdgCOmD/LzQnGWLzvwSD6JRIO6q+DZC5hMXdnfnnuSFJtxcud
jfjiqNtN0S/3le13sjDNWLGOljtkoPCcYHL0tpU3mPcKAjBB/8AKPQ6cKlJzuFm2fTwe7z3HM7Fs
Y7mZ0u2q7j/Abb23u2e+njsefXgmYr1l+f/ul57tIFXCRcPuJN6i/lpfe07QINmqYt00Ka1iNgon
xx1QIFKdogHx1+7DcO++Wu3J1RR7WSFxiQe+87nrzAUJsfHwbQdULvmCm9wZDt2UulZRTWNpphWL
0B779HFxxANMa0KJAtH22XU3Ww42jXxkcyHbwEdv1L9FSpbCXdXgRX4YF7obAnMMnqQecIbabhH/
YDKyaQTnccG+SQ9pou7HiC3lDzc40qm9xiZpGA/pGgUK0W8m+ernHlJeOOSX6Q/VI9L3ue4sLnxD
1Vg8i7pjOGvOOYng11rpEwq960w7xHPaENSuCooZmmVsWjtAJZY3fsMR3FV4cSd7jwXIsnkTOn1J
XRlpfiTXDYQ1AbPTJr6OUI7+SdYe0K+0/TMfPqa5nyzngEpi9PAntQTiPeIoHEiF3Ojepa9Rpn2d
5ZH2gUd+nJGwp2UZD3hEU7xqtZaYyutjWz8LwE/m6t4dKFdFPRfb7OeRAkkhRXossdRXyzNCFCVY
jv7MWEaXG9QBuIXAUnwXB5Ht5UmJlH2ueKRR4XnvhzD70BT8pvhGwn+NADGpbA6RUilko29ZKR5Y
oR70HiEJY+GIx+X+wFCXvzdBBJKnEzDS9XVhMRVrE8PFBFJc6wZ4mZhYXtsRfkDN/FwFLARVLsrS
gCid0SwsR0sBKvg8IXwFvgrKIKr9xskihsWQw+uQTZbFE3kTnU1iIdvGzXJ0hMAsCZeusf+lakuB
0jE3GFCaoTTavYsXT4jIVoPB9qOwXtTUjaxxp6UnU1s/RGfQ3oq+zIQKYaTFe4wba0ihrBeKfC5S
SVDbe0LqrZjKVXhXbciLXKPW2ew/t1lfXqOp0FnRki5leGGgNIZl/iY2R9kRHWiZaAAkE9lG9oUY
YZY7whEuo6yJHB9HQiLx9H9I2WhQvLKIDzbutmTVu5K/JNhuGdamRL7mkkxTCw1JWW2hmOUp8LAV
fbtQqmmZZ54sho/kMVrls828ijjftnmGD33VCX47h7Fp8MfBWAmLMhSd0DXkIIaZOiwjK1qppBoS
yJlbXjGGLYcz0VbCwSxsvxWf9+/DO/gvUCZVtR4hUPgdSyFXV/vvIk7frGAZgEz8LYNOIA8eYh8B
XbVNs7RFO4Q4ZaLDTXskbCWqCs7eC6XC9/ED0BYAyMFPpWBH3jrHdabzYDhcO2RVwtOSxwCuC7CJ
TJt1K9cMGg4s7Q3q3mjBkC1vdQY/9dWMf6CyhLFt4qe83SfuDp34+nb5gX1N3YZtEQ4Xy5n89rMp
S5zzW8jGTCKZywl/vvllWhxKJnhPMqPnbyY7qXfddpURjSJKlvnC9qC4cZLR6uy//hCKt1WjELGE
rN9Cr15UevquNDMjDdYBXU+V8oKajvccb18Ggkif6k4sFID/EsXvSe36d4vw0g519I3g6c91tczw
Dn0WRzhwrD97nPzZHl4uvPoY4PrGK6WnTQaCYHwXNi5P2UWGAUbvEiMrcbVtC25ba85oOHQmlXv6
1zSJ/woNhQmJeen/J214NIVpXbKr0x4e2iWVXbgPfXyLksHNp0SD1UMLkpkBSlqb4sqmyDYvMbCu
8TksuuGFOqvstBeTtauPPfLY2yp2otiVTHADt575mk8An6G+nOtQl8nSc/2ugu+BWol3kbX/a+Mx
nNJRkzMmxpffnrqpZryn2v8A5+ndS3Uwjk9xUOW7lbzqZU+EhB3CxcSv/INMhpNJizbHh9jkIxXx
NjGleDEL9cz0IbWttwOwmOCHFuyXr5N0dg27/9PuKv59NQEaiB2rT3sTAJiYh0Bngn0RMRXNChtb
+L9Gl4nEEtqleNdmPSUkvN9KfljHnkWuztBF4pKTxoMG6/pkXRBAF37BorqoTlGgE9g968p3qKTb
2bXuQIpgcuQ0wHbnkC/l6Tzx35VjwiIRRsXcEsga8nsm8JeZ7Bz5FvoPfI2iP8hZrsn722P4+x5H
vkq310U9UTeYvagZ5yxDVxqTgSydvrEft/pbo2ZUowUEZ6wSEh0xv3npFhe8wv3GOE7gb3EbnZTB
pdXAd9wOMwfhcAanL2GJoGvImlZLWcjBIvcn0rlPJjAl868Zg//V2+FURwY0IlGUgRf/bnxD0pJs
BptCSk/yGUrDSKRf1gyqT7aXboEE5XiL7ahFgY8s/3ZrvljVeeggzKtqiGpH6cJ2Ln13oWVkcz9W
6Az8nJTPwA3FfmkhOC9P18yCx4MoRBRu8TsvvI7/e2+Be2M1KHKmfwsJQ6laHIXYLQB2pR0A1KC6
cQwdd2GogDYa23MRhxuZ8rFU3ENkhC0WL5/heFkinNf9lWT/2LWh84wV6TiCv7Y5ZhIB/epXAaYA
QL+cp1yvllzN1SyJKrtNdGkvrR8Q3Mrv86Mw5NkDtcdDc+r5RF5POShocCldQBR6UqpBRe+1cPyP
LyGZeoY5K0dVNj5Rg79GBuh1ySFWQ+oOgZAQzoZ1j3FguVJJXaJ+BlbFxvNyPNFIJNC18W+T1pUr
dF6H3AT9Y43YAxrxGfCKVAvwtkpygg9svSwOHB56Pr3c3ef2NVFBmglvKA6eEPNBTDw4KQccwomn
gKPsHQr0LzXaZ8zgaxvfAXbv1yTq9G1VpgavvKcm/iIr/WVYCUO72XEM+++vnRLPMg0T1xg3pAdn
DCPYOv8sDlKHVT8YrmhgBzngVe4aWoTOAw0JCMIHM/0jP+cbUGaAiDVbqieaGab6QIhVKdrSpnAt
PNAlqrklqS89JevPjZn6WoPIi/tNRyw6ZUa1vJyIS4nf76eEXpii5/oLyi1Idb3Go+IRgabSI4qd
cEH1O7QR1JxbfpYBVrh4tW3pENG6xaIEr5NvIizgs4nqKxZap9LBkYMZbDoSqe1KBmGFcOyju1tO
V2qIiZFdbU6xUvbKFyPGNo8yvsa2HzvHLjmpz2vssvqBswnMOegCeYQVwjxK4lJnR/1lYLlaHs67
w/ilN+vU1mSUFWk/XqhHLRNBMc0wM9TQchvYeAVR+CIOYj6VcpBIdjIO5JkZsJamhGyLHxe7ABOf
93SH0JKS5pdmwfcQP+C8Ej9/XYlw6nHAwD7vN3DS9Ib9lGSeZa476V9kZokNErGOxLEVdbjl2adI
pYBeTRiXxXzlKW5woN86wK7XVh46BRmRy943D/eAkkp7tJDxrJfd7FJODQZ71W4IANCfck50QfCA
VAxwiGaNbu4FrSg4CAkz1a4GzPglLbAihQMwkywuVYJUo1Nk5qw3P+oXvgJPhMdmvz0molbR+AeY
wWIX3Q3pizQPs8KCsXczGvnPCQyb7Ua3KQnX0Bod1VY12YuHancUBIG/F40yWJHF4byvA/HIoJ6d
V9xZzGR/1IMWXuC11JSrTPZ+3pUIp06JkWsIa+oxDVYxQGt6fgoeHlFwKXmQRGxof0z0tFuUwsw9
uJpnNGilTAz1Sk0FoR1a1/xX+yJZA3Vu6CheB3ktN0x67SqFDzTatwKeNZ5FbmPq8Enxo1JTMToC
mSH4BqiKFP3ddo7Es101ii/c/26nIQgSN9d6Y1DNJeBlHO1F/r621TkOGXO3vvAQeP5CKNWcsXcz
1Cx0/GGI34apPK7gxzyMGcBLosS5UW6mRyPbqqM+eZizs77px8tEFYfGLIKHXyPsAFIfjFvB9Tn4
2JscR9EYqKFFxXXPFmClmf0ngIrDUhkQzkBoELkRRdUhoslDyUq2T2ajUHrTu+xFg9hILLAQgaNj
iJ4TOfVz9YFWQ4G0/pqFVdavtvDeh/RENXlzNpejiGJcipsICfWQ6h2up+tbGaIOldTqTYEgcQyx
zndTtFUt8HwfWtq5xWu9h+9q/iHNRz+89kKWFjHud1/rUI8zgj0MK3t4z16BmW5+WxcLR4t9Mc2j
MFHqXsj52Byb/p68BykeoKQZNyvsr6GPCOjNLG2K/8zEn0hah9b/TmSMQqUEt76VKmvERQEWbP4q
GoYkMvN/9Cb0y4pzf5ImRTZFiZvgC7OA+qNTgAY77xcDq9bpVlnoD26+wekYba2jrsGMSn3HYs6q
90V5Fh6u3+sR6l/Cz/mC9rlROLQanQXIRXHYkBGDrxovp0HDfLafZuJvFLxOyXJI4lKdgP5wsR1i
P/3I2MlH68pZPFfCboFvCDDD+7gBbAMm0p+9P5npEOY2GKZ6hMcM0VWb97wurr+xwCsvc15dNOrJ
Ttn1Sp3nnb1+AjU1ptiuyPjNF4TVPK4QJ9m8G9lryUiY0EOAAdYDSYkAXrsJzuL6Q1ZAX/Q6c/3v
rCSYhHLlFwdRMSPifGTbf0ud6jRaZ58IdKXYZreKcdvhMrJoWtmMY2MgEP8ixIjQSSlWVmer4wnK
tUPeTetxb9fOjilW4tRKnNf0CgrttQ7S4P5TYPbfkoa/YZLFPBTP22YKva33oYwnxi4GLaawTmoX
pvKTIx8FBMCOM9lrUv4T3COzzeK1A3VQHjvtJa6dtEhvMONt5hmZ7vv+kr81uTC0C8wyKV+z4hY2
1rXYqI7QM9bGyCJdgsBUrSFOF2Y1AIc3NHUFRDAZ6ofbfMo2ZwM9dA8B7a79cdkHmSsC7CcwXxou
5kkZE9xHjTaypgqcJaSEiXGCBzDsxcitQFiNE8YHuTeXuSLSh4FAXpmFkPQnpZyhPR/qCBwZ2ECs
+7gA8baxrwPAKsjcGb0ZJdtL0MxudBye1G/xUE/oh8breFtJ3D7RmQYkebl8Djdg4OQfMIG1JrRR
l0VuYIj5DilE5QxPQXZcLRcuA6UlSek2Ox9BbDUYbo0J9decjgiP6NfbavR9mOSa7Zw5yg5krO66
6TbhO/xplJpuvlvVZgO8pnNyed++DNcy4LgCvzHSOZQ0GD8Cf9uvHmf5hL12n2exUhjMBU0vesGh
v00rUH3/R7diTl3+mIbvw/PmOb+skXkba5qDSB4MUGEc3IsH3YktZdQCo6H9KL4ptISUMW8aBqHK
1sK8FpgysFlIwnPGQ0hJoFQkiQQlSLhN7P6LgRaozIlU7MCFt/gublGZQ9aneoboXVIDFOq82P2D
Mj7cHJMwloTQtH5wNbW3n0/v2TR7j/TeexgSd/R8t6dHwX3tX9SPzShxgwNQiJLTeSk7x5GjuNHy
xBU2lMsZLVlCJlGKddThcG+68daBXGM67A2LrDPheu68zD6miDaYbv+31sN4Kp2YDvZtI0K8YQ/n
/yYAxK7NqndwTDvnFzn92Aa2Rc1UpLxxeAnmzb29UtQqZQTw4HVtpDRtIuCFF9x2xpcRqaEsn0lP
Y0bS2F25aMlp1JHjfGsW2UAHHc+cxXD6M3SBHlTAF4+0RmBte2Xg+Awo1sUeL/43q8hH92uVVcR+
XKfICBK1UBZAzcLNIhteV9ahxBGtOfthXKjOP1OKMacEfza4+mNP1KYoFWtdzwHuwRVP9W8oP0J9
XtUp+MzRvzAOOcGldeOzMcaJdx0zKDy3aLtzUQ0+9LhsZpse1q24rYFoqit3DeQCIXRa0LJ+fApB
u0dAZq589hGL50VfxHCIL0/yzgGTC05eL30QwGR+OZozD6iKgrn53OFF0pIUXADUNpfePVuqudeg
0Wm+SeFB9dOJzPx29c4jZ/4iZkTDEOsN7JPdUd3xVltPQRkiInHrVZh+czMhbpoYmKDIXsC7RxUK
BZ7xlFp5awuL3W7AP5XVpLREhjRp9ca9XB7n23b1KwQemtKHkaVb9ieFPbK67IYwqZb+PBdUvLod
4+ZRuxsKkZxVeufqJx+Q8i1J5AZlKtX7VI4HYHFOAMVu5jLZAsSwIg3C4q7HqXOTZ3jcyrw0Dw7K
l7VpEfxoSVgsunx4Nh3ClX/B8XFd/aeld794ZNGjeeBjOoEJ3kkrayES3FFX9vmJA09Nqa0Rj3Ow
Qr1d3q+OBCX8VVi7Lg+BIT5I4g==
`protect end_protected
