-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fiVR4xrczJzCiggAoSZ6hop6kBl9aI1cvZx7vxZBYnYXLI5CEsG4xegxE23lQbhFWQV/vdTwt3K2
3VuubXeLcM12nAzRxyWeWpWSx3DHBW+XfkRdXY6iqaTxpiIFTvK4awALqO5xDpzOcU0ppzEdDeZR
bdrnrbaSuMsd3E4l00ygthiRrXuyJKzV6CosfslPcZBNmS+sbhwff8wRGP001VPtmp1ivQwUvdAR
9z6+gcl0y0ykfae2r+jMgkP7bmShEVYaodjJyJMDStQSfqG0bk+q5/Mf/0F3+UD1B0LnUC/8fwHn
hrdMmgZo4BgygY1DDZj5kcyITel6LgsptxPzGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5104)
`protect data_block
3fbGEvr8I7wwOFiVD8grof8MWGE/6hyi++nGsZOQk5il4Ygp9OZ6jT2TRQfN1zmD7GYidhkMbLuj
/ASVAC9L5LvSHG8QC/AxTCn71wJVo6Oxdutf0Zrfpvbb8RN15CDNSXRyLeg79wCxYPB0daIXV7/I
wnrpq3VCYNYXqr+eMEw26GdEgxf0Cbb5EuuSB7cZWvQeHWj3UvR+fV3MWvWZoQZz+xQoe2cKjFmC
o1T+rHOXPrkBiGD5vX3pkfTD5XqQMLuwNbkGFYuZMxWuU4ycmzcYMvuIYIqvjJ9FoO64u0y15d/o
BgF9JIZaij7i+DkqcAq6SZCFlRjadHTViRRWaE/IPcth+acsaMsVRD4RDZCQAFNrgiKr1RVLwIMr
5XkO1l6OeV+/wZCH/v5xL6oBfAiDJddM9ngliO48qGjgsfrHLX4xLz1AJRdRC7xGnfsmd97Kp/sS
WlzWraenCznjFfYQ1jFI/M90HeJSsuCQSfPjp9gwr5+khHnVh07cOnrnWULvJR0S1BPMm2DWz06r
XJM8jFhnve/ddxOC9E1eAgMLmShWu1HBdcKiAWgI1NhS2BDopjMOQEJ4+TNdGcE0VVBuPePug31Q
L20YnU95Pk7uH+wKG419/XnLq68kjn/0i72stdgSkpGJscR7RurqYFYy0faeSJMNcz0Yqz9Epyef
H2u/U0Sg95ep5bD3rX0YOHu91Y4GxO2EWjuAgMC4zIBPD3kEfC8GIvkjggntYOpmZiAS5JC4ifiy
tanp1cEEvInQ+7ViGIessagLiGgdh8n9YXVlGNaWJghJRcxVZvZMv9yHFci6LIFdMoUJfeuqTV7K
sTBBT8X2c0chF1axZ18PDAC+WrMef+jHkvl6ceteadooHsIv5CdYfYWjPbBJcJR8qfYqiqEaZODs
p1Kzbc1nuMp5B6aqt3pzKa33+Kuw5P0jLsmITdAI7XDVoGgm9bjeqPFFGQZL58MoUicUNLZ1hhQp
8mbGLMWAV7rhXS+jHoKSS7vIe/+vENuo9AQL42bvGn0Ep3HucPFmh/K2fFU1DS075LKvxd0Mgerg
OOzZ8oS9c7m+5ZvQM7BDyWJyuGglzAHCCJpYay+6RlqzlZujaJQ2lTQ+PNCIcbikrUomY9dkE2NE
lfh9Wzg+MI7RfwUs2heIqLCxLWBVuaEjNSMr9rWn6BHvuclVGD7HgT4/ZVXfBw3ZwHihsRPcaBo9
iahvd91zDf3t28lZNTQiOMqKe+6lZOEsocS6b1+8HiwZPygULdd8dvDwCTPAZ23Sa9B3ZGCPOGwa
N1BmfspP6LLPBgx4OO6qoGv5ocbq0asjYYIodLUveut5Mn08VyEmY1SiFZ2GPJeDCdDu22+Rf4Bl
+Okm71NOf55j+MNu6E1qKYqV1wXI4HazCBIpIvXqiurW7R/VetoO+aX4K4Sc6NiLFT28ad8SU2e9
PmxmVKOmJH2vBkvookxuOMA7d61toKLVLjsZf1urvTlv7e4qzYGSu2ivAGi362R2QZm9ur1ZV9F/
BO+up+5BzI9rj/R/kbB0CWja8WwWRXylc60JU7tSuydhe88nODpW35lVwYxXmzuKBDpkj8nXVKsl
EcGyXHtojVb/rCsTJOtHP2Ir6s1vTlTb4NacW6mM+K2LAsTRvxjNKL+XQon+SbTGjiqd65W/fPws
+2VttOM9TxrfGqGU8JhE7j2E+muzA6RkCpexBgkVLgICJoxaIbOB61T/FlhmzrsucCIFTnUbbjHX
hbeu1y0iBT3GiZ6HljB6ZsBCQHxTLbzzRfHZB56HRqroC9G1UzmeOv9l22LwWmDP1suUnUY9Ry1Q
9Bh1KNudSpu5UXShp+kPddxQAQgwE7fQGxcum5PD1Cz2SVnso0G6T3q8t+4lPQ/L7WtL3FmmJvNq
B7gbgEbyMmVcc3cNLTQ2FHtJ0TP5S0SnY7XS+5ptCEhOldF3DoHYzWOcXL+yqUfUY25dQLFN3fAK
lBdKBJtKkpVjUK0CteyTIGfcisVscor1QpRwHKzbjKoozgKkjwr5aRWDrIYrutVKRUH52oTDtwjw
JqXUsZeFPMoiMHpD+ZKodR6jIaHLmuYkPSqM0orNFdUFo5vDk+JENhlhCeri109bOxVvwE+HY7b2
mah9cPusRUJMr+m/OvkeyVEix8Am3Z1ayJ+bnYd3iwzlqObx+DT4SIuF8eRXXS1UcnutkK7zUlIY
DJHuJrHdwKU80wz1O65WWlcHkualHpRd+qMogXZQmteV89OjuVBEVnyLmPeT2xU/8kiXf+FOVBOj
VEYmLsV1z9PQBKFWpC7Exr7YNY7gBnzdThlctT7TTxWiMCtR5VfYW9nd8BeECkZtT//2iaYgVwXa
80rxB+K3GlsYzNX3ZCb8yMsgUDyj8yEBjv0R3rwy0X0rV/mEy0F++p6pU+yYIN3sqv76NDJH1unD
6sqa33GGSxwgiF4qMBWttGX65CZzVhRn58yciF2FlU/wqxlZrUf/iDe35nbspS0ekQLirXoSlckR
6ir8DewpgnqCuEhNKSd7k1xgw94kIMpGyea7KQXCA6E6EPltjGXpXFrKqdu6WpE/qDUsaEFGEhSy
CqgQbjBa2iIt79oSkq25x29XuHYn9T0fVLWQBaq8gD9qlx3r1MLEKXbgiy4PqgnOSY0BtMJsjxnp
1k/4IELZU+FBjMe/q0NO36lVdbG2ZxJd39JUQGacx5FjytplwmEJtZTfTrwlNcNgccMX1tYzLcaF
XvRYx8BVfadFjj/57ursjJ30lgaSol+4ifF3Cd/FJsi0sDfLwlO9xnChvEb/W/0hw1RsIvic1TqM
16yxP0a6sHfzE4lJT57CIake8cmB5hlQnCyIrLvw2DnrC2mHu3WMRdso3JkeB6tD0RbtUka7B23e
O7faFmgRNdzXoVXpYH0dZlujDIhV/zwnbTLZchphxkmNWYU4bQMxRv2lkIwPqfcPqixvIP77NwOA
oNr6Y5Dq9HzAwncTrtKtgaznjvRbKQKmmWWbXujzTQhX80w32FqOYAlYYlNUfkte+BTIkGxH4OGG
MSAtKEqgkCkOf2q32Q7ZkFiTCjoaLB6lvNjvwk9t1qp/rOLYomOMkE2M4Ijsz+X/PW3SdyrJOHE4
hoiKOWQmn2I7doMIRWA/GB9mmfiuRv7jXHH0kRdF4Gg9TUkWu6LHPWFAlqunQ5f2iX9H7sbFvUkh
JP68rNbieKTnnpeVuUcu3PTvNzeD2OwVsU+AJ2BY+U8WcopYpe4KwUFEDSP6HoNiIPl50noxkcH7
dTu5ysLrYqylTw0nGbupUj0r/Lmx6kGbb6+U7mqwWkjG7dS7azCk9DvX4RnQTGWjv1lNjq7efgoC
5iTtbrC7oEZLbHPSdn2Qj1iNvzjdzkarBFlE67Z/5r0XBNPahSgw5Wgvh/2GfaRhWczoiKw8/1Mr
jKLxCihyKg7ApwXj48tuCFPH94ixf7+92RZCKFLHydCS9v4K3XYfUrKv+mCVckCrwzsSnzpbAnAq
IZndmKqCNewGz4Xbjl+muIbY6UC5wOvKj85i+7lII1iW1Nm9kZuZrz3joJH0UzMQl2SuD+ym1sHR
9S6Z6RZ0ql9Si4l1QkOeRdhMyx3QkXkn767aHVBVwZOT+lKeeN+LOoabtBLvqNAC4QSsOMlvjuVr
Yimmvnvn0r9JlywaR2aVlbEsemDJbCi1gsV7wgK5nfKymtyrWysjba6UGaBx21owKJStuQPw+Msk
KV7g5RUbpW+XVRARAL/yB8BHggYR1SznBx0/NyvobWPEpdvYnJYWMbId9DAriN5paNTB/sOt7/R5
q1JZiFOX+ErhLPnY3/G1mP7TbVFyMYebSAaBVX1tHZt4KcXjsZWvU6ok8T2k29aPRX20ScI13uoa
wgRoBBeampkOpWFfDaraLrbGeqCCyZ/dhmMDEGrOCe3auMa99yIStqpwmE6EAA8zGiDRTo3pwCqB
z6wXldzL69Ci9Wsa/UNYM/qZBIrmbL8opc0FDudeCAY3G5YW9alH+vmOF/OsaM1KtzlbEMHVVOF3
hWxsLNlkeElpF8k8ROBonuh8svftg+9jq3pgC6SMvzXrYGecc/zxVnO8IsG2PT8Gig38gP0psLOE
iqiLQgkI/VKxg993dGW6ThaLjvcJ8/6hmJlnah/4pG78yXqmzs3AnS7drt+iKxgP3pGHAii+hejZ
EchKxTs/SYTKrDMwOx5I2dxQFj6M3t9LP/+g3suPS3kH3R0FTAocn6nc6OJFgIEQxe52W18grLY3
Bkvdk9HF2K4G8ha6WnPPKvq1XgJqyyRwkPY/mT6PmmW3XMpSgt/368Zjdkoauz1LZIqPNDdcXaCZ
NzHAuDyOPbxkFfsbOs0qTITNNb5bFHXFMyfPFyBXg2YwyhpoRDUD1L8mCyLLq5luAEEFBWXJQcRQ
IqmK7S8F/2DzW+UMwSW6FiXepwyEJz3VzTL4ryZnsDcstrBEDecbYWqc54ErN+XSovM3iqPsDOsP
+FRu5bwnMsmwcv8VYbGzPeALW8mVl3JAw/L9XlDjCV4NZmTR544fKxmLtuK4RrjZ3HH8wcgG3ws7
m8wbPh7Es2d308Qv8EWK47nst6bu0Hjk4tKOWjXC3/WxWXJr40Kyeib4tKkBsaLCoCM4cIDWPeHd
067NFn7BVeRmho8C6j4iIpzI/B2EW1FBOya4c3InHvsiEA/kdua9r6HKRmEdQydAq8t6nF0FGS+S
xWcgWveoEOx1gBkk1TpoCzLMK0Mh+/dYHfiEk6fxw/wUV6HuocFr1weDv8fNnWSMakA/FXFod19d
5wHF+trGlHFyWQjE59wdPidn3HEf4/HyvHbHxH3R05L+4+dTGap0ndHSM6pCwN26f3jNSsDc6LMD
xKcK0nUQy65adjBREmRs+ai17cS82ibFxkKCOEOESCT4HU25mHoh/jw9ZmJChSeYbnbq1E8Lc2lO
lK0qO5K0Rj648oCvHWSUraMk27Q+NbOof9QlY7BzSbZUtVUWI2MCzWI6MBh0jqCxZZc6JuaI70+r
e2ctWCzIPBNL2aaz/CIOEY4nTViQq+hqTg26jONItPLFu5mmp3buFAF5Uck21MboI8XXkC7HoonQ
/dtDHzGIHDZD3EKAyPlJEWprKCM0dDuJIcR6lA7gVZLCYpJfR1X59LYZ2o98VZHykUVQQO9n6x9/
YbKGRIz4FFN2hN3OTV7cO1TioE+zBD1g026wqpqoiYpVy9Vn5+Iw2r184qx6vkKQ3JiuNBveIPyp
5V1+3qoRG5A/DezfJFIpviqxkNfh42BsDzg0TIxCsbzETHi4MVcjLNYIRdUbGmT3YEwv+0//CBUR
5gZlOqa9KqNOFOXV4YNR0h87Ry+thu6aZXBgEXi5ZxF5gDeyED3uuF9DQUe072GUgaRVoPIIsqKA
jt36VcdxsjZaorThqtEQJyxlkik2D9FTx+N5xFYb8axeuMtY/t5bEL526BATzsnwveZhZbk5lImr
DWLVm9J455r+pFjRCE+fz4dQPQJ6/gBl4XjVhmjqzA7oCWAv9W65aWeT7AshYlez1J77FiNEjKI8
t3LdOpRLNP62PUpXeoGkcnryuzoAFgQbNdb1NX+iYi+lrmryZJoBobF1Lz3Hz8d2KJJGsJ4ocLKq
PGOMsY5KJVffez35h2vhC3ro3gwanenFkJSCi5pNangMFWpymxYdfcFx64YJXdscx1yvBlZrqOjk
6XbZAko5UopwDKefs2QwuomY0UHbEdmR8pRRs0KiKgnoBkRsw9dKanVOfkHsQlklbXmlVjzQHCFy
OOxSLSZsbhWOmrpxblR4MJWsexdlBRPmVxkawLDeR3Kcp4CyGJRNamEWUKVnXkgG9BW2O5fDJMiO
H4pAKT3Vh5WmLnZFbxr4oTnBhoM/zcK4Rxk2V2wu6iVkLdLW108ELCmx2NiRAJFimXYgJGzTFbm7
UaG558Yh32BBaSOOJZ0o3E/+GiPdV5rU6wBFD8HTfAWpH+GFg+6voJvzmfsaVWKmIOAgdweu3WvF
C2iaeLyxt1P90fcnSDeq/vNaXvhsBQ7kMoY7U6O+My6v7Frmx2v4HOuF4ziyveJdoJ7CJxUJOTyf
oF9kdnzqsyI/wmRNAWwVjy6rzb+gsuEFUkY/P9tLniPFBeuV2fbu5yRYCEwLkGS7QjkCn5/OtRaG
I8Ftd0EKqnRhZ//cD2MwLmYUH5BGbfO2Rifo8GEahFOq1ZyRzsXrQrGvKTOUuEIU+p9ODRzhr3UI
eF5BIiTVMyIu2uhcKbTkrKCMj48/fPlGzB65QtVjkwg1y5/19Kot345cR3oxXmNru5mOZMAAI99O
YeI8Y55iZ1tkx4mxBAlswat5Z2Ws8YcJ2gP5zIrz4T7v9oaGoPlKVA7y3tH6getMt9DLIwL2YIry
gw8fYXQbTDeEPlMx8HU1HpCmrfFE5c8pTJI8rO49YJZDsBs/ybGd4QKjjmcRR8BV4aExFpl8dS/e
/tO7ZxipOCOKC/WtEd43Mgz6tMdv/qyivTlboNBiguRsj/8yeT+6XFu4J07MWzYdE6qnj8DjHmzQ
4t2CA1IHHISe9Kviyzg1YPww6hj1OK6W+hUpwfIOrM3Xpfb70u6y3lYbaaQhO2m6CSFdfSSdzz1O
fIRQgHRnMRtsBh2n3kJMqdj0OpRlJkbeclTzbHfqKnfDvM9wAm/jPDTm2fy4cdKOq+jwQ7ZtssRp
N9CnDvumDz31qK6S5TUTlkLUvdMs3UO6L/82mjI6AM7f1+3Fn1Y2eJGCFhiIeli1wFqhqFu6CH4f
XgLnrj+Gz7S5Zv1CdwnMrRbyhA5Dh6rIP897XSSQCg==
`protect end_protected
