-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
bM5V64MX7JLoRA8Vsxplz4MpJzhCU8DbhOjYM4mxD/skxSTlkBo1jNn6OrnaojCo
FygLvYYxX+EXPfdsVkyE4iu+jQSbNVFrs0hX40NLna0/birpgfVlAVOc3AbjCydC
EVMc549J+KSDXIUqIO9K5X39xH/xryWATD0TRTVqP2F79DezPIM36w==
--pragma protect end_key_block
--pragma protect digest_block
Zpv0/y5q8VIu+6A1VneU7ISd0Do=
--pragma protect end_digest_block
--pragma protect data_block
7LZxnZaLRDs0sd+BGdCPu47bxritBEsm7cqgcryVKRQNxtwyLq86PkIWPBendipD
l2eiaEUcpxlxvnY5dVgioEPSA5ztACCLOJ3/kay9ALTwVACYRdpgSr7nJTrxsPrf
cVXz/6Z/q3pjvbTF1yyYXcVH9HxAJHj/LjSVDNKzEPhomL3B6GnRZa8rD78acCKJ
JEAle9slK60Y54sH7nRe9w6WMmB5qoaHqTuIa4oz5whiX5GhTV0sYIrc97PWO4Fn
/GfpIYHjQHD0xI3LKvqKP7YHrJOtknprjbOKE6tFaAAduaMWPoK26RQLB6FncvaA
B8AtPSL4HC/LDzq8s6GF2mGOoN5dEmerpYcydgERFnwAJJOkZr5pKnG3DV9oLfPC
zV8uiUTeqAJ1rcfhHfiZ/ekJ6IxFOdREg7Ft/yh+WQl6xpekhdc6nDJP45BzfqFb
kOPRHuoOQqyWcsdPSkCCBKJM7GfVT1Akz/uQXaUIGvUSr3VfPBC28dGBs+13HaR+
JcckfYDsbQ46RAdtojarwj57LtyOv+8DlIQIs4UhJYBCBMgXjI06IlmMzyFc58F4
jdQvhsibGo3raF6q+jZhV7rH80ypqHVxtjgFQYytKyEyUKb+chChxuoUuC2KgTrh
5Wr2I+XEDAet2F24aVu8TaG72etFiSpZDkb2sTtcebCG2ZKQ+ev1qVaHzFmwkh/x
f0We5gicEeHbxZEtG0V85RTsak/47aR6bXy+jpStNY1LCfEKgy2SHocvutSg5Vyr
JpKejiTTpsZ5MjWoe/0Vo+jsRml3FRpLELMxFdowg/kk0V+XJRiJ6dqE1Hq1fTlu
6x2dDjP8W0AguHOkN8VzEKQhuGY2ifxcv8UiChlmDW5T0IBlNm4qGBzSJNtoP1pr
VtGJy3dNfgzjnCSnjw5M+Ncw/4iVzR/84ztxH/+zOvXSiBOZs6nWdZq4Nr3IjS/x
nRhamsQFjvm1+ntI46LcReNDtWKXRGqHNGavMB0jTz5AyGuquk1fvskFfYny3UuW
SbJ4ysKRVTupOrBO7CVmm94kQ6r4YxN0rxwh4UvJZgqYrt1QFOl26zVMkOFX++rW
PMIUxE21aEheZRR+FQH745w+g4QKtCTdDmGtI6EUL+ziXgr42evD64TNbb+Ao9vI
ZRLuZCCgXQr6rGbS5C++j63yjZOdeh8cZfh3+vGpR8cAkBEGTUyA90sxUVV0J07p
lFfgo4yq/Rvss7hv4IANdii+CZDamZNuiKF9X69PGPJ7XV3Wr2jkpZ9hR3Wz/Ko1
RnqXBuwNAwK/w4ObJFuNLRJFw68EB82MXfZrG659Pguzte9T9eiBxtsaYvJMsu/I
RzhNjb87tncfnF9DabNUjlhElyoVr3MYP/PZmVwvcLHgqEukydHin7/ZArRDGImV
6FPMrVhnTaRJEZVVSr4+1K8/6uZpAmqt+8SQdw10zIOFA880LhiO7OWKrRHMO6Zb
v2rdiDpBS3x3bes7pEbgLz6B/gyYxeSDkQeWL5aMw78Y9TZvgsSMUmW545WIDSHo
RVP7aOUnMEZ8bdVaXvO1lNcCxdQXAvI8nr34c08Iuy0Rf3JQ/flHiJ/Ug4dYQGm4
unSgogWhFfpSoa5xyfzoqeCA099dd3iYrufSpXp2QZqG3wK9y9Q7q/SK+1RXPG1N
L/qBxup4hCXB5PjKL7KxDCb7lVM/cS23rC+LvYdf/VNd/tFEhhVulhofmbiT8Jtq
FEokVOMa1f016OlIUnWqFGysuFkpk2IMDis+HGE3cRbtEJ4AgFXqIFgHkEte6udS
j5NOJTjcTq02JFDJjRJY8eoZFyd52c3WQFyAClFraWOj3YYtY4GB31236d8yreqW
muCxOEp9h5PVa/HvpREZmCGncbkgjCvB5iZ914FGbnmwUuocFRaKr/+S6vpm4YHN
pnj2stqJQketzXbd6yfrf/i6/DTMhdtOgZ94jZYSE5UKxICkWcKEBuN0ESRhySAG
htX8hUL1OEn1qBKQVkRKL4ZaL/yhM4dtQlLz2tKwauE1v9HWx+0BHIB4+Y9Ur4Mh
8cBdRZWhSMa8/0IE4S+Pyf0B5vddpmIxtrIiHrYWqx+l6n5dTXjCD0q6XgVmwetM
+DeNg/a38kTRx9ERz1az/0wEdDnM+lZyOOhtC3EE5Nx3BKTBBeWjDxIGm3VxnFKE
uPxvy5GKkS40PHiSzPCSdBnU2ipKeY1eNA2wGsGVqul43JycIExCdP+xNJiStyme
Z0a2H50AMYcFk5uGu9gswyioY9eBzwZH08s3aI+90BgOQ0YHG24iIs5GGtQhX37c
uOXks5t8D6CWWu09GbQiHheAA42ms6MXQBjX+r+yOSTCf8bf71SE4dF7XV1J5Lsq
OUBJRMfeyoBUfO+Ns7f+vjDQwdYCC8tjj74onyCy62U+1OHidAHZfOWZE3nNwhFH
JUzuX9DBQz7767pC8/8tWanPFhYkB8gCPLT6xZfDd7YhIOVHHAM5fyjSb3/fvmRa
6NCFjKw2I022aoAgb2OybMzCznzW8wfR83ZORdtbPMvyDOtspbWSMBTWhUbrf5ak
eRVUEDHLEw1zGqxde2FLQYdRgyiAGVYs9VzVj/05Kq7UYHpUg0PXoo5F5Ve7LsNO
d4oTRShx8x/p67BD1q1MRijMLQUE/pjnSm3Oe8ufhhATpzIy1G1aVspTcanB4aiC
MunDi1Qmc3wQGvrAXqy75Uklf0QyhRj//k589kEYtvTo7lrBtMnC7tGVBDNRfhbl
CK94PbrrPX931dCfTgNozuVcGArmHrg8F+SnxqzpapABZHcUfy7Ikucb98wVMWfn
0Q9yBZUQM3cDI8PDcLLD/56nzeIeHmJsGtISeZxaEhM6iSZVZvFwo53ocwZ+u/89
flsRuV6jaYGRh2YI8CKY7Xx25qmJf7/BT+C69a8fq+ffutGnEOT60pI9/BbM+7hA
6JzckuCWfIdQR2dpgxeu9qLd1zyqDbVw5S573q0FtOyzWI8dv1ZGLYs9g2d0BwYK
AMn5H2rMcRQMuDkF2mLkbTxvQHmkolWCJ1j65n6EP+r5OiB4cvOkILX0mz/Z/I5y
C+MSB2hPm/KRdYHm+L/NDT/voQ7EQI+3I1CLInfo7dAt+eX1WFuLmLxpRgLlH1pv
GhhcIIrpuMwGpxekFWLj4fPA16yJLM+p06dIdXE2GDFwAq2vfEVBJqc4FZWXY0Im
CSqraZrv4I4FLWeTa3IboopVEz1LZiMF91CFVlzBGyxUpoudxdqFRkoCTKPSWqum
c6k0YpTf90onxSO7e1KETGcI2ugdz3PZyEKUDWHaJV4qVOQ+NgJ9MwxBtBH+6n05
UF5rMTlzq3VVtZn9wM6pDeTm8ahUFhDMbDgeAaAIwH1HsT/erWF1Wi/HRmAJX+df
7Avpvwm301C1IqLFhcn8ACFIWkT1bY1oSvGZp/Qg7tFdNCCpYz0edKrB+WPj0Oi/
4v7TNq1k5k2ZFCpGgkYfXSmRXlEORGfbw5VWASFSRSiV1OxzIINQNTKLNtp5V4Xs
V0ITRM37WABzHWgPDC8LTOtWbgYIaSkV4os8pb2hkTHMWa2CklouluU2BxEtr3OE
Odi/zhFmiUxwWc/mDeMIsOcuY/YBNoEin/CHMPPJNpRe43POPgH+DLASJKsoPwqW
kEF2TFgX2aR4X7kzUKqzkCTA2td8xg9ynOWS5t0VmaDn1zI0UsQZCcBKhCKFOsyj
g0O8uSPlhBMUrTNBRF0HshwOX8t8VmIE3DLhGdEjShYPuxkamdL/4f7eQOikwcoD
iCaZDM954w0LG4cbIQb6lHdqzk3lR3dHB6GeVNkB6kfw1xFolPHi4+FlVglOUWrO
9FMuyQofWbqoZtxDCILvp4i8cX3VUmSLwUMOBV7JILDYFHdvjq7CG5SHjWik+Tgb
We57Cc13jSv6u77qsdlYetJCi1GNcsqUgcYdBxGD77QZUtpry12ow7oYvhXA7om/
WgnD17GOwA+UX2jIfSHaBzQJo6gqSxkRVdzkYQEybQscRXuJk7wSh980fX5tub7X
ppT4/LtcxcmQlihpwbORxaR0jtFU9l3HRe6AAEeGyM8gEJaXd/ypTsVU+QAPNAZ+
5uGCpbra5T8bLAMa14IMqQ0EJ53lGYDzTeS87nq1piTkVVCpo7twWoDsZnZ2gOJJ
EbrQdLCKjrmbUOG/9i0wgEfrbrddDllUJTSLXHeHazaINlQ350Kn2OvXM7XNgI5U
zX5CvJb/vIR1VfEhBRaN/CDnz905VBHVT1gYy32vtR7YFiQjrqoDewCtE12IT/xX
xgZKtauRL+swjmg08DuRtLwsir4nRfAABiS/bSJ1wzsfVmWVnvX7hORtPQl2SfxB
LMztnNc58U+9cm26XaIFe9TmXsLUDre2Rcxe71Am8wwYgVCMkh5au03VdXd0Eqi/
a82Fsdx8HPL82Smfr6oaufJY6XcoeQFYCDSXMRBFz7hPmMa9H6Ixpi99ZLvIwFL5
yBM+WWgqiwY9nExqYjONdXFltNcXPLkwTAeLg6hlGbO7qdEaxeAiRYcE1Tkz2VCi
ZfCPSjceHvYQh5YbvePssPSRt2zR6gyq5eVOWHRE6oaqqU0/EPHdfyVoUvum630v
p6i1QNoEPdBkH5P8463jRxFUMmgsWGexbzBdgTl+mZK24q2RFlYeltBQmGrJt5gS
KutTLu/D/agv5hREc8xCvEOLGpeBlExY0tidwjR16b0+QS/gzBktFsT/RQZ4Thxs
PsZOLNLNzIUURbki8c4chZQrZ1fIMMiWXl1pKWcNbsKJcy5099rwik/iLaSeRSvv
mK+TcTczN75fEQ+L/dKp2G80UmLbdl+tMIrs2ZLSJLq3T7BFjdbkQ4G10UJhnhOI
jexk10Nv/WI8k+nUXP1+ADGeAkUpKYxaWf86BEvXoZwewdnAZknkbeevQBhkFSu6
zLzM6EPV8759N54LRTwbz7zMG+ksTFYUzDKEkWWlBcZgcS0Hf6ActhtHo0anApUq
fBnDWFKPtscRgLwlldpxzyrqP6kwpmlLtsqH972cF6D+OUj8SS0Y26c4JBGu5rJL
kfxU2v1US2eAlbN9WRih81HZcyOVxowDHUZZFGs+i5q7RoIyJMQqDf2Fk/z7lhku
NgxF9qzAygQBIdHacQt975cS8ipwXfg9LGMVCXL67VrVI6Ou9F5ri1YVBbufyLjb
ssHD6Fs5N5MqEDDQz8ovfvs5yD2bLUdFviYhKtmTmhTKEVBuq6Wp2ebZx80Ngtte
thEJk4VPm5jUuFYooHe6CcYFTT9vgeUcaPv+22jKJFXdHB5EgC2qzREIY5zlbXUE
WgvcL7G2hiliZsrW+VQ4QH1QHYPR/BcMk7cSC9hg5lpSHpTeRHHn/7G7gdyZpdZs
Tx6Rlppi/5bqc04MD0vuk1piwceFqHTLXakOA7m4B3cMHH3Kfw5zkCerx9XN1pyH
Q0jkCJGxCfoNzl0s4g7FpC3doqFgr5TTaaDAQRi30v5BWnC2EGGve1VviabWiySj
JxpXv4o25frmlHG3nfyj9qf2dd+133z0ubYGRR89af1Zi+AWwhnHjVxk34hQskgC
Jv0JZ1Bx+GIOwFEj7eJAG3t2wtiE/iWSGC3/+/KJRur/deLfn6+xrrvG7sbAkw5v
vUeTkzR2DNi64ckbVRv3EKLIf5drUWxkb+tK7Br0xl1pQL6xiYbcyQZezac6PXHa
O9j/4GxNq2a+0noAURXXsbKWvm9dvz4mT+zNl+43Rm71IgfV0DFXGdXcJzIg0XwT
kL12uUuEZfdNowzLuXr+BT6/XOWfqVqouy0EPY+J5H9BYOnzMjY97Uzy2StiFqw1
K7pLP1uitJTpP7p6VJK5ux+VGNvJ9ttb7Rh6vjOqXSiQVWbWSvMNlcoD/JjN1nt5
h9FuNh+wc6YoCJwtLMJ/ll9IPjNQhl6ABmWsvFzPNjCZui/TIvT3xF13s9zRh48B
cE+tnkC2aBJPjE6/22NoG+3/m1sduDR2riIrOZfKXIa/4/CTE6Qp5bVm/f3huP2R
JSQQUslhn/8Tg6S4oM7PlacL97vnfpTlkcWw2tZzzhB1AlWZj8vRmKgQ9oXG+hF7
A8pBnX4D5vAMuTFGrvkSd/STQLwZW++RzvXy2JXnMrh6VTBrBnn1MbIP57w30n1K
FoN09r4bikaHwZf0tn1hCGGgG8N85aiwPmkJeyS4luzTzdDGE+fPVl1eDxW6bb9W
rDTSnaDEnP8YI86C7hzJiVM/rDKP9VLUopyOMVUd7IvkopPx6wdnmLzpt1KBpLCT
JPJCpqFZx12k3xLjO+X1ubh7A3ZFHk1yxCfkwn2wFBWjndmzHUDk4J+DN7R6kKr5
dqS5XfKFm5OMI4xgqCXWQ8tGiNemzJTWnrmNmsXSDUknZycjuix4gZkbX2EvuE7s
mUSXJGAN9790svraG0AQCSJe4qLqoQYQbbntITjJNbdXXh1RUcX4gKXaoaWREAeQ
yJqZqpAYL/FFOkjdJ8ZDZ6ExGEiqhT+K1JzsHY2p0kvBfXAbSZBEGmZnTSIgwtZ4
i5ljZSf7460Vil5WyHF2VwW0+uP3aUFIMCdgN+0QOq5zkf0ZRuZkf4D2l9nPtRNq
y4gHF+OpyV1f2aBCiaSzDN3FYMH5uvILdC/Xr5H1yEzceWC/yZgc1z2k53IPCTHC
ySjHwh00nsQOpmO/nDvPBgZE+mRAmmCYTuXhBzvGBlA84CtFwMuBVMYFjnSQabWJ
a2vZOB22qQDT1+DRIK2n+SnaH028bZKkUbZJI2jEwTstwH8MiBA5CU+1iFydJDeZ
4cNz/5eErL36kTc+gul+IE1XQawkBvi+2MEf2uCsGLZL7tYH4VTL+QtLEGj+/Ji4
4Q6HUWBVPHhlkrfGc1ieJyFksKOvD4EHeBxInKncskiYfSEHBjqgnwMbCjGeSYBn
iXMBgQFYppdrxuVjQChFdIjrggZVCRSlLh3HmxHfRaYjoP7VfXpykPRawPWK4Ssy
yiiR3odkyYbhVYSw1o4rh13YOaGoVHl12B2/cBVqZR03ZNHR+S2f63csx5eKbOig
i/NFO1ygsHNzGOGxsZ6wy8xvB8qMXiHSNp6uV78A+3pZk7YE53JymJo8Ts5unxlo
/pkBzsL3q79lVKe1hKC7+jnx5VHQNM4KeRkJS0Qa+GebfFgYbzRnmKUlyU2WATgo
aPvUfxH4YdUltj0B0McA46NySS85Hf8au77nb+g9niAokEDmBLnyTQMGipo2j6uA
oeVodVUJjDvLgUXgTzV9vdHN+Hmk5yh/QKAG0v9GLOBxoWdsIDlzI2LPoSyhA5hH
CoTiIwM2roZeCwvgzNyudDE1lyFf4TvZlcRS8O9Jz9Dit/gQtk8gtT2sC7kZ/GaU
RK9ZgSisMJZ2kDLbOX22QrwxlqUFDI5789jPcIVWDSw8CjYmlUteRYYKYZOHqL/o
YPhDL8GQmzCzhkxbiga56cT92kOvpgSMtVcDDCYJ7/EpAlreF/UxSJ4HdO4qOpxD
0aF6VdeAXjuhK/WknEiFAVFvLtbCqZk1zK5OCscOOWaP94Ddfdw+yBFpxvaMhSL/
M+mdrTAskgg6HZAnMa+9M1JgMhc+fZ14YWO0ffjavhGLTxqJVZ6frJLyARaM7bEL
ZX+g0c1mCsOQK1CTR8Hw4IWR0Y3huo9Z+jKoGrJlXqettNzWsyIpcO2Re8FWkVlt
NYo1vlN3Cf58BOdL78MA6ucCLMg9iK3FpVp9JwPz+T1OlUCBu4HThsExoMMwh6ut
BNyiDcEoKrnHaJdWMmJbo2SPC9+Fc/v8cLo9Vv1lJoUpyA62JLuf6E5Dsg9lbU3L
6Hs3mxaWs3PS7ZY//Sd1Qm2HVB/vMv7gxqYSiIxOK1aCBFXzM4vw+QU2HsvHHimF
lYweG5yjpnbvEKXlQ/w9EhPLfm64AXwzCU4tMcWH2EymE3n51CI/e2/dKZWLlLgT
cUnjG7zumPoL56X+va/UgvwobiOysIPHvrAyydq+DtkoV8+93BR58lH462LztrbL
WtTi2PBNNErcOpE48Erwu7a3cpeC+VUmMqEedRyKzPdTD9PJx2HxJO+s04B3zxTW
5spBLC51WCRIrC6lWX8PX14urk8/uVJy+QIUYepQqXWcHagHveSX1DESiHqETr8I
1TGFRRw5Nir1HWpMERWRsoETUyGggEVmKm+4Abl1OfBr4J/CLsxAWusDIO2DzVvs
4g9XHUH0+BEjr8W6b5eaP9KCdL3pahSUxJheVGpWXdna6iSfCzcFAYMh/N2nAT3F
JDu9SJ7NicDqRbOldSyx1uoZFf18iVWGugfzZk/ulOLV27daJjt6cFUOwySMUmqP
TYXTS/tPWNehBmcVDBU58Pi6UpzJKfTQBPiTGQb1hiVtzKJj0lrN/P1mHfaS02y0
9a2RII4nI9YI34FiiJUHi28CeoWcMc424OQalhjl51/cwVINs5g1mqJpY63XCRXg
m6cQdRYwr+M1CY2jcomj6K7Jt9wQ9VI6tnVxEH69gkqLOShpx+4/Nj5iFS1LrKPU
LY/tx+XDkbUWU/G6X9q1w6XNR/Sd5D8fyrCMOWxP4HDXDOkXlq83XixzCy+NAx1S
XrRGi5Fk8y1OPkt8sIfT/YRTY9N7wa82x1EYq8BzixO/cexlhWxrh8/93fiQVRse
FdeFdM0wgUPEcr1Y4zo1I+vmY5nFZLCvX1iWuB2jt3KLEpCSYDhNIwMMTMaUs7lc
18k3ImortBwAmdarSB+dLrnKXPa4CqB+FR/2h2OuUQqankZBiOgiARQPUy6jluaP
vLbnb1kn/k3Bcdq5hJatWDLinhmAt6pebJUbyDcXC6wzqe2kyFH+bwB98eu5oyTo
1YyXllZgi4SPHhPYO9BfE4l/Ne7S7ZU0tJj6OtGx6fz82+z0QvTNwILQFW2tgK8K
cEbfUzm4b44V8QNVoIhUU0L1/9lV+wJC5+8vMs3Eux9MUTdHdzplMuXd1VAAYzAD
FQQ3HSOituPKgbZGlnoPD+7NsIb4TIGlLw9FVv5aqF2Ge9aRg1fXT95feLf1icJX
3YtqJh8nex3NGzXuKcOb/KdWR+x2FkzT5gedVcRTGyDPwQdpkJ3tU3o4ptT9e/ZE
g5GBZwzx+8oBeUByFd7fGd/u/LmDuYKJ6V9ma0V0QNcOqv4bIviNJRfscw1JxEm3
7qw+z5Cr+GVOTMc+6b6RDewWpihIFKncwdPf6JYligAAb+wKa23eytnQwyj8cpxB
8KNXmLpIlLylbEdEjXKSSSEMbjRgj89xEfBW7Dju9uXQsaPxnDTJtbasGpORJ89x
7yWlZlKDEN4hgBMVkhgfEJqZL8deauQGNe/Y6lPRFfeNiP1HFgdEQzVORZiU0vLA
PRiPtlhn8NYaxM1J16KhSFfz5+5phgBueTlqjXpQ46oIduWi5sG6gDyM+j9e8egH
eV2KHYkGUZClZrrYDJc0pFy7lRaL849mF6fLid5DvL36Z8I0cqtdAlUcZIbQdeaA
c/nVSf2XziT3xhMj+LXYTnN+slMeLWsR//a+/faQwIWKfXtQIUtrqbP1ZiZPA8tt
nOFLJd0+3ZQj8SIbBQTIwUAXXFqYJ0iPRtGTe8fxWcN8oSYkBP0Z9PSXJkbRBFMU
5+z9IxTUQ6vQ1t09yDjCzGJKN2hdjIHm27ZneKVvnJErDo61A+z2NARHeZcoNQmk
SqeU+KkJiRwserMGpFKTCdC29XXEWjXOJVQRn7ryUbQywLB/lJUHvIro/HEoDWZi
Ikq2rsESiho5jBJMEvF7c4sYFw4X9GVcQK6fs4TNPBlB3TuCgRj3iR6wuq8wawgb
YSZLDPJWqYnqrDYYIpmXur2FW29gXktTYt/i1WEVVaV9lwk7qfkqROLJ1x1QrZHL
9aH1m9zy+TeYclTbmGUxwR+Sq9PZtcEGBZqBYPDwi0PBB5C6c5k5WuADe1dwtTJI
eslm7mmKgXxGPJm4yO6z0lJwGSoivOgWJti+L6Lq/HoGWyUbnN2XTRTSmPLtjiBg
804rVHVOgzTstDcWKnwTX1+LP7s3CcYVVW5gYXlVF8Xi20lwWXViRsPPAtqV+Ug/
WVtEwZVygDGuGYTxcIMc5CtkPh1SNEEV/pXWOmUkFlzSVtcCl6x7yxPLkloUKY8y

--pragma protect end_data_block
--pragma protect digest_block
hOMFT01sjudCjhWexazCmJC1AGE=
--pragma protect end_digest_block
--pragma protect end_protected
