-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
inKKrqjEydzFYJ7lKRMq3g4/J3noDiQ7ZMOfg2QFwhCBcQ2mD31k3QWp+tRpthuMihZUAxcSu84S
YDENQCsOIgMkqUpCv1MjGe5KxEZfbh+bJgEMzHo07DOv+UV4NJdD9XU7IcGSvR/s02D5qm1h/+u+
4V9HMZTbt1qhKBylm1j+WkwiXacJmbDJoD/dkOkWM31j4/xSLV9WgI4KddiwE2gp8C5STZLPhxQn
rNziBUoQL+X8Jep1tukJBSX+W/nfSRn5Iral1BHavVTdtHofl2odV99yN86T+o94Yq7IIC4eQsh8
jZt53E14x0PBNBCyu8EE5jfMjU7/4cPujRhIBg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10320)
`protect data_block
sLnCW5/kaiFKINZnFW/JRfDwWfoSYckK4wrh1dVPXE3FILvxdN5ReHV7FmL+css+FblJcMd9bMT6
Fd164Vz0C2uZzQrB4SelYdEA28Pml22HLq4kr5QwH8xnnhIhbEFueDEo8PYJxgiaSoctB3HzRbCj
ApUpITiTJHdpQLIJzbySPhVAIyfqdxQR5B3SAIgMmhxut5Tlk/1sJg7sSnXQD71ALE3eWiT3JWDM
1w//W/Cc2T4HU/SZdEGzAL2UkQVsVn5Mx2Qxllo9OtB9qHWNyK9rmoSRd2sH2Cmq/ds0VD7GeaU2
rCdURSbJtyF9u0TZIUjSQHltXWkpRL3MdbnZKug8UF1wyc19O/XigGTn7tqnNjGn0uKaH+N/i+gT
dtrt5qigKvNjISlm4DrhFN/fnXVhsZdqngGQ6Uq4ohNyQoRRQSDHoZ391xZvL99zIA+9BW/4FbKu
oOyBfuv61GGnGqmKXh/p9xa0MlbSbxUUL257DwUYs0uwM1pACL0kBzm1Mk0wJd2Y+aAR9cYzWX3s
1u9qSblj46LpEzX3s8zmcQSer+2porRdh2BMorCI04jG28XOwPFG4KjGEuwyUBEIOqRj6qOlAe1R
6TQ9GYGC4lO62LS0Q3DqWuPvdpfTl3wHQntGjc07G4MSKgYUq+bYPdH90T/jGDwkf58tzFE9pPLy
FEMa/+Qci7Xmpg/5QKU5WG1D5g776+GXnftMf7rufAeCoXB3ffP3IpLGNs0/OwQkf/i4QWZi3YeY
hnopiHsi4qSR72zpAbcL0e8drCoufW/5i16kt9SoHESXOn5dwTgKdKYJV0pDQIoHMRWxzh/81Sai
Fynrf2jn/xf6hl+c0jochlrByX7kq/pqpS1lCaRDrOPqYFRPRt88iN+c98j3nP8aiRN11DvbCI+k
ntbPNr9VLk0lEiPRtcpiJfDkkldib9SvNGUAb8Znvz2GfYsxLPV8J6+Nzp2sse3m44SqcCvN7HcR
D/QyjR7+yqJjz40iFPdK/CEjndLcC5F2z71XK3mf+usPveIEWoZHTy/KF29ptviFH20CXfYAMBCj
xzghEC+m2D36boCnRdnAWmrzcdsckl/kWBmakQ+e9ST1BJTVnTTLDNC/wO7tQw1ayjOZUV6CDCDf
7dTVowGWSoJD5PiIGddm8/kmF+sKAzI7oyt4ywikkCnwXlh1ql+Je4YSnqF4tnQbemAQ/obN+ABh
E6DlI87nFfIwyENcbukgOPzVkQgbFKqyJ8NWbWjho5unS8ozO2Li8G7vcz2grXRHd5feBkqkNaUQ
v1bieduKHWHai8mAe96gNb1VBjPdVIvFg8Yu1Zv2qpz9NjzNVjWgDerq70oIQ5aCG8YqVeJCa0Q5
LlkEAXV/fVGUd0X9D0xL0iuR9CuwmfS0iOTSw3WkKxyQlJ8K7oh69pnMdb4hk+aXut/WQ7fvWHDH
QU0PW9xr/aUNYCB2lallNXoBouaj0jtmK/l+xoLUA395gABR+7XerNgPOsY9W44SMaXzll9Uo3dS
KVeXH6ZOxPsWttM4FOwOc8QiBSaPtC/z5Dv3bTHxoTiYH5LxElhXOFlCcyWahuhMGX+LSu4BB6Tf
GQmtaHfe2+1QzSAE9fsEG6f0ndgeZvyaZL1tlfg3EId2zCexX+2Upb2VZby9gb6qhCCLszHsEHjt
YTQg9eX5FpJ5c62WwzkDW/n7JkeFGDYLwlQno9OdWoUYeds9qy3T+tIzI3VAVnicabaClT8FIU/D
K9LqOw9G4wqP3n9s6Z1pgyq61fmt8RI82mYljSGv/Ksg2bvGCdrNZL8hZjsn5twWoZqggRdQKxXt
JG6JYqoNMVGnHHmPrlyVGIl5YufyUAp/XaLi0jibMtlCJykdsXyhJT/gP9qPM0wadJQJXV05PWEA
1X07hpGzsVypD9+OpxwC+vgkxXwz+VPdmFf2ZhPOS+YaAnrCmku1HvBezw4dGQZOeCqMY8ArTfwf
f0XIWto1x/+RO7QZAa+zLWK40YTahdnCg+vSdW3XrhEqcPJVi7RPKK+739dlDZj5iMnMjx+IUS9d
eDmhyOYAYI9IrlF/Pt8Jf7IaBQVfTIN8mgSqqFo6h1e96GpiP5Y+N4yAEHXjDj4/YlggBV5f/8Hk
5wCPJoWK5lnf7K4+3PAf50iLmlpRkMN+bDq3NFe6X5ST7EyO/cDcn1V39g3mhchpUCFT7zrLpjPU
gC9rtM8Qn7oFEXgykp4YFeC5eCOUJIgwrKnfBVte6+rIx5OQCVi6VpBqkKK2cejYfrExdsmeIm3a
L502MUHrKXPZFid/8Xmieav9WITOLBdqhrIjT5fqnjUk8uMQtS32LPpaW0GjMOKTiitPaCj4NfzS
c5YkI+nisXNgMvm6ewA1PKAnYWBaMYWr4wzkamQ4Z0lC/aYsNtD39ibmgY/XwJPki1pQpt13Vfv+
CMv6oCZXn8R9z/co6yldHWmJG4cJO8PvFMDSxZ1veMerJy5EKd6UVoVrr3qTTKt2D97XDshUAaHE
2J0mhqUcPY8PAzoVlMCKT+K/p9TUBpw8+LKZfCpA6KZ2nYC2wmfx9OaU8kJM5Ck46UtbL8En6e+g
EXarvLMF4siIZLLcPOreGjuBcNOWgUPG46HG1x/KGDTqFeO7b/km+0WCF9WvrmVjaVZQosyihYyx
Qq86UdM9AnnA3T9foz5HhQUHzxGVQWaM7HAVhdHui1l1D8E3Z/JG/ewT8q6eFlfuyJJZoOB3zNX3
s6gEXTmLq/Gp5/rYycyhmsUuMHolnmpXUN+Xm9Hih3qwakQDZK0FmA9HXk4fB1a5DX7b83osGpBu
pyY9C2AQRNYZIaqa5cOifMx6GNE+TQIGz4F07RhzVljOaatkH9+nC53/iC2BGqTRIdK1rF8O5YqD
lUG9n9u/X2idowZFpWoCdXsxbBmBgANfgxz+nYnE12UyrwlReTXefhacSTz3dpAOqzUmiUjV37fb
XjTWMI3iwJmNf2qH9RSutkIRZJlmmnbNJ+or3IplAvFqykTSU8g8oCVAap70fDLwmywOucF2+0ue
9A8Em9XJmLMj4Ul+grfHS/hOC6bHEfu3unGhaY/wwMN7+a36szPsdZGieLbP+J7Lz7venPL9zJM2
LcNhkXSQELOXD0jO3vLdScH7zEL0FKEGcoRNMXenvb/vu0PNZiL7CshkluSMZXYqCaIXHNN2J7Uf
IXzt7XOVFWfrk2v4+Pl+ORex/NjGOyLP3nOEvfQ4sKLtyJ45AeKfI+FsXEKPGJLhpHDnPoZb3Rlj
henZdyVsTkZVnnA03XJcmTQQ5oCbt6neo/m7A8Qo/wR2A8mLbegLmoBZZwOHNG1Vd9oEe+GTC242
9iwD/m958Bs51Zw9YtoCcSUW90EpjeRERWKF9jtNCfIwStHu0Y0oPPdu9ZA/+e/3QyBPAZliyAD3
nXySu0Z7aXfQ7U4RdUf47DjNbEHJ0w0wz4e+TwSvLCjJiTFjE2r4pxZSI1VZlxcNz9IWYgqodPYb
AYJHJjyFPHUOrRMj7meqFfp3NqFoy8yznXMPUMKs+zlY89brmhPUiaPvb0G3hlKfgnKZ3N7+tjbb
4FD/9EzzO7iRgX11KI2fZirsHP6rixLx5Q2zI44fUxWYdlIqwO5vOFoHCIhBLIfPSzJ3ke+WBEum
aVaTUd0qwewO/9tuGpp+LBPfOHTioSm0a9rTSLSb73xTHDjaHArizQuJRxK1jabIzgrK+v5HUvZ7
vH+5BFzOq/vtzK9mSicYatUKMYl9JpkyQED0hsWr4joMWh9Iu9eNKrhvOAgGiY5mioLSjqQNqRhJ
Q8deQ3CWwIhSvN4XBrdWANji4VmxSLICUN/+IB5U7I4nFy3SVWeS5OpYUrr+1zEVjzie79iiRWUB
OFidU5Upto8R62MtU7EJ5d0Gj58/QObCQTGecBCm0Rc2Y5JplD/FwH6S1jnGH0L5tRPlPe4YcWQo
k7UkSNzEXJla9+5X7b4ExZOBnVqeRicdP4MeU+c5BBa+6R5/1qRpYqRUsINLVnCRrkActcrgnLg/
GkfJob82unnURR/Muhi58aI/X9/EiJCfStp8zyk19cEhrF/QCbP9isdtozLT3122UjoY4Ph6kcPs
Db8p/UH9Zwbwt1d8VQWZ2yOBnKr+6rFer5oCB0zX9SBqANNbQq/7QRr2vWOmS57S3MiQpMXZ/e8U
1gdKvLVD9OlzzXo1g1531/u1Jdeymf86019C2LWRVim/jLyuUvx5+SiQWxnp0uHMvxqn9WRxGgIg
3JQxZL89r4RZrgPLOmb5sr4eOUfKkdqAm3+yyEsNdmYacX0Tf08ZFF0D60aELhWb4cdONqOwJuKz
KyvNXhjnNXNb6JuHMJi/UGjv64QfJTyYzJoAKOfLLJr+cQeYWKTjF6r7TsFGnPocXVtiicuYT/QF
aOVDNZOR07v82JGpZSpki4bcbOMIgCTk1hkBAnz7+KV7e6ZmD/95lj120b/l7bnJu3cxlSRPoD3Y
PHlpoZwqjoXl1ses43gK1WRsD7eIySjKOETbjEnZT1m6DucHqx/fHtBUuto5HgCEbYZ5fytCoeyv
/TZHaLgM1qMgsPRXnRxRUrZnF6HTIdMHhbQqe+22nABXc3mXIbZh6vfxatE4sGJayeIGI91pF8Ci
fGJgW3foYtWfWkMZ9E3+/Iu+hPkqXIlSwz1XtUeCsTJb2q58cp2VLRTCCSzLSYlfWG+4gTeLDXM6
BV91W+NMVQhR7ZoibT5eD2Kuu5GtQjrbh7hHHEv095thR2/5i1sndTyB9CJSxDAZ9Yst2boKSqpv
X+YFX7x22+A+LxUIEUNa2+nPQfKNphJSJuzucwpioyugEsTvbmJLP+qBO3a6qnyxjnFwDYR2JCpi
VnY7OBQW/16xVh04/jb9Z0vfVQSwHFLuvCvu9vG1VvqnH9goqD1Tlu0RwikQpas5eusuvQ3Obtl2
4Xhm+DNmyWNvQCJH+ZBnyMZVAftt+1SC+VdZMtph8S+jbvjcD+DQ3ZTL3fW+jL7NVDO04muwycJ4
HAzZicrQN07r68IBieaWc4Wzf9arXajfO3+PPRtPJGUwe5igWFc+p2yUXs+eOa4RUrUkn7MkoD15
SufTUDuq53UOWln7KxzQfgAlYRv41cyKeSxj5CoMS/hn2wXROmMyTEiCJ9lPaXCddZ7A05MPeZHa
QgbQvLzj377aAK7gZTYx1bnN5l4oHvEUstwwvTDRZb2nPsKse7sDm3YyR7oQHvJiNlSFRN7+YfFI
Wbi1oCLeGDkQ7Abksbbez6kD913qOASJGHD4nVTJtbvMVxZAbKi88Mnx9wNQiEwh7qVvMvrfiO+y
ffwQrGKI16OXtKdzmb3gCGmQGqvzp34enRPCGMwGq1To1akFAq+Fbbd1fmt9QO+Jlqvgap8LGWlr
DGC3Ka9xW3uHgiGklfgCwmuV0Dfdu7dJsXpQC6RsXuKFdkwHDra3LpWQiTzVNl096Nauz4aPbMCS
xYAnK+xLOIle/aM8cVQi+aF+2Jvg6S569jS10m2O8RSzmEnhsNOzsY55eUdd23XDfUb//9h3TLew
/24jJUHBKnAVWrE9WZpcOO4wXNfOnmvgYzJkAPwPury/SczQql65ZooOCBzETFKlj/eKtqnIINGL
vEMq35RciipAtgwOBEPz0vYUJfxfqbMYCbzQzutihKypYAsqKXyUBJze73tpXfsjegs8Tri0+akK
24pXrk6d1AJD+fV3MvGbOChl2wfqTGqzqGcyGu7EEC/I7l/QoBPMjFXEOTYayxq/e/M6nkfitdN7
cSKrNBxcTrUsrDQBk+QUtZrSiTSN+Cb+zly2XbmbYow24KP8fn+4gUV53IHoanN2z1SV0BkNJ6oY
UpGLBkZ1zQRIOlssSo0a63feh0+CDlqNF18zX9qL64nhuU3wmljtSPdcL5ZGXSxT4oBPAlPQSYym
gVXFely7YRRQiUe7EHYVgF5aMXMnbFGIp8g9vTSNbwKsFZADf12ezmbm6bJ9xa54/V/9OUe2p6wx
4CKnrY3vrJR8Py+FY6AT5B6/7gnotez1RmjrVHOgU6ktBnStmvqo59FpBxNbwJE8Cu1kTDhfiyGz
gEnI8vF5bDQ8ZNNFja89g3RfSv6XSoET7Kwe93f6LFjOmHg+CHbj6s/3oBa0rJ8NH/JrLmHLn5cl
AcKd8jKVmWgHyLAC/xR73rTYn4Acatpztd8ZwZl1pjRAN44OsZETX4TzumXKticOI/pQk0fM2hCC
MESay1ebmX4psCxDBPQ/8k/JkFrjNfiuk072HeOJFCFdbXEKVERm6Si3nIdudzUTt3KfoVjjyP3q
WJp8hWg+THvZZ0EjNZDV8cMCwkJbcc9khe04xJaqOaea4w0/YBtaHxAQ9Yf9c5Aq1wDo8yBpJhbI
38ryGljMw8TRLfh2t6/FYLvpTFN+m0V0XvLQM79qnr0SWtK0vpOPM0o7rB2myoMLVSGXzPPWfndc
n3Yg0sMz6Pdu8kqkzm9MuWybBoYsOmlCOblD3hMXAfG/WzrUOzSZU5DrjGBfdYKJXWtDKkC5ft7N
CyXFSMbMLNh8qStZr1TNeEVVzxxGs3+A2cMB9sxTeV2xX0QqIK8/c/TqzSWJbGpYagKZ3Mv5w4O6
fgUn3QGmhLenIuJgRpLkkEQTuWgXy59QuFnXuAmWiHYLmKASYnb83F/SWvg7ZMMWZLIvpNS4BX2n
/Zsko0sQU5eI5DKrtDWpbJkhwyLwm+xcNB3MWgAaWFpBKE92geYyM8p89iB3GsFwYI+oCHLfFFmj
the00O1z5FlCmmvUCdfRpOswwX8yc8Fu+TA8ThDiW3YydBq+axdiCnfWtOHUc3bAnboQHf8zT7r3
cX1+hMYW/26zS3OD5NuTjnnVgrRFDXz8OOJDUXMdv6nGHl0YVgd1WRa3fnhOsmkFt0PiVBPhXx0Q
IxFH7+Y914t06DrUdyd3rr+P1Fuvu/+BPByRt5/h0G9tScdsgkbVtKw/Ol/i9mp8yrw8WISq/sO3
ux/Iinro9ojFllFTSYiAmTA7vbiAltYlAFPBuaw0KEU5YXVAYZlpLALGagzadhwGgA8kg+3+vnqZ
gIacBX9cmojKWfMP4jHlbKq1djm3H4q8TqGTsBodgQwaWK1DNYT75Q1Py8wbMrZW/bo9MwKujgVO
UGS4/77xaqlytCvAQFp3Ouu2bNLGb2mqdypDdLlSdTCXzs4Dlt6mOyI669pbbNu/0riei8Imxodv
eV1ExtrvyetfE4zXAglznhUnDUZbSB+/RSOy1pkrkN/IWyfTpcbzLgmnQSquSEtXzohMl3Hd4X0H
vddVQELAQ+NS1J+rX4MZWS1is/lqD65gwduoSstje4Uw4phOuS+zyn/DXxkvcLOQgN92MKkptvj/
+4OGHrsfF752eE65PtmnSGv8OwzTGK/zYwqCPdGc5RuZiLKkTfT+K3hjKnJ/jumTmF/13MKzm4Zp
yILv0OXniO0xA37eydUHcDpim7wrYOeZ5nrIzP6BwGRU/X39CgxsJE1jUGR4sUz1ygO43v+2Opgx
SXGEn79oWEF48wwlpA7595Fe+jU1je62Jcd+fVADF9B7kK8BgMXwr4922AMjimoPzVqsr7DIXQIm
AC0rtAik4XUTUlS93V2oTUrGEYIaksYQoGQNbvUVjU4bdpJNImzNXPRsYry9CbaQGZDAXOQuzvyB
Mj4XLWWDE6GA7/9eH5UxH1DyVY/N4exP7Xv3mt9vHzoWX5CYDyxaB4fh1Pefi7MPZtaa9ly7FS4b
gBaSbBNgrrzuEMpd72H9l0iPb7q80yKP138GB2+QVxPZVa2n608zqo4ts9TrauSitfFWtJoG4Idu
VI18zl3IpV1vZhvnDnDZwxflx2jpmHfLrlFZe+4duFVD/3GhpW25zktxf4IgyndF/XpzIDCBHo+N
n/fKF3hRweb1Dxigs9gv+cqMzw7mX+iR/NsmNOSo3nd7xuL/r6Mrk/w8C4Gj3e4+yPIAvCCTL7Of
9epy2OsiJlRMCY/Alg+ybmkmdUbH4OkgUKEuiEKTDkquVYM78u+3OWr1HMPmoyomjb0kPhGVfVBH
/0xRfqRwHf5p8yuAGWbfU1NBhoq9DV6CKgITUtAtJHoLJxpPhaJiDQz3MiBQGOvTVab9WEdkpJ9P
75u6bl0Rt6eQkImRyUJbpAY/QPT+uG+xzyTz5IcUIhsADB/RR3I+n5WnPV0zkr9+7KmsYFzyhvEd
XlAS9o9bi8BmMf/TBpBaPNsQ7oslZorpKgumQX3QsTsN6G1lgZGN8YLikC6RAMYd4E4rPp5wadl/
0N+5cWRQgSQssDLbgIDxum91yPaDFNAKo0Fnu0nnXrmhhR7fWcCPwEtq8nqTojRZz/l9mKgFrF6g
NE//hX/TZErjZsMWi9xIoYizybKIjVYM9pvzAalpO6JgtW6FgYTcWdwM9vuSIH8PoP94WrUCrcKk
JWRZ99hFFfIRFXshCN4qndW03FtdULn91WzKhzv6rpzbzHIfQ1zTqxBB2Rxve/Ut8pspRD587RJD
jJ69uWEdrmJATBP76ByjKrEnX/G5QwBFTGOKbD3EOB0NY6RQP03alCeDN1AOh4XlKkLiGKGnV5SL
4/ZajXre8EpYYudldpGH49R1763dUzjPNwZIyYrH61NC3bOluxALfAqvFY9T9s4CQpZH7/uginx4
zBAt5YVVTgB1kGAbG5TtOkmnfgUaMhAtTWmcNebR0YOrpOTpRbDhsU2mvFCF+C5P5ja8dZhXXdyt
BdnjdATmyFMhg1G8epWI+ymcTb2lleY0D3/cuq76qFSkzRFw5RQ2Fx31XBpFBdodJnviJ/FQzHIT
eZxXDG+MT3uxi1Xuyj8TWVyVDDazEdJjwt8w5LNahDv+Odk2EYae39X3cq9f1LJxXClyB1EkOFfI
pjPxixaq/Re4aLKtVfeg5464WXzhZaRoIeHWhSQWjlL4ftUKtga0Wa5x8lgsHuOP40Lq91L6rifc
7Nw91jmm5GNL1iWBgsXrcdaeNGYirRmAZxK0RM4fEKK99dfuRX4639n5lZf+YoehPfSCCL1sMt44
K1n933Bj9iwIEd03EEh6l6pVbUUr9n+ljNPcDez9eO9gY/6qx1jj3x2y8UuXO/bp2QguNJngLyWY
tgFJoq/r+NlIoArZK/fR4pc4YKAlr5Ibz2EV9nYy6MvIqHO6fVk+XmxfXqmKSbwH9Ony3tfZfMSm
uCL6a81F13b/jX61QzHfq/M8KkeeQyaAuXzAqHFjq9xGybEuOxPKvSDpGhYyIIc0NDoTApu+pNH9
ULqVFzkAr8RkqQjt7LQ+uD/jXmCSiatb/UQTVLo7LobzcyxrwvMRypayH2bw1otsby0n6wGA5p8F
HwS6aHQfcj30MLnGoDRi24DtxPFi4/wql5gFR1/W+ti16tLAXrOJlh40NA05phf2aipUyawVaWbQ
nX4jS5rNZOA+Clz/3GxXXza1DZiG+WhtyiLjdoyQdVlLi2pSYgmn136cgUtp9GLbUSe0tEEZsOZh
xZpYG9zmy/cEA4x9a61901tibi5fMQeTVRdc5gA2hrSHNj7Nzj8QHQ/hxTob42Q86qc9PxevYDBe
Pf4T2nq5tJA4hBnVqNgAvkJL9y4O543yUhT6Xvbq5OUClmTdNOYAIdtrNL+3l2e2eGkRHw40UPCg
ucdoNJVa5oRSf8abxrxcXEAcYkWlMweEKnFw5to9+8pfeIioVXSS2ymC1DJBK0wkQSIJshcga9zz
NKSjzTyFOTqFW5NjVcx2tJ7jtrzveuk1JFt2pWzqi9FdHGXRUHZ3+zTGqJHVldFSTB3s8HowZLgW
dckx690On40VwdJ7woXbPFbpudijdSx6+tO3N6kvSolBHFKEEFLvv9NUHJGEaT4r4tlkhuolfGPt
hQ9/eydGkqsGg9rsdldY/waqUHIyhQidLndMpQoIacwcWHyOkaS+qaXCIN4XjcWlT6k9/dY95F8g
TPYrynAtvCppkRpccflQ2Q5g72lRTwmUULarYcYRTcUJPc8rMoqNyGp/4g/ARM9MQEycpuS9T/lI
FUhO5fv5AJiZDHEg5Qud6lEigwSfKg6+Zv1yNg86ees1E/tzCMZrHgesCNOkd4K12+eWNi7AQrT3
kzBNe9LylwnyWdpieXQA8E9i9qyRybHfGQ/WYKWAZEQGVbZtW7CJ43nBx4Hs+XZXxfrHLewgyGBA
01xIiEfoq5rWnNutG+G0lD+cNXtDlAlxcV+F6bkGIQd4H0fyiBYoZYfMLkjypGry+f/NjoqGCujG
3rTdTyPl11JiF30LjrVqL5nENkBe5alcDFal14jOSmfTdSJvHnXQzN05my9YL6YOpe7ma1VOYJIz
IcM8pdmPuSuu7uW0gMnxAjvD+CPbsNUFL1d6G/rAY4GeoKUgrLAW6KsLmLQZ/44+smauLdS2EJdQ
ruspqlcl2Tm/MCKc+itu34XWo4AN2OziLP0esUyIB2r1wC1yt2EsUrZB8vcwWhK71s16dlnXKGgp
Uc4tbRU0b8MExxnwI+I6A8zDXFSIpfYoKYZfkIr0v0Q64hNAr94IhaK1+/O+t996YpneOP7q7UAk
yhylC1Q5JWyFKDoHSJareyjS5ufx3eCwUCII/1h3D1utNNs91ovTOemGzJqhXcDbzEuhuFXX9y3p
l+6ppJSMCXkFvkkRBlixLElUL5qweojvzIdmKRyR0CqP1L/6AD1Z6v60znge1wCimTsG79nSZ7pD
v/xTaivh8A/O5+UVm1Zkc6Z3tHhGXWynTKp17hVOD1k30wEtMsPULJ9nS0BZC9AytbCKdhqiIPFO
phhtr8nHOCdgiU2iNaccv36fgQvZZMhtOdVZGYHS1OBlACTdnx10q7rclH9M9BdbRiFt8wFwHFBA
cVR+sfu9WVIK/DKucBsr6Nsrd/C4pN/ImxwMbkUvzEdw7tZSlPWHREa3Y6sdwFSnczsTfl/7n9XT
JaKnJbFLsOnwTVALBKzKOXK+QyLsMXQkC6piPTH4mvC+7FnL3IBVM01P1IWjFmpSj2qJAyaRuWQ+
I57o9+GfCPPaviA203hPe6Ht7fUbYSPFd0WfhsBD0QQehUlVFXxZKZzjHb6UwGgTMmV//SpwV1Fu
+CJ9rtQ24yGeMbAsu0JbFZlXBSZ1E42coPZwuIdnmybYOFj8ZtvlnHMyy7paYSF37tkwFkQF87Zy
2AZ7flLlP+qTHKQQjjDr5n9B02j6zOQHbBukmfOzTepJxiznh3bR5aaWZyY/No0kxokIfFEP0/Ti
UAkm2fvpqTs+GgKxib9TSp9O6toIGCaxNiJD8q7Ho2bWA+5uvd65auWITabAitAS0vW5mxHvLTsI
/+H+l2aUjM/1jf9y3zrmzveabfiPSETfxPB2PVAn6KoWu8ErVs2LoRmXXz+qGxERNzP20aAhr49O
0891eKSvTKVcKvOqB6JjhmyIIAVSsNpW7/cSALeSZWRJ4BIaKMwMesFS2RJkT/NmRKvCRgdWwTn8
pXxDU7jmsOCc7n/yZaTDnjDacqQz1W/88bNTk1HtRHGUlNb3WapHeHXOexPmKgMe5n3jGA3iBWfp
TxCvE4KEBXZ86yr1y6v8egVCalrNgPqYwhJell1vlpCpaKccYwNRz/rOKOLE1ISIyk1ulaHoqi0f
DJuTPqcPqakM8Y2UdCgMCVUQfTJzXoJbWvA2rHLEwA8rGhV9tizH46BtcxoM57goXPWvYWhOS8ts
F8a8wUaf0COn0fivQoi05EBC8eIZquOY5mdneKh24RcqzVZuqNVaZ22fIiZLG+iYHQkWEZ5qwYOh
TJUzlHz/HrGFX9GNVS40DlEQuMv1Yr2p+lcPw7aFneu9OQHDipkpOwFZrXwtzDxn80FZmFTYvNBD
vUOviCBvGP4AqvMuGeQhnuJrw466SZ2Ge2yUQ779/76jL8qP7StbXwfHI90K7E1xzCKFmc42q3nV
FdmRWXhUDVcGCbUxYQKbeBilzC+3hmrhB8l4QB3VmbQoqpc0D/GdM/7O0isNh3PbWAnoqFr4g113
W1rElPwZaGJKbGT2F3MjdvCS1WOUxA4cuCNacs6X31TmrDj6FLBb5g5lXpWZ+jy5Q0R66y6xQDI/
i3reQgKuMDfWBWhh4NaJQC52x5RHHjylATva8ZnB/Is5MPTtlJsglc8qPCNuGrJR2X0NfB0atYCB
xhP8JWriGTtIKiKWLB7Fyt1O/eG2ANmcWS+/epekmezxZ7f3w5zLMKtpxF37aafbcFyJr3FM5bil
95eDTbo7nlgnkvHrj/5t4fvMVQQhWLH4G/W4Q6Yh8pBjKYvXYvsHMXK92Bqhx1t8JfW0EQcONd5v
J2Fh++KNHUus6bC3sFhM+m9ob1DEGB/glcISMASAiJm95bMR7MbOrTci7UgOoE4xh43NeM27LnXi
wY0bRONu/fvazNbAun2K0ysRqffn5WJYSDS1SiO7PjrTMCyAtvg9S9VD21G6RTUHcBzfkZT6D0i9
0i5bX4FThF+JZ/gZScaM2behBTz0CBvMUtd51Za9crxEwdapZcJ4Kl6zY7g+CyxDzN5wwFOiF3v4
QDXPhZJV9nQD0lPfzpjFTGoUknOF1YuO8yV0EXK+dcH1Y2pJl2Q83jNEkIjspxFZrrjZeQSwuKPA
KmInvRco6ih9TW57kMauRStBL2CG/yg1zhR+u4GwEfXYKdrveKdpA7N3s4GL7CfYmHtcMxEG157Q
lrMfeyPw+izZxvyNE4bMJ0LgHMpJfo2dJ04RlsmLPvF8BHgNBA5k3xotAp4EbdiN+lQCT6hPsGHL
0ootTP/CTQSLRUw6YkbBx4SAl6BUnAdc3lZS39PDrV1evFWni6PN+DL7zM0uEDZUkFkMQpiKY5Ef
6CkOEV1VKzCyatYzGyO5CgIK0AC1IavlcNw+sGYRoRor3LLsB4j8DVoexhScntCP/pls8jqqH5x5
mlX85PpjWqGbF8Vun+YpkhyNf5jtH7CuVmUqURAFFxqhVkttK40T53eIJuIQb5RZLvMDaKqBG3eH
XM9XaeB9bL/Qw6Vx4Zq3f8j+WGgmzShl0uEY5db34tT9QbP+VLbnLy8preJKLTiM39+tnOGW6Kus
We8sTZVYAMGMADQRNM1/JdWdFj36cjzllHy8AAigrUZPkMOAn/8b+lJGAlVHLS7t07V/piUUumQV
vsQMia3RsiJkJQP6KGuafzcfs8K1D9jxeoJRDycxen6FUFWYx2Fo9qV/H34PtFeoBVScifj+3pCi
GXqwauzweQYgvJlTk9lnp4IQwA981aweAcMNkH/5wcMlD/LOHlvRJZLXjWroEXPBOu41cY32tO6l
SBjz1m00OiQNWettjnfePS1xFkVsz2EbZZ12DUDiXElptKWZLnb4igpr/emVASqMUfviVUiX3uv4
CX+44XXyWIXhh9QIIVHuch7WbAhv23Sye/vWjm41+XSZ6SOE+nOhOMpeqz1WUKh6F0tZPG/dgE3l
vtIc3pVspO0O+zH2Cyew0gP+7amQJvMayLzvGgLNI+jOqhVfBRm8KBESRUxm6lfNuAg4VOMsMePG
YhplPjfsDry6g+DUfGKQbhSW9iyyTpCwOlMT3Rq+7JCdLF0RFqU2WfVGxuvT9D/wVQH96rVptfVu
o7WSDXbUQptHlTh2eYxa5jSCP/5g8XqQctPVsQ3sayTWIgnxBqWTlyWLBlEb0WSiwHGHbGTJgipg
pqofRHhzAS2/YSOEzJdY8WWCFF9uUgeR/Nww5J9KhcLacGbaKDTr59tL8LZLkLGl+LbAt19Tu4OD
qtCY
`protect end_protected
