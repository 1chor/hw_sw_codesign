-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
O8s1IoNOjxSYN7aMHx+/HcN7L83bQReETX5c80nOzusk0B2cX2ZrAJGfZD9TMah/
XP71IPLzrxex6VKQCzagZmhxuTP5VvBKV1X9e3jPdexXGQt75uC3GP//TRWK9ItY
eGDTYmEiGZ1Wm9jz/8ZV0CCk96nJnO9diBNPYPdGEiA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 39376)
`protect data_block
YvNq8t9eUgIfugo7izFs6lt1gUePUkfhXXHitr24NzOW7B4ZbG/qInNh7x6qZrEl
5qIL7yyswd/uvmt9zFaBqy832b0wdGu7mSYqFMxvmFlk/6O9jFKwMPHKgEMOFkvH
LOjDFNznYuXPfLYuJ5EzoPuYTIAKe1N6NrKcz7GTWSn082ySTI1XKtzZ0prPSU7V
iY5/5PAjG2QS6PgHLmVkqdPLH4RfulQgDODzZEDwC/VnsGz9aoxWhjxlylpr4Xyu
ggA7dKCRTjvwTzghiRUF0wC6I5is6NN+LmQWQzrqIpi6TICyyMKEJV6v1wjyJRmh
36z3BDyk1+Y7jdwX/rRvbmNelKFonb4FBTFvri9CVdtqt6GDyayI7GL2PqJx4bTj
FhJxf+O4+qYkFPjjfLWS7Frr/insXH3JMbjkWCry7PCQLjMK9BIjUxsKM8iGbFPR
hI3Tk6y1wRC+j1RDMaNRLRQOpAukJIlO81W2ExCcnEOgGvnuPcTv0zVHH1Z+0jKc
xODVwTlRvHo9XsKAKf+BwtsIw/5xKM0/atPZZUK6hUX/4LFL8DvIwAAXciw5cL6t
tNj/r1S5l1nioQklwig7Cz2bL99eYvQb9kocYep/nL6X04r6MS77q8TP7vTe9G61
BbQvtLy1M+i8m8vFkDjHBJ7bkqTfn3Aqxl6C7S8tsn9u28N8pMy0jy766jcXHRJt
7rXpdI2313g8dj2rzrqOm7E9IXKI5Qr161RKrAbvT5jcDgyXoEhsr7iXAD9USAOi
Hc00fiotX881k2wbn7ssHtyx395oFQ9tZT45WfmSa6p3nkD2M6LczYmq0D+z/P1M
xAq0reL818Sj6BpRMb/xYnVtL5pv2EAGq0To+IaKOfW//NCju9pM8FiMSkMRKoEF
6o4OxzwugH17FeGDAWyOXSptznc/lfhAs3W+GG04LWgx/g+E+ha8ZEdQR+WGpJz2
QOGRlYuDKQjOzBGxQQtkKLHG6VRlYn1/t4hDVym1/P7SZFDTH/3yZ1fQRii5YofK
5qnCjyyQU3a6xddnDxvrI+OFovb0ASLdiQllA8t5aJmOUrJGJFmsPcKmQXl1nzb3
rNsD/jPlXVbjSRdH+y9Q9fXlvgyXiyJLloZWlnn4SJhbLc1K1ySGS3JgtE6zdTG6
q1HQYu0VmAzVdBLC2cO62hPLFrJockOM2QLlmtBjVHOrd1eQ2c2Q6UXscY0apE32
RWxia7CdS0l/9Qw+XkoJKfoJtx3d50qE1cqiozuT55s/Ov/dPGawBPBkxm2HT8Ap
168cGzxsFS1nwq6jZuINXK8lNKWKl4lMHo11bAJAOYc/iu0ghsxmWulqwGi9NBor
OFh7jwJY4WotXw3OFv9CiaxGcwkW7/J17UAlcDzDZcHeh9U6d6fI6Qz2wLevkh5B
H3fqYvgzZUFWPVYiacZlFbKNWU9sn675kTaBgDL1aDJeAGzcd2IF7DgrUxrmPSLE
2Dxb6pVSExwOxv1eSbDBdZI0SBoU/XvmG+pMP9WlIPz/nPLfIdmUlc4HSfD2zSXz
h4rMDynY1Ptm82UJ339OG2y96Mpj5w9afZH9ZE5+uiRrvv/01nM0FbI7Jns4zrul
YfKzQe6H7Vbu3cke70gSwwAr09ieTS2JsN7tIjlxrm5c6Zj6PmktXD5Z0vr9Gowr
PNHCmbwItjAGIXp2NP7eUFV+vmcKLmSOqU42eJtpZSrU7i8UWjO43jtBoNmPslPM
3q6rq+uOw5BjLbANd9wDfO6VLKwpJJ0ElyEq4mwDJG7VZE6XNk133t/b6mJne27r
xnYwadlJIabvEYcprRRJ6VpqDer1ShhnY3MZHrQTWbpaGpBSp8wmBLDThIIQXxdO
xIFf9daeAThN1fRctBHjS+BmX5FV2mcO5401PwubbNGvNQy5jJQH08b8AWjC4nQ7
qcdbpZAUU8jMF33H4n/V43z7zbVcFOply8IKDHx5iJXzFWK69KYCwHx6Dced2aN3
ztAMzL3oikS24fPZIA2P8GPFGT3ytR/eSdAzobqvFXSsadKyBdWzF+/KY4zlDFgy
GQzDiOcQj3pVbHKXCANSw1+a8Hx4N6WpoW966biuTOD8zsxxQvJLfV5p4q/7TUNk
FGtwTWVi8UGpsi62C0p1Eebbtojpq9MF6tsnEVP2v1iabUgHAA0vKWkVwUxtmcas
CAu/lkj5jspL2/+g31qqPYJNDnV9xMRdCQfLJkojIbPNGU6wOoxsl4ZY4XUcLFFo
tB6pVEPMsbEVIkzXU9dGwYanGcpG0K+iXtE9ECLErRAhgXiC/ChaSPyrtnzCU8jA
wtLcr58HvEO5hOR716/v/sdqY4ax9PqEpwpazxjLtYMhVNycWXoP7E2YFB8Qhfr8
4vO/mI+2prN+VpF03jwlxK6yOB01zo74eogMxcN+XTU5Q+nPuYRWSMGjtblpvjXA
oQ+Wif+XS+Vh/hold0INK9kDsD/5Etk39dC+7XLz1Kx2ljdvCIJSRTUozLGeI3OL
heJEyrJ6AzagpZJl8W/aZNq/ro89KZHH0VoPiehximnY3ZO8ftIJGEF6Xe3Ifwd3
sOmSVOqLDjZAJULuzOfelSZkD4mVxqkyh0RW4wqc4Ck1oxQgajpGDqD9Ec9fcn/F
DXx5g4FOG5AgOag/NCyF/gGHVo/iS6uzQRouaQsH0+8QOCGiUcsA+hMKcAl6o8x1
F1aUDjH28zMLneHbXIACjV+QLVgUXF3iEcYm9MseRBjKqnS9jzx7lbTXwuf6cyEW
70EBkOxavWyrIjboZccExp8448UrnnQ+PZpkhEc5QjxX+zCLBJHVdr3JfrB1+JKl
eF4LdycLK0cu5MDkHNc7gDPpStdZSTZiv+w8BEXJridVoVo5WBxHU0kHdXBb4kLQ
egsB0kQQcSD8+vP+ArMGFsmhAa0PDtfKX+Rhnq9PT1kFnBJf4++JzqI2DVquc6zl
xkE70JkuTEJ9NSYW3boDFk3ybIsRJKeFPa3cMO9+yfffYtX8O+HtMErKdnaDuetK
4A8B6gwFc3rsFjqHKnJW6URNj7HkJqOh/xEzOvVvA8gFZe5BBn0TiHuamKN22yP9
EWU0D+Tm3z5yyl97ZFKabrzSu2ACAR4pCSMMVMnsmCzYwByPGyJeaGfVTpfP3ISX
kdRFUQ4HiHeO6tfDBtHeqjcLp36Wxb4MdV9DO2UJtd2xxLb6FeREegP1UULAFHj5
2UyuitiNDZw14I6I5dswTNBS6x6F1FpXRs8PwC6kIjdSEQpZ+MtvEeCPGbLnE4jh
MOJsteg/7B3xFpfk5w3MXWUIfFMvBer6mioOUyzsmkNGbAJ1Jqa/ggccB2FVduWZ
D5FupZJGSqV5k8K/Ns9JF/VjpZQfW2HXIVyPgKjmZK26Urvddmc00PFzgBJfkqzk
x5LLy3nLA/I2/y/rnQnOasaFtTz32SiJ81CA9IhrY5VKMrOPpHFoZULOBo7QST6o
psNFn82ftnHLPbkQ9ja0coj0+/wgyZefirAjoPSDtOnLPMyquRE+Pp5MX4Tx3LtU
rpjlyiuMFUrw20PNePiMaK2p1ID08f/DUkyf7hNTEFhIFMsbgTf5meDO7jxeyGYb
okGETXNHOyDFYLHSdu8364rpatTXNKEQK8Q7JnKorABtAqTejJbVqW0leQ/n5kQJ
Owuia9NoBf9eMg5OzXKD6Htbk71NAfavlH+JLl9f0bo67nU+Oc6+ZxTY1ax+hAcA
ysG2Cng7Zss6y92d3utiloGOddgbaX69lfC8q03/lM2S7Hvi6n5MqZFCpA+UmdqZ
zAhxi1mm1qlTEEmkt7IPjX8h5Da//e+iBkraK8jYm/DEmO1Fb7IJbc/fXB6DXSuS
A8VI+RCEukgV0h0aHIk33unNi1zr/9Euziw7WQIQBnaaZGbC9drb3sYxm2XqpoF1
TVfiOatO5Gz+2aKCPPPqPRl09JU/Jqc0gQQ+FXzXK46YrkJYiI5epMaipSPD54u2
rNGMUNtvFO8XaPzD4S6oY2fhuutc/m6WmKhgQaLhyTgJUNjsaWgqhPKnGbz7d3jA
W7KVmOols1LRBd3SjG1YLjpg/dJKTjFrzi3qc205gaMw6nVs74pULHpMMYRu0BXp
tG0E0nAxrcVdvFvZ4PdnLv1cAy7EYUBLjdpatnPzivAWQuvbpidmjgwxxzZhg/A4
8M6QYkhB2IXo3XMfGYnW6uC4rLzOAODfgNc3pqofvRviOJgpH6GiLhfdAmq50kO2
roE1GRbGkDUCmL7HPwiwiP+9XAAxM9kHuz/swvY5XQvGg6b3NrnvxlWapG2ZKLXx
XE7tfm15l8Obz9phh6OT4RB+ruFH2yYSiVU/o52k6QyJKO5FQzH/RTY42Qt6uf0w
wR/niq99QUvbJAq1Yssvo7ufBvkubW+aa2lYDoD1npObyiKenh0p3t3bBao9bY53
URkx3PdtsWhZyTspkkZMIFJmpxtda1Ij0KaxhyzRBhbqfTn11FWn6IojvvIaAwRb
YQqKOb6qhtjDjBiYRDZ/ba4Gb/uF8fX+wwM8gulTDPsvHyZVPQBMQ+sBkY4Ka4M9
epyUZC8ufMWwAmT+XdLx2OQtOdSBv/xc5ZdFPTjNWbbpxiSkS/jDLCcnwZsNMVri
65c2ym8jYskqHs8m3CE0r7kL1Cha5cFhty1pQSyYvXKwMIy9jRKQLrnaU4Uh2K1g
YjUI7HVQRu2RJ7nQp3HqA6w6lrqHvcpQAPnP474YY/Z273tufSzjpn+FxZPzQi6C
3rntdixf3IlZGtoNAX/d0/Naz90meVQ65aC0/FL0EK5QEIdTeO6zY4UUUknTjWGr
vcfSkGQ4b34Uxo9k4sDdhdzoPCUI1nA9ywkYrKjiDpgfxFhR/O0OBvipBhxG5Ggf
1YY1ToMPWkV/kjqOiiu6cHmNfXkbyHNJwDEi8jlL7msMhSkJ1txV6Mo4obGpiygZ
sL5mLkdaE8B1X6CP9ySdJvoQPUnNJAP0uf9A7cltVhsk2B8D2Le9ZyQQtpL6vQm9
jqk5x03irdPJH8HWUJXM/ypHdzrr7rVWZgdlv7ZCnn/C0ig4VweFYGJVJfE3XHdY
vSlagiRltbiDArDJSIAkPenZDmb9OErMeqQIzWQnMgPzdsn7T9v1xIjy6Fq2S4zh
Ju9s8Whn9iydl0ojJAHNa03xk7WLBU44QKF8ur9okfs8cyiJ6PUWzJXz6T8hMsMo
3IXVVqMHxN2HtroYvaq93EK+W7FzsbfYUzETSLXgBKsIOIERW8n7RfmAOv+WGDkz
X/m14NnLIdMhxB2aLaa0RgxCR17dkRuBSjX7MAwOAZkw84XnQIgbzGJv9fAAGUDO
0iigynNJMisajq0sJlePerQUWhE00exUw6Wves9z/v2v+P30Jcqz8Ouw0QznXNkY
s092JN2HIqhrfbUtnu52erWRiOpMtpN2JCl2ABLrr+fIBZTQWQOgF5+IKhw7/+dh
XOweoQi2n4VOpFZ7pmn3m3D/BYtU9Av2XmIAZX89r8AytRyZW+6NJidT98Zz38sK
s9uGadrHpCtPTMgCBjNFu2En+FQyq7QbSE5zsHqmltXUw6qwInTLSggOZP2s9fz+
VDvlyNTsuKg+fS+Ngi7EHgTs81tkuWWpMrj1JcvRjIv+ni++jgQSrAgRPiBLcD9H
VyC8wFx5y51JGqX8e/bxDYAJ3+yS6tlG1GaN3NQdfUEtCm6yVEmzT50l0YfzUJGr
n/bF/RhWyNxmzOjuSowTiwTr0/kuDTwb4U2dKpwJ2q+7X3tX+5DKN+lCX8kv6x8+
IxllJDIcuOvVOsdsOel/FBkqg9UYkh5kr2x3YQAYPQlWi0KW8OtCB4Y3dZ8ryzNK
IewNb1pC27WfYpVUDD23pYzaXt86K7Ret2QEW8l8CYEcf1sl5SPzKkrSXZNPEFk5
oFgSHn/rqf6EbmXD+QlJE5OqWaJXi0ipdqPz2XzCuPmErWlM0Q47zcX2OlSq12yU
vUaAygml/cl+PHv4pWo9MmuB+As56nPzS/DAwm8JCytR5kNBz9BBu53SjcNbatFY
VjOSeTDUhgnIcANts/HxqCqGoNe/f18pllIh2i71UIcxX9Fz/Oq91RJCzL0y6tru
y+wzUFkCoOsqEUWoFVvAihNwndxZktDjpV4YS0RAXS07X6a0lnbHPCpyPzXdQczK
sZKJu56uMv0HYaXWzSUN6NiSJgZnWtKXcLxrJOkwtd5UR0AWkNuHqRdJ9/u76VWQ
j+5ORMKX0ZHGByL5y5urcUNMdW/iirSYjYvx97Qf50hQ28NKlw0Hcbz6JC0VxDB8
oDJfgQLSR7kHWa2ZbZpfAxrI9/pDS9ihiQAVzUFA9nIM9Kk+qoygYj0Vff2LvmNH
bKbgwpNKe5tUjszZ/RBTAUjMv/NzQreZahuoa3y6SYQCj4uuDZY5pkNyz6UEjFsg
Vxmf8TrjEhy7K+q0WyoumARuSE6cg/VCviQa6btCtEUMBJIPo4DXYalVkk/opVk7
s+GZTHFIlKPRT5k21U/YxeTdnErLmFDej71qKUjilKXwyrTWihzuxAdfHY6n0CY9
RKP62m/MQDYCNFR5RfhM9BZfqPcfZvI/1p6FRVuHlbdjG+o2oVPgK5jvQpkqAPMH
SmOGzX3+zaD0VPPt5UtAl40uVbWfcftMVmyJ7zCMKllJhvIoXOF/EZmzTq2yam3Z
bbSQ9icprZz6WM1gGOYiUbh7ZbX0dVnuvpn3taRvDHvR7QM1Z6xvjDZ81veoD2vI
KoAGBjtNBFRjEc0iId/fboHh7SH9urFcB/j4lxqg5Sk3k7TwRF/CBCp3/lu/z6/z
9tAi4QSFlQc2x5byUT5cvq8lnU4jnclhABy/PTWunXnVBhQDfiQ+bR8xVYcZXu/B
dFMFRdxDEEeTefm69UjXhAvpEymKr7dDjtwdXufnINB4VDgb6HJk67r9TYKRh4Yn
pW934FRqy6Ywi9O2F4v209NOhQcK3gslrAmI6O1bjeh0yjYMhTeh246b5FO0pGvN
MxWNJd/blsPjQRlrfFfq9jTFAyFXuwg69OEFbybAmnhTWVG83izKSz4GTYX7xHIB
5tcI6MSxbgkq8Xy/fohEFno6PSWjdyn4XoMUW/A/Ii+d5BTxl3lqa3YeKF+Rl04T
ne0hggsaWdAzSqrkxMinxQ7iEF1mi9v426Zy0b+wcsuJDNCLVV3SW0sXbGe3Gb/W
6JD/GqsVr5a2l/mMdN3dIUOG+MJo+uaHhMiibhTvdh+UlZWD3gNjKmrr8sj2iIcL
aWy9PeCgTg5AgS3VdgF8h8Warn/oh3/StVN2NGaOsK7V6/gHROcO0cfa0YQU1Jc/
GM2HKLydrjDa6kyOiIIxDYXTLlvqkrQCBYdY2r5tW6Xgd0CXNK3AsqJ0Yf+kqL5z
xiZ2JzgKmaWSiyAwOZJRpCyKsZaB0lJYkAo0TC3rb5XWYPc3HIl/JpRnaTZ2xUPQ
Mvf9z43V5YLVTGa+F/PNPQ96yVHJv1cGHDJVnwtZVupG8zQPpyVb5TIt+ivPU+Ao
jverB/otD6MOGZ89nLK5PafV4VTOL7kam6Syjw/RlzFptWqtx3yMaWIboDO3RYOl
CyzDj8KZx3r4AkT3gAmjmclx+h2frsEAiL/d/hPzJsG8uHqKBgLFJvaCNKnqaUjP
/0iT5ouqMk8oXLmEPdmfCJ4Y6zaAq6HaukGmamZio0q8ZdM8oiciivKlJreoVvJx
WDr/uhePIzGh8pw8CbNPbJajVVF4j0LmTM+nAX7iAXdbmRwevlA2KihgwU7jkQE3
JCscjAsHHj62+v5uB0mTOiT6zG5sWWIV20W+E4Nm/zb46aGGMf2dVeajUDqlI/OG
HhWHV3Yu4MjgPQKIPTlhlHuiK4eCK6u6dtwWXPq3oDu0ygRdF4UQQDnBmL7W3tJr
+/wBOUGLQiY4CEdisxl4LSarz8lpPZwx0vMddAaucP5PXXVxd2kXxqE6QLVQpW81
9c+STpytXhJJFILLkJqCQZUbjQR5andoKIywMN4JbI/Dg4WfRbRsq1cxcASEsHF0
fj7yoeR3J7bM8ukGSH58u5PW1qxhCbWgfRUoxisA3Yrqr7NwNhTe1quy6yFXJd50
G1UeyEBztge9SYzxsQ1b6xXJ/7jtC2E6TH9xhQITEfy87aAUNi4HEOiuFlEcDg16
RXBsriESlDCgWNyiZuscTT+8LhaFBWXZU4VEO6WPDdVp/CGx2pcEyhD+3CAYX/Y5
Tl1tOcTk149AIlk1/s7aaakp6PsV5JDj9uh3r9hAO90xFTkhNL4Qpzmge017yt7N
DYyFxob9sfpAnGF3Akkhs3NB4JdqjuE9gu1/s2i4JRgB2AWT6r0icHXklK5VGy8J
PQ4OxBMdeu5zg5b9yELFrnCEEebqF1hhZtosj5Xgc6o+93+ADSDWTaU/rSoIodFu
Q9CPTTWPOkkROfACrg+hFMU68zzPtk0RJXUWX7+3cEQWVT+Wco1QqUR6nJFd+3ld
6Ja1SaHHAW5YJEdDGYNypstUo273tX0G3ZySu8lvwIgaTW87/ie4y/5ERNpcX4O7
3i17DCaTn0iZFr25qWHMHrcGKbboSLxyfEuDdvTh2lE3BQJfUk3gdd0K+a5vG3VE
L1odsvuSsnZC3OOo4cgKuPJubJtU/Unu9GkAyGa3+DPdpoYQsbBDkFkQyAPLmC9F
2UwkDUN/NSeMhIWxMGXnRXLJTpPWumR5+qYZONzB6xEba1JP18HkFnetF0x6/D5D
mqltybXGAZIHdaf+u+6oo8R4AsOrmjMneFKJGf5SGfQbMah3kgs7OMFwhVvIwXyu
igVlyc2sHEToGrYxz6LREHg4dLw+34/r/6TK/Z3SnYRmTFoJmaxH6LefhBACtmq/
s++ryLKqmVX1eIDm0X0UKuesmiIFQNVsEO/i7URWw/uZoWHOz8olXjZDh/4vlEpI
njZwExFUlrHpn8WeOq4b2sVTiiyIJCw6V9EjbizaLWptFpFnJSf7IiqQAMv3j4Qn
RbLNzTijBBAR95bYeWkg076fR3adwgeGjZm47vlxgUSN5bYRJ3mqq8rlVul3+zAS
D83N079tA+WNQBkRXfvOl5dwxaG/GoreLMIBMVeCwuBlYuluezPxWtkYAGf4flVD
IwrRplTOm0pv+PJx7I9c74XygiwTyU5zpDhRJRtKwKyNQPJbswA8o06+TtQblAQa
F/2b2gdxrPdNPaL76ngfduS0ClWd9newKqtGNghHLXGalla+RD278Zb/eSjrd3tF
1a9EqtHORgmq8Tv1f38HI/sxkVY/Qj5PQk1wtL71rKmRbd+ZWEZvN3It4pWpjG2Q
m/6B3D+WZl97yUbq0MzIDPO+No0dJ2GpqVi1CIFX+7XOCv+eBgIjrBRwM/NdQnYr
nowlPzwEINDsUfdX/tMUfl5SLn5kSopSvQj+JcB6Pd/L2hPwzQzCQP6+UNanZkME
ndhjniTpm+PhylSON2TjX/PyUsvLLI6tq1dwECVLp1dhTD4LtLpKW12N9ImWBu9o
7O1Ph1EusgV5wVm9MogKnW27xIEw1Dhy9+kNXv50egUp6hnkMBSAn5KxvEIDxSTH
JBrADd53quO3FXp0Q7DzJgaRmmWIPd1f3ZZhbhm6mD1CcpGIEwo920vrZQCw4aQ+
LFZzjgWnxRDAeUWjnwdSwFD4Zeb8Pl25wIkZ6qvJ8eM7F0PsN1Cw7h668/Trtus0
qLlgAJMQ8BBKpb5KrzY/QQGU899yEzOWzC9w/FQZl6T1Psma/yu/kqyGXvGg/xW0
svUZKV6c6zkXOpgRJnon/FxDvBEiYxs8Wp8XuC7gNJXn4BFTHQYJnoWqnu4RbRUO
0EbuFZzXQor3kguIWJx+C/dRyoU1UCT2JneXwlX4lGZy95w1aH6WzFhtGq8I1fUn
fHrfqeUFENEbr9Il5pHoKwOvXIkw73wfFZZYgJ/7UAOY8zEt4/xZwh7S/alH0PDk
LDgQgboXk1Ys/hCmKI1d8nC3yvbo0oFOj32R7riLqxDGh3AP3xtMvodoEJGySM3i
7j4eoI3m1CAgIre5XCVd1mnf3Qiuub6yutYzsg3FVAeyNp3MHojuRL5uQc/q4MgF
BYzN23A9lXIrOdd8odCg47RvuN18Ot3ESYGT6l4pOBSd0W/RAwJIROobQQwZ3U6K
gYfQPPaEao4xCp9KYNy2SWxO2+1fq+yXPCBavc8Jm3ouHycjkWeigtpXn8HTPjIr
1+jb9Nyw36i5jxU+adSV0b4fgcpff3Zmr370Cp+FXc8NaaCe1rO/YLTqhaQd13dl
E1F4TPuveVXjRjREmf+PII0fjCimKljq6RqhV+oErf9NqBH0/55P3CPvHkriOU8C
H3rB//AoPMkpLXgI1AsIWF0rpeEviqdYkAhPUjOiY65sqGpon7P5V0FG9hEukYrp
JKFmuQBj4gHsPxQmND0grEIyzL39CGQgFvHJMtSPSczIGm/cZHKJJvpTbvTghFqe
JQO1j/EneadTw1N0sjy6WgtLLh/Ki494uGxK0pZJb3E1/yMwlfcPyredRD5oQYsw
O6KjUbSF/gZSTC7kf0xylHDIvRdK/x2+3uz3quY6vwbJsqYsg/E5p5glG1OszQ7l
Vs27ZZhLWMyIOkI+mMyFf+VRoJjdEoQxIrZNIjcBreOmDrjEIoiZwZjFTcQahWlM
nQ9wsWLCMVF1pzvvC9ywEbj7po1KHPoGOa+1578jeo8/3KUwC7EAPKJSvWSKqaPw
WpMbN7Gm1OacHDM4EASsSOg/oBNq6+czWdadoNgI6OUzyT9DLx6ZCgXd6yhS8hEf
oJF82MPE+o8bNloCmxfnO4qH3qlZhEFXJNukaDZD5jt12YhhBvOs+pYg7kOUFB0N
CQcC/1FqUXE63j3guB8mlu41ulEdva7lQOr0Xtdfb0TyAfg9Ww3B6OPV8fhdF1oe
Sg1lHEAwus9BTKTfTbvhcZciH/waqQnhc89X7RphXwNZ1+0gEADUiPHavpoX3/11
SWiwemNNjAXxxnm8PG6T4yMCklm4uT7fKOAfAS2LBBJBZFYzA7Ct+OaDOQq3YcVp
H9lecGfUX/AZvI076tDL+dwNrRf9zxzoTMTB383ktcamMtSVsmCfxaD8FHlIq8rd
+ughMeoaudccffQ1NONB90dAB1fCUw9VtLw6YzCIQdBTLX1shhFy+IxwfcbXOFGa
0PR2zVRjpLO2JYVj2wsYoD2B5N0vngAV9m1ZktUh5i/ZKW3arvGIUWHDG9ekH5M2
O1cg/CqPNv4Pmv5ZFEH0XyTI1ckyYyPjaZ8zBil/uMC/khZ4E5+Fe3KP1XemdOdU
bDzg4AaELCfXJRqyyWKEgBDMBZR/KEluNORGoA8Hny/mkpjw8rYIbAF1TR1B5RCy
4pTJdC8Mmvuiqpxc7QAkyIeJx2G79p/TPdDGs/3FKfyjt5Id+E02m7JrqcJOaJxK
MFx8hqklW7Xi3NSguglpYvy70R08LwCZdjjro1YTyamCsNmmkUSPcjWS41uA0R5S
sQUfQH/pkqSag+HxECtMrKKDKRjEJ6GxHeA/2MevJqI1gQwCxX8yNmEGoaPD4tDb
pSrSO2jXruQm3R/Q/C5q9pAfXrCT7REXvlCA6n8zWL+WjHyxpZ9t9uqV3Pr712DG
P50lqSeAqyOZM1yH03E0W0f7v/We6zeK1rpWV5LMLBZyQmUUeQko6uDjR9xp+WUY
SLJeCrBjF3hT1O/vBgs+dhRwqg2bH80EiooviO3tAZSj+YbQjeeegA3iUgInLDus
RmfHMAMAkTSjEaMIlRW7TTD3XTutPCjr8Me6er3uGNV0Wyr6Jciztxe/9djJniB4
IbpmuWlojhLdybVFUcwI/c/R/I+71/oz3vttFUAKs2dEgH2M4W20MMwVT6e5E1j6
4Lh7b4vYw2QCc591gSv1z0JhRvnney1eDSysjyTOWz+gQbsASCKH2GehupmCuHLA
6fh7TzmvOE43GXDTRvvQe4yms0hPZvQLFzu9sYhWDvI7cIHFzT/3BdvphYtcjJUG
sWZLn5M848jVjxSPv3Iy62t2lVfqCAoARXjxXP08YsDDWenw1MDA1aeFgXkSA5G5
P0hU6n27aduE+/aRQ9Dz+6z84Ght1ZFm5SG2cCuDL3oM3TscuZHlHf4FeaO+7MTr
qBRckPiGR0DEUehApxr/44HZWeSZmqqMioBQQmBBAnWf3QRsbGctivHcY3weizVi
KqMme/6Ft4rhrlRCpK/SIcgi+s1o6HZpfhTURXTDVBYzXJ2I36ogWW2I7L0DPENz
IB7bdcUOB42OZwpYnPM8uFP1OJ2Pyw7EEJo3f6WfNy6LG/V22m+Wd5dUNY74/qTU
UF27Vjf8JY02weCIoRmEAnjTbPoyWDkMU4n88WXguMZ+gWvCpOspQpk94ZxbFmBD
tYAn/+eadH9zoBT6s6W+jotK8MwyF6+Waoa1aufJGJnNFflMfW7srhSIM2iLATCG
IUb2c8RQCkFeje6v2YwBY1BkgyQoFtkz5MkGlH2AU75V6o75q3FxKMaoUQKmVLub
38JHZMdsCjRKI1fNEUDEQazwPskJh0ZPmnUWtcEkAGBvPx4/JgAEQva/fZ9d84CT
AGlf8isPdkeI04JlCjsbAdpmJmUZuTFo0U75azjfd/Lh+g+izf0ToivT4HYy94oE
7vu8M6SeAQGD8bxaARObDobEOZLtAoFwXM1QptjF8cjnTN7fUF0imDkckzD7KCmt
8hbicqXW85RnfC/QuEkMR01Wx1JTegF+lxHAt5Bv0Tim5quR4yDXZ4AQXXUXFYbE
gcWoKDy/m70fz6ye7Ecux1o49Y6Xtr7dFC2a5bpkAiIDOzndHCM1qlntkCiFzpRz
wyIxd8AU+W4E/+YsZo+bzdcFXAxjDtU5AFNr4q3fNxmok6reaoDVrFpKP3rIxw60
27hFOSiUr2CH6v52qNP+HttdPInIAQNf3tZLDdm9KYjLSgVuX9XEs4RRKeKlh7MO
0SBnR7SQwlE068z3IHaOTEsIe+PNsM3cpGNdIwlM9RzxnSTdJo7AUJertY4D+R39
r1R8/ilYIVnC15JFE9GzQ5k69b7hoEzlRz7WL1GdYwkK5Io0vVdLtOZKHHusCZfM
336W7jQwynIIsqLoFZeP6BrsbawDn6wZnyWpRahiiRFt/Kd6lpRNyBv8qUGgEWFQ
Y12IMvrXPegzISOxhHO9RHCxiqS8FE/XynFP4cWSikwFtsW09m/KZK41t9RONfNb
Xhu6GuYVtloym+tDyihwLes1iV4/95TwVA1UpsXjJAX9pmCLOSxCGJF2GYWEkNRn
xYJPzYVhrf1yl8T9fm1Hv2KI3lx1oTyn+k1O3TbUQkmzJP3ksBefSYVnOlu3MKBJ
CZ5l9yLJtShnrZKFN9oBDm/gDdTKhM97mTqiqjq+y6cmtpewMONvhDnBjg3SgPMN
gylIuq+c96qTsw6LPeXTDio50DaUHvXkHYNi2FKWREnr2ilHr0gkD3IXZZACqSD4
raX418Ven8XfbJBr7UQ5N51PPOgYNyhsnh2XZiU0J7F8SPy9c0OtGcSlq+AqLp81
qjsA8NsCy86nhREfd9R0FMyZS4YpzA8F5JH0tVN+rnI6l5VUNACoB4K0qn7Jzo+Y
+ZC8yiyJXyVsUTLWE04s3Ev7m19s9n597sIM6I0zwNS3+MIOLPoFlY+ZIERts7A2
YEeRU2lQShWoHt33AYydLyK96M+YDvtFjiPHAunH83FS23rFGgBV6D1Gom0Kzmou
d9jmGVThZ9IySALgfpD9RI0WjIxdDs2CfsWuFtXjkKgnz1Noqo4XSBKPAUotv8Ey
yvon+4mplNCYhjrT/zdWseUML7lTxgR0HlQJ9fZ9iUqjDFERhUvrHDdytuVjfJf4
gRrNZjG07OMvcAFGwjmWz5S6n6B+wMOjX36s8yokFgdzkRqwbU1kHljpJP3DNLpf
BGOX3v39esoJ+IDeEsp031Pg4x1bUzilsiWy8oktq04rw3u+1Kue3+brZ9VEZXHI
JValqGJVtRw1zjBU4PePRK2qj86zPadN6e89JU3CE8ddi5HHJiPdl0/iEOh4/YuI
pnpyMtLiYbt4bxQQrlE40V3LVbg6v3aINx3TfHKZn+jv9ToC0vaCZR7NuGXvwr1o
HH8yFHtrMkvGXWdIRl5D0DHChana6eAAPelayY8pgPsSiurNWKvRnEvhhMZCx4ZU
OpFcm1g5+pWU2NQ9srzbXtzBCSRbCc3vtuIi7ek1KyxPQabGt+7AcNqRHLI06mdJ
V2P1Wx6WlT569mqYA8CqfmL3eTlvl+3sGT4jsaMA/QKQOW7tkGztMgCRFGi0uXc4
MeuWUGffK4XCgKae+17VGnwP17IQSYFnhiQ7j/SKmKpUQUwdNiirZi+8hqfkVpb6
4zybVGnVTu/jo85uAKfbwm2thCrLpz+ZnAkGEyOTeXNoFYB+KryaUeQTuY6Altql
eeb+AMpS7qyFvPqnJpDwu6rhIxo9/Xq9fNZPUdl2B0zdy+KCUxQgPxvZE9hhkG/0
qsbYP44ZhYiVqCXO0kL4ZtQcJ/8P/ioRvIEq0LMWSoS+5b3dShd9sHAiCJV3s3Zp
idyoicKLNWYNE108kHFIzai0Zhel/aQvXj/0WVmSmZqHCPh/QG7oXC58EfcZ6uAt
7Lumxl1arR7rMnslJRha7/flzPsYPoWuRn51ULoc+hIgCLyp46jqT/jPQp/JzSu1
RbG+/LPWFe5O05toCisdQIK5LW5qba+mX2D/Niyjn/oWVGBMeuBlG1FRkOb8zgX7
zGY5Rottde5Zawx1ECaBQpz3TCbmsa+lKuPrwrvwmSxzPwYQGzRb+cDSCyWdOkXE
mgEi+whFQ/c33YlY/z6DQd4RXAv/api0hI8WARijbN32M8B9te7fezMunqzsUyoZ
kPHJPVSdJG2D7DGK/I3YjbjCRQcW301XgxdT77T5a37r4sieR8kxj1mDoUuJGanU
CqqL2NHLecTK0k2g/b2RLkqP6FUmkPzqAQ254QMEEtuS+O81GvhR8C9aGswjA19T
XNGWSyMqkA8xG8sFTbvqXNVROGSBIHhr978DyGWWyEXs48J4MrgwqAddCip4Vz4d
5CKaB+TNrctxnFhK3aoJorUa4iwQCEFVdnlDpSwzEQxBoLFNHbYiQwAPz+urdZ20
Gz73evxvSXJng+efjgO0JWY4lACJsSFthOIFJ3kWTqQ+igduRs1iC7MLh0e5WTJ3
777YnuFF56Wqf2tTnA9uKlkrHO6VV5xOw7VbxlJ09DsUx3d+koAP9AVV/78/rmaZ
ibLpQvkCHbVgUJnXJqzbyCrfEmSxFCsjzkpzpX2nPoRMGu0MT/vA13zMm/+vH7ih
zNZ8Ef0PTXDObV+9W5Ddsagg/jJZRe0Owgh1+TfpwthYiP/1PmGzdPBunMfqdMUN
RDZJsVnC1TeqRJ5aqHS0hvOytkNr8FwSX5DRTX2MNaSFr8/UOFEB5d3/74q5zQ1C
AvHB4TMICIKMp+arDtrhU+i2d/HHpdZ/60y8TAt5vrtK/81eNweb3FJ6QDs/L0Pt
lDo/XVedBE0j94usUUdsx3YiCxCWLzu6IgwjdIkvp4tQye5QhG1QWZn/hytukc+G
BaacmW4NIvu/hiIX9TBfLGyN2DH4ZEKhjssVndiqGZ0zSRpl1/sASmLpnnlkLjRv
zldd1KOFZFW8+f1z8Oga08aqK8NgCVV36qaRiW5OJaD1nyZzb8waV1N7um0v57Jk
Is4vvGRFt8wwRwotEUCQx93SyEx1fHWGHtfnxIo8fs2gOsBzrZsSYUVtq+DaR8vZ
rkQ5bR/Fk8fbasFvCHB3xFgaEAnwU1KE+bbqKxhcw2JUprWcEXwxrEtfsH72VADl
Z+j824sLOaQq1i2MNOGR/BfrE7NlNnNUy3RasuyeL33g0v8BPcaQ5iKLn0mCef6c
Yqlol7q1C/irGW4Wwwx2CkeW2NcGfgijY3MfI8Vlf42yk6xkSzVLv7e86x6ocWnT
qSGykDhgAo+JRdDrgFAnbKd8448xKAVeIU77llu1yxn1pjLr5eDq/znKr5Lv4V2M
zUpRZCtHOU1/2S9hv+Hgpnf6ZxtAqZuULkKS9stF1WypWApe2H2YLkvcUIZl9BYZ
W9afxJCGHCVYPocHEQtx3a1PchtWj1DjZB5M+eo8n5Uf0h2axmDZWfD3as/d35Bi
0np29Cg2kJQwa7q4d6zrmWl6F8QonnKGCPZ9+IyfEiYAZ3WdFTiwuGPTeviVJ0yx
TqQePyXgBuI9qI7T+TVuzJ3oQKL1FnJfM/fWCm7QOqMV8Y1OU7VZebeOv6P5LUsz
cGpyh5osmvcLv/viVv1GxELSX8mz5k0dWticsboR3Li6PbgjjSHAB+tZC/NekTFE
LbeLdT9rAFXZLbEORkFfksXWCU+4E31lm83v7kN+X/5znZDMsBd8W4mk/WrFdZaG
u75G3vPGoPfrhktVWGxCyO2h7UFpFLqIh+Yj7uF/tWzwAjGGpGDEl41EizJ+7PKX
BFwD7YuYLZFu8IAweM+GU+EOakriuCYQpUf30rPqNf4QdNrr/E1GPlS+KGUo2s/+
CbjyPSfWmoDNn+j6uvccxrwC5P64ZXMDVRm9U30AIbPyTZvP4Mtsha+aY3Ok3//E
D8eshDvD2hENcbrs+VC29flpRrrIdLpnQLle9tAxnOiTa27MGE1z8PjtuJD1Eyhk
VhmDZX/7fW/f/eQycBB06LKz5bkk8CPgKh11g75Ii6ws3cEStlSTKQwZ75ePkeBy
jj1MRAo/HW7MAN7LDoS4rlaQtYkHUQ0PAaE7lCWUxbQi9V1B+uwzzvAzeRev7iIk
MnC8bSrs0hwGqluE0nC8xvnFy+mjhvz6BMdd/Yx2RuBVFXLoUrvyV5I8AHan7jl5
or/6ge4+Gvv6O96mNZwb8Itkisk9sogY2vL5wYTCHyy4nmt16mEz38YonmTGXo20
xm75zdMNIpr73k6AU+BHDTc4UcUtWABpcXN3iBu7FUs9xwmZNRo0v62QZiGCnXCr
pxwuQs6xFDz9OGlM023IbLubpxiJzrPL3oV0uepEr0QG+l/ibB3d61HroYv7WKcM
+ISqHem0bhfl/6O+x6CEPUMyBw7CS/K7ki12jY+nopB2qt9BpUDkyq+dS8lt8ACN
P3lrDfsv4UH5OX44lh0osnVmz5BvDEEeUi43mcuX9h0orWxGxyXYJoj6/dCrmL0c
pE2TAv2Uxgu1nOMQABthcum6/TjkeHU+E0KY9FTCvSjMiCyh2ckyx1Yjbv+ys/NJ
oan94C+iovI727lAQPHSSQzsCraXfhROVzhpljzUJgAr+fQKH0/UM5ZTc+R4SaEi
c1+eeGg5FxcZlHCjKjR9QUlqznK+8a1x0wz8CuDEVJBsCuGBZOVR7+AMjittyHmF
oZ3WlqwcFqgeIDEIQZ0gbgzs96F6oAwhNiFVdazLjSoa4uffgZIAN5C8ZajMdtuq
8ephP61HDlJBn1Pxz17iwE8lkbkxa4TX2tVGzCEmjONR/cXAEHvCqxZOyYuD+Dbd
D1Z99zCrWCBJTEF2ZS3R4vqElo9OZs0W5fdGkrBtQ56TQAa2IeH556H74vjgQzSb
OjF9bXx7bDHhZZEHvZXSorxl0u/A3ClkixjnsvWvNUbOEf79CdLrpR8WtdSYZSav
q+6YJe1vxgVCEzGfmzqkjZFVFGbcpjq05E8cBqpsFPHUSFWG2g7bv5KY0M0MJx1w
SWYkJux5T04rOr1nnh3Fojl4wAX2gwX44RMMx1APYC3jGaJHJpbNm9flOLWVsSu9
CR3O+BaFEK3Ip5b/ZNcSj0sYFfhtaYPWEt0dNh2bU1aqdszYfFdatvLzt1vWrO/l
SQQbGWpbGcyC/KAbHk4/WnGvhtROJ57ZnMvjKC1xzegwRTN3+yvwI2jaZ4o3sYFV
pFEL3DpV4pbNx8M0843HJShJjkmG+bGMjmcAX1COOZ8fTzF13dFfEcDft9cs1+ZC
0BN7Y4S5RzUHBpmNMgQuti45qpUTp9dx+xXJ+z7YSVR2IxzgZzhXQpltxApJfKYw
Dh0UWf0CbZZIlnAMAZurYsHEeNrYj13BpFWFrcGFqUEhojZAF3YZx524pgxbT0Az
07TspTUFJTgk4tW3usV4iv0+EgRl2K5bwyJ/jDGZoNa0NoWpnz52mCl3i70zRpUt
AxVkYXu0SRArs1eOhzim+AMteT+bZvfR1TX7MdV7FgsWYifU41sFEzqb6m68a7/q
GAqPw/kq0aKs49+IpX9Ex7jhD5cq0Jvc4edPbv0DwZarj2Fas9Y1QvGaiCy8lHtQ
GSqn5B5c9fSGNop/zTU2pDCicyuD09nPjsFOC++fKIMmARhj5BqFfIPJ+KZvNPkL
lTKRZFtJPcHGSDZoIbTR7VGgktsVAbyRwHGFy58JAdSmpP532FSfOCWXMOOd8vaS
cvEXPLEgNY9EC5lweBuWaiatv99BwUpPIcygm+HcKHfxKPHqdx2rFfhDgIkOcffy
U5o8FMyVhM94Ixfezo4+RAfsNyLOlDUEua1phjB0ZwdeHrnmX5uh5mPsFt+GeCOp
bHAkA/tMwW1e05NR9faZvsE5T5CjvGbDqt57Iin68NXyxpnP5ZypVZevFadjfGrh
Tvl4uVavxaNxYmZrcY7gPLRYmIdAGAaRrXmzlSzXnS2J9ZtM5dklVzGjRCilx/5u
2atHe4G+cnSNB/0MBI/MkDG+WjnxR6z9HD6U9/7z5b9GSmbgQAGqMRl+AZK0AXAc
BjsM4TKtx+d8qS0E8dRkYhJYfkJ0F/3C1xgUJLvTr+pFecpyb7FekKEByvFTuCZ/
0vBYWR3TR2oC0DdpDaJ1DhzAyDjGKckaxyfvVbKs4kVj+e3n4K5Kb+oiDWPNjLMf
AJL+htwDyFN9Nwfut9ggBJSsPl3XWZ1Nds7vT80kk2p+BJDSlqmr5gfU8b3jZENW
is3iDN7PAY7bZ6FcejX0Ikjkc2gtoHeOWdqM8p/uy2anzjBovkohBtFiuSZksV92
aULFxgdT8Tq1+uUHo775q/rILZHbNDHd+F55JRghvWfMbMyNO3kfGlnQxyyTWSNt
1uhulVsIHZdXd7uV1AAlJmmz6qBkAuFcqcSc+EgM99ke/2ajm7PK1aSXK53rnSlN
BXdKb4ogrQ4ctQtsB9KXlD7kj3fEYOpcpHFMypqvnPnTCsdgBh/XQ/SmtSLrJQGX
EbAMMTpYpuFXijIOZo4DNfXZoYBBHQtPEXtKwRHSI3bz5+RfZT+/rM2x6oxAJJOC
wu9L1og8oAg9GhaGEqrWwYC6lCFgHmkV6A7E029OWjZl9na9QQSBLxB4dmNlkGXp
6WL/jtrqe0rrWt9B64k2bu2o5QY4GlfgT4wJtQkrTAZ3ZdBzczZiISVsN5BjmKgi
RJpmRJtodZUESZ1z5udvCTw1b5EuzQaEDkvDlgsXm0awIincqSsEEubdJuk3MEXT
y2Wk9axBPCY3289viFCbKWS/gpFXXq2qIMnqU5EhgF0tFHoz819iYvQzgp+P2w6m
IN3jhA6R6qd7b8pjjZAswXTJ/zY7Z6zOleaCdfPX1selN38qeo0L3RXCc+Sf3pb6
nvg+LRu32JbWujqtn57JW4YG0y2zna9qaSPx/q6NzCc+CMZq81+LxFbIB/hkh9Ug
9FO6eV+O+ZWW1J/Ui7VK8FTX31eqBjhVaeEIDioucQ6p/7Ad1GhhiX+fQsLAYRhB
aZmtcukKLLuQk2/9bIFOYY6vh0LV59dY6Wtn5Ip/ouiZPcFHgcRGlFetXtyNfb8x
ViC/W6d+2Qwm69t9qVu12KjeBec9VEVzouch6aSjWqDAJRn2rsL5DlWPev8/qmfY
EQcSaj05jsOjbQIbWFp7Qf/6fZgfG8/SiM+4OJe4wjs0OAUIx2DclVyx0vriqvff
1IpKCIb3Gg8kMovNT14bUx0D6s8JaYMhppQZ8SvlWtaSRyV92lbzxf+MFwkV5To5
rZLieu0i+1pPNaKi0MupXS7sEi9fp3XknTdjnK8i0wIHPM+8xF3ESWjV7PRxw3Fq
qGTkpuzHg6ghBWjoCC2zfvM2NGCDpDBLFdc822xHv+cg1IyhQ4VH6CfRvgRmUHQe
Ud7M/oUjhtwJ1wUoeA2kB11wSjkehQMsJ47fR6m4u0d0NTxo13/TFOm/o8TO1A/K
dwkwBibFsnrQWSEck5FOa31S5q5FDSS2gIk4izlxpAcetK9PpJ8y9a8j6lhOWchB
gvV+pk878tqQSkiEBIbDf8kOv57MOg/c/nVHKSB8N1mJLnAryaAmYc/WSu2pfWCo
6nxSwWYwNuohD90VU8N87wUl4cfwO/ezCyU3jss3tPXnRxLvg+2G6KXw6Xn/qNgd
5Z1W8QI1Glw3bq4Y2E3EIVXfee0RJg0Bc4jWUcFhu5ewYWGMTd5sIJ5So25NIqzS
lnd+jO3Bga7LCTrUA6/PGOQfUMhMXA0RfXu3KDsVoZuqBnyJ6pE4c2is9ZzZv4zI
CaIfRq29JZoDY8Ghc7tB1KSeYE0kkt7J6VVVUlpTdX2bpaHFR+1/LqGQsGLP7zcx
JQo/miX7YtMx6LqR+k6dGNqAPSH2yz5UltCL0DqOfdgr4MK5J7v4OI5NaJ7P/mZG
eA0hDMT33BNBisXVGsoW6qpus9dx3wRsDgNZxPAP+T2XEROE1VIhp0xXsXOryTgb
BMAgvpVfovCFtuJzw4V7pK+8CyORRPricbQK0jZlBnQ0Tv7FWX7WenWuugHmhM/J
3D6ckJmP41Q0GGNGWrLjXv5Po9xWjts1qn6wSmEBqjS+2Is78hqfDqFRjiaZnAq1
1kUny39vJR3UZfWT/3xgrajyAFRBJpWA1wiVgg76bdhlMBfwPdcKMDX/W61oP2Gv
LbARwYXkfw2w6dTUxvRekCc57oMy0XP5pFM6Mc+G2URF9YTlkd6og+JEpm7mvYuW
1ZTvd31/CikPYxJk7smlq2Us9hQwdU1n1uzTGj6MpPk4IhLovhNRd2hJyT3bm6nV
g95vXYwy+/x3KiPjJ+9EG2GOFHwYpD82qN84OqjxK1WiGVcGMYSr4x0BAxyhgOcc
sxlmzQ7YcIBiKeip5Y+cnrW6Qp8zMnkGjx/e7SIw4AVB6iWQMUb0b8Oi8r7jrkmE
jjvC2VRJGPXLsgMvmkK6qf9qF2ygG5+ROC54gHk6UsitjHhdMFyM2lTp2EmeXaF6
69val/ijCf/F7aHjsbZfpOWawhkJ93eetNsIlYH/Emead85KmzUdBoKZYf4Yjbgk
G4XnHHeoaNuSuA9xuVTDvhnU80ZMa1Pu8BTUdqIvsHonxGj1ZOWwy0BK7LjxsDRB
F7UMwjJMj78hE4CaZVzcL6ycOg4r7tlw6geX7cdtZrMtNDurWXS2pQi1pV2FpmLk
P+OYtiZVXq0hnyMc+iFjF7q6akCtJ2DCrj5Ogc7NLdRrpNABD9y5fGaodGWidMNw
dyNKc5oaK4ZTR5xkAJuY+EnOHAPigB77naIdXA+g/z+3iwTat0pL44GNbTSZzbTg
WWwsFIfTSBtYzE1IDixJAUQQxRZ9ZwkD1vd2s/R68TxyZaLCJhYzTYzuCGAobNB+
yqF4ROAJadABb5mTDJ3PmJjP5gcN7Z9gqSU5uL+qYk7fVjutgGQf6/69V3V9PwHC
2IfcRuaiENr6Nbw5pWFIKRmjiS79r17dOiMg0H5WUzDiTPjqnQNVhX9kxrjJG79D
uN+vMv7jDOJ7ktg3Q0oHY3EBiJ3aQPqHRxNnV79Zru5PcbMg2v9l9YBS5e8jq0GN
ewQV5G1cAEkW+JkFqKjgszjSNef/3nm/ADriaG7C2WFKgn0726AYQeaTVvi6rGvz
nd86KMGbCj4ITed7vJSAGeo5B/rFdfrbSkDdKawBLAnmHfb+z+1LJPCASYboG8Ya
gKyxwDcdzdDrSMDXSdAfmWzQcNj/tVgrfkYG3/LnGxRq3I9NVouegwOsBV83gzIY
OZAvfWKgO1zIakrbDaL6XEiV7VxQb2VTC/0i5bg0E2DnwurneGom2hLpo1Iu5ind
1kHz3A40/V9MdQE+Sk3GuFJ5wDrkB97pnFTEBibWELS7bpBWjBaZIeHwrOeLnhHu
OP601uRIlM9K48eNtd98FwU78waj09I+9Wp6EMgJ9X0M22vmzgp8Q1z96BqKLc0T
Sbvyn83FJT1oR37d36chXwul1PP58mknEbLVEMkA0uXzWb21sSbny+kK5uehCnQp
kp6uZ4E2S5e9gbSusbiyC8rabq5ReztcsD1pUwT73hEFMUeJdhOzJZd8NikWDuKC
ANGP69mnvqZTLy8vKGnprcfO2TuvccEgaACpyNHK9uPYT+zusPQwj5ZaKEiZIKY0
qf3aToLjDFK1plsqUHyH6AyDkyIKoGrfGHEWuTU5wmLRKJD5iCvZYUQpOFF74SaY
Y9EMnsrUpquLdZTV0Gioo5ePcPQyMTv1VR5QSwaX25iBt20Km8QfgjEXXTpvYWT7
GA7EPn6xHqKbEc3kl5s22o+qTNPxq/9AnSdtxUg9G2auDCDdSEgGPvqAvOTbP2zc
ie1x2PbqeiEojSUihPW6TV92JeYRYGSqHGEE0vRekE4EOG9y3bjHdXscGY6AAHoX
kdeAB2ja96STbTjWHBy5kZsAbJPSvm3RXrjOu6IMFWbl/33X1Gkg1dRmdSe39Z73
TjwDc1sTg415gS+gbV/5giB3ebT3Bkcrvv8/xQne4shLNGBzBXXQxVqf0I8U/dnX
6Hi6d8Oo8INpfvgKPLGsozybNyaJ1yBUokzxyvnvGzTJzT4oKUAglOXyvx2tEGPD
EF4pjIMoqJ0QdBHgkLlNhJemkZmdY1OA5m7FUKCs5VxrtJ5frB696MJhexcRVaPY
tmwNhp5ypjO+AITnKVdHO+qi1Ihg1o1cy2nHwKvTlDEgAqurupT6fJIcio5v6Rg8
9FgPylFI5OWgOoeiKdDcovgNRBgwSGXEL4u5binp5+vqEMngSBifnlMspa3OAGCJ
zQ8NU7JTVZLX+oVPjg6f+NSIKy5BrqNISAua8Y2BcQir87mx3mOcpVYPpesm1QP8
/wPpZsahyDpe7vAdTlKVnCK1S6ect71Ssx3Cfrztg6H0Fqno3yzDSLHs1QBLm6RA
avDif0KXn+SQ+eMnJkH7vmn+MIbG2kw5fw30sparzpTwUvBI5qI6Bnc8n/axghy0
Yfn/bnTjsWc5no4RFLKA20OFhPnZCpTy1u9sn8V9xffE8ucA/Q7m0SlQOSA2FHz0
GC0iqlhvHt12+T3kLgvfkWxWoB120HiEaHj+/YSBGWho+ifFExgj4qUCu3MTllqR
6Oi3QnetwHahJZhaGFI99vKc4B+BpYeewPdsgpu5w5gdjvokP36zefmYimfZGW+I
6d9Zue0JGBdPMYgKbB7mAp4Deoof99WC+guPI33yD47o8gwmNA2WI67VmXuPMWNU
0xBZXcoIb2ek1YEn/Rcm8mXiiuFHyhf9UAUeoDTcZ02k2PgOTbOV/suUmy7ViOxW
8mYmd+vVWHOpQlLk6G0XfsSMHLXufj/3fC4ZN9tT7rV19HhOZHIdldUjLr1BbVBO
k3PFdCuDYq1eemNP/ioJ0Bzld4V6Bx4lW4kLKTLdliokdC29tFOCgtjMmyll8D6P
bJSdqzc1DU/no+citaDOLh6lEkZXvEENM1gT2DaMz++KdyJFwvM0NlfdFbOr/LhK
6eDzTRIYf1cXUtXqsh0vfmtyaLRZP2me6DazYZqZ5HAmz1G6k3thTb5C73iEhMNT
RN6wk8+zmVFwBbZE5AClsNNmccj8oXr756eAzQfEDd1emW29UWEBZu7rejy4kIag
9IEj2D5W8QmXE3lo0HDvB7wWdxXNtmuJNJPjPv+sfrJm4/JIPH2kkUN2cGk+0td5
tG/k92o+0+Ek6VpUVUtKcgXbskabbIRhhNwDsw5G1Gu1OwEUT3JTYZ4N62+hLsX6
R7qo1tX2EWZXiLqgfLNNv7Nr1Vj7vmvYg7rYIAnyijbk2k8LduLU28tMVjm1rcV7
7oLphMWec8mawDjSaethoPrCgkvaa5RrjMuuQpxuIiWKT7pPyh3qHiW9NA0vh3y4
LNejWYhkI3++oAQAT1Ar2bAwo5jQ4y0EcnGTY7GgNcQp9u2ErxHioH7JnPWpphIK
jKcBcv2Bt4ftJlbUuln803dItAputUPCUBQVhkHpppJ27BPI+snNRt7pvpbHUWdD
i/E1Y6QmLXE4JtW9MlkxbdPBJKrV2xTjwD6wZqPtaXe/aW6hDOPBrzEnb/WnLyI1
vcnV7jSEVOML7AKolMXgYHPyBF99OnCDA1mBmBNQ2kNjuFP1rFNAV2re+yJCmVVK
8iHVuaSgNrb+kKeoEJRE8YVo48XrnEWtLRhV2F5B9yoC7ZNtSArXpyD6zEGOCcDH
MCcgEcZHzneSf1H4qgHTqOF1GHO7JXwbT95LOn9gpT5jXItPi4Yiy4lbe/OuQAlp
F2CcSe9fAjdhLAIbkS2i7HzbhMzruGvnI1jJR6hTutsWZPTt+HhIGlvf9EXcO9Fd
HcAhfu6aTybg1tdsiNPmfNy4IYkiEZJqL5EiN1S0a6iVxP7QlANPnr9UFd0xyTJY
986N/UQOBwjmRotxeqOif2ejQ8vq5CScO07B6bXaTif5kyUuaYnAaKle/XMEX9Pz
xI8po1RABpSc+8Wy3ib1tnwkJyRpaADYwsi72a4txQFiFwqOPnx73zbFYBPUwP2j
o9ypKuTLF/8bzJE0pxckqhLiAwI2dQU6Wq2NBneCzHB0ug21sWvxgBkzTl654cCR
jPN0329mlqFjjb/qD7UbrhuRt42YH4enI3iC5CPyHIoBudVvNs4br+8DyMPuOQQL
ieUvs7pPSgSyqlxDExTr99gh4koWnagFHPJ5FDEUPVJuQARzRBYpF9qvXOXQ+InM
5mopLdkHGhVIdXfsaFCI0k9aj3ak5mhcFo2J5WAx2zwtkStJLHjgVMIsbkjRJ+8O
+0OlUMZNLJ/VTRFbzSvuCDUcsglv3R4s6WAAnjcsOiS4OcFlb7WBWuXAeUf5vDz0
EL+Dpyy07PzUzXp3/AoZSt5BbSVjWb7NfOcA6jMoD5vRvVr/y8f6XsiHOXxwNTcb
YLW691hoKlGLBM6owZ3X5aaJbNEefT6+hfLpk1BwWX93vGVPCOD/UKDFrJ5jAGUU
CBugK4qsNBkhWDrHNjtdK7gCCVMGkfiRk57YOs5C+6EfgeeTqPe2LDU6g+tLHMjD
/5r+kAIyO0hF5Ax1f7vu0tkfrwTTcJnTN6N0x+1vWAmI7vv9120pkgroar9ldzDZ
8b31bnMX0hsmsD+vDB54MPxjLpygnSNZURTKeZIUOxp4Mq3aYl6DXomhMdQKS1ka
oqotkJK4AAJryjyvc0xG87iS0l/2pKzZ+ZRbbxGcyhggD5egx3vazVwEtJN4Jh9h
iweUybqTk0j9gycKZ/MG7C6C0apKCCSTrmEJFReXv3WbNc0vEHo7HGviSSaBS1yO
GCLf0kgOuaverPcQ4Chn12nA6T8By41MJzcgOhJkjXwhzLwVBiGKwBxSUb2Yh8xd
q/F0o2vZpMO6YXnsHoX0QQKduzlzEuAqDbvwnodhrqG3eacyTw4m4Q20gQPQOn9Y
S2kdN3ZcsPPZNLJw+tYbsHk2Tcuq3Cv/9RUnz/88qnB22pi9s5bGAWY1qYJWGp8G
MpLB+TEzIMf8YksUl5lpk5usk4AvmOQ2QLSyti90YdLQ1wHdoZwwE+LZw27XYFbq
QvzRyGTy50ymNeqJeDhCWuDD90vTqIlOXfRhy7fXcOVPm8eTxN+CbBMsjevQaNn0
ZN3E5qIIZCaeyCSdgjHV1utbnb+tEfnec2ca7OtxHpca7mKhUEwDHZpmL7nCP2Wo
CbxlT2Zc9F17Dx9Z8Dj7RzpiKiRx7GzQVXhaeEvMfKmcO0V+7I/qlcqQdI/E04Mf
gXHkxqbsu4v/aWZ424CYZneMmbZjRRipZBqHDgMNghOq+sP2ukCwusrWq4iUtvp8
XsLTiLsq8/nE8tBKb9PA8s1kJo/is2J1N8k22TyXIOytLhWoBZ5rfzdBe+Ud03cn
s6wJxNxUL3iFxIs0asbvJoLn4zSCeOKyJncxbs2mvytgfaUBjfLLnBvaBB/LaqSw
9UZ/cELtRLI3PJKaZIzKhiJmBgyQ6ylFABsWHFSSHL36926sBKiPW/XIdCaPFa1T
2UtagYu3+GUuIMUIY4gl5XR00Iks5Rr7sF3Nj1Pn6qwUlKgS6EEmN3Yb8Ye+s+aS
fvznf88Y0UEIjQHJV8hCYtwkzvZKkFv2acM9F3ZnjjCsTJYxhJnAghNuzXJyOOEk
1JpRDszfk6hCWsPzHMb+2yu6kP3Ua2UcicFioyGwJlekzOBFmtYAxnFHFW5k96b7
LgttQdlFGvcPw7nVA5v+HMhd49dXkFxJUPlA3m6SJCWDMss1aj6ZVMqJtJV7PhSk
BLqzJuCqAcKLhT6m2zI+cHNkdl7RVCWHDOPWsv6WAJmwgCvwhN/15okpSNdwfZPX
2CF5Rxx3sByG21foMQb4b2ZyoWPLFsx0jUw6L2hhmbjSgdHOwIUJwcH0TO3+Rbch
tb6D3WhsCIlQk7IIXd/c0104mIoMMk05h7YDftcue33PFwUCec27HH1rS0WvccIe
tNOmK9sIFrQ2F95DrLIFMb01UN4gSshtySWvAlr0LZC027MUP2pQFis7zfRqC5wP
TIgqL6kYPKPrcIYVw7zAUKciGjw20BijToGeist3EH5hN1PwAjPo1esNFV95rK4E
Una+p6GZGSiLmaJZ396iUCoJXcLOKDplobtGykrEqSvnkP6oyO8uIy+2sxjpLQ8W
r28KTmvy08RIFJ+EWYFDa1AaCTpx4VEhEOBYD/ClV58kmaJ6cEr2Q49wMdlHgCqV
SFcpT+uB9q15Dm2jgooV8Cy77doAYwnndLutjkmoEO4MGhkm6GUkO9w3FtsaCX3k
n4UO/1gvkT2pVuMB33kbNCqZU8WsvI09mStMQPpLMAjUffoqPPZkKO2lThaJCKhG
hEZCy+T86HohXqoPwmUUmHcm2uWNsIBKhIX9vyEqZBhQ+Dpi7XU0UypcgzvtZYJE
MNxzdi/tFf2r0I2jTR2xrIf4hLWA0ofxICxzV+3Gu7qBkns9lmXupRLczQ/jAxP1
AOF+p5zxT/xwtWhlIW4sKHvXrY5CpdCGA3Um3p/Y/KfGKVFMEODsHodQdGc1jJJ6
88A62ndSMbEQZZ9GWtFQeXXT2BdUXMHAp9dpp7cA7tv3gvOEBuBwPe2uWYpPmmCK
wprbNIh3UtIpO0pvEZfP9vqnjNHOIyabXie3z2OrB0LUcWH26GZV278+dR//1Jox
s/S+3kVoZo8pzKeRmC84B2M0Rw7wThdAqXweVPy/NZJ1FEy1Rh+lL6ke5Cyi0Yuu
j6zN9er4HmhfLNnS85xWwJ56QesI+Y+/MapMZ6+t94kuABay2N3QYXwXVZQlmLI9
T1itsBwqMqWLwquQqCvIl3fW9+9BmEYMZO4B1DtGJ/ngPKZuCTpzCkjeEyZnoHDh
PSWvNEowDeXtkCk/RrJfYUHPv5WhboKMVbDrK1nnkBTkMeiX9zBJJ4C7XhVhdxed
m6+RPM2xQry0l65+Lx1WMwG/kiLYCtPF+WlKoB5X6q05DWiTBHJ+5L1DA8P39YKv
REAnErTfszQ5wHqPknyTJp0oEHgIZyKks08cQjQ0Q3LK95t9HWlSo2fKgaKEyWi7
qP2oN6mRc9lTmnynMJsC1VEu0RsukuKlHWd4KjgxI5xyz/eibY0vq5C6XBpR4Jmx
k6H/r+xDCmL8Oj71cXyhllkJmmutYqdX6LadnNJIms8STFy9uer8T8ErssA48eN5
vuVyqMAULNbVFOFL52HZWiGstQwDh1rrWgVjXB7MF5Km1qtGRmGkpo9CY/Ccf6Ki
Pk++khKJ82fe1cYvmChF7O4BZ9U1+9g5PJRgfYoLV7zYByj+J5mu22QZTTHiHm6M
MAEE83cBFyX28d5kCPVyJ717DDM0TcDkkSEnEKc0W4WbLlrAfAPaYB9M+GKJtetd
n1YP2JLjG0/86q8ziO555RViHSq8o7+KxqKPHufFB5Pwb3YlPrUFRoZkcVwmBgzB
RHghuYlMk8KYoHVpS+F4tOIiFyQk9psE8Gn+xGkcUbHK1357RJOXtBGfLB5Ky25L
SCvFpQZNYstLrg8L0DEoO4i811ecP6/L12q8AJjFvUXyHndjg/8YWAvdVkkpB4/H
1O6JXnQEOiWbdP/pOk7NXZxUHGIYTrtHKF0cOEVaWq2mtQC4MeKtHLltQiOhzztN
R07bLzcOz5ffebAFk63R5E36jvC2Pmt8HTkrcMjPXBxrYprIoRrt6MyQetfop7AH
QeT4F0ofQKEtHo3b9Fp/YjAIqU6fl+CcW0exTNr64U8HG9obGSNvvqGZaCJSNTKk
6Fjmaz6bua5L+TH2ZRMXfqeoFP3vfkLfxXPHaWyfJ0tSs1cv2UO1k4AzY/Id9V0K
ILUg1UGoOO+qdq0W3bS0Ur1jOurU/ZjsBUOCh5JieE2OgIg7BAxa5SJZ2FVi+lLl
VD9s62LRxPHmsFJ3hBizZQvZbbv05wLE4D+/C24EnjRRQs6HqX91pmsD6nBB+i8Y
hpvhuijjZbKEFOlUhrGdXlMHtMj1j3aiMwgd3P2Ils7yy1gq/b+O2CFiLxjjQc0g
s7euEAGuw5/TbBkhVKjQ5+yCSp28UheAk0E4NSLoNurqpP7L0nW5JoB0WGlLicfV
TlFBG7AQdyI+2CZYEEEWBeYAhWEvQe61iTt8oz01hKpg94wj2At2PqhrNZXF5d5G
eTRNM7cvt62+w6A9n1DAi6QSSiYQC4s/wK6cnSdjrmn3lD2zVvQdwY/xB34rszwL
sabd8/rPbMGei0wtPXdRnD0HCtDYO8m/jXEGjTRyhZg6mXNIZ6Rs0wk7pdLvxJyS
t0g+/cvztBnjHeH/f6G3I7z8tjH2oZfQxeqTua7vm6fDwXlSXcU5kYjslllIbSrl
Gt3i+RGaNnF32l2bJdg7AcapbklUja/vrd9EDXOYEqFLvKxTy0AU0HyC35aKgYM/
IKX2LpHlRvzyE+1qU6ZUXHp3XNqKqcha1n2ajeM6AQR+MrU5EjNI1i+jSSuLyUPW
TalXRLtyKQBn0WjIb8gnhihwk53s7qmkuuZQahnbHT4sHvuW36AFxAIvEIlbu3q3
rpx1H+f1uq6uuaa1CgroTTht9B1FR+N1IlP8xVjKfzS2n8FCAoTtob0z8WKa+m5Y
bC8duswvPpuQycGtyljwF/uWRGPIBrGKS0y6SCOTg+0+W+eUAlYyU+gc+/Uz6hb1
ZvGrMEoBOcLYxMgdY59TLphKs2QEoo48GzKbFj9J2qww2EwfTlwS/qtBdinsf0Vn
xpRMPY2paOxe5UCheqBsdA0b5owuWvltfgKhQx1DytbwSBLumiprTsshGoAbSuaq
IZvPNy9wyr3bTECwJ+tFiFPYPLiv9nGsDOhmQwvlMAVhYypy+vhQuVq4qCX6J4KV
QodYmkvUPQcsAmt8ufGMCvSq9PST9x5SEyf6x/RF0Kcdf3eWBMtivUzeTRQUse6N
4Rj5gUmV7SmKlyyjw8JOSsUKOs/pipezDRzy8cjXsUVU1tnmQDHuY4UqkasrATMN
kVfuK8w0kUYY8ioAbpF8YTHuz9HZGOACe+V/cYvBZ93uwPCRHZCnhpicl+fzqzTX
hEtYjHk7OnDsumNvp5TZZy2EHYHNbDCPSs1kCuSWJPiN2KGZeroWRr/PVj5+PVW3
iTury0pY9xnieeMngtUyYMkQUOefnUWYZzs1IyEaYkFVMCPK4EfinvAld7TaEJvU
3uX5HDBgf6NwQ7VDdMj23ITB0lm6+PmWIxL4fkH+r/keKldOJG1FODgQcrWBMek0
Uh/WKt9RqZ4b63kcRIQ2nh/zyhDMHnq5AJNe0CzJ+ZtgP9U+s9zbTLOpZHrqeyeT
JaNCDp4HIohabAJXyEnAU4OZt6QcSkifz64rU8zz6k63s7XCa6R9Twwg/ko4ZQfA
16lEqfW+cCZkcMpwjBj/Ixkbss0IdxOjvV67bqDh51Z0Fqifp5qmw0NioDkCmXox
LD/fn8Y/QhEje8OrpKtZMQM4cB88+pHwZ8w8F6q2C9OlLjQOdTM9OgKi+taF3tjG
Tnc5SXF7LVvdk+SltqJ4QAdbI5zfWh7lWWsn0bceOs3jvAxUo3rdZr3rzgT75z/C
xIH7C5A8jO4A9aR4AuROaz4Q+CNP/2kvg38pItrRhpZx1b2TAUOIpQ/yIdd+Mw/E
5MgpfEAlgucyL20mlY66qdUXsGXNpYvpHENopj9p5ffBImzNLI4G8wMlWZ0dBV5f
4RNh7rIvWpzbAng+t3t7pvt+ShbJk019ZNqr+iYt4iSsKjDgBww2DFMdSm0EFTaG
BImr2VIPXMa4Xao8BcopbvLjY1SE4wkqmKdv/V9xpMaMUNcofTYeNInIgtrNK/dK
OduAVyWRD37j/1X3P0T47lRj1zhPeF1FtSJxHibdIpOcM4bTbzqDzO5XGAPzM68A
JxJSyRx2p79Gxq8cwjXLthqJKlUsC5CqR1MhXWmByLtWq4yGIDpaGNjH6Fc4MDTw
uly4wF1iOVqII6KpHu2sDzeEhoTWqP2cYmY1F1vYLcyAtq/A5qRMUveqde9p6AnP
U5bVzUukFAfPTRMXVUmLH34wgRfEM8VVUIXKw7VFcLuoaUS0OjqVp8oOnWQhDkFO
aY+tFKNam8eioCFfp6tJsVpmB9KVUPwNSsuDWB9aAgK9G8Qg9iU2LV0pvx51KGwS
NKUAOzw8M5NpTKqAStYYGQa29BSVBtGlA346JHYwOaiL6hjQg9G5hQgqwPKkORF4
VoCEqspPAI+zL6J93R9Os5g/vDDubGUsHg69JnCKnFNuICkLQzikrsmU1scDeqJj
8NeE+SkWgfncIQ0GMUQk1OwoR2XvhV0uTX6nSnFjJ7A51QBt8ylX/6Z52AdGz0eU
Pzjqu4uTEUmQEsE8imT9nEgHEuUV9WbP92w1GNJ+FGKMZRq27JOnwCchObs+JuSh
4IOuidE6Wj4zzeVTWZ+iOB0QEhWhAxa1eoHE/SE6ZCT4yMbPJGBsYNLZzRpczKRV
2JImFg81ZGjsrbUnphS5x489JGGm8FlcSKDVeaARkVWUoe+FOe8tc++/d709T2jQ
LlLbUrWo16yotHjP4X2aPw5rf2OO3TpkACmKWj6Q2tkwdD5mUU3P2K0KKPB8w6aY
0yQ/r7rzm7DTZOq7CkvimBVcCEAjcP2fPDMcMHYEDAvwmPzZwpNl0i640gJixNQK
26iaxQOn0FrBinPWj/rMbSvxY2WKTJMjHSnnQcism8pzm2yv/16DvzAQI3dY6OhL
heyN/Ml+eptctVTMP1GGw0wsOqCaiz4YSRhbSWB4LOhsL7gAsgRdGXY+CZsF1djI
josxurbNeqd0Io0TZdIUqzIJRVFf7Yahm3btPwBUUYSrJrfdhJitVbKld/27pXZD
zfTbQEEKzk1zHejKlV29TzINutDWwl7XbUVdI6laW80l6Ni5C0cg7jRHTZZaAPqz
WUGMT1U+SYl0mQtFwNkoR/LOdxMCoWknf6Tu1c2kR3NFlQWHy3/GEwBDaSgFsm84
ZtYNSo8E+IifkNFey+hdzHzlk9Xvrx5wEwNQEnfN+Nv6wKVx4w+gvFmWSldebJL/
ublHdw1OTSxAsbFxMoWcHWs2gm9bNbelsJpKuWKdZosv3tZw6zILAzKuVRjeAeMo
C5HiLeY3nxBgS9eVBwmt0p8N9EXp9RUxMlMAgWwJxOLsNiWIo9ViyWXE/gXv8SzC
PixyEma2wpBYaT815yMW28mOuoOr4GDG/jQ6S1mpvxw2J09BvJ2+PLsIZSnMZOJM
sOtv0g9FgRJureHiFKni4BDJJAK4m7sNIVnbOP8nHA+7g40Cvdty83Tleo6OchBI
pu5lKDkdtAIRJbv+grYLh+ixKeqO69rA1UkxQR+9Ou6Cll2ceMUb/VoVHS2POYix
/kjeLrz23/aA9OLczBy2TXU/Kra0bFwDfwM1WxJn8CTKuYI9gFCLYjHS4Fvlmyd9
ptf0hJDXoWm7wxQZX0Jqe8orCl4VhTpGpMxPWcUgPjmXfH543TAfbGVW/eXAAvxA
x3D2eNvEAxsN8uO5H5iCmrvI49djXSUiqcANKNHvvPY312/Bs0kijaUFSZXhLzQI
1yAk+SJiNoU/U6hHeISn1gO0iz+eeag5rY0QAvg8m31wMFg2Z0N0g2OiH+3eeKUw
tFHQSgNJratmVK+3DWS1mVArciLiEeJxtCM9vdCPf5rejkZyg0v/vBCmlCgDj3VX
V462Xaws+bnf4bejfXoLw3p8evfJrdBnMeRr2NuVCHYU3mzKj3jX3AcdrSMhrcjW
I+PilK6luD1SnFsKt1a3X+32Qi1rp+j8wU37XAEjY4BP3F77RlFTPtAQFi+JHhP5
qzQzIk9xd39Sry1Sic8d/GOyLRg6E9vZvSqa52mH+IQIFC8PUCooEGXPLFLQfGQq
qLQjvLc9Ew8VQSnHRWTp34WjGPGU6occHBbj1+ZKU8ckd+mJ2yDRItvKE0zPMaL5
NLdlOph/BoB7EgSItBeVhLdmp3RRU10w5YCWc/lYdMJh9WHWNMadF9L3GzjOqdfP
qpnuKN6K9DttmlRvhvrT66OgPxRc+R4zVSHb57cSqBPQaDn/M56IbEWOVLOiJAtR
X7nTMXW4VrPVxu04Mm/rgpj9wAYxbFHU8sm+mWj3dci6clDWMZyGBa+4IZO6IEGX
CjsAl+gGcddR+22uI8XDP80sRBhOseBw0UjVaBuAbEsI2XC7awLJfbua4otyOq+B
4s/8NonVfN8oncr3AzZhVV5Frb6UuspehEvUbP03zMMGNua84ar1Q7ykU11kGZ53
M8OObMzCUagyy+7VYkqOwIxRpRB+GQK/qN6zbBiy6kkq9i3RMaCI9Ay91YBOFTQN
PTbhyD04imdPJY8IIDoDJs2KLiYTosGJyHrcXVe5ReRJao9ufqaFosrZ58pngoQA
TlgESm+Uq5P0cy1gxc/gE/MIEI2BgLpWpBTEaDtNk9ylef1S/Gl753dnCGeEXDwK
PNjSVXWRB1BtmwrKxJiNdz3cqxWEugR7SGV/aQwVZjqpxwsAFfjbv0swVep2jMvO
btpYGdaowgjn1M1UXL9srjrzdnhavvKNSHBckZRIzF6mYYIW256+xJhi43lMKy1a
PayoffS5cmXOP8wtEzkTjM6YYT7eMnkp+H7vnew28xXWzWG6ORIbrLA1dpfxHdOi
yJLqt/6CvHz7PRuZEbswEQYsQgATghGwc3Yx75rAPwe5uCW0TDKDwOtYVpFUucXy
K/4JBKBL3DJGrfP73x6KFo8SQG1Vq1fmbmSlaBAV9OpMix/+RB8XGKqbIlXh/2d5
o9uT46L4h2gfO3lV2EURj7hY5zWpoya1O0xe8XPxQxeKIuluA2nOBqRF2Ds6qy01
p40K9zTwAmN5p8vUrv0Rg6DLySlxxCmZasgaI2GC5cYfQDJNfP1tBaE0k+fB5Bw9
1+qnVcN5kMx4ph64hLOmeBnEt7dh3xuq4SdJBpQ1y3KqaaD6a9T3oX42021jTwK1
n+Jy0S7zDN/qeZu6xGCmm6S453Glhld9R+At5/FtKU3fAyLQC+f9PxVvnIjsg483
Yi+SxM9TDL/BC5HusDXCL1AoQHV+kt4pd8rY3h9ivHzHrziIeQR5UNilOxpyOeyq
1ZeeQVVcuwrbCJYVr1fRtqxjkCnDqVLfUrJd3bl6NqEzw5zjXx7PQb/RishMXOCc
FX+/g184gcpKKrUEtbRm+F0johmgiPX165eRZbv9foJJC1ZRzWDlEh9v6PJ8dCKC
PSJ0j7O4oN9n+49z21mBDOJrO6OB4M6zmpxVn/7zlA6Kn8DnOeSICO8rQIwgd8GA
4UrlExx0pkC6q98IfS6mQXDe+ZqQirsQGEb6qgfOHpgbmlvKm4MrHrHgAj8q1aYC
xfUJ/lptiBJxbf4Gb2dA6iJ1GJNhOcTzZZxTB0Smwa+1S0/eGmx50kwsSU49qMCF
h1m5u263UZiTNoRvDpmPrO/klkQcTO+8MVx6RkdJuUmYZSITqEpYmd1a5flSQzWf
PVQgLing9LaBMgx9BrLCHx4fzpW2o5FKTYEAfB3e9kN4P7N6bOQj/wD6VWQN7xe5
fcyXb1Yt9JtyGiV+vItK558dh1nx5amxF3CTaR0me9hDnZ0mPExT/0C7rhkz3gJ7
5XBV9Rrz26ZSaXSFf9U3KzZ8wl3r/0+1KdhCGILrudeyC50nSnd6dc/hhlXLHHgW
Kdtr8uUcLGbRN1xDPjIeVUy8+EJkYnik9CNxaq02cSeQU2BCnhWTtHYbeiUMmrPU
eGsfPk+QythGZyOEoECA4fkD2DOy6AuiQ58HuDaKjwNB+hA06wHEbXUwShWhemtL
fDLjHYU1ZROxaaK2/EgaHv9MKBR+Yb3QM4+4YWC9P8FD3kLEeZswhhitb4m/ONTs
vaGui9Nddg5jbzX58d2/h00faDbHRcbjYgNh7/8MFHgZy/Ucn/AUqdcYaHyzM37v
dc2FLsTyobKhslmkNq06KOfJyEY4BHeOq5B31Tv3efUXzB8opcbDYa8aqr7TUFFT
/VV1kJOA70rF9eNhckHCK2+g/b6uAedoICyaRmjK+Uz2hFSjyUiZNRXdPmUbeo1T
2qdy+RhayBZOztUBmgBMNtmnF1u1wrp4SFcUw3vDCmilbxMR4lrVEHovYAi59Mxr
bmobpQQwFGEtl8LsSKWWXFCQ8Dx4lxdDc/WQ2q2ifnvx2wQhV96mEW8u/FXFN0pW
IgevIMCLuv2ZuIpjEstjCtWpVtXgD2Lxn9o3iZ897b2CpY4j9Rylk7utANNU4hTu
tXCntIJALvV5+LmfwJDKhGUxxHkFoZTBWAmxitaIjFQAPO+5J+7iGRCRjLTz7Vua
XfdWSdFRMP287H4ThzyuqXhU6mmEyEt+r5uUSbdYqvqLu0VK8RkGn+6LiePdMWzw
a1JgMvgYsYWZSKCalbJfmH1htk/raV35Vh/NtWW2yCIbPaRLAHZPFbA9dbL8uFUd
pHEoYGIdHUjpGIjAU1U9/exgiRXUfSRXMUQZsBhMF5FUmxPzXtHfrS8zypn8WbS0
WxB5urysaeKa7kvcxs7rNLqC/lD/NkUzW0+gKwPQi3+QAm3lH1y1eYatUpI7n78C
MHcwUvQhKRZoUXgL37FHu31K7SRZ8Y2rv6UpP3qSf/WzNGw25U4CG4tFvT6+UQdx
HXOMBH1LOZ1E2P7Azirick8XCZZy3nyo3y8sfY+ufXAOpsYvdEA5tJucGRVrQHcN
pugwsk5VtqsllfBrTtPnyzMEvmf2p/w3eDOdYRTsUZptKHg0pav+srVCbRkO0wZy
eb11AuNH9ecNz5RNXYZpuw9ZkCnS+wvxHkjc5kpCmwZyASqx6+Q0JZig9aya8TZk
81sDjfBuTg0WUkMLRpGo1cTz4372pqsW1MjUQoS9vRv40NDPY6aqY8+Ftn6dSlXb
CCCOHA4dQbcDiETDRgDY7qCMrqDrrn1whu1PzMAO0R7jjByWPlyleleDYApiUJ3W
T1+um5BbECZMUGQfubbIDshRjnJIeIvma52Rk2egqMz8NZUic0ENwGDNLzMe0afi
AMRDDTBDkn8Rgi+a9tTfinvQEyV0xEG1keAVkxzoqNcpSZ4CuVbR75QTaZp5t5mE
QDcoMM/JSXDvtHMJKvSrERa7ZAhnBNMmZviaLGPxAOUEGPlexZbvMMTuHiohryAx
r9vNorvIZZrukxR0iH7Gq0LvIUAy5C/AgbKyrt26aR8YdMTkAVCVcw1vWpgpCLpF
LOW591Wfy8hu6LV+LNt8SBk+hWcrkDNv5gcqI9Y+1FadOsprCw0elUQF4GNLpnc0
H5j5j/ORYuxfNDHwWBejECLYU9gPo2u6zzGBY0W+FRjNrr61gC1Zvq/YuhzSNbcu
YxVUPTjkozuZ8bACehKBXkWnbQ7Zhd6ag81pOyW14bsh68zh3k9XM27pc3r64Rdv
twkzU/KpNZoFcQtZLNW3PQtMibXRS83hp00uVAH2tKxIN+Fwk6rqAZOGgwTzQ5U2
7DfXTy/vpI1cQgoUFcYSSEr7HirBZpkRuuev+AWywF9n3VGAW84T/jtgaPKA0O/c
CxXx9e33TVkdPj560gcl7dKs+zwZfjLHLv1J/JBieCfgLgAQlMwY4FwWMAg+uVaX
dz0OWF7/VLbBhLjsUVBvIp9n2QoBWHUvQOMK0ZxN2JLHgtbp74J5m0ITWkjggrph
Wpq4Yuq1fRhQIXsAn3n9t7/RzsNGTZ5ug5XU3uYPCk7nnehkazmj6HDPPPVIycbg
kDrrFStk+Nnf5bGRGvV8X9QL+MlfNuZNCxIQLZckiTnUSnenoaO7q9ViO5ABdl7u
xYJoGDjHzsFCa+a3jTs6YCEKq0IsG3v9PKH07Z5pdT6cqXV8N2Wuzp+fRdoBmpEJ
X4MkF1TN+dK0JiNpvSSYsA2UIU4Y4OBS7shKnzBQyA2Hw+O7IAFm7axmx/HFyWt5
EI9/QhUDq7YagEWtVz277w3L0l9a2ahiy0IbrYcc7djvxnBnOrYZ0vWzeiu9FOSt
op4cTeAe6uNiOBHtlpMjAAxzSPJGhGtatkitN16qRLli3Y/WjnbcnnmR03EGL5Uw
GriLWBb9yAtG6cVOGr4JoBTWYJjdtm1QIHvwhHVKDEElo9qwfnrxWubo+CAbX0IK
58XkaMZsy4fAoiLS+1yGyFliErfX6SRmGqOOhegKckyBqJLoKVLRQaUcwmQGDf2+
0WYtYHQ7oDanBogh2SFWFnlLP9FFXSrt0yYuvrxhBs7YO0SQY1QtO/kzikM+4InO
S5Pnr+CCBEqXPnNqPWLCbY5fKNhLPvSf2opqdgrW/DAaOwJ/rRfJ1QquAs4JJJKj
8bSAfklTX9m3MbIpM1l/lRzZcf6b58yZxWT+YkBTmWU3UY3fViJs0k3fd+I/XFF1
gCRmdIRkp+565lNpyYMcIo9WYzK/KqSRLgw5ligOrrPrBqGF/7Ib46K7VrgB28xU
t6Ex0Rn7odIq7qqLZn1fqHFyx5eEDuskB/3xij38EumCRj2RUc3TSCKCyNxJvMUg
Sk7oUxbJXHrOPfGjw6QAIoqE2ZUc9WtNccyRHqKHW126+2d80Dj4Toqvryqt5Bxu
4/lWi073x/UX0zSWq+aRGe9TQ2wD/vXerD4pvaObmQu6qpRBT+slaE5exA4PZdTZ
oC6UEaL0XAIvcEe1V7kjtkYs6D1aWeuJnWep1r4DVwymDmcba/ykTDXrCwvZbhtV
fdZ3/Dt4VVW3nupoZEi/fhBOb24rnngmlmLP8eGDUjQNwTWpvRWJ7GLL8DivmznL
BhWLfQqVPYlbjEuSjPlCEMhCNwWX+Vbo4jtXFr8bzCx1K6n+175Ds4V6/jN+6eW8
EADJ3ZJRVJDuw88g4J+V0S53TgzvlpeTnwcMCtRpn0k1QF3OH8Ta2V/wU3UH2F2g
9oTe6ue7kaRhwSdi4VYX5aJRJKoieD1al0BV/wmfltYRa6XeHuTc4OF3FkJwB7mC
ea4fYrsXFGciSs7KHbP+0J7/LVT5ABFWKBYwXs1jrYZ/pd4ZuJMxd6OZO7Ik8TCZ
0F0gE9A/q3JhT9ekdO1ooXXLc1cFxmF3ulggrzCgS+rE8N+u9T8TdvA/ArvulS2K
5OmwB/eBQEDw4B1A8K1mdHv/PVu4VVjdHurkgAQPmJ+amk7RaBWikObnrG+itMAc
L26h7J3Q9qJPp4KWS7uj8lo589ZKmuxk0YwC7q8oTdJ+uxzTTFhxgEhauVUfJ18g
ox6HbHkmF54nPW4xef/W6mM1CEnbiP1VGAI9vZVS3poROSEIypu6B2eTT1i9FS0X
lFcHmiXrJfiruqSrDitgtePedSYKJevce7ww9upVj5aQ6ubLsnshjIZdCTXiHjB+
L7TY0nM8qElNwxFzQVu8rxYYMHRXjcZqsGEL1roWIWlqU78RoPviiEuHaafUBuFe
9VLeQ2dIxb9gaELKO/MsrmHPjEWRXnMUbp0A5wPOOI32P6ohRtKRZISGu1rBHv/w
puxwfDL8rqQKseKjNbyM5mFXY00+AugXhhAdcWYEkP2Ba3OpbrGI9/iciBV8LL0N
yfHqxCqMhCJgYI/j6jvm5ETR+Jon5k9qkTYM186Fs8Rfanmr4ohWkuAYAnSLgg3o
78fP7cM3s5nPkz6UA/zJoooectqnJTvhH+JNH3QMfi58gQ8X+PTnkFQQsIXaRXjx
SzHjqFAVlM+8wrpglCkE9ntBkXvUZliR0ukdGD9qMulrFysodImjfu8m40GsNQUF
/09P8iHXX7Bj4ewF2duFvToPWJoqeAvSQynC55dClr+yMCIoMvGY8OizB9mkBc+t
EY2wUJg79TyZgHtCLqR/ZgpNujos7qTI+FANhkvRiIdQ+resw1LuI5BYp09XNqce
PzmXilY26OmfWxdRwCAxBNNcxu5/xoklgdIRVSkoeGmweFr/yEIqXQ1XpQJC6mcR
bZwdqmyfbC9/AJjk1IALMwqhws1MidAIDQz2lbyL7hHoNmaHp6jzcP4bqsuci73/
VlHkLsVrblvmb36jwuvsP65YqbE4/S453Z/d3aJ8WZ7zcTcHKar0y8ziSIjkNqc3
HO3n+VtIxeoUUQXK0TyrYsUF/TBYi+2dkco36AiYJGU8QInVE32kwCo0r7B9K9v+
+4pFhOTZYNe2rIq7idwxWYkgV4qzzqHgSOygO9Z4b6/op4K3yn1Q2wyVnNrqjWbV
FTqJTApBm8yjLoerQN3WDNNpUf/TXQP9nx7UGF1E6T3wszFxM5lVRiYEAPSdW0A3
f9xweqma0wfr+2jmbtecPPbtC7ZP2batO1yT3rT8/IMCAIB7ggk4jDGLfaidbZ3r
t6FFbKiljZYbza0YWlfjYPiyZzjgP5XHvhHWLbR9BzSz0TD4eUCSNZvFbUy8/Kux
NrCTMyIh959b0l1lajMZvo1bvaya86GpvSMoErtLm5w6Z7EoOZlpu9TZ9jHTxrRb
dXMoK9xFBhQ2ZduwMzJ36Zim+jrKTuumc0HmFiNTskXGfbmQ0dn1yW6V1Tz180VZ
1JcgaB2cuhRcKlISYOfSkODbfwAwPNao5mrCrE0pjkmCCqPkR3D5IgAtV7p6k/l9
h5PS80yinuRy2FX3NymJLcnKwjZO/ApZXTj2+o85YNeiR6Q/FUl7PH/AWmYiBUX1
0cCg0Sa0HxZwnmMOtkAdtspSs6ao7sneBhXSLvBF2edYMZC7B02mNr6GIo/KmL1i
WYNQ9giGXp03pQ+YFWS2g+OHTkCLXFc1PYbxVRSzn7m99arMNsD+8+8qIiQqP4xL
98sPm8WTCcUtRMNN4qjfvft0UJssBLcjhbRVNIP2kCBmX3KdVsA+EpAkJ/N+6/8B
xV87apzRtDJyOmHOnJh/kj57yOQ+N1XOcx740IEctkzrlro3K7grPoV5W0m7Rcvb
1bhFIjHONbqA0dIUgcz7VKhtVrX1GIpYMdXMkacwTfSfGg81KFF8Wu3vptQxcbVG
53Hej2JTh3dWXeCwtSCovZARzI1RWlq3Wv72E0WQqN6PCXNtP8KR1/h8v6trPaAk
ksnUz8k5GWTsPUhLVStnSFNHgWMPpUC8kyQYQ6ABALBEsz8Qr0RmVuOaFCsLOb4z
HAieuFszDAAXqRZ/SaQctreEw+BzEOwPng8LFvyHAc1315Wu6IDZ9693GfRNbbXE
VUUPZ5Jqcl6JlnlxhsFHnHrSHHxpksBFenzeG8udJw56AN3n+zBHVzl8DJVD9uE7
XuYeOHOCtL38ULOuIvVVAa+oBDmZsPcPY3+igwsfyHmELpnH8xUk/eOeLsUYXMRL
3hhLRRt0m1spvBIz6lZHS4fGwOvjXuyUAmTslqJ+T7unL1UNHIRXChtNjoAWbADH
tbjOVXtnfbNGdq47tNQ/+aMHOAR9xUAXXqUfhGRMDhkCLU1aZU2AX8t+FGbxfd8G
/t6NBPONEVIdFHqixKBpUxwVZj1LgmdD8Qe0FyZXh18i0KsQ2o9UUCT6MYsiO5kB
sz2crKeByPFcpRDyZak3IK8anFf4LytaCJsX35Oe5SOnfzOyscDo4DsjuTQYsFF7
tarY0LguHun08T1Fe0raoFyi5aNbCh+BmW3QZZxfuAqGksm3kxffOVf3ZS4E//lg
jYSshxM1taruccoT+Dr9etIJgcSJJSrKbWidAJ/ni/ycB4a1mejhlioAWLdQOz8U
yWkianHKF6hAQDk/JQAyNwGno1pXh5AwrdwTWJbh24b+09gZvo7z3Bv5M1Y9mt3l
7HKhto7pS5XF+XYanAXnTFw7m12hr53TtuRkW2b0D9PT8zOg6VR0jO3xmWWhzFxE
0PJlMOYYzvnhenEXkmPnHRRiNYUXsjG3Gdh0vAHAxIwowMP2qQqStA6snJMwa/Ab
GRb87jgk6ViOjFYx/BjrnI/u0V22dF8keuz5CIMA/v9gjcZD81AfmKYlhiSWIJSC
u6fHaVKSbIt2sF+HLpvSWek0E7E1lieyVKnIYPo3Wm4gb3RF6rnCvsz7qUPt6V3W
S4mBsMSSjEms0efuhQz+oBGKexK3IUsCqZBmxwuNlprIsJRFQVmkLfaqQ7BnHkF8
7RhajvNJrrf8B4eyaLSZ68K2zySF1utPzpOErb85I06xK+Izrn/p1pObDY40Oe9U
kdCpvAW7G9ocYlt8u4fgzY6OayfRHfnfIesduh4yQ7WgBCWu44Gyyw0VUVhID9UM
BFqQtW43ggxcaYdmfq6uIlI5hrRBlRLNCltm+v9nsvFKZyj8P17qGGeWiGE/r26f
gjtcIO1RuET52fGYhSC+pJmLQev7N3PK2F4wUNPb22rhVXcLznDo4AvZRL06ewzM
u6PhcZy23DMwhgVl9JK7vE2/PnOiumePvpsihbO+r8vcDe4jm3XIYKscl+hUclCe
DG+Bu8WoPLUhkorsHPlm7mbJhHag+02DKq6rQkYzAx4gAsFhnZi86RNT3rRfzV9t
9ufdQdPVHbqMMWJ5Kw0iy2iTuO8KWIU9PyFFEy0/Ghy7Mz7MWEz32aGSPpy7G3/S
z6ZCOQK84032PZCES6vYvfTwPlUkUeIEV5n3z+H3d9cN04Zzf53NymCtE30gF2Y1
19agTFyj2iYtj+JEEHTgAA+p3cW4JmKELPnpoEhoCz9OtEDOq4qNv4t7FY4xWRIe
1We896sAsx8ImDiObMPhnlHmQzot59NTYQExOx0YSvrEyQkZpXdu88lnPHZNPjZ9
wzedmLKrMS+yPJy1R903swN2W68N65vRf6Cy+NghiUG9NA/bF+k4Nd52LkQGUne+
wx/wJBMh/Js3UX8NIAsytYOpun15Y4XFg3nnxgVsZWCXnmp9NSoKLmtgo6UArfzQ
u8wn3p4oMmw6451lVObXQJJ4J2iN7EQvColj/O5DCcWtmFLf6v+3BqYX7WVWxhd6
MKYmOmqnya75VZlAmvQr0Rc+fKKPzAl9gLqtAE7+OrE30VEML60MVRxuXYNBCOen
GssCQiowLTbq6/4ZHxAYKnwnpsCaAia1qfBKdsqlVbnbUBbZLnV+3pus3/xBO8fA
PPL5GhCjdJZ9zbiQSZJDCh5FrIg5085odUhjoSzLukYlQgbDQiXY2l6MItDdJRPg
TGrxcmWR93x9DPfT4MFiqfZ/sYsTRBmTOvE4tewGwCSx9EmDHAuFYLnRM3fydd/K
AYFC2O+x0BzJ864iEIEFSanNuldPgjo/28V0C4t1AKwv+yBQ6fLUT/W5uGG7ITz4
//NoZNyqmpLlTmBfnYhLQRCu0uc+Ek9g9uaBLYdfDCJ3PASja/29j0Gm8JPSk45x
9VjgYAjvS77wt+xtGlWhdykfw+X8X8/rJ3DqFmbYejaaQKaYFQCpEm2xG8hsnnj+
a4s2ZMnIP68PTNSjBC1mrvqUTmRiw8PlOeKQXPUkp+0otuqh+GiTzmZsqOuKoGAe
/UPUwt+JbYbBkkOVQaByMOK/2dLIDutfSQfP5fR9W8wpOro6xq5CSPWCYwg6im/S
Cey9EF9V4h9RDoi4wv6JbvEBDmNr5khjxLlqAqKk0JHCG8sNG2/pg+AD8jAiB5Xb
g8PtXYgaWRxIYfwrJ470Sd34DmNiK1tAEn/73XdfMJR2Kh6Iirnokrwg29eJBDVG
R3buuJL4YzfZ0z/mR7nZvY5ZozvDuYbGUz1l2krav9xyy73fd7+cN7p7RuVOpZNz
RgWyS8I4ANXlygyHFF7aAwUqP8bxXdClHhWtp/W0wHXbgkZVFRK3jH8lb59ZsQ4S
U+ngBhYdBOjM+TVTZzceD7X8YBA0l5XofyHNYk0anFT/4GdwLl6x6VsdYvVZ93qB
ayxs67WjbQfBlzb93lrl1stRGp+GaK02HzunlqmTuMxkDUGEP+PVeFWeTgzmoMTR
kLyhh/MNAft8gQoWeBgiztv6u9MHevJOe4r18/ccQLBZXpeSkWC0cjYX8XKKihy0
qM3oGRdXra3Qy1RIKTvSPFgn73kHBWT6Z8LTxKqdkKMNlrYRxqnbg1i7YXzZwmfV
2KEy46uIPm28sxovMk7wvhrcTyPXzaKM0tlGboDO31ieqfZx726OodG5QCv8d3mt
M3tBLfwfZceVYeIsdfiEZVDJ7JQT2eLqTrA2rIgEnWS4quJ1N0/4rqbKchLvH9Kb
C6qsibUmRtOhxhihUkVBz6YxLhYTJr/Rv3na+zOk5yF/Bw6oFIOMawZFFsG1IZZT
E1Jgao15Kc7jlYiqUDy2JpEItIw4jDeRqaJJ4IfUkQVsEhGZCLmPLmsMKvXGtZCk
oFd3jS+u1eiYAB+Q0x4o/va595pbuNhox2v52topS5Vfj6xXCqgUI9ZrjU9EiIBa
qRfH8DaYDF49zPpamAi3nf0GBlALgtVdgLReyVbP+/M6ji4tUWHReMVM8xb4qgpH
1G4bH/4fEP76oC3ZfxN75ujwEmP2gNh15vQGl4sX7jqyQMKTsJ1n7LgxEwuI7KAt
CcYoQ7R11ScT2h+n6/Y2tPNjLhGmA/1x7z/NCYctMrmYd8uAsinvsXNYC7RJCJPH
Ww5h4gCMPqik/Xguz1h+s9zcU0+8Dt7VctyPe5acORXCO1VVvtMwnojZS08OS6+l
zikPVersOGOGszfT+JDzIIvLq1gvx668+h9Eiv3Pew2Dz0bSz2EB96Juu2+bDzqf
QRMq42lUr/RlNuM9jn/uii+je8cETQ0GH0curTPZUTZMY1xlSxN5AM9a3Iof5g+5
dF08kCNis+ByWsOeQVsTjBfScxO83GsjlqSRw6oXOXQfRG7N6rg6dqIeBsh1TZT4
ZeQRYx7WvrM2neWmzYYEVpUWrhn3maiC+R/XY3YvdeRZAlLtO4Y2y7O7f4sL+M7u
MBVIVKZKmTdt4n1mEGGHsGtUiSzWAnlOj4sZg7YPXN16QqP1d7MpN3g9DXozAaSe
Obs6xJU00qlKx+dhDbMmTXjeLzOY+i4+gWuT4zhG3ylpMBdEAq2Yc7eVevJdxjDw
Ju0xq+r27FaQf7OX95IFrsTxKeugOZgBCB60PVKvDKtm4hcfx6Jc0cqQhs+NGfJD
0vcuCcu9TiZQRR9eAoQWcoGkmTjyTJw60pcHorj/beDK8V8pKiVaXykK/HlDPuMM
g7rn99ER3zuEl3WaW7WBoCpCPK2RQ4nT6E5Wp8xSljGb33yxJqKbaw8uK4e/zdC7
YoZy+dHu4O2LdWlFbmYfg6B3hdDAWiyyLJlXyK0lPJ7uTvM97ghNKMDvOzc2fGAa
zFfluDZeslMu65a1OynVFeA/Idx/Q7OpqzB34Glm/x9nxUDejGzJ0PUGE/DS2BL6
zeEzhNXUTCXXtHawpnJ/PXph1MoP1pkHkiU912aEiU4le48xNplkXmEpIv7jAAmv
1eMnUVvRFc5br1oPjPM4mAaTb4kvrKoL9H7blG4QU4LAXzTtGBINsR9d6y/mKOGy
XmNolNshaiCJG78RBZ13nN0OKsCmhf6lnaZuHAkif8KuZF72UVY/6abTFuJXu1Xy
baUWL04gIuO+OJyfL6/jVcrawdF9vZU7/gmOaul0EM/7q5ejoUnT7dktvr60RHpU
XXiZSLdwWutFzO+OCVW0AdGDlVJeSlxIPH7X8ujanPJKjYQNL2K9Sh40/bjgHaUx
5vlZOi/kuKVPh2vmOLc8BRD9Mqpm24OWUsZYZhdyrj8sZRsyFtM2s895yGWRTw0e
qZHxE/DNyvtbYesNVYvdJ8CiWHjTj9Vq4g3tz9lNN+XUgZLClufbikdC8Fhm8rAe
QdukJd/F8oZ8oxMe2249xqsv0bWZthZSt2Z0ZIHvVuQNAIPCP7atR6xc43KxAVg1
N0rjJeYgPLlgz3BC/mbyykvWirppsCdnQm1r1NUs2ojneVJ2JHAKdI92OHKp0BjH
p0qXJ18/RU0lWS7tOdMl4tsIsXi5PGsQ6g0a1lSpHMWxLof360BGf3CLtZzZ6FY2
/42Xv+945n26jI2v0TQNpXgiEmEp02J0zrNoQU4kebX677r5gBVfoEWSdx6qDFc0
sMa0JdWr67zdB2pfqrlr33ZRajf6rZdWNIWZXuHnhJgAejEmwba56rRqTauQDbxg
fcuv6gxG4NUMUnuJEHBvrqlONRgTCfQmt93IdyuqrSi88PtZQ+UZmAShQpWopKvQ
+0POuWtU7kyRMMvICNeBfK9Df4fpBmaWPl+InlnYzKhdVgmmVL0Df9kK26nbL5MD
zUDyTmIHixVIXRmTAEYOkvdhvCxRurlurSov4kk95A39MCEW/4nlPXYr0wT2Hq3L
rxNsB0J98f1r1+8KlP/KgUOL/jvAIVkGBbW4EArnNjf5thDhfXn1H+D24CgWX1rB
21wgR6WAEKJhF4m2q16Ms6mK5mAajp0jpDGBnYEDy2/NP+AgW8tpt7h6rmiURdyx
5irCXajdfIvCrIwTYCLvwRPGhGdR1pLVMjjz8BU8JqOtIFd2LYtsRNC+/ilSDVrV
5biQ2C9Lg2PP6xI+aML++elNvpxU/pAFDFggj03TbONuTd/Nh2eEARm9lTW3lomo
xf7lgT2KBTsavw+WyheMYk36kKsA/+pvXxOTLmnRNZaKiCFWQHHGNpDCM3slxSYc
HAGik3AaFsj8+1Mw8Jnzj89v5tbeiN9ow/7f2sp7J5sprhXtBncudNbj2q1kA+el
KBvP3n1H+dm6klCuzmkjplWR0vI+sssCJyDF1RwZooYghBBoU2u0XyLWg2ZcNM1H
MnITJu0FZBGVWDt7EaysRnJSW+TjnXY/NFWXYweM1QBWIfP+6rYAxIkK9t0RS+Kp
bPKAKVrGKUyay/RPQa0M/t0BzPdlx4KAweLbwbTJAipa+JJRcssexArfhIfsM8cX
LC3dkUm1+u5Cu+YYeE2qqvcoeRLCPayI8aHlOXivDPUaZzYOtIh4B+8+42BWl/1Q
8wlX/aA6GTlRSx2IMrHsX55q/45s0GKIj1NMmJd+YhcqE2Glw9HFiVtFq37iaQ7q
HnZeitUi/QC+h4TAvAbnZXR9IBRFTQBMhuv+HnzyH9UG6W1ORA2ddKBKC76TXBcV
3tjfm+1P5ZrkZOKvz/Y9wbSB0cNpn1G8sD8ndpPVu8AczvUH5LU/s6CMJjRomKQR
2wSvUnlEjWdKgwUeBC/Sun6yyy9G7RP1CbO+iU51n0kD/zNB76SuTN8b6yyyj4r9
DwsG88YpAT9G9D122FTwHmLV80XpR5K1dknd1aTUJYebE8sp0ESPUjPB5Z+dGAVl
45Cf+oZ98rlYX/TwEbZyBdj8apxiU0Ue67TcLOBeGm61/nWi8wk4LE+PlLX6ghoC
a0pIFrbKufLFrBpvFp1oRWZGGjnRjJMPywLek4AxwYB6DbvAcediDrN0MtltpfFF
JCVCjPH8tLzOo6quKgaj3HdFilUFhCPc+vdZghRopEZ4BrszZlYXLylXXg/Pz48X
wrlsUgF/tHyioENYqrE+u+ZXvkU7OKDdRi4IxRLqGahLPKXszxYvwfvruZ3lBnYv
7rURVSgWSAi0orP4zPfUgjL3NajydnUaJgiRcgcKk6GCjW5NS9tX/e0snoxX9msw
I4TnjUoV9W7mM3NmcbwzE2qyxQIfkqeVbr4USzVJA4qTLJFmwTQxklYqZX8aQt+x
yxDNiKZBRbChRO/asZgOmPYzo3cD+9qk9gId7h0XsDEubU0nPNM3ueb3noTVnPBv
d0oY4rWnqh3r3yNvkqxypNM8P3i+tWm0e7C6EEynRnB+xao5+8ChOyuiHbjxiEsL
1qJUXpr4DZDeUP5Y0ghFl+fELoPJeKJ+rLT9mpS3qC6waTuGN3rSuVUs9PxEhFv6
a+NkUOUPlY8Gb+J4sQ1wZsag3ANjn7MZqMZwk173FA1tWvvCVNqZH5mS7fmpvlLH
gI449ZX09efBu43CiCTiADwO0kw6WJx649HMCju9cMnhdSUfLCojDSI0FiRfdm9e
X6cvmD8b6pGWZkFtDutja09AiVlbBc3Jx41pz8yON4L/kxT/S/Our2T5KZFGebp2
0bocK2BB/OJi6aQc+2PqnhpZQcnc28Pe1t8Qjkey2eY9fjnkxIHxeciGDBhOYc7g
A3Oinb3s4LOJuuCSpBsZ51L6FtpKYMstY1+sWDXKlG12d546iw479NUj8tnMRMRL
gKJfP36plvU6s72lMlNBnfTVoEHVQqCXx2lQ4ZXNvMe5BcI6Bj9JuW74IHbkq7tN
/g1GDVBLJijkf5RkuVAMLNtHaqe6rK2cF3niXvMoAcot0mZkLvT9jST/oShoRY3T
YKEqJikqDywWEqRBK2mwB5Sz+ssUai/SZ3P7J6/l0P8Q7TL0+SPyVYhLyAHBxHBX
VImXhmehRHfxtHqOqSN1I2p7q0gQPKryoT3Qgv6cqplptL894qwqjfXR/EypW8XC
T+pHyyoak7aRy8JTrY0Pkt1dRMsWu0rpvPPoB8w8KvNxfp2CwRNmK8riSppDJ5BQ
y9bR3yC7xlZ53dW11v5xH6K8FOUWp5AZh1H6FxPda62V6Q/nsZ11ooiY5ioRfE+h
SFkTh2q7OIozKcE44sj4NnA8I/8pwls5o4aHgsgGUnUeH9XQadvHX39jp2uCRQvy
u4ozjXZO9ebvWWWxIfHjnVp0OEFWXHwoHWLNhxYfw+I+OhrqvdXj737svDKWbDOj
bu41T17t/YHGdV38U8SF7s9Mp1lA979EtlHc0HWNtNXI/ssDuBcmLsgexfxNINfZ
Cl6jUDVy4ezy0xiPgNAjL/DOUo/5epTCKlpPtvU2EuVZaNtqAz/hspTJag84APwE
U6uFevSrRJ1pL1LvZVoSfA1LCurhQEUQWoNh+1h4stTYyVxsQOt4MK7TamKbz4Vn
XfjTc26d5em7pzEaTAm3umLNs/xdF0NE4Qhc3XMdvyPnvGybzZfyyMSJrY22bqeM
y7cd2mzjVxKKxY9uf4yKT+e1spMIWYa+cg/q5mcj9S+fKJTfEu4l8AKBnXpYK4pX
wUcGMi6EsFrXPUVNk2vb5qeRxVxEr7gaJ5kdihosfvnmCAO30Jcs77aqklIYJ4Vb
51Jsw3zht/QzWZYHmfvVfRrTk1Gfz5su2166QvutD1yCEPFPFxQA2iO/quNXbsFS
Hp13wGA24lcU0nuw5mn2LaY92vXtyo+yEIowGXUHFZDLPXARv8ck9XmwPKjJVqXf
M9qJHhtlPjlKXGon4PlACnIIjsQe9oKZTh3QkUbq6Zb6WOQMt9xmlbsz95mKSESh
qaXMYDdIsLWbZmexOV3tKg0X4Ilf7b4ffDNkUvLV5kuJ1MtW1al7M9APIBMmUTFZ
kLBdfLAT765M8/hsqEjJ3TBvbn+y7MINnHqnoccsiiNkSVI0/nK0LAI4YM4MlQdH
WW0qq6NjZ1xKyGPXb1k+vcyadTW6BXrb39Fzpe0oQBZbm+j93K9YCsFVAgoEH4Jl
ljc8pXTZ1DNoRw8fyl7nCNa7G1jySGh3c7XlLTYQ3b85nYOXCDjhuZu06x1nkH3D
oEUEWKRAajnCT4nZ3RULJglwcELIuHkx4Rhs5kFI4UNUzl3JWjwFSDBe3itM3E+V
IUXQRlDa4IkxSb7TgTMDQuzrWt71oAnbomh8BDDewjuT1xBnb738cmxUEO7/8hHF
VZ/RxfW1ng9RxT0KN0i0pW49irRFHi5jWZvT6Y+fA3nJMURJrXhg1OudiB2UhiOR
28YMvOSl3qEmBMs9xN4Kt11RFhN7rFDr4Npy0+GtTsexwmV9W6/0Rx0XnV9BbXjL
QMMgOwGISOxUMhPCwRrtBNshKU6GDSom9AbVSqasrpcVWcco4Zj7fUZZJyfu8Y6P
jtcaw3y00pCuopN0Y5CCM5xSJi0MSeOeWQ4kCPYf3FLN1zXQB1ozEl0IXcEiSpwh
FBXUawvQ51iQd8abeIhNh/32+HnO+wrvUYUsylWFHw5ATAgbn7cImgUJ/p+eZGjl
SXUz9P/V51TSq2J0R2amvb32t4VS4+bTQAgnWvUj5XLq8tqXJ1CPPO6KBPIv4C/a
KZII6szOlV4Z1347ETjSk7b2C8GcK4B9WkQDiCPkiBBuOxtdhC27LVbffYMQExDj
/jN+eKb2zocAkJtxGHr2wDeUWyyeZKakzHFnLffseU+1ZElMKnn6NRC2AO3U/lnu
/tmMGTkE7u0L1jxcXdu0GYw0KWOINUxe0v1XEfZr8iPRDuYHdjGFxXsAaGDk9UiG
xN3Ia7PxzUqBV3cf8tULCmKQ+sgJhHyM3YQ+5Bj0qrgkBjD1q7iMfQeN9ukZjzJ6
uQMVvdkJAShOGhjDEIBrMXQd0BVzHz/ykhX2qKD6rAzyl4kn1L2MkVlnrPG7oMn4
fOrojiHhGjISgDWCD9OMizoZOZqEPkQIIxh2ocQYp7L56CJhg+JcMs1st1f5DKym
PTAcaboIMSS2LKk1YcHr7rXjNgstPJaBBGsTzDFynToOnbo/ULZWEPO/u8BkYZSM
6Q7ItG0dZjTAvx9bcKSPXJFaGeJtBm9oj4pVrBGI8dPZdIXn8+Zmpg2pXW1hQsza
zHE6fK7M0EdnQFaWgGTWNRYW56Hb0Ro9JY3MqUcRuMbMu6MLO7V5asfdUjQJcuJ3
vkXQfkWXUq32alSOCclPLdQ1zH6OVPujriO+viEIDR9MQDiP2mNsUyi1fmtrof3/
kJh1i6trVJZ5gzcne5XnnG9jvPxX3dGpMQhMWK8LA7ESm4wDRsdCbnwlRxTVBs8o
aQeIp21YA3tfMIRGIsPTxqQsc2Tv4N60w8AvGHoPY2STScddRkaNpaaStqA6L+kX
vPAsry1iYbQpvs/YnaUmxwPiTA6AvsH/T5XM+wrXiCM+Z2UQcw4IVxfGZBVvnFHI
SGQl6baS1JNYRYsLphc6nJIF3zLmqsz5F8g14A3JR4Xh8gmftF/oIUxjZGMcmfG7
KgspemNPkmgOtsnS70+yGFs+FmsDPvX6P1ElEjHqZPqLgfyAhK37lnwhdRFbIQed
PsS7Qrw7ael4GHxVdvKvHAwKf2beTzpgSP1sbKWuX84uwqr7XQe0wsUvim8cY6m8
LXBMELFHBCm/p7XHojDKmkS1Gjoa/uSR4oFQt1YmXOjxxyCng3Fws8ryF9QGxzS0
T4Da0kyiTn2IdaAcZUN6uoJwJ4WcS1IIvVcsNnoVT1fP3nJQd1k4T9AU4HAbbjDh
hMHCSdo3MisKWBNvcXf9w1ewB9mXstDQlUNi7h2EjCEB2SvEN3k7jfgSx2J02Zrv
a6DMSsol81gMIm3kf78xcZENqNN9aQbvwJqLBp3k2mKbn69J7z8IiB/Y/CwOhBrz
3g5XtVW4kqs5+zIfEAsKw+B6SsFQpJV2YUO4ascV4B9Qlx+E36D+O22Dqi4/aFlP
frIfaSRhqXsBaXI5V3fSxL/fhL0dO5BxfPe1GdXLfHO7i8eKEUGPO6WpMLR8pWsf
nDHaEyS9uAyaXgdqsQ0MEHjKdtsSNpkeASuRdVAszpT1OVbTnXqEh9WFdkQ59NAG
fcz29h6KGBwo03O/0/h8peAXk3+5xyLRY6gmlsMlptdjfiF2LGucaGEsRThu4PdP
4EbiiK/7FDtYPRBVe9GLrkPbvcfMFhYhA2lXOFchnS6ACLxCdXM5p0Y5aEM1fmuQ
iJHbH1ibWNQ1RdNmWqNYus29j9DYeE2lQa1NlsW9CoIzs5FJX2yxBPKwz5tfAyJS
HZEkluyxh4hDhVF4r73sZB0eJnFuNYPxPPjH+UdS1mCBqQuj1k+ye3uNLuntGyJj
kN4DJSLIOA8qJSjbVrZSXcn+qOZC8cGjy2n4fnui9mP19TBlOUI2+I5XUq5Na1u3
Eo/BB3H00GRYyfQMgJ0ipDdQlxAGzaidwwJmNMEYNU6wdGJ1gvsBGc9Q6ZdpmllG
b8HfdxMjFRwoh+oGfe3CS7KhT5kii0VPNvWqw1+Z/sdP/upYF6E9bnZIePHycyyc
0EN1GWE/Rlp7vjsx6GDHc6J5wnSGAic1ypXrnmnwVI1vNykD2e3WCwb8zeQq6GuG
53FchHpsNrqOrwQZObTA3q9bIt6R62c6g2MEsK3mdAmlM2rVBHjEo+mirGt+DQ6D
Dm2SjSGq7n5H2+QgKX0TjKuirLAlAj7AprROwUQcMlVFJThUezISIL9+rfh1JOFo
RWMhw+a48fdYITyY2T6UrD81PGdB2eDIx5siZAdTIxUWEzd6O4u63uNuvBKkQNSe
3rLlR7fl3KBvtIDEHaxSGoKAxx6/zDqTIfxqUlZpKfyU/OAIyhEZyEA0h/sLyo97
ZBJr3/WyXDoXV5E019hJfl++ISe/R50XCxFM4sQi+3Dn4scDGIsSn68znRq5DOSm
ahUiCwDXgEFxngz8A9XQx3tI7/BXjhlJkqHf0o4XunXvdeYJvzc3sm9KhylfFjek
IKwINLj//pczZxR2Sk4VGHmhQ86Pi9dNm3F+xNQvEcu1jf+PCtbH2kQAlL06SfzU
wizYqM0BpVk3UGC2yEz+0XJZ+UNXegBd1P39x0Ox+rBfs53iCqyQjKM7n9Ei/Ln1
D+7Ehyh0/YQ3EbSa7BKIcQp2AauPyhx8uSzQJQRRqFa1tl5Mus4lWG+FCwaWnqvm
QAuJscG755HRsVEJZEmP45d1bpLcM0JmXl7HD0hRSoDnVnXnRPMkH0s1JCEG8Z/F
FVmGizOFGEUYTS3jgtfOHgqiMSH7K3ryrAsiEfHHkX+jkFdddO4EnvVL/fd9WUlv
4jp0trdnueYXBrRQepwVQlToyCIBej/2XdvZYLDcJco+t0huChdDiKnkYxjg5t3L
1OJOpQNZlqutBuz02yD5W6YTSTXKjK4nSTPvdp9Mcld8sGD0lukk6SNkE/uqOSfb
TyBgluVsMFPAeucmeZp4Qpx6sQA9NnaqwDhwE3a/CMgEMGd+Mh4zKfXPmdPrX/mQ
pnyi4hV2oJqJVASW9twyofCyA47nGJCgTD8Dbr9EopiZESeOwqiRigJHAEm/9I60
+IGnVV81fB4T+JVO5noICLJQM7Ji1Pz84SUKLclnE5FCXJQX80dB3KYqobqanfr4
hPkMF4zAswfQIH52gMZuqRnT5GhYV5D1uPd7i2POGY/1PBh6PCqUn/gUoyj+8rxc
dxcIDSMew2aDmvx0Onj2ElKzfr01qmky0BF55dswSsxhg1+dIXFet1LQk3AW/bY9
03DoOkO92/nJtdCV3THIP9NRa+s7I+CR4AcoSBZiDsVTq01gQOYoUyF7Ure80+GH
FCdAzUniKvtHMGpYumjLFXLwwlzNOrLG7U4HPWXrsnBVCkwQmiXIYd9fgysY82TV
6WNUL03x6Zv3qUDFPU+po4STfLiGeyIV390kkqaZpfhbeZ6nGhUVrsfcDqOtFvXM
Us6Wt12xPxfvjSS2pj1lSQclQ23Hd4IE4e8tzmP5DBysC3qf9FJI72G2llJVwnIJ
1ci9uf4uyCFpq4Akc5qAWPizSaCJaYplSptVlGDkPk1J5dDx7YfI4lBY4PlZMq6Z
vbSN0K5TJurGmnpH5OKDXqp5sy3lMK9m3sMLvaavQ8lbOzlS5YwheVegZsqJZhat
KdVNO2G3atPvGVEzDPnxA+e2HQ3x6/jYsqWs6oLYbw3mwVDyUk4C6xpKTpvXOJhr
EihjdWKhAlL6AHzTF8jdCuo8Iw4V5PgI96SgmXDyQcqYJN9a4u/D107h6UOMaZRZ
A7QQV4HtuVzilUynFzzl9YbCOpoq8WrbLbMV9cnueQntcf5tyTgRFGFQnd8+H/4t
/jpa7tYFDgN5SVosR7HllRfZ9f+6dCRZ9F8c8MJG8utecjOcJ6GzZ7N55CdvrTSd
fPy3m7gZ1HsBqolGoPy1gEU1F8hvlBa/iGeTLjFJu0f5d/eICGFNwnLddqOkERwd
WQ/0WcLgeBpr+fXwDWg44jaPhPo8M3HSENWJ0SzJUfxrhc2JScsjsJAqidx05ip4
x4/cVGRYuyiGnhc32sqUC85TVlNpD8p1by/xMZnHhHL2RFT+n0fRnG2/wrQWzcXZ
shP86ep2sIPIAB5Vg82O3mP6Fbqq6mVMjQk+fgC4jeUdjlxKJ8vWiTTCz0VPtRGj
qb/NCy4NAyCGFyfjNtblUg==
`protect end_protected
