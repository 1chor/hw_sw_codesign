-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
E7D5E5UTPCiMv4FoPZP/Drv/gm/ojYwGjvU3Bu+aRNKsjof2tI71ovOO2j5AaweJZrO4qzlO450t
qlE+fBQdlUvMzpu41C1HNAxu3vG68Bf/1MZIZHWsjIoMAjnK/bQm6M2ovIoTvgxpYVItgg06GsKD
i3AtngRcIWMYJz4CIHdd+eRUozL5uvmsv/rVRo2ZjUfrsqgKY/2QraZh9pYOIrB+0OtJj1tnzTzl
ZDu+pArPG6Z72vnAShkGCSIrG+HCKM5heEcnpMIaLQ/pEFuOGIJy5G4txcrKWXIyKicw9OZk3Krx
Rng7uEvYaImAajo60flUVEL+ZCW/1HVDYDAapQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 79872)
`protect data_block
mG5F3l1neLiurNmCsbrFxPZCQzeHFnmeHCKLRZ5mL5HBqDLxlTPujTVfXekj6DsZDmFiyMDxr4yB
z4R2hIU5CLzw77ejIdeM5VMbQ+Fg6ZjIbb5dYUFpIP1HM89f9samKaDKniQRb/JpPhYzib8dbFLn
By1XLIWsecP4pqB0qjGgqsiTwd1TjwAIDrhVS1qFWVNnBlj9j3a7zivxrpbbMyscPfQwPzCiAPQR
bACgw3dQRGEpwOE6NL3kJ8CLL1nk4DRGHnlvXYSUNFSn3dXfGH6FiCViHgLzx5vDpDEekV8aywOR
H6Kg8A9IukPUQBWRNHNSdZENZ0uNGV9uZB6pZeRvpkYp1vN8YtB62i/O4lWHHCd1QXdMGjCS5X5a
27Jwl0pJZ+NXu9mCme9wR5beQ8Pv01O9gCMmvIg8KCzkN8esK9YMi1ABZJp85xRa70ZPiBVSKCrx
PlJjoXN4+1bBzHW2FCCdMjc28uqYRdDV3wwb8KqKyyf5GxmaASSajQBjrZxzlGJmxGlogLFhUJDy
GrCp3iumds938QXkrLb3FMqCFVbS9cI89uM7OyoTSlXSuAZgBvPAjwVM1mdREZnw1KwGAJQsSkCz
/bM5mPXTqN/JKTxtn6ZegqiS+gVDKWzBOrL2jtInCkFgTVSgsz8hd8qj2WNHY5aomqNqq0mQQbRr
aLUev49LG5oHlKeMp7bej1z2dBfAqhVQBZrU6pyAsAvePKKfLRauwIwz8ltcBSGPIXcxWlGGHvxA
BnsLjiOmzD69Nvx2c1PuJGWlBDIvtCjiRqkTka3rLXXa8l0hUdu0jajg0ghN0tFfFs0BfGBf7NJk
t7l83A2ckedGfYmaSiHCLz1iJ2xeXgswNhxC4CzPz6a0gQ+Y6mXIU6fLdZS0ANo+Imd49nDbHBEt
ee2xWA220VvRcvAyD+cDkq/2WhXwLCCU2gBLYEDjigisy0ZugqNqC9OhMgSzmmjrKqwXxD2BqF5B
Pr8luG0nfWB2HFTZZj2eHzt/JAKN0f4k4qk+GBcNL4aCS3TBWJrn8r0YarYG1erhPOr3wfKeIUyr
tQ2v2OX+a8TvCa5jCU5JjufcyDG/s9tS6mg6WCTFAcTOlo5GZc3nw225emPHa7NnVtASY3EH+mMp
3lgfwfvgBGPa6m+eOcUut2zTOUsAFAW1icDj+DBKZi63dpMt9U4bsR2I8bKMIFIH2M4rJX7XHwY5
lQRHX4xspmZlDS/3ZvL9yiD1Qj2Y3TtyIDDlLVBYJjDGMTxlIpz4weZz5Cc2+6u4UIuMcpSrpacM
DyET3Guq/jxCOc9YRvlq55XSND433R4rGF9CRtqot021DqOfl/pR9bWI3ymWWT5FAFZ6IQLzcici
iFQ1HOu0H0y9q0W73ryI8kQjcd7yv8LsyDbNjKTomWJdjsb2XQ3QuzN74/tDkhGxZw5FJINhdllZ
Jq0k/NaMDaNr6wu68osolgBLejlc2kp55CKRB1rSkyeh4B+UCr+lkOrrYjqvdQxRDJPzPwdj0Ca5
eqb6NlLVGonVWInLa+HienV43mQV7KVbVWrFGm598aC/0l/jdtZ2DCd+XOFWGuR4iBhqs+S1kmn9
hz5hLza57BzXljFhhBMVYEIt0pCJQWkMC2Il2A5sKkJxsCdkEjfUv8Pl1HPrWlavpkxdCU+ZliIf
yE13E77SDPweoLMMkR6ad2wii2AQcp1u90LyRSv5izA2ji1Tv1VA1n3EQso5t3WSxViYFJK6mL8u
6M/VJdM+RKBkuNU7yNf3K7EkGFO5KAqLfKYL9RvuvYQTDupN8ZK8WDrWxXBqKzHwMb0fP8vfApiW
/1ZKXdFii0oKtZ3TX1WdQ0sPD3eCj4DCImuLpU1zKTR2Zg7slIJznqpSQ1QgLwQffHWMDsLoPShC
fX5VfpmDxjg7RxxTC/erY8BjkpuSycA5tflWqzosAR+x8wcJBF0EtitPhctYPEDeQf+5qydH1zb/
khyTstCMeQ5E9DN+NjsrptB5tisOtEqL3IBPnIfK23JxsbDa4PlSy3YmZRHdLEPBbgxJ43J6UeUo
TD2l6Y5W1GwfVN5Df5wHIgUKUe4lVU455eFFRJ4iX7wLes/0yyWdSbAE4KZDPzVS0OLU4hXY95y/
CdZX6jm8rLh1ip/4vavRo9T0r/JqpF4dWa4gdLlUnAlEDmADsYVNJyHsQal3kPIYxkeFOsM4auZd
6G9MsQePxq7vanp+9AjPwzhq7qiqdqdXtwGzb8EAHCDqNvRHJ/XXPtpPI5r6vU5O1rEcSNy9zSEo
fvrCNnZuAKU2bO2O/n60VeKJmwVzOZPgbU+kiGSjq+m6iVhH8WyAOldVIMXVFPA7GJq03HDDSWa4
2m++P1HpagCpnpskaYyDKeUVAvXrfL1+QW5RRofZSvpXr01PsvOFGqIuEBWhTuUyexsyoCoULF7E
gKGhCAe9wIdRMTm+0ir5IESHmeF0WypzLEtJVeGDzN/c+cK49C2o3/Ztl57GugmTnPZaqZ4RcUqh
a9FfhfsrxNmNKI/bQK5Vf9ZynKE7WdMpnuau8rwTjzFhGpLE9W75gBm01FTl9i5s2gSDRvnlEsIC
tm6DDxTj6/rZbzD0JB5uSE7p5itc+zwJZJz5zujvOlGeNT5kcQtk7tmF7eHCv6zKkKVRqQv3F/5s
b0CUVtRUX4+dbyhdsCT1BHu1HG4IpU0EAkMzL6lS2lG/90nMCZDs2127JFa5MdouiVrI9Iae2jeg
1g8ul56gAQsH8X7Ke5+0J+TDpbwiMTz7Ix98/XoywFkdgxBUWVF0FaJK7MrqB+5XgzNLakFPtj+Y
ut6eS5QXnZQTElrcwZRnlCGyij5L3pgKf0mwEzkRt3Ty36n+5OTpPvLAEkAQ2VSgz+RNc52wLvUn
bfHRe5205m5NG3kNMz64Fq3Csjqo5+6O447IquFuZksMtQ3STM1lIfFli+kGpxGDP3bV5kbV+8vd
zjCyX6Dun6KO39DeKyFZOKK9J1F2Er523xOoMgtODuY7SHbXNDipiXk+YQ61FFKYCv3zmMo7Hy2R
pN0Y/7diwoPp+vJlklWvMGinXUqF+9W5PI+GVNwhbdSkJ3olqiGhgDq2wy+6DlTcSR6RKRdo32eC
uYjHoVsLSUu4i7a29e7E3ZIGKh59AFRTvCsbs89WYO8CDVIY16xQg7X8XiGGRu+G6D8kdnv4VigA
KyBiXN6zv4qVrHN0qzkQhixtoESblQWnhgrwRuDeo/c/AgiFcj/1xZ102gkZG6VqSv1NfbPZqeAf
WFPPYYhh37LRe4H7R/rktcmF7UpfuOnV5XJTzopt6uPutToMCbGriwo4IB6QHIkK9rLXNSM/OFpa
BM+WNntFvaQA9MoToihdMeZwwzyHelP5m2eishasNUTuoa6DNFWNv4wAvyaMXzOE94g8dKvkNzgq
p4whfW3RkdplXJsEDD7HGI8ydYgImzp3FOdQYWKKCPV2JtK04BuJzuq3yl3xL5nOK6KomLJvd9lY
BrhxEOHhWRC7JAGHmffSc8cz2ZZG0ettYPXsAQqWkL8Q0+2AzGg4Vczq0lrYj9Gu2lHNEjBs7+G4
KF9d2mOCxl3y/xgF4H6wcOr2r8s6KOEmCCaqAIDtoRfzCmbway64Vup8p2sN2Q7uEoYp/pKvmT/O
y1oxan0MRV8RYP/tvPcAHAZmWhHHIh1piYUPzRg6WglNbMyMQE5gknpDz9ee/JskqOFp1vpMuRkj
YVjRxTIfi6uMrfPYOl1oGa11MpiYW9LjYT9mCEsVpUyDLIPpuixwUhDHmaDnLqjyn9T+zOvRLysO
6vxzFff4BT6Z/maUqN42iBLrxyuPQznxShG6i7JFQALLMEepjrAmmp4xcT//aVFYTqXqhIQxuSso
duWdY+U6f059+QHuLgPv10f0iuCJqsv1SgGQFQG38V8MSvYSzv51oFDQgtGcW4Oi/tPJ4G74m7wt
+AQL3k0LgRAwXwuRe9C05ipBGEPeUobehEmP/5G63JzEnlhETA3Rh3+L6u/83/dROTjna8VTUlAM
dvEMbsrJlu3BHmH8jf549RDqCIDHg3rtMpcGIB02v/UfV3i0JY9LDdVgpNVWJG9qGWChRI58+ROm
qbgfMRrlkOkhLH3x9xxLiM4xaplVTb5xHlUNlUjhDUiUthMf4dvU92wYgXGUmV/mTNx+idSdP8gu
YcXlHtzJBM3kYrnfJjzNI8/t3xk8nmhxM5YjD9vklmJPT9FirTZEqfT3MyWwRzxVVtAZNv31ZaEC
fWb+75W1bQhppJHJqZSZLs9aBeE5W2HT8D0/LBfR3YR+KU9J9Iis2qsMN9q0ONOmSHOjPOn4Ks7u
2ou7MaqXAfGIOrU7tevK43Eg2yEiw5+4uU5cxlfFVp7t61EdSiq0Q+1848/t2guzuSSwDEgZg6GW
FaYcTaBuhDShlCQLnfFyzMegwi4nONBVQsAs4cetrx3oCLGsYupTUal5PqYnyyCxF6tk4wv5idaM
b+MpAE4CUtG9nN0/K7OVZd389IN2S/kr0Mo0y4cQFYXnl33D63tt3xgrIHYRLRT5AKxy/Ldo69gA
XnIT6YtNGoQ3IH7lE55QoqOGd9dZaYUBrEAmL55r/kS+Lu6qlUTgn01Y1l5c5jlho+W7mMDhMR+q
bVUhqG5f9KvJ3Hqg5RtuNwGMgM//vW1GdLZjy0e2NZ4QZesLsVtqNWnJbZ79utUoUxouwWyHo1t1
9uNHagd8BI1y93Jr3qIUtSC0Nxn8ef0ev2qP3EXRC74F5eRZXmPv30vnj346p+EDXh4gM+wsotj0
XEQmlzwtLCpVkElyibYJeU3aH19z0XiqocCNoSXeJX9TmvZHDYSQlobD0e5mIwz2Hxt0jSjfPtQw
cIKC+SqTwyWDRT2ytQUjrY7HFdTK9OG0BaK4s3jDVd0HKcxxR5+XGSQwFax5kpQwKtezdBRosSyD
f+HsEDQeTMv0A5Ik4nN1wLjAbmY6b5gIkOk6tPlulOykM1WoSa+BNYezIWtspSwy3B6IsbJ8FXVo
HpuGtZrb4l9f/2qtry/QASRgCf6fZOMSVpQawow3XdD7CeKMywl+CVNLNcnoJqkknHs1/QXk7t5u
fURU2w5Y+MFXAtX34H+t342dfhmKEQEhVPeie5FuXwEI7DhJpT6prbqedsVXJDYgZOKgrgkV72Dz
RhHHeJbp7LSOXDDuFAPnO44IzWrMDguw2vJ+L7rVq0Khhzw4Utg5r+m4awtLcj/gQeBhzoyiwRr1
cRYLt8WXix1KeQa1f95Rt7Xc4o6DLWZ2olsci9RLew4rB68JzggxoPgTLDn+/0vXsDusSmGKuPLx
Gf069aSqmNOFpKh+7K+RNze5QNyGOls/0s4RABvJKWKbcpU/blWVBa6mgBe+eSa/ixLrrUAmSgub
TWtg6XcARe69eYMYYpHa7YM/9mITZtemiic7xyFfDzyN3zke3f0jc+uSw6He5VmMHIjPPKalUMM8
H0sxyvnphmu3Wld8w5DHAmh1KbxzDs3SULQ1+1Ihk6apxAAEzjNgbKfhHO6olUiDLfv6997PLvsX
ggQ0MuCKbgs2u4mtAiUymgWU4kqL+lRvAupK2pxlxUxXGFCV2Km7vrsUiSOHF4uD24eljzd+J65H
6Zdy16D6vC2j8u00mHjS+A3qxv33ywTb2X5W+xurnsS6dkP/+I873nKtvDnX9tVYNWBzhPJSiFXk
zM91ZyOQBuuVBVKFWatQqJa9eh5jbASsYCCnZhT+pvDN/rViB6SsFa+IUjgkHuH788mj/J8QWM4u
eCcgqc+I7smZs3BMN8RNtJQS/2I6Duc8Vbx2TAO5SsDle23ONfZY+UJfOqzVG1DIWuSiYUSwCujz
5BPpEWoEm7PEt9vg7tWoKWqjgzp9KmUz0NrWoEDtmdjQZQTfxcp6D2xQMEOIzchG/2ZdswMFB0Sr
4E/KwkmdO9hdAG1+7sWZ2sbbNWX3iOuayFg1ZroOBfeles6iTdIUrsFQ0i5J1NlULrLVaxTd6r5h
YB8Vi3rRbRGw6ZpqcQ234YQuczde+aOtJjp8IWKvdu1bIQDP6qH++YuOy//3tV81+EKvcWBu9qxU
qu+ELA3L/J4sCcXT+Mbcb+snjCktpaD1ULznMEE6BV+TFTGMBTtFEfL/OCT/wYRkZCgOtBLc1AvC
QlBO4YVNj5afPrDK3fn7OcQKTzoDcaGSo9jNETIFyOrGQ1AESbXDv4R8JdZ36xlfugZrfoJ4uUT0
I5wAvI/BLdfKSk9TWteq6vrY6gNsgHjKYp7FzRbd5bQgqkfg58Ax9BFSh05NE9+Dmg4YgAwd/+IN
ZhIV9YZN5+7lLJM7RbHsJJ28Yp5FWtNgP6gd4BBQet8SUZ2agq/T4boCsEjWMBy/z+kCvONRNStN
FUQXz4sRSR/QmRk7cbDsMzRyEnk7CzmsejTE9GxqKo5nH7nHaZVLq/N/IU5Q8oWrI5HQRU44uE5x
Pu4+x15ofrQ/luADkYSokiEyLA4ep7hU1RB9+1QzL/z3xXpO9jDUGh6pAXafceWURvIUEeCtCSxG
S8QnyCs648F8PRZ7cHM9uZrOMJtcoY+/RPAJvkXeAeGzPhwwE0lxVyLnwgXDZYGa2fDX8eTD3XGo
3HOs0pgX7lFUowQCRyrBu60dIT9ms00VJ3eDieosIe7XmHoB4wLzk4xsfAr8tL3caX+TRr0rxned
bqC1GkXYIgc5mB+F04q+PElNUJSP0ma+z13EqDxaQalu9+e/6ye/y7FEzI26qRr8HpqEdhQDSxXC
V2Obxsrt0Ki3nLtVL2YtYBNpK8khYzEXbQNf+fuOUAX/u/kzZDJxLF55Ut7m65rDWUqZ3FLHqARs
noquwySl7D5aLQMjb7x5ixdR+u4PudUdRiO3fBjbe1LrXihZL211LJqlb8JbByhoVlrL8/A0DUZR
MBfMsqxN+5mrkDyEqHNKTXVa+qNeAQ+nmcFq8BpOcYSol+WSDbqddg5pUQOfDQbDcadvSyRDbnuh
Ds0ttL1xINtS57nBS2AzVs0Auxj4vcc2Scg68UPuPYg8lzDPpGpS+Xmr3cEt5HOXSx2TCtvgxt+k
lHnqTzUW7t2YauYdi8WbPpIbpfSmyNR4uJCHJ97rXiPR3c3V4QYUwIYgNetObOulYx0vVRlRkhrd
rLJAkcvCS9f9iJKJnfVwo7ZAVmZAeigmQAKDJqh92lb7T6anXrPv33ZrE2zyt2GEQXx4PM1j4oFt
C9NTq9Oo6v+N9qFq7kJcHwSxzio2Al6AeCv4C8B0k2JxgVd+KG2MW6BbdD94KD6T9QmjbumjysfN
7BLXF7kC8X83GyQB8sqQ0XSMu7xEsSxWbMTRGmplHrsagH+KFrDO47dnZAnHYz+R3S6zihvlL+45
zVVWvVB1YkZA9etGQAwhs0Y2wV8GpKyKLabYnAz1cZabMVXFnEsAptm3YgCQT0e5SWJCkeRiowZ/
ZUiOdODfWuU+0UdOfDsYEp45yaRQO8MQlRyL2K4fSSr78DIjKOVvEBlZoyxbSdkA3vxj896TS82e
Y5hBUIh9VBcX5cU18wP1gOhUVlul9cIvYGICFr9icKPjCb1Is2MtIShpIA2KKQrBKsT0zT81UlwY
C2vVvCjoQiRlb3BSHU+oITWmiY06ykoicJYWxXhs3ACJF/EbbxTltSLHtkeC7kCy09XbRFburWmb
dT0z7LVASe4Tn1Bnmi3o52F9R2EajwtH0j+SJoz6Ynw1iL1pzG6C7CjosBs1PgigHxYmokvZCPte
inCUhlNzPs/xDCFlHEWEI70zCWLHzBPAh9nN2WjjBZ6fu8C/iaQ54HrDwwlkwrLxUszmLjZIRs4n
uLQvMw+krmU/IUGXNQdZQASD4slqEqRyjYzOwof7pHk3r3RTlhrFLg5IOzgOLUio2VTfUd1nocCH
eAdm9x+xdpja2zeHCRC+KWTl2Bq+FOKrOWFEsLW32FV2x9ygvKnp2u3HqGh9BRWSo+6KjtqMLQ+f
THdoz0F6sWkAAoxd0Ez/fo7X+eg3kXqzdySQ7XhT+aZhrkLi4G6QuNgcoik2Dy1zllIt09rk8Db3
/a89vat+27rcg7mqoGHDV2S25MteOyEBOs4S44HQ5Fb2nT2kWmPjng9lkIbx0pOJDPPd9ry6Punp
po1yjFvCfi3DVW74Ite9yOas7UW6VSsWyT5ksPo1zVf5ck6xBiSKys9ZlBeSmOXD2NF/3y4gwFso
NMSUyrAJykPk4b/8H/J27/ucsEK7G7YWVjIcHdQZipVmyNDq8Ygz3c9ijsFHksUXkQC9Y4Ba6o/B
Wm6arFZGS/fAaLccWxyBBT/1emytWAbayQD5WC6Qw8I15x7zUXFTMp0sTpc0m8/nX7p9k8bTjRNe
9+C/b61+KFSBluFPOC9cC2ND36RZ4YU6Jtgd94HFlpLwb8yh8eVbvI8hWvUxcSfGtsPno+BnabSQ
PCCpCKxqq5oOWzA+5oh0sZHfU2mQ9WFMINZ6TxxsWxsmmmo6CfEPpWgQuu0AMYHc4bNXAD13YQyz
Z8NwuOPeoEzU5e4t8tSUHGFp27XRADO8IjKdZbNDOAUFh7c08tsw5SZB9xSmq68uAp5V/jZew8mh
awLcezbUs9YhtKlNdKE5FogIH6h3/U42EPPwz+SUHk8MDUq7GzR3gGlI0JKEM09FA9b9jiRkwDTn
nkGguC+S8eDNYiXtITyW9yo3yH7HT0UJeojRiFi2wjzTDFyi+DT8JiTA1feQ8deji+H6nbIQwkPy
wEVKkj0Tzjh41dk9n2zJNigJ79zM8huzKnfoDHHPiTefhZzuKHwb9j/rx7gPywMheqUgOvtIZSnZ
cYL+Uo1grhQa/gPQVDD4OM5pjTdpxvTxy9YP0xpDXHeBim7a3AG/zMBI1hW9moaUzkOYcucA+ha+
oAk8IhxlyCzQf2bzWzQc6phgmviTVNkSkUrCLLR05IW1YMTQ1h3BFiBR4naSI7gMREocIvnpZZGQ
E/5Fam5TQIm5CujY8YPozsjaztD7CWswztjH6KCZpEATfGxlEX2eKlAu27IBu15ZZ5KuTQwLsSh3
ZKpC69pczVJu+SLHPAHKiatw9W9Z+3ooQrh7BGICSi62ZP+M0WYY49n2qanryh5t/+MvYq893lzM
fVDd4/k3wXIjYWttlOHtfEq8NEjc766hwloQD/j0dmgIiya+rEjkhlzTrTgN8dOdB4F/FWFo2vEW
om+wYFiinNyiJ315JDSD1mInaDinkzIiZKtpR00ibpDDu6dY8L3ql6V18ckpIutUubs2HzzHn8yp
cK5TFevwIiDkXO8eBX53Zw4cic41NVNGm22gIX4hDD+AnZ3k64XEZsAmENSsF5mMlO42V4huYiD7
PpPbQ2vH/hP7Kt7PbyNfyySeviW4f73ar2pDdA8qEgBQyGlmKCXkUYa9uqhD33MPesSRev/t3XjA
e3FS1Pa6oHAxv4Eso5OKqUfDOZC3lelHwTWuvkUjWvPWYanO3FVIPeOEIqPUM0jznLbN96aiyxpG
rTlUnRncLMedeCyyMOVGySbp6H5LWWdtu7V+G3HkPTqAnLEb9RRUx3HU7Z3rBtecZVl7JnlgYizV
harmDAgznvAXo8vm+DJXdCL/S6HbCpu25GGuCn/2QbQFnJU3qbev+X2BAZZkicg/37Ib9Kwk+6J5
H52SBOHx78BS3QuLj/As5YHNQt/fXIRteGOtVTU7R0h+0tnJAkMCOKFnhLsYQhRCl+gBS4JsVVDV
Kd90RmvMmVXg0BV+C5IUz8fCYexzobZcsgAaScOq1dtcfNN2V4BrioLBqANdfPFcbCkGTyyfbiny
ZIbRCNdgO6WbnZMBUaEfGmXM1xPWpjUcIRC31K/k6TaohDMOXJ2vQMuGuuWhvl/5CtWlDV9v+WO8
7LrGcZS3k0ODlOt/yDw0vxtmjgPnzP0n9NJ0XY0IccVGrC2qQnSOoFgVFcgSYNQzuGmdGop8gNlg
Dl98ec/jztEJmD9uInoa+1VJfzuA5ajldzrXFQ+lbI7/ZxTrf5Ghnh8Y2+w+4nlgO9RCu+LPRTHR
GnoUt7+lHeE+xXP4GBClFhisd3CBamjUNdF7C2Yb7sjHmFhiorveT8xud+dbT97igCc/TUe6ZvQi
xv2OhKQUesSfFSdRtX8Qp9+Oq2s7Z3OW6YZx4aS96h3pzQB2rvEhIzotmrqIFOcxQJKR89sgZId2
DTc+U8YYHaWm9+3cIsuaXXuRZt3o2NZed5pe5E+jNIPskzmcMkOzILEuIkIpqYP7yTlYW1lwbMJK
mWOsirZlVeNAhpxgAqRMRFSRj/C7RWaKe0hR6zrRLHPpbo3R+Kp9ZT62ZAK8apUDW3SBSQCzJFHl
xz0KDoodqPRNnqlyNr/OyqU398P4pI+AFffmxVFZ0A+S0u0hIMATJCEMfo/fG+lFlqDRX5XOHkR8
lwU6yn1dAZdttGrMF4QPbQiEsWn7f0B7KrCZqS5bi43lK5OUn7mAUate0rZTqjL8paT7GklpFSl6
6eu5mJFqTfhNMcxbgjjM3MudJwPu23gX+ew8YQvPEcHu3KgcKoUaVdJ1GoITNXlksscZLtwNTacU
DDaV2z/R81waxqJwwoM95iQaZ2iGO+WBn4iEZYSHQDe+h3WdUG1Hp6mhhCvXY5M20BLtIW2RXN1d
C2zlwH3JZFAuAN65WARa8hHtbVSDQNYdVE8p7YV2kJy28NmeMCqyHKKqewXS43w1tS5yxRJwLrOu
UHR/VfVBirVkNKORhUZh77tH1JG5+sxSjG0dqjutROxR3RIn2rJTcsyBCaO1mjSlVUqPM9NMXMb1
lvYZYVrnryf6g1srSkn2LU3WTbbwC9B+8ZKgiIjzZsLTb/W1w1BwWuoeaVV1JX8LVO51jpTtNLky
9fMGQKzVOYdNO8ERUZEAoYoZzyDPPM6LaYrZjVrXEhC1b4nSn3m4o4USlrX1hFVjonEMTfHl8xJ6
O5gJeoheyeitru1vzAukU3TC4FDEU9FnGNZHYmrM4/dcuOupEwzaXWVP+Vme6DG8vjfQNOjBw0AQ
7wJe84Gi4MXpSjcSfa29ajBGqY1BIvUTepEQHP1oNqCmiTT6Wbf1qoCkIt4vYpX71U8tummZMqCT
1SCMNRQOllyjnc2QWpXziOA14E8aTUYjLC85l8iwN3oSYtZ3P0/TEisadEK5vXtAst7hklsCgh+A
vXOzIiMWaUuG3PmX3AUvDEYRUlHokLvqZTYO9ybJg5FzV8XJm+hdpwKTkcswvJYOxX9GctYT3Nh0
Ou8aqu3Md4N2lLpwqZHWb+CXRjwI2WLp9UZ52pZq2YPGM1DTY55lauiWJLKmkciVT9uUSokr/2Ch
Jp32fJxc+6faeHUkk0LiUxuOUcsOGOtbGlvMwWd42e/UYMyIgJrc+mEXlVrZoR/rPWzq4z5pZZfg
qpqmmKjmfdflkqJ8/xVEnLKXlxOjTwE0nE2Pe1G93iXiWHQXb3dBq0a2xHmnzaKm4SA0asaMMRpz
HnEXQyuIxLKo3flqtmUUFEjHIQMANLUij4+T/Fe8IRaC8QjLCymF5im49woj90jNiRklvS1Tm/57
sw8/SyJqGvX/LqDIjbiBf2Bl+OSxmVQ1eZUtfHSD14jQC5eeKrdpH64DOjK2VmKI4IHkwn1oEFV9
g0dna3YxXSQnwBbrmaxo0Nr3+77L5hVKWNUaqdyG+bDgDcHLrCuW9nFP5HDKZJz6T8BZ+1sx/vwj
6Ex7f4vhxV8RjFabcE86Lh9o7K3VZmULQETGoiDlo9eYYbSsvjZVxvozXls1/uC2atifT1mZ9b72
uLt5L17Tb4cl3s/Sa+sKkC0NXorAm1R2CjF4rjK0kaC7PB2N+XyqsD6WFTzs1lUGcJ/FxDgSTu5b
n2S86rPuhlzB8ukQzmROfCRCpMPIJtmAoKabjYYAqFFm7YoqvurjFMfM6XfrPh8DXwSmnIty3uYy
7Azk1f3jH60Yv3E6RC8Xvrj8qMXWZxYZyDhjYjZ2hxkpeULIeitPVR5gycEaa7HnInF1GG7K87nK
cikomlv72jc2c3lYL3IT2ZyH5v9SmQfHUKz40BQ4O59b0ZK7J9Vr5ARAvPdneuaSRq3Fa/rYaQ7R
bi7dPekrXvSov19HuIoyBo0JVI6S9t1iaXhyYJDtrqy3s59UswkxUEKCZn8LwP4CSk3MLaCcqh/I
v4Hk+ZLI8/z9fUNsA3tp7VldAEhulkoc1pkGDNBDw/fKDk0UT244/8NZCL559D6zQRFcBhCDUbNQ
rwwuHEjmZkqloNRDqsQQ0DWcAkfeQLnMsX8fT+I5RwKFzlSQ4NletO5fxf9zGlv58JW8R3R913EE
jxm1KJsr74gtNCD/Mnk+PWS2qLRYB2f8ymEa6XyanKt3Bwa3F96oU2ztCyRFXISx8FKVa2kTSLDw
3IAuVEb8uBg9h25Vr855xcR57f4kkXzvfFYr6Tn2qYfyFACm2k0ocj2dDIJHlCaVmJ9TcJIJZZqv
MxvRpc58/3aasAwdrrvcYXe+dTcOfsl7vR0i55S4pGcuU4H2NZc6uEG5nh6WTGTAtEdW0Y/EAOvm
5DZPy/XGMkOLkvZfDWv60Hu2Rnq24JLStf4K1e4F/UlzXCxKh4LUN697svy4FbkFJPD1Y6q3Wrhe
2TgkmteWQsFVxps6dyLSuCH4CLN6eOcrSDq58fix4mUdVJ0IEaaPwgetMawiWLTUH9QNvkT6Mzxw
mvyUaJfLqbXMRy2j0nbw3r3wURgS+XuT49s2oxJ4wqXnLW3X9HsTy5s3rj6kFxR3iF9FQIBzuFtU
Cg0r3rcIYGSMw9Jm9VnoDx9o0OyqNq2gyVb/CbMbinFPPvVuudz/KuOjR0DxKM8fmnApyeNKDUCn
ULJ6EuBGHqJTanwCJoirpJLzkI6lD1DuZmgZowNUlAMxCxTl1mblF1MLCCgzrgTjnfet9HwnHp1/
2+b/fiMXh3U2chFCSp6WA+VhohW75oTnv591azE2oxZT2NuLfrfgiPcd48rSdOfafqcrE4Y7wG6Y
dwsOtCWoQqnkazAgxPVaTix+sE1jldKi6JR79W+0NOv9lQz2yUD2EX8d/Eds9iohbHHjmdPG/UJa
7BbQHF3rbNrcpeoO7hXkwjckSPMmuXxRSHk9cwlpjyHYkeQ75yO7u4puBnEnVCILtOcBHX4Se0c2
KxfxVRwzwrEbltgMvysJNrZx87WS+efmH5IDagyPS9mVuTxC9kZFQKpkJPYfW+YxmY0JRDwHy5xw
W5p74i1CBzeIS08/DdQRni3rvoIk4nUZWCj7tW2ZuyK0XC7poT+sdLBTCr6GQ4Rnc/shlUn86C1l
Q67mssJMVAax5j8B3FW3TswL9lcyJdYiL0o0gcesb5UKPZtEMR3At4mH8EAN8e/wlZt3TIPhJgWO
GPdIbGSRMG1wuWyCPYbGJIPxLYIJ4IAfBfhu8SK74Mg2Wlg/CZTKsw5m9rk9/hqQk6a4JibWJxpu
KMGjMmC8Erwx+D5Td+giVf2ymxXiGflVqfg6/5J4my15JWcbm9BAJOVy7O8T7+eQVL77KvfsIdOc
SoXoMa/G8bW0F0qUZ3wQrFOFVjq0+sQrAc5zJbzpy2tbO2ttg+FOM2hKOedu6jclH31yrn9xookV
ycvzVUYlatWD+f7X0p7mMxpP15kaDoH47I3UiLEdT1Yn2z9adAvzlb4XUiIvL3jefntraa4mJkxE
ej4HJH6StyOYdMnAfyLglm7UcZ5UjX3JdaszaBnClzWdJoJz1UXxPCaeH63SaF8chtbMS+J2w5ha
zCpBqnn9YfyvDHu9RE44dkLzCUcExpRBYWrA2zFUxckY7EEpuPr90dnEWaiRUA2EYGWIhhcbhTES
Njz69cs+FkvWiEbqVdeqfU+oCnpkaLpYLmIdNKL/mQScGZEqKovQlWWxqLNWh8UROhtj5CSUdi2k
RohwrPyMl6K1TAFR5IqU1LSM4gp7a02Q+MdwgKGW99coemx+aFr624f38LtJ3gkCn+lS4/0dQ1nU
Jn6W592up9qbX4E08W/+EeYYpsr3dF+3wHAP/ugS4alxTcOgHqud6a0NAwTQp1jVZp+XODaGQD+3
42/GsV4K+GioWoa8eoW+2pcMCbktJf5JUA1KtvHa2rmelI9uu0zxUidiq41Fk0FHTJ1faDYGElIt
u8SKE9vulVsYu+nTV9FQiWj6bbn4F02hdhqkJiZPh7I3JzorzsT0Mn7xR9eFfQUXH/198kczs66O
wGrCqUne6RdDc4F4eeDK3BTgbdwPPH2kLBI7DVVlp5Icaso4/qapF/G3aaDY/CfHcC6RMKeboJRI
qjfBDIq4bkcJzMpC4aafawYsJ5EuE5ezhLxjnTfkNBC0uh8FNxn8i0/xK2Vphoq2rEMdbPaRi/Fr
JGJsWey4es6LSfKvxCUHo9gHMceH93i16pEGPa/gs4KOLykqxWdwvVafi8imQkECLNCpMoURufUT
qTRW4UWBFZeyWYaJpL+8J95pXS+UuCf8nsChDff99lQ7M5YyBaiIsST6vaQpx5z0A+y9IzVQKQ1z
tlatUTrJsDYLtNYdf/25b0RVT0RbFTcUXY9pmgHa3sY3BSy61Kwh7pTJD5jbLKj8/pS8j2ywcquv
ppTySNZv/D8aTFO5WSIPcEXjjwaWZhDNX7IDJzNT5i25qLiLuux3ADEmhArhUXudr3IznVQcFhZh
/lE7sVPKRiLan76t88wz9r8DqLgV/BzB8dFZBTHeAlhtWqWapchRU1Wtb3kRp0QsKOBXRtX11hpf
TyLAUdQrTbK4EVblxn1Do7CUP4NQ9ARdNArw9zeTdObkC3WnhvMRNsMCOD/FTGTzlQYyO+8YGmKr
+Ewyb1juRhmvA8OFpfhpEMtZiLmw7rE54zUGM3KmmDlw4C4EsMqKE4erGGwPvp5BYZ5JhcOL2sv1
dCNuSSOqZr+oKTaCVNYYENCMGSHU4cu3LyxK5Pn21+LzeMQ5aWaBd3vj9pbwx8BFhu74rJRcGCav
/DQVevjNpduVlLMn8veInFtJOeEyFIVfdOq5IgYWS3HWBuAU7sjNJOwJowlWBadiWoKkWO/tru/P
VaPnw5oEuGYFOF5bWc+9GNfLD9VDU0R/MFRdfdmc/Nd22pp7a9b5BEbethGZ6LihdivwScLqrL7v
l669fO6rWItNG1MW3yVCuVpW2vvmWX8esNjiiJVBdfW9ABmkiPn/nTCxWReOEmns/Gbq9QEgZ7Pm
stjjlfp9kgc/Wi+kb9Qb0DF8b4HBqieLjtQlReKd+jrvZu7+TLmO3lMljIHxixeQc18QqFtTR3mi
FTJTsry3FEA9EvjBoHEpNTl9xiSYNSyRIBMOdYIKE4+dVdONVAyiSvBfWzRQxypvDS9HHVi5fdok
eaWCqNDPP1pyQI2gnSL1pcCHlEFozNyxgINNkEVih3h52FIfb3iEsshx3+Tx5o6kj3cwxS5XLo3Y
k1yLpBr5YDWX7YqEd7aqPcpzR1/zAvVzk21eBKw8GAzrZt6CNTADvxa5U0BtBOTcj2nbieoEadI3
Tz8aKAO+gRJ/pZ0EMduM8VLjkr089E+3TNZeaaCjwNyDJNUc0H8aAFcOyThhYZqW1FKSpBJ/eUyW
O4mm812h5JcjgWuCt6DACd0CDeLoh6qFYIdEZb6UmGzhA04PUHR28B8a2Toi201T/N5w4fl59uoW
gEr2ZfMK14uRCmJSlh+SiEHln4V3mRGgs5zLeLgdDQGR79gXtiK2HIcbsCtZpsvMTBpcrCyUs2GI
e1pGB9KnTeIX0YOgW/VYJCW1iNRBo6GFGFTOfQxu7irluqmXMUMT+xWr5InWjz4PtFPCRs3mLlSd
EmAyJQY3rxPd39B/TZPP5TIkhMRRQ+RJs17iPb7wd8vgeqc56aI1f303kX/JEREedTZOs24atMzq
7h6CZ/DMOoSAKryza3ZqV5A7jqxK/5ygIbGPvF0eWvJSl/vrNkTrCDUPLC90C5/Cbmua5LNXRaiK
ZuA6meMLjZGP/vzNh5XfFukIyQb4b9Qt/OcfoRtCXrGKR9Mvmz3R2Vy+PUkkrRjFjKwJf1GwTVW9
Ew4PF1vCQTKIXmiFtCMQX76qlmN9Jf1U3cRncZGzRg8SbNlz9tL6gNmnGN8IgAIy3Q2K8FDQGo7n
eTdUurIqiMBWP40e0e853yheODgwYDPyFWn6+MeLqfmGOYgK00/Y+ojRN1vNRjIb8CURT6BSJBOz
taLRVzAO3Q7ePleFuGHzGQCVb2PanyvEqKRFb8/lNGmbMEOqey2LwBQslaUAG7vTuc3nS8b9v18T
dkWvrQ7iAUCmfDNZHeBhPQXLZk7PeDrdwTBY0pAAuBRx9w29KESJ2ZGo41VxdA8NRPgf1zoxd9zz
1ibkiNV2omk+ToyzZIMu5Y5S0Iel9JubXtCB4ZBrnYtdjReYYA5qgv3gfoTcYU46Fr5mJcbSr/Z0
zyyZpO0/y3KDGaeleWkL7c9eKounDOxDIqZCGbL3I0JdhIviiWJ6zPcA4Z1XRoh4rthe7d2N+IcY
ietHQVsqLqoIfH+Egj+9vwC0aF0WVLDYuKkFMEIR8Gz7xbM5zBI5k2oqy+rcUWkyjHs6hdXftwsQ
UgAcveuETTwdVC882AMLctP6aPx6MAYMq+CMSyevBeyuI9x1BQWsIRK6vLUIDf30OjnblpeiXIce
m1MX4btlDaUc5S9LJDI9k+Tuz9HNCeUwYwMbtGAP/eUN8TdMJWzDAlb31K5I9ARklTOKONHCkhXz
TbQCvqOraoWaWxnBBnffYgH6a58bMxUASxxmkYlgX9DzyiLGf4WC9CrD9l/W0Of6ds2zuP/JHn7l
U8mSF1knBJRTHbuplZYFLgP4h8mC4pbYHbhOHUfQakmidos8VrpNtNjAkJReGIQFr1ONHMdRC66Z
1pl447EGpl1xGsPLzf7kN+0XpzL1Ay5ZemPgByG7EkAuGDgneKWUFB6aCkl7Cxnv73b+38dxziC0
w7tVJ1ux/6nvXbMoLmCoydK2roR7MdhMwQfS/zQtefgigCqmsv1DrCX/z5Gnu+3E3IEEizqTs80l
O3GkigfUuXIyuQhQBav+gYiQ3LmzGTjpgCEdjcMOjcyCkmkkzNfktxLqUzKFFBWnlaU6Tp/jQrZl
Qn2Ec7+meprWicDhHt3IvGDhy7FX4uqUQtmv+sHYFc25OHUQvI/bQui/Kj08dMFJIJ2RZScsI/2b
pT13XFxFK9B/FXS0QFkxGAXtq0qGI/zGffrCpAnNgfkLH1WigE0e9xl1+lCz4P4w2vlWpdE4/dG7
pc0leijzex077H7gmyubl8bpSVdhPWBa9DKgdsK35bqpEgSpn4h8CmO83kL3NCkaSjK+uA6EvVcD
iU/lHe/gYnLC4YDTaldjG4CVMJ/9ZGMFYGk3VrhDbkiDhrw3eh9Q8pafwD1s81z9Ot4qGBAEoWWY
d9+W3r63un6qrmI2EoGrG0JlD+RCz718+8HB3EPCwcvD+YyT7NiMjT/wWJWewnULWFPcIZvz6F5c
gAw7ty/7f7quIUf5QkppuMWBDn18kdkCAlLWIC/UUaIenBLYcEGKbNhLESZ4msRWN0jYOqCnSUNf
5K3+DWAXKLy4oF7CiCg+dKNLlz3fsaJNQqZ5fw2SdS0LwI90aubhqiEjyrMVcGbaU7ouQ4rsadM7
qZpV1EqBXdJrYKHJitVYkhLuGqI18MpuzLaQoJMg0mZubxESgYoQ0L2eoTCsruEjv5O/QGBmQUe0
DobsG6F+BW5qg7MNnTSBZGbAyKCD4MjoxVxgiJcRhHaCWU7EVMy7DUKmP/CG9enjqo6KcdtV13Nl
0N+Jr9dIS0U8pH1HgsLQUwJRPInzEmHOPmTyFMsVlonnqVEoPTlH6W/1ANMJETSBLBYcdgphh0AU
gYI5I415hrovk91d3vnXSw2aWw4cGWaHe/srnHrFzElk3ZbqGycVAyVMAXUcyw6JIKMR0dzw8uQc
PeMe13d+FEIFD6fohdZZ30jV/DHXQFVi8DXbVXIGtnuGrHfuJOp4aNVWg+5i9QpjT8OtZlx3LCpa
f9dOc+LN3oYGCvyRMFJ371NSHzpWoBGVpbqgqcKZwJQY9kEFM8cPeWecy6EZV0WslSLG7a5Nw4YT
A4l6FEWmNu53XmSGCAxA1g2JjzwiWiMPHBMrAP+12BEyMdu6XpLgXJ9wQWSMWsU4znoGAyLmlOJ5
4rii0d0mOxl+N1aTU6EOhdq5/qHgZOJ3K51/jlDx0XZlSiSXfijJRUwmQOBnNntyJ+tASnHHBIMB
KV85EXF7ksNMcRaDDttdETnFYF4amR8oOO7NZjQi6zkIhJ+6YtKoV67Bh0PjwFszbiYHPXPb4LIA
ZWWEr1Yx8Ew+Y6G9MvwD/gWeP4O0sMpgV8WUsaaWqokY4uzGfLDC8BrJqbcrHSCGGNZYGTwIn9Y4
XbuaQ7AIah92Yafvg3/qXNGziQz3ueaQCkEA/+xk1RwkMChYw6uTx/LaMiNlLTqia5envdrCMH29
RbMJxpimiE/IcIrzldZxk5LTA3EkAPmj521AQn4IC/UEOaNV0KwBI9hUmzr607b5k+SIEpJ4Kdiu
P0V6GatFVQogkPIQsY/Qm5rv+U/DV0Yh4vxs6LgPzCskEAuKii+g9ZdiKTyeeyr8xsU8TxGGpwPU
exrowebtNe7D1d7kWXGNL7BKE8Z23cT0OOnIPjUFuPHAK2dDBrTPuPkNh/yERFdcumAjKADq0BF9
IMLX53Ultu2/Q27L/OP5LbkOj0vmtIhVQCq4D428JRo+yyHIyndSrCkKQyjyaYg9zlGEQEnoOTwK
BpIvwLexbTAW6wvdjD1DvTQtY0XUJ4Y6xsy2tz88Q8FHX/CyRMn+TKeJJGv56sd+Qj96aqEraZnN
kPkM/j800cclSm0No9Nf7FViKa+l9W6mpfDxx33KyQtr8I2+X38QtQlQjE/pMSLaMoAR4gwc1rQl
JAZgVhl+Dq9pr3KYCQnHn1yhn8M03A/FuZL3ODlUGuZ48M/CWUYXyjJeyxgYMlawerSah/ELvPiY
8M+sqmNovFJtoP8ozw/XQuQ3tk45a/0NUAjD7ZW6Pt+877pUIMuqS55bgWtLuPxu5sMm3Q44bMEC
QC87/zC7+PdbLqEsOq4iYV6lVm5gzPYz5OdvCwNEeb8dmtBxk9Mswg83xRC4DYfSdt/jN4jtGI/1
ccsMxsVt8v7UtRl96ATIciuzbd9scQkKq1ScLD6v00loowoAXRG6yV0OQ9918FBNOkWebRYuJKFQ
lIa/EcIXDV2oVE07JMSXLCMKDbWaeCfnZtzeoRfvm2cGnVueDCn8pZM3EtiUkpFkYdegKYa4GFML
xsZbLUqSRrZNfD6d1/lN1eepLi642FX9FkV/PRuLp6d5xgTqDBYo+wgkD46E7mZMz/gpYXpURxOg
WJfmZEYmrnHXuV8zuCL1hWw9gk/5DLJouxTPXtXcZG2bODfPDowLtSiIFyPkNgbHh63K//DPdphj
CVnIbuM5y+oBvspFuK2sMI6ggZF8PyWF+ZZue7XnTb6dYesUDyrI71PBOFMXlSVoQMq62qEpDp/Y
n4bIZACdYOBOv6AlHKUADcPiPkYWw1wnZ3vtIU1+BJlLeWLCfzknS2xVNACVn1ASWbrdEqtHswr0
AcAtrZQrF9WtoipyZfD5TRPlHcS7zYJtPNSrR5cjuJDLDrjnuF+vONKHS+h9wqQA4k6xDNyvjq1M
99OR/0mTvSjhNDU7S/wMxiR33HYY/8GsM70kUf2kpgDMLGsHqMjya9WKvxb1VcmaP2j6Tf5dBDvU
/gY/7cjBP7Z1MFUXILsNYNjU/oy4WH0J5DdrfLtfeaZLXEmnuvRMvBiUYkGlJM+9WJPJxGl3s1Uu
MMKqJHnrHCvT9WuLW1Dyw9KH1YoP1VuUOHLAZ3rxZzjBEAauD9RHm3vzwmrzXhkREuuK8/A5rdex
iXCf2tWiU7U9HEU8JD53c3E1jP11OY1KyyOiFE9d0SVEHK3Uo36OaozWHEL20mzxgeUYZHl3caM1
cFMqJ/N4dxNfvdNkiv6WcgMHfoEp1ntzNX0XAx9zg2ADCxTrfwXbekpmJ1SDvCJ5o3KopCuqhjo5
y5nehnvU3U5HRI8qMejYNP1A1eMmJUpmFaL3sFXQ/yw6OkqHu96i3qTjktziW4S+2Y8qT42rW6FH
+imTCjKiJ438Odm9UoMkdzgX3hOFNo8urpKF68HLRNA+Ct1vWGvaAzarQ1Qlyw2iu8NeMRQ7ZILS
T56F02RyzoZKHMnCI16gz8PePhJxX9H+mLAgqRnlO9PecevJTQN1Fk7l9iRiG6WKCMsWu6uFS+bJ
EC4tvW/K7MrdZO7UvIDFaVq8+tHCvsAndY305ZuQ51i+vWAHI1P4/XEn+M2Pm+D3ldrtqiNwL5gL
YKkQ+SW6i/lIAcxOciyob/sKrQCqi3Y2/YWS2e2/UmgfYHoOuvgtNEx2qFoVuJBDb0fj3t/jmCxx
qoiRTAk0BpDCoh9l4WjOQELDT80fXENDaou2IUjOIt5INE57kXSuIczf9kXtxIc+8p636rOUuF6Z
v1kqDaCLIvg041DRhhcPkA5n5gaWipiEc69a6aHm42LaGG3q8lOx3Vg6dQYIgV6UjsXtBSHL2K13
WUyQ3I/dxSyUruqQNTBRNfRjwRIszNUx1nI95kYRmQKlaMLA9FYjg+QIrsz9Z4qsKk8H0vNWZ2lB
+4cIbp11gvEZqBfDam5NHZgNvXEmpObxavH8OO/AmTN+y6vOQNc/s7RuzIyjyt8PiEHuotv5ccoq
6U1QcWRZL61HxtqjZLKcTjJ8ZNt7FiaOKD9L16OXiOnY5jRP/nnBWTgQLrMByHUOFq5G4l9uRIP2
lE8c8ShOgyfHpS/QVzio+AXRjfh/d0HhUymaDs4PHpq/d41qMcGMdrxkSGDMqxKaDo6qJFdOKVsj
lVQmM0qHMXWcLB57z1EWTPOKwvl7B0DS+TePt7R08fhwjAXJCDjyu/TwpWpe87nSHAH38ApnlgoR
A7GHOFKDuk9roy8lThqO8LMINb1N5xqC32821T8jnTTST2UGJqe+rFJb8eodZ81wNUuSh4VIeiyG
/uoFJ+ZJKOiJkj96xXYf9fFOBhT226f4uoeLeht31lIbJtXpyvW0PTAO84yQlziOVo25WkkNMEDo
Iar7jOHdgSU0LQx2WR1sZGUnti8SFO7+8uHVhNK2r1BRqyVcOUoCutBPXO1PMaN7Dg3W6Tg/dsMy
dXliYju6uGa1rJS7MUb81xDfFm5n2Lb/DtnR6A9JMHb9Dc0GIg4pmncuwPFhSxabjKZR5dBSUU89
OhMExdNx2yA0r5yFQ1YXgjXVzGDY8VkK7IMEs70JFC+7SlO4ckXkx9hiYJH9wV1FKHRK3jWqJx5H
ZnBg4dIurz9FirlNC/HMQeB2hJSDtD/QLhhYhiMCmPG1J+invfezky5bK6oM8UfiGcUuSDh07GQo
wxTA7BtNJHeY7OTXy55aToLDo9JX3pPbUjge/uD2QcyFNUecf1eeEY7lCSSnrd8hru1NoLCbWd/5
x/2vreJ4+h/nTAw/MSv+32+BMNdhGy1Q3GsVZ5OwN3kUJGI6a09JUL4J27rZejDGneyn46co0dYP
o1qU1yB7OV9p9OtpTo+QWpE1zkFrlL1Y0WoBq2kLxoyPY3lfYvP/GU19KD3swela3ytf1p3T99Cx
BxwedIU980I5BTLukdP0f9FoRStr25q79PxT3ryoeKaateBW1TAajO6wnAYddOPbRc0S1P3dRULV
dGDsnn+YDNkCtS7qZ37AZCoX2dLGCWNMzWS6m1rJw/u35N6uklZI9Tmm8+kFlhR8MY0uxc4lG9TY
AzgvGGGTg3XoXcq+76Vc8m1ky7iCIjLbQisKrRETZw6T3kdA+lyEOah4iyIII7SwST5OXEFIvYvG
XULxN1HQVGgLDevKS4whU3XyQ9lw0LjYgL/m2fkeuH/pigag6e9/Odp4crMpUKPY9+eVLNMAnTU5
MTc8Ruk9nAbmBRq74VxNmthxlykA6j17lyadhJOZaTIWEj3e6YYI4YcX+VNduJiYkReVqfoiwaT4
sTdleI33iqLAUvcGERYavpT5ZaEL1M+PAOfsnCro8e7OF3KnNnxpu/ODPMNYyZvfzIRrJ9pU2J69
GOOOQUYoi9HxKwGs2T2uEpLOwoDY7X05u+oltMqXW0dE1dDBev0EQc/TSpf0ezF7jV2Adyn99noX
/TqRoOMf9QWRuC4+0fuFhtIwRJMQDTGdQ56TOPUA8u3nRt56rlr/Imr2HaUIAzYJREsTHwd0Zq60
C7NnQ/0pWLsUU+iN36be3BBuxoG9exlxSikUJjh3KSTBE1lS+Efx10CB7KJ3oTT3+KWKbSbbRNH3
msetdNDyQJ2hoMx9MNDQEXg1BeyfSJN6CbA/npQc50it+W0nnbk1D1K2uzcfOWa45SaPnPt+yokf
t6Vn3mScuDWkUvwTmaZH8SoXOXwYMTw0paPV24uS8cb7G3qW8EkGFiRhJmiJ2a0NbFDqPipLSKa9
Uq9/Cfl6CT58iH38XFxIsJVPwfyI3cvaFEWw2DEqt1FuB6Cx/a+6X4VYcauKcrQIVezK6KtgkyCP
aQGZwfVBEmLmN5i6SPqp2UdDKa78L9s5GGTNax11Y5hC5gspUkUYu2mtA2rPP+X8M43g1oLRMWPp
4i+gayFUyPEDH1fRhh+mxp3LDXabiPw1BFMLjoePD6me7jdan0B6wKV71WoQtOlHHxxDwhF82qh0
d8g+Y1+c2Pustt/5C8M7g8AIc30/zBcepDfr9hakXIoMsf2ejFFNGzAABRDPgIbTLaBHRIyOBJcT
9VHz0PSbxxGmlUA8utlgrHTrx3sEXLW+R0olv8IlUedq94N+JFAo7+N34ihf8f7aeluM1VDFkF1v
wF6A2t/zumXXOhizFVe8TH7BB2Bna+pnl8NoWlmot/iWcY4+JCVFVlXXFJM/KOHo848uJWWxXd1K
F32Uf+PmJH58jYBq0CJOY+iw2x10ZiEJmkOvhd386bHJppkePQY97pU+hUJh5ccf+D7LU7f692eF
yjMXWO92i8IBNJx+zP5MNPj5BjVnZlH8IjT0KXDPboV81nwj22wdR1UeYOMZc0erdK4HeXeZfvvc
+767Wnfr9FLjRLXiasErbzVoEWL8eSoTxk1cDDhQ0HG5P5rzPZQNqG0ZQuSCBElrGBbx6SHVtghk
2O6kcHTL3aOZQC7h2TFgJEybbUeFE8uGHVStkWz01Ikhb0w3p1gyNbr5vsfA0Zy+JtXWH0sfc74m
AX2dQdR++XjITmFgzFf+3GeewKZG9ksq6fPOjmwdJcby1YbCzF0mxXtusBHU1I3AijqSNlznKe97
vWv3A+51ZyNjYypkJIxx9hRazc/HiVtmMG9COqj9EbnxDdju77+gykEvuCsjx4mFsRhMaZ21Eo13
lUu5Wran9QEA1Tsm8L7fLXE5BLsDKhdcBVrwZbRb314aQ9nPlboAvKDF0V9dcW3SXIocgObG/5Jm
VvHmyw57JyLVhrUhRvXm5C+qdR9JRrmHu3mZ5jk8AIQD5Na8qtMGdEJGZWmtiKwB6/rWikCLg08w
g9Y8sGLWeRVR0gkoYnxEWh1Digei2NRUKhSLllZgbNL4HOxAMm1p7X5aEUAlOTrtPTK/RIbtGbsY
5zRQ4lVieH55DUVmh0md6KZOW2+5IlXvOpPCGlFugMgD5pUbSaPu4h2wPu2+5ageBkku1NYugCA2
QHWJ8NEHSzgbAHoE0cnotJpr8tdCmjsIA9UvG+ZBp748NZmdxZMjgOMPrCupMnSNg4ZKwwGe3rAl
1ffJyvkCCyenN0MeLThadtGJrMlACeXLeawvIYdHqs1782iGcHiBRDInW8ZBjdttZLmoTsS+7syN
fxmsD04hxsjtdOYnfaxb+/nP53Sh+SIZ/ENcJjSHpwQWjQ2XeIixwkA4jIim46keukWhp6RT49AG
oRccHvX8kM6BsSTb+t1SnUZIEDwNN36KmGTg1OKpWJc3MDzwnYtdHFPElftXyYZHSXrVKjr7kQDX
6h6JMWNybSk3qXqz4WVuLPP9+U81pdYNb+sFY5fqnmkE3youCHMCKkmivmrHFSQuOmeB22CnP6kE
Rd2PZhdebnnH58FvJTomhtk9wFUpNGcRaIY5eztOTDD5WFhsyvjjzKZ7Z2c9oaeMaFC8YHMFVTzu
cXP06L+XddBe34yKsbIKmrL9RikzbYklTlY5J3G6WwDZyf/NFSfbNirD0ilNOOiZ7bUrHI5P9qiB
+ZJPfcsI8olwFvbdfpYsRmUT98SmI2C6npdPPRQeFOkOt7ueA9mLC2EYfexE3Vxd6Rx0KVt7Do32
r4ie9CaZNwJtGPzPqwASAdQxSPEKnYZ7xSCC8sg4s/V36vCVJpA3nZ0fZeteH4/OJm/B3sGht8RP
ehjb6LSa3cHW/ftxz9ap4F2CSg2AdvEMT/EqQVnbiseuAoCNNvhWFVJUSCKGvVFVzShr4z2+bTu1
mgxWS4X5lJizQYlmQOm1HSKegYnrEL8weYQj+UNlwr7XQHBCjMP5JkVit5SrkRkWQwfp11es4RlY
tOYr0Nam+k7et7USXqY3c1jVwJxEtU0fgv1bJ6BU6THEKTNQf9FPgRNYUWjUaBx+7jfGpMtexF4v
6zESfkRbYGiapt2YQg8oQVItJNvI1ENQlMG4K5rAiJbUUKFrsgf2Cru1k60xBKgc7U/mlK9jIDX1
FWFFPWr83r46gSl7bS6t916qGjtOIht4M7IrbJWv0ODM5aUtzrpvP7Tsf6bFRwUvECtzKlJPckSZ
nD0LenWKoLa+0wDZaomRFbYzSWg59kHzy1SCsfjs6TyVOFEny+iDuMdtg7UhsL++zYUPu1YcuPke
7T8qp1attI2H3I5VfmIdUMem+5QsYdmh0/7zrHx9IFPtbQiNsr/5PbIrCFaJaG6qNkThUfuBw2fa
3T4bEh/6vBkWOihNVPAXSEgbk3Kn22KWlXRq5ghXf1LSwkaIaSZ1d6J/hwCe11JYi+K66+h/ZWG8
Ple8OY2MfrnzJB8Dmm/W6RsMgLrvCpF/dUOQcuGj7JQKaKbxQs6EF+PWAV0bxaXszuHdsJP8jM+8
0Sg9oN06m1NA4MDzNVJtAIyeKlK5nIXY+xBPpF2DUAatOaMlkB1Z1+gEfmKqdmtvn7zCcX0q/lRW
KotGtuOp6CYhhZQhNOx+k/nYj0Vr+gsuUlwj04nZIk0eJbZZM7SleZ9bwVFl6T+avcwmpQwxV9bc
N46LvdPu2BDGY4JwRyTAZbugw82PdrD6sxPI3G/wKtSA2wIrxyJ+dVMg3woVp1ZMeKqkYqCo9W1c
PqSgtJ+eGczxn6xHJRsXXof5xdZnf6UKEFzDNT3cKB+qflQGgWsIiY74gaD+CEkprAPvIcciPMrY
TMklzhcyr40aDuaezjLmc9vr/ya4sbhFRjHvrZGf3o6/rB1UOqfrd0sP2Oav+I713DptGVG6Ff23
a+bz+D47MfCeYYX2GyQ31fc1XOai8pt2L2tV35aMr8KK51Jfol8WFThCfcI4jdRkkhvEyKnkS3wk
YW1hFZqyn8B7XwYug3wCxYGgGRjDvrbmNwRi42ZUm31MPYP7h55lIR6Or3WBQ3XcEx/hbr4GjpPj
SDhtYVnYkHLj1k8+4ufz0KugW2YTJ8sAay5HQvhd/ReZP9sePaOoHmcSqV79+ijc88GcTN06+ZJn
H44C1qC+EoxnE5z2m1oj7H7yfhidDby3DxmcONsr2oNT8faRGSfV77w27eOZizyDguxjYBnB3uVR
B7A4nwJnq1SgiozMAqm4rEabh90Sag2JNc5korqeY3oOlIdS0cSqepRdit4drjx2y1WP9okCtQDx
EIzN1LVE5Gb5RnWyvZfxIUZeXvp1IDm7SR0Xs6sieQ7q/RwaE7wnVUjDU7PcRNt//i6iEpnEOY4h
y3s4sCIN52cDJudYaOvQ3uzkZm3Xt2tshP9+lKv8zIebIIMe+88zckcPXpLfA/ZWXQnGbj3C5aBV
UlIdIO4FHHZ20RhUwa8jJENWGCO3Tpp6OAZHxc7aFFyFKEBrGSgeyhEKVYSQ6OURzHA62uIX0MFi
isY20VGwc2DyeFY0BSd4cVrgt7mMsItomQsTgatr/oYTdYC9BZhzEfMGVguuBfaAQK+zeQQWXzgt
A2uS03zJ6jxuyCilcIkPzR+MZB7FZLIwoONYbS7tu2GoQpbrrHBBnUGt5sXNNggtO+t7uwTdLeku
rStlS8f5BdgvrNStx4X/svxn6yRXi2XBY7xzzBrlWjQQu6oo9mneZMo0+TggnIoJFSjr2v4V+gaZ
nMsxMb44OelmIpmkcDqiajvmgq8mQGB4x265vb5MW2pJjwMfpmIHlfcStjNjnqk/rf8YCNn/h+QN
hd6JMpBHpDQd9XyAQmDf6saomu3ikDzDHeDcBaflEziOGFeiY+1wDL4PETNMSauzQT8WcKhACTIF
rKiDZ026qab7fW4GxLMg3GniPCifbbuNDfn7y7xfNw34l7alQ/BVW9MOhlWrI62r4N7Fx8i1SqCp
aA2+P0FA8ahYOzAaCAUWAF+HMLStBL5NibunNy3D7m3Dxi5qnA0SdtKSsdP0ZBcFUCxRcDnk/ttn
WcJyHTZ08c5uUcWWlcAQGkhUM965To9Ymp/49aFunATbig6JK+V7kCjWZu+Xy5tJgepNnt44QuGk
c2QfpIAKXA/RghZyQrcC1eXxJwi2CjgAP2e9OZPLUAATfLAfOdDAtNz5OjoKiqcFiDX9RmsqTbaC
Bb36THAFXol7z2dZkq/WxeAicI981dRTXVKI9QxVH6LbbygI6Dev7v2GzOpsSbPkYfWr03JDX/gW
ghrQgpDQXcFdLBEkfd+Q6dmjQyLJAgw7Ed1UZJCq0LePmpPFQzQm17GmcRTuezNhe6JAaGic58Tc
74BBE+nIAa2Rudm4NajKbq+9IIwBvZsp4uX7nqY93qblHUbmIBZBxgovf0Gw+y+7mjy+84jLgVvb
I0gQS53MHdf+KQwNeyujPMqcLfJW3MVK5QJHS+CYRL1ftohZjakUw09AL7SZIFyKZ0kxWhYLa4hc
Jbn2Culsd7/gVV3i2Q18gzHwKpCfVROnF2cpnSyNCuIJ7y/c/v4yXPb+Dr/KA2Tb5lOiSHaC4+wm
8Cqy+fgIzVJGnV7OkuRh39eNow4OB/sjObvyrPjVLYwkYbuDobjHal+XNPhueC4recihR8268xzX
9VdjYFM/uIYmSR28XgWkb+42hJ4GrALB0JHCQY2+vSEjH9SfriMUe1qaNqqgGH8u4saZvVm2HhFD
l737O5z1YFmGKvaViV2d1i1RP2wRc04k/QyOCmf9UbOA0ZyGH0EUs95c7AIlXxg2KUA9Ferb3Sqb
Cz+4CijEEvMR3e4qIPkaDMtR8ZhTLILXv05nWpqMUlQLoE6BYE1Q0uBBU5yr/jG5gdcrREpUbL3E
sFmKJDyx9gEWVcM8d0fCLay2WE2IEObVGjTAD0Bd5KBCp6c2mKesMJAVBG7Z966VM8Ai+0eOfmQc
RiDPLWW5csuxCDYgOAaij7I6yccE3f32v6pssO2lS3Jwinia7CZUv+ZuA/wLIpm0ziQlGQfsPzlM
FP/746Dd0Is7No34LAxO4cN2YQtLV/ZJGNG+vIv3KgqyxRpNFsLbW5zmYj9sC27nvW+zY2yJrlNb
FlFAXE/ZHhtddZbFKkMfKMXFEb8jJ/C/tGE3NDIJbhCAPB0Ko7w96w7lTjIeR/bnRGV6qWwHwKmm
CnuVGejJS/Z6x8bGR0SEBR0CCchSXe2sNog3qrx9XdsCmKJbq2bIwqDh8Sk4c+/HcmsZ6TLcErp2
tbrT+/sJT5+nH2hXx6nZJwjJamTqyntElb+hDKIi8M1ajbIXl4xEjYD3peT5GqtYaRoUzDS5Mevf
BdKFyVn5TI66DR5020ljbtpQCa3YIIDFQvjx/hU+IDrOcMzNzHC4l+g32NkjZoU9iTtbUXjG1BWF
+PeNooh+VQfvbBsHKmV/5hbNGQsLL9TnsxeBPFC3xQ+E68oDuAGo7ICT0KQRWE/VXxQzMmEpdHwd
rfXyatW3hSaE5U7HHhbP4P2aEaSBTin2vFfxkAq+ponVzoHH3OJ73ZnfDPecmLijnu3I4OeWJAEf
DwiU11vxvFnKG5m2q7wqoV2nFctLDy4I8Xlumge9bTl921+rkp1/GTXYgL2lT5fVs1YA3DRrdf95
izw6ixS7BAjc2qf0q1qOM7mpSx2YgnUNP6A8azSNMEHJJv5ffJrdD3RVXo8mnMMPqAzAR4tmaDhn
VMcVGtqauQNjU2XKPVTHgGJMrdAPMQQzoS8FeZzRJMvjrkQLaEMzyoiU3VgcycB2A7fyGm8BCcl/
mAEjVW4iX6aWN7+6pu3Vvm4vGnTgbwLaCfebE8xfXgU62uyLsQpYwAkbLCpM2lFIfoVi44y+iIIV
cLtKT4s2CNAMGdOux4yYQVNGu0sX0Rmyz2IxMUHfkWcTW0Eyv84GypN2vo8WbXoSAJJfB2urQAI8
CJ9vyozI41C0+GapDpMVmmkpbmEDbyPVt2hpgzoGUYtsw6fnbQu/0DtKs2rvWzHRRGjEvP2TB2Qv
vcTSe5RuMhUmR/jtqyPJHre4mttPkomSPesvf5vJHPhWVqTVs+SbAItldTaJHXPfJRyl5ZyGhsa2
TYfCeD27K+ssfL1nR7V8bnAzn52XISTVEc1uTWvLu6L90V3K8SXtOG1Q2oO/NbsUc5X32UxflGrT
MO/S86hVqEW4TF29ImOit502AKWnVta8m720+hQdY0LX3nZ6OnFAracQC0aGNAiCjsELMikWr0r3
FhDYBSzF3WVvHcysu/go7lM7ZsYlF69+2RfZ/PeVurQ+6dO4oK3Sm5dnduH+VB2BX5ZTz6KPPW19
9O9JJ2IuzVMi3ufzdS50jSGM5cais844gMfblHAb5CjdS8BfhW7cwVjGJI21M9i7q8k6cyhvUyxy
o/38atmHISS4LJpiarfbd3Y4iUzJiELk8bC3z/+TnHcG7TDwIU1iQjdOqChKDCe/XLHWRbp/A0jR
5zRanJv09Rq96ZqW68uo+zaonEAAJBLUeXV2Ece3cnk2l9FJ8B7jz1wf8iiRDNns+NgKjpofy5gd
KUMrq2+pdqZKQmY2g1AbkzqzgKKhbM9247QE8/373oBMmUL8e8+8Kgr3+Gbvo6Kvw0yn83QNZI+u
VCAiu+RHsA7xSz+1lQA/anPpzmOviD4vvc9BQb4hvcIolskuWkFD3DvkRQIMBHxt+a76WyV71SZy
+BcrMUzecmROKB1heNXIsQ5kn7CJWBwQYVQZc624aGt8HjsNj7r5/fUTIPau393KQXuTZuZdkPKo
tvguNZPCfIZEhZU1XMKBTVBABGCWIAH/bxsXHtB3Ls6j6j0FbKbCS5Q+FEW6nmnnrVg+tD1Dj0A+
xplsaqCyR+eFJBBE4q26jLqxpWDILUSHtkBGzyPmgKLD+SaucA3DBlUVvXpMMX2OBj8FObU/Xxau
KZaFzLusbW40g6Ro4PciGjnZ0b/SKgZcXykDPRLuikTHrq8UxmsyPdjLpYJdiDJ7dW0/9NjJSru3
WZc+QskvOzQUhj7YysO8EDkYBPCsa237y1gIlHUNvTvemcl5bIqg59mSA64Nvhx/BZoL9/TgZreR
IBqf3RATNJTZjKKb0PXvntNre24YMxqFcSPoBHeXVqMYqVlPxvzPGH0thHT0weSvmqoigP9NirOo
ZskKRdCOsOgaqSrgglN6RwYyF1bElp+Ju/cripFVu90y5ssu73536IcMY8O0uTejTAt1pqzeicVF
Gr3r9BFeWweRmmm0dvghAFFBj9xdFRglAGvdAQ5ydBibMqur5rSqNe7J1nDg0oUDjJYzrv5nBcVc
SVQCszBd7GDpO8ly2TGYGzf0sJNjqeH5rNHRi3NZG2f1DGLGGwD5G+1PmhHwcnXrJvI5SPuWe5ZB
24HCvDg9S6uR5l13rGtSD+7JQWTOmSQtBlJb0KCRgvaNglcPmuu71zEkLr95LW2ebvupLQj4s3U8
RwbqkpCGhZpOBRNYCZAkJm5RkZpxPI0jMFedaZqBHI0wWnib7A73v9q7rmnSzv1OhyCWNzWdvrdF
b15aD/1F6l8fjFlTD3LNOJJSoCV/pebA8SvoEzahRk7rBb6YSG2dZ8u2rzoZGRHSbCKK+fLao/Nn
LHKJZz3Om9tyP1VBrtmsgK+pqmdjqUEX0YzQIANJqQ0P7I/a28Kh3LX0sgSTkPkwXT0z8OMaeP2Y
uEmQxnTwkhK09mwCnNf2BSYbymfOVGMBbDjUgJFqvhfy4b56iU0jkNbB3fkxaEFkxVgbMaVLRXFJ
3cA58snGgGpscndgGk11yAC5Ww0GnnBwul1K/I3u6vbZdzASjmrFRIZGESHE8sjqoCYTR9n0IWit
hIMJQviVPV7syQ1aju0zJEwH1807gCqqbBN1zTCP8CjQ6+/7wSw7dwevrBQqSEijgHa6QKVD8Dt1
RUu8rx7fPFFwmLEq5AM4nHIbM45cdYCDccvBH5jlcBZiGJv4crnBISl22OREM3OOotXmY8GCQTcd
zGufvbYD+x29KYg7yiV+0513jKwQpWK3VykukC8wVGw4gQQ/lNVAq+OpCS2CRsUuelc99jFXiEqx
G55Hx350+0lxmPQE//zoSSLe0qmvlF0q+1Tv3djxPA3oo+nuEuoY4hgW+euC9Dg7WqDwFbPjs0Uv
vyvziKLp6XSOD4RYxBXb0E5nDTkJAutJMRdmBD9VR50f075XSzE689W9Qp9a6fINSHjzwe/ryqVV
NXK5aqFjQwm9e74WU5MOq2Jx/U1gZ79Eo9vR2+RZRL+hDPBqOlbK/msnu669DOP1laGA1JE89ubu
D0M9zRgQmXqwvmZr+Bv7suIqOepW7tc2IyfO3KyNUlfmpCgJFoszdIkuJuoBPO2Te5g1cybgDtEu
6FtASvbNfJLefYSp9tLlEGA97+TBLYYnv847zzL+eqH8N2V+mTKWYbQrDPn86lQjaz0n0bR6oOon
jn2ESgtxgqCbC9PS17BJJk10gsR6DSWkUFdHXgUgk7QBvv8UB4zRKf3lpSq5yxQUAy1KCdvlUFrl
DY3Gw61oGqt4hHM4dA1LTDL1Q4xtsE+5tVSTq8s2TfJ5FGU/dlbJuWGyUe5V6skwgLfiYGAbfy80
HxAYEVLVic+Th6gndAP+cA8Kt6M9TZuxxoYfaJB+BeVzH6WSP1AxTX4aIEd38wqQXaJavAAB595N
07PVOQyWGBhBNKiZ0JXZr3K+i9sqBbHeo3HC2Wban29DJeJSBYuHz2xS2j7nB2BsCCWIDnQMieog
hS2SptjqqjzvW6w/bvB8+QXFpQnea+z6aAXZWEGFCjKzM/GjgaAW+Zrl4akeL7fQJofzUtN8w0Mv
vFrvgwW0ac16JvLUG0KM3SRYH6uiVWI7WSTLb1eRnPmr5xuPsBtIY8BAeFyZV1QGEkyeiGd0kXoB
mhvFrbL2yAf/nHvX3+WkNrNJ4/DfPWaLbANqxgP0ElPe3UKKSlFUbbWWjm7Y4E4PiznHlZKkDxFH
kPCyR5jS9emB9rCvJWPa/diocfyEZc5/k9HxvzZVLTxcnnlP+FllBNdgDBqoWkGPd5zZTOwteHD6
3No1RIYFySwlNaVFolBmATeqcsCN4C8yo140jrXrsQusE9uhD4FL5vCBaCS97FifLdOk8EmXaERU
xesJJWSgZ4c5tBqWXCNfDZBAoWokbTEIVl5jR+u/Fz/PDbOX/9NDEeaG/zunB45xIijHeezV0jxA
C5s8VQZ+5OG7lGV4cXDpCAguHmjUnUAJ4OMe0q1hnPoJUJxsMiyQOYv7QBBiqYM9dkSyAydbZ626
rgvqp/riKGPTxPtKFVVLoeisRVLpgpqTU0f3tMCWjMsSgKJsEpTZiGLEO5DwI/UgpZSg0OCajxeI
0zLQmSoNbiNeNVMxYTce7XATkoTTjWTjkkFokIoKSPRyx0srOFxBKLAI+JMKpH6ECQ8zUOJX2g0s
A3u8jb454LrlKIU3gisa7pJ3vpNL1DwwH4A9FyLV3z8TeUg0qFX1h+XNX7BcJVW668AdsxGLfk6A
GNweWdi6yneLW490J9FtQ1GLNeztDBRRWnv4tP0MdlnlspseHgvG65GLTCV0i71diNCKHZyjmTHN
QH75BD2j4CPd210cVHjBMB0NQheqh8ymHMRbfvHHP490PL0Km/uD04sy9Hcapj995UYIbXN+8H7X
FBxHAtM3DBkqKSegqroSQzNpJIjR+L/z3oIbztriyGkK7Vy9XsxV9aWFpDaRLZN3X2ek0tk4cpSU
Fl2sHykKPEZBlEw1DTSV3B35gjW2uUE/laqr1IQglh/wibh8BDEN8PIgpgsHQ3DbYIhm9HN7Uh1l
t1UALCXdC40MEbZiAw8qZbcNPJLm+Qmshrh8+WVIoqUT/kSSVK7sGnGu/bZULaHhSFCqUQPXNAAa
cCiGJvgVDfSbWk+20TltDC5WiOSDnT6GSK4EjYdTs+6i5EQpnFwnwtNLTlhn6L+NB15Qmg3mI78U
5yk4OGIJSj7pPF5cdIfLQGY4G9K3xrg7eW/9drt1Qf5d5YkuwMuEmVCA1jLQzqjJGXtM3nImZHLm
J9nXGvx8/1/Z7d9TVtvXgYZLCqF+TYf3GR79UC3CFtpbm8zvCIfD2jScVRQOV1aOTFYQtqk3bFh/
2qnYLfDfE78/eT3FVJbSEBwSNlr+qQIx7bRkQ2a2uXwU6ddZKcfTcLZJResb8hrnn6WaOKbv/AVo
MmdOS7YkJA7Co6DiBdrg5q5gHDwWJUZinxAHBGAfsxi12Yjf0Sv84rhQjwWp0KPBzTteRpHZrhga
BT5kag/WJLtlXkZb27TndtosRzE5LVOEkMNhT9jWZr0XOhKwSl9L/e/rddT5b89L1TaeTqRB6Xjq
fF8xE1a0uarFjDrWdlkU5VP4Y1xkvAPACTL4EY8YU6dp23n4/cd7cyqRwVBnUUQ8PB0J4xolUflW
JyRSqZKBe90wuXzdgIriTCqwboR8xOEa6gDBjgcUGwj5TlNGJ1CtzdV083FqdtmO/A6E6So7yt9w
wV46CmuxrnjgT6+k8lGDd/xt3L/udK8EPLF8wWxZjMsSeDexBpH1dgsOf5xXzK3VhF0WrV3fEvBL
9f0WURzLvJ1TBv34VPVx2iBhEhCxsOy/fXL+Qp551b6h9T5/gBU6wzT3XJXCJpbweoyk+dMSaJ4d
x/9Wh12dqqMqZOnwn5y4AZ5w0FwKkPSOwOerun2aUhuTvze7PmTGcO+ws7B+6zm6V5L2bcbL/U5d
g9+Fy1Lml3/v2Pa5Cti8hB3e7viu9ebZRkuovRcqNW05My8Qfy0EZS0s8k1UZihjxgiFFKlbLMpa
QeiKa78fUsv1pXV9kK6R4/cYxgN7LBZlX3LZLWupVdLMsf0WugvZGS5yBu9flf7Ev7AwZ5TsqlXF
7MkbiPQ9YCKMHM41kuUinKEAEnLddu0f+2VVZ104RSTa+tyDjP4sDrD0ZkXaJR0uTNF/QF5k0vbb
xVJjo95XzBIyWe7ZVsr+bOgJKqCyQ/08zw4ZgTXx/c8SEwCDg2WLyrJIbQKKsFdCjvP7NT9/8NWY
xLTe7eJNTgrd9KmQOyrZEfxgwYXGiKQb33T+ugeagY4w0imDV8hd18Fb3bszhN17I2EUZ73/l2FS
2tB0gHWcUTiF8enP7p/xoatyjizh/LzabMWME/LHOgFrRLS76DIUOMiYyy0uMbS83fvbtVIKNAKx
drW88oHJZBNX4BgAdTG/dz+s9CrjWj0epvy5NGV371wDhzpmh7r25szeIHk1tGo+utKd0n60VxtG
VATTunuhlZSg/0RpbX8yH2fzeNgbad52jLiJNilLah78EvYzvRX2SqEEbo7BM50yeVnMDsjjAtkV
ZSAY1x1dCcz2ZT3Lz8AJ6UaPFfpDC/8rdoHTcja6icXe/neSVF4jGUNLSJWQ1xM7Ve6YvBQp+igm
7H+iRan7d6nwl7lwmETx2xmQVHUTN9Q8GNQ1NwszkxUm7VJuUp0f3zmzMMgDhZskSw/CWq8ql1TT
wC3VCiG1Vdu0wOh8qCpT1+XZqYYuclbo9LKe1adddggr+ENQKXPI2p//gmoOcBU4oMMl4zNKI1vN
pjjdNhFawmPsJKwXD75V7vqzFUH5QUWi5z3DlEqG0tPRxJPnOMmKHm/VQeOTICs52t7MzkmXb/6m
5CWBIM+FygqpXGKV37oM4fAQu40AGWxUNIz8RGy7PyOH5oUovvLdW/qNGdjHZ3R1hfOR16NphwGr
9COd1dj19BK+B941xDDz33m/JyEQogXm0oW8KrcmhG0QWlNFU0kZtKfUdvhVGyZ6uZOxC+philU1
FwaEJ4H6EtUrzEeQoim4JD6uNI4w3v547Kgfcfuf/LIY5BndVex8NrsLUPO4lwiNNxZSn8yf6t1Y
B2YerZsJVBUNWOXRk6MwC8WXo7vXv42Cbag7tQxbBGwaNVbGsq8wCSDRmQE1J7AQ5R8MQVchOAgB
GFuHm/xMRzeyPk3IqjySS+Ji/ZO+xpUwgNub04PEhzAP1wyfH+OF7k1hUeji1nkcj4ZlBe0Tf4f5
ZtFCUO2V23tckfQno3HhKiQ0zbQizkTRawcEGfYmEqSuhax4UePjc6ijy4xrbNhfyFKp8MoW4RY5
Jdgy7Tk48JHmdvbhd2kZPhhoEdjyQ2iUpNt4xOffzL2npO65wFi3jqicBrdn6esYJtWJLUgDV47w
SnFNhMQCV2lyK3NMq+9Gv3+RY+n1z08nn1PkozOyMxHmnWA6DrUSRV+5kn/vIR9B9X3KtiYNQAY+
n1LcRtn+e2k+ZGcvTjdFy7DDKGk6UA1QwnOc+2slcufIKnQ2lJ4kCp1ppCmJ5ZgwYg6oVZqNsgI/
o5BBaD+yNT6qL09GR6ilb5qwlSeLDx99Z1ssu2kJLsnXcyc7Pi2570k9uejhwlBb/RUs53a8eMOR
oiGY90/Pxz03Iqi01vZbHIBdOgscUYh7ZZ0bmje9Nhm+lm+E/h9J/pOyCYJdDcQLyxkioZmxoqXj
q5X4bnXYq4yApj5inoHiF5EIcO/Z/yRdAar4eYsoAeZ9/y+cnMw1RI2LCIGpdNDR21GN6ZEboPE4
OL+79NHutuuQNetY0cnpdmZmz4bBiUahJTL9ypH2JCaLqVEXWToZq69Vm1K4vH84G4kDBjqihz2D
bnYxLW1WlInjn2cmV3uT+hLaV1gCDUNFY5ttKlGTIyPXGWIG9BQ6H5wJGshQbmPuCQz880wFO5O7
Z3Fe1jJolfFRrXGEiLJzK1gc9vIQxUIzRjoNLAqPIqgTvW7q/0BfCK3a+vp7UvOQqOUDjUzelnz1
X34em9V7VztjZsJ2tAq+UpUY8HD+t8zGH5ymlDDwgBEYTBtBtGClzt4MqUfAKo3YulCNsdzW1XSq
F7IG8vb2x6mAlkpuAvuIdWE2BrCiBMEWi7owRLZdb6oRF0xxAks6+yxp8OGsUD0ukR7g4ff1Uw5R
m4H0oJ5QdmOuVIituxeEXMlyZFvbzDBBphHH9jI9xwje1nyEOIegPkEZDsa4cvZEHAUIIEslW2qi
OhjaY0gSdHUVfsL4reZG0cDusEFerRmuip+j66BWh4LBmLxINN9iufEnw+3LlLgRVP0yxlgaLesP
cmdf5vAhgiSMqe7V665Zl+qcoPE0UokjJkS2bxIwNuEWUY8bzDC7Smmcvjf3qfzMmCS4tAHG6JlY
+Pp525nPu/Tf9jobYaw2omFWDP4aKcZV6+8QESn2AjCByTrp2Ym8dt4X4FGf4HAxrEDEOl8hV/gG
31Lk9IWcw+eyel4CYOH5bakYjkQzaSKAU/ZPmyDIJokw9hVtm/6HtuDLYCR0Z/6f/d2E1JfnUj77
zLn1ZnBgeceneGKwS7Vt/xFLgTRubCa9/KHOScHn4enF3cfhmhN60+uwkXwrXED3SpOQ6lLRc+yE
XNRKnAcsMQUapbQxgcZM9m4RHRhog0xZZbYg9UkLNQFbC+Mm3LmqCoyeyKQ13mSV9AcsUL3WjyKl
z9SfWb6NI0laAEv07eukOceUUXWFciZTmiIIbKZ0PXf26mv26Q/65HiVF0oRfGnBo0QlQPnS277K
0KLskeKBjCXxWEXU3+oxUuxJrCLKOvy+krFDMdQU11wvTxA+ER8tdh+AoR1RQcvu7ckCzRyTiCDa
udiUDYSpveH+gU7Bkp1cHPx5hNTUwU/5zCAVB38m562X73W+woWjanssdbzvDAejTuz7eFbrllAd
bAISj0ChBylcOQdWPXYsZl7sGvn9lsrCDUawkuhhhUpAd8zFFk1RJFdpb8G7t7T8gJf8BhHFkDJu
DZ2xYGhwqlAPZdLoq/aVi8PFlTI8YVo1WbJhFNozpOZowMCkszOIfQceA7r2fGm6SZfx0Qi7IM32
URaFbloe+tkfrSYT6mKw7gz0sFKKODs3/23P/H1EnmRVqAz2kkRaiVUbDhxaY8k9gmMKGZwnQ0a3
ZDeKMudn6HSXoSppB9RpypHD6HevlLvNxxA0UF3fHRomVip40p3DGvJQ/EHPfIzcEFPzFZZHTZsk
FeKSa/W0aBjkiKWGXWH1qulZYnHR8tnjaXjpRpaxYHWMfb3xulfqulssqvC3rmlTaRn3ltjDGMF+
lueD/WBI1MbUtsdLM32OBUX4Nps9JJFeDp6nsD0qrF+rlQGMsXvWIYcsg5S3iv7fIIQfP/vOnAby
vvKQFUcQZpn+H/0HhAfqIES7jB5s2Y0/3hb30AEGvm3Ifrvc6dYV+AcTEGsLj5z/3osh2VzgjdcE
Q9XthD3BUAcOnDIGGbTjvH8h9A/aKIi2WwEemlfoM3lwFQEF4sIL7krYjTukhTjpjrngQ8CdWB3H
aTiZD7k3/l6OVlmLPkZqHZDr50AnXUf+lhO58+cFp1xBRComLmriAnkmHwMFxSFxAqLHFscwy73u
35cm+2k7t8KaS+SoRftJ258agNqv/wiuexJ+kRDa/wuxN0BOssfJ2MmTDieUI4FBzbOco2gS5rbn
3Dyjw6wzCVTJDdJ6uBQu4m/d9PKGukAYlW19BqrcqfIDXdh7/Qtj0p58qd1ECiojbLxi3fNm9AsQ
lfbnz2AU+dN7bcGM+SOIuyeJE1UMUG+C56+oK1oKWGNAIon2Tgej3GZ+mxORn3Y41cYaohgDCJ3A
lnvsb/x6aVtsL31Q7yTfPRiuBlY9faKCZOdj1EFN82xhLf0IyCsh4JWpGQCALjn1hMXZfUzhtiRb
HfSpXegAJPYBfp1WQ37tvgvETyRt5dErpAB9M0AM+CBgi3/pTnPOkkfFKwTAW4OxM+mYKZSY1LVj
I/tDQzMUbJuzvFVC1XXWDfAVTU7jfLyTnw280PHFFVA6gZgx2+aMfhIePPjg/FqOBoeM4X7JKBg1
J09se4Jxrj/moeknSUpd7mZGafQYYqaSVPHH8w7fnrwzCIR5yLDjNOLJpy+34Te6a4tiE3fR6r1j
SI9b8LCqtwxlsMailbLB4g6qnDjNOJ+Bk4SI4q8IOnjWtvlqoK70+7Q4YkGDjPmF7lIE1sP37R+i
NiYJ5z3eCf/AJJ/bg+KNDetd9lSoRbUaOKnR1U0wWBj2VRsdS26vHuqCoM2HmTwfuNTU1GazzFlI
mjrQNFUDDHNuiNEkdpLrRpDO835LvJ/L1RYRcWCMhPnPuPscMIrxgs9hc/sDtPZ3DY8ex9V/DDIa
p6M0saga9Fc58BjaJ0nMsxjBndy5hjK1r4wQ+8KIQcWMss71K2lTEazyYoIUQ80v9MFPI3EuSdi6
tVBZCvDKfPtr5YVdB/I77wMRMFl+wmZ8XzX+eoATSBtwScH+gto50dkWMNJIGcCvLZg7g1nPOMU2
wH9pbHFxLr3UixDBnZnnsHbXrsudu+fzEtw7CF71IluYRmwa3WTI2vj6x4UacUjsl9XogjrUJFFD
3myVAh2LAXDffmRmv8Z6IRdrIrTNR7ni91dgc4PdzTO+65mPw1qydZo8bQJS6PauF0skiOWYg2wz
pD3MySd+8T0Z6/SKiZiSFTRp+KMMq19koSzlGl2tPX2ssjJ9GO1Can5OPMBmkyp5bSqjKPFbc7Xi
ZezIXyFrvMZ7iTMe2VHOPGqQ82d1mPCk4nfz3OVG85DazXWHlK+vVT6OIPRLkho8lJcWjZcmthqJ
3W8LS9aIA7v9FU81QaBKzo/pxNA4NzT0DjKdVmRdFi6MlYHlYzkd98/2HESz393xO4oC46riR/sb
cn1Ag5OpSsl/3arLnoF9EHv4MMFX3So1DOBGVM6mueqxi0RhsGgt8RTM2FQtOXtrXpknlR7Wb50W
MDmm/rhl/6cjXXkTSa7NRfk9D+HTBGoU7Sf28gdMNA9iP/9upu3jL6o8yevHcFFKCijpiWvgvL4Y
nBgwvprdzy49RP9r9KVyGyXYWwDnTo4UPyV/hZkwo790h/Zr6+fzSVGjx0U6Uqa6rtWF1vwZXe1E
4aYm/Jgv8YqWYNAuJPNWc8c4JacWBRoLIK5g75+EeJOD0syVjQ4Xi4G7dbUAXRkPFLeRpd+Sd1p5
Xakb7hiM/kC5QKRItxV0FR37IU5RrXNCNOswiWR3wvQgludX/Veau+q2PnwANOjiIZxtL7QwxyAd
gEB5BpXee3cPnBzstvZCcGX4Lk7wEIAz/wIhjvt0P8v5FkkqyvjjKhHrtFEZxN4wq9EIe9BnGbej
A4tpA0w6S7HtLSDOKVrDQFZW+5DvanEoDVgBboeKZHO6pRT+roJlFGQqXBTtebYxIuopCLoFEswB
1JKvVtK5VAeIOewjxGLLZfgVeKl3wQwaZZchQaR+cWe6UXdLNOIY7aUZ0QwbDECEkQWbktYv7hmj
g08Fa01X5dfwhGN8TSG4By7wrrbTO8Dfma+ldfwIMbbEgUh+KoGesY3r5G/yrtq/jlz+CKI78S8+
NkaW/xCCvOeNyn2cRcukuy07dPTQ/W3abJ61TcBPoc9m1Cc/B9smSp1DwRFlosWPSam6C7ttJuCH
hdKHvcmqxH5Pau3t7P/10z1Qjgo1t7ksBBTfKYhVjzTjE7pxDIkv/2fRkn1g18Yi9pe0st+aVC4T
kZu6AY4PSTr9xeh3L4osZiEyPAu0asTi3cqVkHa0xQ4y00bijDZE8zsHq/t7KuC1uxQy1XlLgWMu
yeOklJUjbHV4drhcouzpWu6bYvh3KmTfS22VOcZ3ult2UrTWAwcvlHX4/9KugWZaw4qTqyhPieka
ss/Ynu+4BWRwrENWSjSlQdIxWu/bo4C/HyApqUgAEiT6Nwzln4vabe3u/OvcvPwOZeVcwGax4G+/
DyRS2/sb8qD74b0bziBwnVfLQ+kMGDcYD6NBgWz3V84OgyT5zLyCNMPH3C/rhybYJo2hcscrJfc+
hMWkpM9rkUtAhk8BhtGi4XNI4RYvnIJXwMGMgpXXJL/cMH2+hdSTkMyoHiwCDAJHEhTovrYSAQ8O
HPptTH8U5WgvQ1pqbXJAtiidAERd/lJnXHRm9WDmfEpL6LKfBznVSLR7hK/rctacOz29fJcUapOV
PsczJMPeY1V9eIoUmZTN/ArsUxR05k7sNVnQ2rht2oNa4S/zMUynynNh5HyNOzt6aHhHaFhXng9/
lUh555I9kKuUUVDLOHCvIpnOVnnq/7g7Q2phKvD8zSVHx3oa+2miHl4yKAJ2AukafDmUnrw89Yz/
nFOZjHJQsp09so9wa3namRmRaPPBAG5YQGlk3C/OSwp8kzcqQtt27G6dcXGM9FeDiSbTNnjUyvO/
yiMXjk8MT7/6eSQNV4s8dMyrADDb3AHlwF5tcntfEhQj1lBQ1TgIW/iN+RwnXf95ubfx3slinHha
eJRQJ6CBmr9oaJ6AYkry3lWTRiDzh+UXDiUs37OpsFC4EizlgpSiBQoVBJWMX5t85xZYB1akQEQ4
aqcnbkgmZ1Bxfs+5EiB0dt8DVXZq4ejJIiNBy6S3UHiifHSnJ1X5v7opczninV/IzihEtChoQvxO
urbtqd6RMWgZq/Cwl55WhGgQFUS6fojN9PtCE/x0Bsu2Y3Gg/eAgbxjpIP0LNdTb4w5kwvYGmYEv
ME+i9fTThKpfQX0kgNTAJR11pO/6g7U9i+1RmIeHHdsWgZp/KRnmlu1iWsREwtUxFb74g1QBQe4r
skQ+igEsZgmiuXrpulqh5wQ40GjjQ4mVf3/djYboEXxLBcwDzG/Yjw4kR987D8T+KicUlh+a2YOk
DphDUCS9v1N6r3CHrTthu8pZtmrLxpv3tXYCm94nUhoFDBrEg466mF0jAz0zn8MKejZ8uHO0iH44
N420d5uBkMDQ0Onl4MCRmAz4v0c/JpkPVuwFOdDgqs/Yr7H+q8u7NtAU9WEbTwNSy4rY9m6DnD8J
V7FTBfQBRW94S7vat2CMBfry/47IA0y/plSuBfbFfrvueGyEg3DSrDOV+gyfb/Ya3oV6wWhNR+4a
MZ8dk3kq5WNh6W6+nvFRLwSsIjqwxMInRQlpY6SJ0jNiYrXYeV/7drSx8g94mYhOUh9S49KY+zUp
zEXSIlkyLlJBMDEPmoh/l7iUcUL07q1QJZxpBSFYJcBtEP3AAMveQFWrxHVahpFpsCj7wIMYheFQ
EMh83RUxM7B3UcDmav7ipU2Bo/WvdmPX5dlGIa34bCwa4WJrmVFlqxdatX9ggMSOsFDhuEkDHC2C
XxT5KfZJKxW297CUWE8GydLOoEpAFs1q1nnf5+XeWKU5h94GypKHdSI1QSaYdgVs4lbjZZGd08Ib
kbobQjNhe8ZHf/1z5jZ8K4XP5L51vwSVL0phzfBm//4w5EG1DSxijXPCgBz96qqDgAWLmS1DshUZ
TjXTPQxg8HIIahOZ0Q/uUSoTI6OwiDnlKoaYTjikulWvhFY/EeTwdnyNb30RE5FzvCMOHL6mKJfa
9D32tXx2bWL9sgm+l3KHDcGRet58/Vh46YhFPMRN3y/PE/J6F1/6Hj/Nng4gppoBG40tubXArovg
KPQ5IWmxfEZAEbZDFIIlP0S3h4ET5+AXXJ3zojG7dYtF8RaQhCBFOkst3aWMSrJr0rAe9Hl3Q3l2
q/ES2tkVyDqwd9wHp1sVhac1zcvvNjEW1SOpLLNWDtJFCfdtlxBz/5KSyntP2ZlTcE7X1cPACsHE
kEnGE6rxV6el+49S1BC7LHRohrqVCwGsU+jrocvn5ApCi5Hk02vGeMMcx2lfNY1Z6Ge1zBwZcS9i
CdBYql+8uoL1Ck6a5nR96z6B2SkvGqxXVUdmw5KilW+wmtnf6BDn9gofE6FSa0Cu2QeHzGb58Res
bQqln/gfKDpTS3MILz18TEoluw0vYj1eLmss1ZkfqUbYvXP1pfSZM4OGF/hcDC897RpLXZEmyRCU
E0O30veAIkBc5Re6qLK2SJzIMl09D67mYSV4E0D44ZOos9dr2FYEhMH7YfTiEOo1AqEODKW1dbYc
zfXhx5ZSmdvwcTdQe8iM4MKX48e6pCuAIiBoUiibqxrQWYZg4x8k3td5JvtxprBLNRsmEJk80P4s
vOTyBZzMiTkKdc4darnW4sdYpAFgX8AaL+J7E664+h3DPked9MQXtNweL2vFxKa5An/MoBXRlich
BI7/djcdMJv0SSOvMYx7XJBXXtvishrxfz5hFZGeaaUZDVKaZ7oiNLc9c/zdJlMKKKATTg1Wf7LI
uMQcwTG63p2cAEVPhOd6YyEFMpaYz3qB0xWPOz0ycBa8/JyBdqo2e1bFh/Nh84ldOyBL9c0OK64K
AOwk0VdK3cNOTnMC7atnW/3y+++Uuf8nzfxTPG6NSeCyFAa0VALIyzjV0xQJsx74qxNXNsxTAh8M
Bp3XJ+1EApsZC+CbuJG0+wW0YKBbUyUC08vmUYRTlDehrgpt3c6lFBdSDf0kzoU9x50FuexVL9dL
nWP4qXFVrjYBp3RBdSKDvD8CiOJQwyR9PWE10gEF262H3543W/rxX762bN+MP67vSDOq04rebJNR
ixjS1VwKV7I2yb6vQeYB1EwWcpdgKsJOrB9KO/f0n29sPG98+IHtjcLdoZwU2CwMokNjCirEpdsf
iGrs2AiMPSNpqE9KtvE83wcWrKnv/KDlFFsMqvmTxcgpbPTbm00BEF38UCdujDZNU2+mJI5xdbTv
uu3FmG9ubJyEYkwBAYQ4gzMSpEfpoipMflA0HAPA6xvFyGuCwQuvmEg0zDSLRNlqf/3gKjP0VqAE
cw/vMeZIZcgKpzwcqBH6id75Ustbma3iHDOK8GPzat+Jjm9wKcpljze7GcBw0b2xYUM2i0SrlGd/
1y094EI5jW7sg2urA0EQd9CT2js/pI7KIaDfUeBRYv0j1ABMD75QtelZCf2HYkTldWry09g308CH
KSaxzr8oy9hpdbGwcrRdkH2LI+NHMX5cZYgu62pllydOjLba2ZM/wUDykcmul5SVYQGqROeNseTD
0cFDxxUTyhFPO4fKsB1wkzPtZ1X5/lGUmyZTav9yF98xOWM539dL3wWU4HfB03eEJDBE767zYI4g
WUdiiG34Nc5woU3oIWM25Pqnro+IlBTJf7tYUl5d1owv2v7SYCHNvh5Crt02nz42dReNXjDD5Jee
+IbL2Uma5Wue3i0w5D+hgihOJiZfX2niD3jQ1ATh1jee8ZjYR31oUP0Gdxt5fQn5qdIr/nZ/BtYK
ol1128urvOLkTumhjMeZQK6cPqRfRMOHFtLKn6kHZkrKWpB+6E2RdO+Lj1TWyFtLSa59LAQaQv6M
aMgZl5dnw2Jg/nTEivGcOdC1ORaHTiFlXoMEH42NwBtdHRM7rxDKNo0HSwcIff/4JDA9lmMCatIN
RCHB3xmGTyev/qUcWnEF9w3EKXuEb00ZAqWH9UJHnG85WnHz4SKRXXhcAV9Ajp9ahZd1F72v+d76
WcBMc5gr18CPwWskn+hWSZTG1zedOqkbsbweJKWKhezOaqIb9mI4Fy8iOUnegVwo7/KFVwfRn+Ru
6Ii0qeCtx2SeTA8pLVIs7ca9dTPMF/0IU0MpY+gurYLjn3iQQ3Esm2+co3zwm1Np8+xZHJlucu4V
ZdfcRGCQsizWNz3Vz4wih1cRsaY7Xpt22B0vV75lSWqz0TG5ByBmTdh2qePgAmqPu6uANFh9NuQr
ucKfpKyvn/2WSS/IB3f5YKpnpa26hGsCR4NaMY090E3HIT0Pl5SxS/+scfoWiH+fpRFW+49+mKh+
/wH8G2bhrUhfaLnhPaFSud7H08xD2V7G5evlrWlRYNF6tsF+qfs76vPLouwfNpy399Ka2lTAnQFp
RdebFiDmFtxuCfaVulRlEdoTrPq0hbmCGps/+ucYc/vZzKkcJbkli19Q6SXkaPMu8CWgCA0WHjdP
mCK3F39NMrSLvS3JcGNp28Fw1KGnDPg/h/1bJ/nk33BVdKUh00cvD1qUruYZjXZQkp6CfWS/mmqg
hzODPUWnycDA50lU8aF4iMevXCTveEI3PShc84r1ue1JCHSsk0y+ZU1i1bYZr8hMTCNWSmeZTkMv
lBdseOruFM4PiZ4hce40c6q2dxjjnvvK7nggq83/XPqTFDO6DKwES+QE8I06HiFB3ZhHoH2S+Php
+YuRSLe2mPPnUYr+iem1/gw/h4inJBE75q6oqwFz8pUsz+TisO16JyhxXpQ4t/NF7eQa0K6fm0g0
72z0bI0DWZJkfAGzgppMvfz2BENnq4BziPu+HcoG0wn7bhzAT7rv2Gf19OLAq9MsGF1RwjjozcYm
DFeuwAe+3nOwgLUq/6zTzucg/J4kvw9RVW0cQz8EttUsH4UdBPL9BCini/5AvHw/QxWazkcpFKCD
wqBF2T/3pmbJ2U0LiA/sFRM1H1uufg7avJUahCPDUO1ccF8niRFN2+zrtEgjhAYk+jwXWml2GfBb
vlyAZnUXJGM7o9dwnSNkcsMQC5MyOTjsLomE7mY0isbKsLfMrPCHYz7XusTZRBbqXe0GWf+kapVC
MplKJeqoYN069h70xFYijWH6C9lfNNGUxCfVG7kTSTXfXFH7A4QeinQ4tN/Dc08RaVfp5OU3F44U
MBrQ7CnHGc3eC4DIsk3z8KpaCuILlq6QFWcD2NgtMdG/IIC2sSuY4IEUwNLyk8XnMRBsRy/qw8sS
YGfmILr64RpBMxr4eJv3CYLakExNaPBeE/JoHPSXN8hxWOhyhCsMBgWX+TnCvav0vE4ofitHOygj
ze9QLCVeI9I+NPKE+atBgnlYVquyeJPy9dwVIMi6pEn1jVJaV1EEwvad8fzELF5FYrcacrlxt3xT
2z4Wcw1/JAKfQm1pd0L7eG59afHc71oNSs58OQBvGFpwVuSFcYrn/rumm3xzp/yoDzD6Ai/xTnOY
A2mS1xbOEJ6wZ4NSNoF6ZgNDz9GhTpg1URRrCOkMyke/1f7pP/C7gBiAYPLqSjzjvJkoD9RPqStq
omObx4XVB3fMbrxjoI658YXqlFcQpCUYKHWnP3tocdOr3D2ow0bQYITEOeuSSUTw8imx9F6ON/6m
JoPFBrSpOxYwjf0u4IOJwVaP7RQJUmljQK/bALZCS+KgFIrh5lyp32bVa5aEImPsYAOY+d+Avuge
z6rSaru0K9xxyzJujo28YNtkZ8G7HtIae6uxvTCUCjcnW/5nIBXjhyBF1OOcC7Pi3SL4RqT7EKBB
M0lP5HLpF7TJL0hoZsIEmepeglbOMtffHJyGUUnSk9K1yj4/TbfpuRxmraXB8zVtmZ3A5jNUL8+h
NLG0W/eHlmf2MlvD++Mee1jLqzZdesMkUHGq1s+IMtnFMvs8Rs6kCagKH3YbqqlnePYP9lOn6L7z
Z1RKzkPybt0P+gKJNcHh4ZL912QJZTeYOmQ/NTTvidB3ubM85Cy5eOjDRCaJdhcclTscltWAEv1G
qlpE9h2mq+bKW22xBuEVClakiEaBs8i7S+WcXSw6/65wlDnyDDzDqIdFMnmwl0tBl+fu9D1UY5/3
/ogc/6ALTu1cxUCmw1ZrNCsNSWVqWBS9Y0HwXyuXBg3CMN8UDezs/ssKW7y3Zf/DVkZVQazZwOp3
cC8bns82gS3uWptQEOLE5JiqV3svcNbEsR1NRlijNXmyckOWoi9mqzqmpE5bEH9tl1OlkH47duOU
ccHS0JnR5sBa1uO6zoXsL0V2TTRb79nGbgYnhBTLFrjJ/rLjlUZg0yf0rX9o7iOTPqnnXNYJRgHZ
rh6isnJ0+NED2fdWyvDq9V1r1Hspn5zuJW7bxdnwSw+HUQbP85v6Go/MqPWvUFznB+LXHSwijeUT
FL9sbvvLsQxknjn+VtGn9kuWbsuEJFzwkDPVWQ5aLG+zg7mYhbZtRnGqLtTTlhWJMg8Svpz6dzAU
XPPYm7EjooZDFEpDfqpzQcaky0hbY06R35tVzUyucBRNe/+PWT9nidO7pOUdN4AQj9FFxhuJixTw
MqqB/PS2L4SgThhQnRx3thq+0HQocluFcpt6G9YE5TAAsCwuUjtFmDCKJWlcp0sJw4I60SXJW1aE
6TDSdi+AUDzXXvvvtZGMJHHHJ/KWucz/abJt3j7+CSO5/KVR8KoB3IIifnFyQYlUl6+57iu69HkM
HnXWx13N5waAXqT/vHSukDTzdQTGVUV6/GEeSXdHev3v3t+NP+FTCq2Ea3fYv25gf53BUjN2Pdkb
JwokHobb4lFZnEGE0m/Fr/bOZ2JJgoZlW53ukk2WZVgxgtSvOncgTx9KVofPVmyDWxmSdqfgtID0
BMu5+mO00L5kxGo/2wD66ydF8lLgHGdCD0tV0a8yV5nEYUfUDlb7F13FklWcXAPiaiKGSrTEuTcj
zz1ScI0FvgVqHTc3NI98r0rfNcCgjDXQsCvlvQy+euNdfw1Vf/mbBDIYGr1RjEgyyVWN3mOvQXZF
AI9oPzZWIxYNq5SQP99ASYDByI5cZ5pJaplT7NmYUJzxxgNKouQH494rPFgJMPowjHNrKzZXiJy1
KRzyHBuoI/r5Mguakmeik2o/S/Kg4N0UAYFcW9xqPb7mU2uT0Yo5GOft0+G2kU99r6CeYYeKlWoL
OvtVLAib7mNRMXBnXhcza0c2ZOYxIz/E5PXN56kiBhWkQBEPMAJT3uO9kuojcXxUAvzY38a6Fo+J
4n46n1gDXWAPi5DWFYMn+aNIcpS+9FhMXx8F9Q/HpnRuBVBaei3lmZsQXliHOmh6MLU306Q7w5mn
nTCrpeRHPKtJTHQ6S3l+Lw/ngKxDdcdfPnxCHosNQg0JzPOSilE9YFU4jWBqeat4z5udgQvM5eav
amuyflayb3g6G5smMt23YqkLA7pi9IAMUOZhDjTy4ULHp7JFk4QT9tiX2c9p+puRgMJ4egVQv49p
g6lZmH11YMtU+hvgQfPSLGD1aq5fPGuKM5wA23+Cenw1Rz4fllxuKCtxXSogOjERmlwmSeRO8x6b
bFRM81d0MdohntBpJbcC+nuwg54brAWY4/bQfjiTTLhRIZHYCn5gV+mfmPO7siK5+72+yTer9pXq
mFMMVzCK0HFNDGYab8220W0noXn6Lsz0jVi3mKXZ1CZybCJduC++Wzk00kmAgj4CGScDnBMyY6Kj
4W+8nLj6z7gTREWKtfLrMteXtA5xHzClMNyQpPG9MOGymHf+WgjgEEbi9vdQPvodeKXOSzMGt5Yt
zyIk0JBwF45zO06CrChWcyZVvpLcyJCk2G5QfghxKs+2NV6F1+LA5W3BlNGuuFQzKOyGFP7IiSMW
7+fQXH9cFRSa1tH0mSGydZa3Wv0W2vf1Si6B8d9RWT50KfQCnxC31SEoyt1KPdwo4SiIlpuxQy+J
qcGEmqiqLh1PxvO49dFDmPYI5M5UyGUfOGDacruQe3ovWcR+B3qu5Zc5RqaNCBG2u48BVN1bOOuB
0rv/08rwmy9YFDbaDypmncw1xke6GFC9dtvK7M9Y/d3Pet9O3arkhRUe28fez/JuhWBoBJRq+vc5
UDTzokGBkdCJn0AP9tlJ28gVcjHyyO9ZLJvO/Q337kpVSfbdeepEWPK51U7eON72+3/Z8l7jVQ+1
sXcgbBwLvcwLwxVJGm5Nb3+8cs41I9Yw/s3hxJA+HdDkMFMB9gm/Hhxxal7kGZnUHQIqkN4Q5+/a
Wxfn0M7GzxIF1UrvJOALBx7KScSG/eBHivIBjTkNajH7XYXF4TinMfG3w0q2es2nN1wTtbIlb6a/
wZDRZxmv4br8dPyWG1JQgeshjpJ2muqeCBoovlP4k6udlnFtG8g03pU3ASdcyV7kxzCSV4leSXkD
1+pleX4kWBlNMH1ZqOqXeaXco+MvwgrkHKscXd4iAG48ZP32ZVS6H+4VBInf/vPpy5DS/b+TkRIO
w34M6IDdwXwUJ+Tc5JHY8GHKnfI5ZzYy7pAgOYzJkoRGhb+H3JKvYYXscI6+lSPY8jHidWyqFNjX
wBSRGELmy5nd7DR4GpYtDWdcD3tYkXwxIhP4WMTnMELFfypWkrXh7Rj2L7/ASHrWfWj7swgPy4UC
SnqBQZ7vO4oldm00WwOoRnCWmGTs2p99OUTcEQOlMkMOAFcElipZLlzrEqXKEhFOY2Q0+FZmj994
F7nX5Vas4qUxp2JVLL1OoinNBcbKSdlT+79WEeRzMU9vZEYdCHUtWOrjDLT7EqQSqjqaX7tRQqTW
PNkiaBY4bgcnLOCK2iJJO5quo9Lv00/jlHHzKHGNq5TfAgIHBQd4z8bs4UegTNM7xWAZFc0mgBYu
7TDaf02dFT3ajljMlA6DQJuVdAeU80CjULA9xdd/ReqcKTgrRq4yEyOEut51JvtCPUfj/769rKAL
ZQRaEREbWMQiR1uDVy2ygI/m6t24vQqIwfCRnynCXUC0FWzTg5YGCr6SnnEIXURUhusHgFDwwH0/
wXyE3xDMtLn68OuhnbM5t9TlBt1FaklswlraC9Z5ezaMlhZMI5ZYZiGM9At8RBLMW6ml6jtxzVEe
MRiztLMtPD+10ExNgdFu8dZACHtPlJoe8Ct6TvccFCbmYa2oz2IzRgWdlVE03dQNjEQXtzQrQ30k
Fh3HYculwn6XfuTJk390W0Pd+2afEpgcWDygW0kw3pxA6L49bhOcxLn/7zwtMv2eT+JIXyG/LVHT
anP7Z8d04iDwHPEajnm9DN60ZHW7b9h5vNIODKTvOatx/K2P5juDgWvJZTSSKL4ySr7nNv5xchDJ
mlQTPIKe3Mi27jNWm2jayFYrzPM3Y9kcqYDPiCwEZFSsHzQD44n/xrFQxZMDZdBZI6zdPOackls0
jEsn5FQUqq7nQ0MI5CLo+LYyvuRWuSioKSOnpa8/Ic4GmRVRgA9xD42TsK8xLYHI5gbF6c54DmyM
S+0dvrLiqUgULvTHlJgc9mzPw3w8FYuFGFJQojtaB6WHeAnHjoPaJA0jybvwedsu+zJqHcMl/kEl
F98Da39Q4/aKFbSpe1CCMbvjcG8nGegfgkLUYucoxGNpQp2DfMDP4QKkl/xzpyU665+rnoKByPUY
bW82fADj/NzZxWxMl6Lu/TcoiVYUPStSczCyV7RHdAZul6lSweQLjhui6gi7s12TJDl1qSxtWzzx
jPllyqyPQQyuj8L3fVc4d63tgv6e1wqZMyh7okNNXlHKIwsgu+LwxxGqCiZXYJKgKMl5RNpt2QkX
rnIbYpqE0+3N7eJbG9RGCPXbZrGRZyBv3ozX8A4PKfKmdXQKSfsZBtQu9T+/xU5a6HxIG1jCZMlY
83ECczNTR1xRdHKnRfzfuDVjbElceYHtIegj93pmQWju/3twpU8MyqDS9aiIte4KHxXPtP0m45zG
idRM3JkPusfO/2ULh1/7GfL2YJyCAEW9WUu3VQQ4Tqm3d0y9ZaJ2IbERx7ZzFgl2P2g7+MemaiP5
bviA+RpgcgE+rOsW16pbB0nnv2SQ0HyO5Z9lnEH7FZduqtM9lTpDArTRIe6gjBo2Yv0xGuclNwFi
80GZpjJN//iH9RxKLbPCIy6qC5oRorn+udpUCAz550Y25u/cQrPGK9s2DnNBhSO9zxRoCCAMWkrx
PTpAwxONDwyW5fsHA4fgf5QrX9sNhY4Zt3cLQDBpTX9hBFj4OpoPrgfvpEoiZEHiZ9jIiz5to1Wl
H+f/X65YmbSHGpxvRQfQupXX/Y1o4WKeCf2nCk1vMMZMHgR2K9N0zc3vpVZBv7x4FUrDpXcZteKo
K6S8gCAo49hINZ6niD2Hf8sowc73qfwfMRXZqziGrxaWLhxUYa6Sh71QNOnBf+piXUwVQnpzllaZ
glLjf0FM3wkqIy3BHuRK2vOvnph2zDutdNE4XBMkdOKj7afm1h8vmZOJlFKTc0xWEPaq9m8fhtJL
kCGuXn3JlLh1umJAeQE0dQ+qARe7p+YEnaYWoaPazS4WbkijdQy5WrRc56wT8qqWw2sNT610OZEq
A+HlGMdErv5l6DedeZ9uKYPdmOY44DJcV5TvVHu8o/6fUc9ldiYAJPXsCxbCiF4iwzSR2Vsv//VY
oIPDzAcQD6w0AFoOSsifU9MUNK9erywtz/LDFtiY/FNSNwFXS9ggOyEflPlaOASKVasuGHT9ssiN
dkjG98esa8DsaBRHsbRUCm1ull6pA1ml3v5WhAyRNJ7wF1s26D6dQXUdJqifxetZj6yJLyZ9sjiP
5VjYNLE+rnIfavE2iv5J2rahgcDyn1Vq8Izj7uE55UM4tlDR1uxBOpoyasJV5ejbfOIgVBGaZmny
mD1N+i1FrzA6w4u4C/XyKHprzhzlccxbdaPV8JLquWI6kGpJS7SFJ6BcevUQ2wGKwSppUcX8M1BU
Ex8g19ytxiS9wDXti3B5vyB4U3M5R8BlSmJlXljgVOeEPMDG5eVT6K2ktKnbxJ6L+AekE/Kzrtmj
+GsnNWM8tUJIXGFIqaRrDTlhzaYoFjbaH/krAAS8//ws8pr6h5/xR70v4T8bLqL97Xfc7u9Znqjp
3bbiVcnzPqbPuUFu3Z0inoGxgoDMg7G+t7Dg6k7i5OKTuR8VUNMe6A3T8r2ROPr2CfTCL46deoS+
rKHi+y9CgcEmQhRTCHKycFyed6dIWUdMxdszQ0T5oQon73QUAKpXXr8iEKn0ZvGJrhv0o6iXwQ+8
vr+a3ZxwwN0q7eyRzv4lKa2wqYzl7CxyC1hJ6liHeV2FfCmaU1HB8lY/2UOLewgIueoJyTnUR5DI
HiISZYdOeiwFWV6S2l/YOwj81jv8t4VaOkS0fYANMCJBP3XmBji8a+eqPKrWPzTFfyuAT8eFyRnJ
+69f/aLJsTKdbexvnO1ePCR1XEkoxEzk8yP8TjP4VgdVGHy8ct9rAdCSE3ZYexQFN2K1gKgHGVBy
lFJh4unZpwe349E7ihgQLHUPj4ACDcY0LxFaFQ6wzc/fspd/K/jVxNG7U1KJ5NRI698DsBuBCT3T
p3NMwp0Il1rVX4eCeuTIc9poCoVEsk2DA1nxfWAExeLOXVcDU90GHnhqfvW+P/uXw1Pu7Y7zkhT2
+1QY+NE9gzlVw3RJ0SixAuCisP9NRIfG5qqIY6XAaXpdEvswq67i6UDRBSrZyqXQp6idIQ33iW1C
Kyh2qcPnqf23EfWuBYv0hgBYJ925tiDkdxHjuKbirfQkhe0DHa6uE6inwSEY8H7vnF/GTphk3C8y
6O7f01SJKA4ctMbmd3ftcn17K5jqKL08EWSL2lCi6u7NEjMaq5oeyrvs/79cTSSffRhGA57Mt4pY
R7Y1l/9sDwWMuJ0i7U5PDqfFXdOG574mIUGieHbQpQMkfelhWIiv7X5EFiyON4mEowTwTUy2yIOj
BWOrkm0tZWYg+Bqtp8HiojNcHL6HkiOJRM6o6oAfKivB3cHCz7r9lrM/QF9k+wcPe3ZocGMELaGx
1Efu8MivOOX3tUmyZ7ry00B/Cu9SVdAlZ0jaMOv0PAYZ8cWVRP8ej0LZ0qQ2H0Z4l2lcLwwWJ0FB
SYpgxfMuW1cZxbOMBBllZN2/cmx6uaZUZVcnamDg4mN8luzZAriCafcp6J77A54LY9wM92raUesM
7/ZVeVXIj9T/ROx7DuUsYMtBDHX6bGlxwydPhch0QstIL9rCgXEoy/ayfOQuZegq1WebbF775EYv
qikk1u6so06KMgoqViaM+y4uCToCMzBwYE+YlRLR9eKRAv0T/FAhooU+jTHq3Aqovbq/8MFKdwcQ
3bGueX1cTPoyWPNv2+ZYScGERrLDDErl4pCtA03MJ7HhCCH+zVQ+dtkaZ6tIh88+3ZP+M5+lgOQg
ueBeUnkssxHrW4NkXMGJd/f1w0eTb1JdmRg1b3u5TQbRJcmQJS6ruazHFSgm1R9JayX5Bu4SeltE
uSAkaz426KENkV4CbTc67mG5EhzAAFORBExZOVz3q2E2LjsJ7m0XE9KiGN3wPLJVpRBy+jkI3l4E
A6+ut8CNw1VFyJacJeSHtXoyG70rvVT2nslp8+H61ovl0SZoh9aaBz7pstlHVf0VstUlDYNfcxO5
+aWiJXPftzVpaRA7eMvFRrGJXk6ghtxsoBIk/yU2DMGtuCwLtg+iTKCCqayGA3PdZ8DVmxLcXopv
oH+VqjeK02PnmEU05EuwKp52eRnD5uzGLuVLl8ggxDpW5lVFrvoIi6CLvAKfab7jhuGEybtlAiZi
3aRxK2GVqfWtihokIVeSi6LkpV19WM7DE48l9RRGo3KYZFK88uf70XQdVjy+4mXnPkL3v4pJgTIM
EjwUQgmm7W7xEZi2iwnGIoT8zFXT3ruRtRFhhAA/LbHpTztCD6nzzPnrlXDvV/FMZCyaHWYZsSW5
lVl2dQN/m82SlSEkgaV6MinCj5HoEz4fKDGHB/Xk4C698Fye0sgLig6zu0xxwC80S4nYSI9PuRWp
MXFW5t2wdFvpkw3nSVUynrxDxf2aZsQz8sHHLJA7VSsPFzSOPUi/aiVXmxEyLM51K5SUbmfnC/6x
ARKdg2GZ11QL+ItWrTr7mQt2vb5AQkLb9ZrBhMkBZuX0Jt3iAgCLzjoOz5eDQ+JrQwQVx6Y+fa87
vq5vAD06g6mwkXfVcCFkPBG5Tqb3qXwoBo7PkjAjw3XWIHgHbG5zfupVLFJLsKPeK/oSSwNf/oiy
advCIzitMvAUgLfmv7hARKS0lXM2bL7LDLIuYhS4GeegiUZCDKku27VmQ7raRQLgum2uyiPoeCMo
/hdUZ4tfExi4iJWzgg7auNIXVB+8zZjX39KAT+9jyqcyrO0r/0WWtV0T7Z2Bq4VNWz74pPjPSvhd
qiGjrqGg2kHzDuuHhyKSsCjYAV4HAR8Y1v5aSa7sw4hFxcEduWU4Qr/1Cn6zaQJ7Q+aLPDuTfWbr
pcl80hT43uzCdgfo3FMIUuuOgm1RPsrVohGGnVLEACxbtTQUSYu6Oi3GGWahN3b8eAEX8Vo2i/Ro
euGAOj6mIHQ16GjbYzJgCC8x0sSzYCnwKf8JDYaWoEK7WCm2ht4SuRpJw3aMyc4dWvqw1AR7KU6c
2QS1boGpfC6iNFehnyIqOPMePIlyvt1uvxEaEnEpuK7/KMNaQFtT7GYl3teNKkPX72yTQxDw5Y/4
qVhBDCPFZukIBMZDBd+g/me0V+D/fDOrDg2goatiZ/MsgTuhPkXJaUl3PV464c+qLanTIrdl6gCE
tWVXtndLPVnwVFWlP+wWnFSmOGEkr918k8Ue3JYyL2gCpHHThEEfxVTzrKKVPXdyZp/HjxkdIET6
VvWagpOZr8ni2BMiMi3Z5BEQ/vmRXO8pdBFY6pTwLGlQaXfRep7Z64FyRjd8TQ1VsTEGnXrDwTyz
RF4U9tPvmJXDboSGRfhlXzrINH0GyhTuUKL0xXIzqXEyPD8NlukvwzzjecAh2wSHmwoByn0btkIZ
bT5rY964YlPPOw5pNjavLCVVz8RkbdX/UsTu+V1MZ/056KXbVAtte6FFPji3YsniM3MiwSs2PkSj
6Iz5mmB046raKG/FdTk31cSWuOWvBPfx0YOgIHKpDdYG6/cLrXL4wQVa7UVwPLlhVwGqJpKtrLFK
Q50rTqmEQqBFHFgQauwxboHHFTBYJWrBBON14CaKYTGqrI679jOjyz+1HyayhQ5J4XNqH1fVheOz
ijMBr3nMl+gOk7yzZTHHnc7lptYEKzjQxII1yYAYKwbZcRNE0b8Se6Je1uzSB7z/ObEI41gg5U1t
remBSWxk9ivboWZl3y/K9fipEJvEdDM2vP8rMA7LM6O0uBI9i5VpOWdsMEhOCCYKla/Q7vA/Syx+
O+GDdt3ytydYMOS1KrS9NN+1Ma8otTqAQxzWLJysj1MvhfVvusjXE6xoCWRnLjunBstvtMCiUkxL
bisqmmllUEWPwJUgn9nIrth5qY7oEqV9x61FLQdmLbQq5ovHv4IXfV0TcLopkbW7WSTqGCVcSaNt
Tp0XZ9/yEHmfGhStCdwT5hU1aR5dLheyF6sKQuQJqjeLQUcysZIy2lxES57iDYhmtQS/OHhM2T2C
dFQYCmnnpM960lMJhgujfObMgNgZCRiN4G1AWwmJaX90Xjk63rLPd4h9FCb3rLRHTMH4v/5U3ySB
sS22J7YtrmcLkN8zyuV0eVGas8ouAiHUvFyZR1lRPdupzqiizaJtF+fL6+LZ7iRcKspwuEmIM/eo
OrXrXlT8WpggbgeDzmXwY3OEnG9Cte0zTqa2n0D0XhvQGVEAXvjMhpEXWvv9hF6H1mOG3sVnYdzo
X7pwawN6kqCbndHry4yWMUpTPDFkZipDPH4gE6YZ5EItsVZchV6CV63DByQL/00tMsJZlcb/VgNf
QSvH+hcg+LXvDI5swzTQb5cxL2trseFhCgoUS8hwiaWaXzbkfd+TbzXIhJ+74pGb5iFC98fBtheD
PCOGLLmfLor+Qjm31TXdeX5nosIJunT5y7FBhKMJM9/w12TdKud5FnAJAJp3G5lkfrXBw/3d3akW
MSgFNOdR+AqGBcATlAJ6ROgOQtfOQduhDHlbJ5CILG+qk4LwQqW6EYh4vtD7b3fIaRoM9y5fgueF
N/xAmMWdc+KF17SHUgrM3NNmht4zFMknbBCYV0W6+QdpOYhsk/KuzGSxvu/oLOMX3wDYRmD6sXv5
RrcX26ABIPDG0nCvMx4wn3quEM5XRig9eqMpGg3VarUJQEwDNBiUogu0Uv5Hlk/A6uwruxiAjOTu
1ku74/nQX7EerhhsIhrXGWSpgR72qRswQoobSYmz7hitNnKxGb3as8yZfljFMg8lgWAZbgBSmMke
lMpHWpSpcGmiCMY4CADHhewQraHgpC4UEMNrQl8GRgCfM96QtKG/p6PVpVMfzQP4stvPalL8VfLg
uIGhUl1iprLqmWJOlZCdxytE5al8KDQriKtLeHfAwCVH5RXH9Xd68XMY8nZ3VfQAivs5z45B75Aq
RCZj878FpR3V5guLcWLewdJYsYyTHxtYOQ1bdb8lPPnryyUEGsvYtQAAP/ki0dgaFWa0JDu5fzRJ
N6voq5wC4ny7X86YzmRKaYBpJHFE0l5lreIODebT+B0YIt/r+m+uADrOnUDV745flcWv0Py4Q6qP
zYY2wJPhAFo04obsPaq9nSRPgQuaFkNCqFO/DAAOOtgV6irOgw1dW7QL6E20VwLW6lWEmTStkM1N
PbvLYWvDupqbhwKVhKUihoKQke/6NWBu9x8xgK7U0bMfzdk80XznZAcOjvNamdRefMwIOYi7Rn/s
SKkkPw+t6O8y5Oj4+IN/MqHU39DICmArB/5wi/REiQAkeIbHFhce8zcoaE1JUM4zbbevpjgrPYbF
Gt/dCIXELP85OEyk4APnDxB16/qZURsL96jNk3MY+6fyRwq5SGFV4woiECSDB4bhdeB7ckC2dyrp
4TkpXGMGtEveZW63Mlqb44rhdvAq5rOcx6DpLzqbCi/YDiRotpznpLv98eE4+ZmIJMrxP6X2dlbs
cARY2rNrvRYIZc8feC+nlGhkcDeF5m6uFDzTEoTlhx2Ew8awr9+/a/af8HX86IBo8/omLFbKwcIY
u96MNmDKuTcaxToM/h96IT8ELqR717VUzTBg5SQswZnZPXVskq9zN/414wu69DsQy77tdC4vG4Ld
npGxd+fwhTVJ0DPeX7HjhCEVvOVqNmuaRJTwjLF0VT94E19J4y28BCt8p2WQhehNDDInyUEBRPBd
zZyxs/debXuDcS4cH3BuxXuINaUjc2BIdOrfrEb7iodusFKG1chwlM8KVz61EzOyHl7pCqb8gFCu
U387rKrSbJ8XO39X2noDQHlhN+NMlXj9hD+V5JpsJmkrikrzL1dEtI8J1oghLAPiPsCLoawzjTVB
ZzjUseCWTyik6NRmATbSF4sBHjgvTIMBiEKNP8DAJXVg5R7qMHZ8bAXmEGcMlI/qTMSSfRVxFrIa
P93iXhaiY0EqU9t3/Fm0TxABO4sN0mLimsNLi5/Nl7PoHdnSEiEBrhWAKNpOGO6oMPhiieiqD86B
A4DKQTM04sX5QT12bW3xw3EVBqrC0t2gcAO4vn9AEdcEuBZu6GDD7/HZpgdz25Jtjx3+5qjulQPO
NYaHBUpAQH9jr43BYMxNYPze/kI6tvsktU/I7iMErvUftALsF5mlitsTLsBkpmjARwYYQ28iV4oX
9ZVFGjGpipm30YY0nsjG6RRtJ0D1kUezLmlp/KGGp6a8xXSDmS/8i34gMJV0h3El6XBD+GUygAd/
wEAOT1JVpSPb8d+2iu6KwnaatG+xuXeIKgiKfL1gxs7aaRJ6VeOnncPFlCuOTUH3NlKjm2Gzfh2A
1hbZc6nNAe9iKqMWS7foOpOIOKMJEmcYoOf1cHSqGtQUIJ1wvvUC46nZ4CCdaYGT9SFmufeiOVWC
rT5EXzghovSaempc677SZK8yEE1MOQIgZsFcpGdtOWlW7R4DaTyh3lk1vlft7uIX09g0Zzw1Fd8M
+MZOuu3VQnYV4BwgkvygL/hUwJF82kOhFTIfmbAtI9PPhi9Qs0WKcZiJCWRM/K0L8ybWILZze0kc
SPWWhKMV1WFdqKxEIqsbz4hRhVADhwYI8BARqSdWFGB5fyDX/B6tV3B6r4P9KWDIFj1oWTW1DkvY
JbmPu84KLkcvXQjoTXJGdp0k7aeVb2vOZ+pJlFulY5/+12y91y3gFkUWGW6p8LJNjjYKWqGsVdM+
zMR0rfxeF1HE6kIA4LnlmawvbPr2dm4tIsIkqu5wQfUJKF3dS4G+HORcSoVnrhm2cbQw0ZdLkMl5
+YAQecuc1DYIK9U/SXhdDgCEmAS6r9fHmshjPDTCVbIsomV/bc5oe+BUym38o+iYo+VsaL84OgIK
f/PQT/eUGbe2pS9RrlrMix3Ipd0xudUzEfk4uktLxb7/6CLGgwYF8eWIBRS4POD3og7LHwcA1kT6
yur73BmuIsJFdfMew02TYiVovSDWYZXFcCzboOM5EAPUSvAICEHtnHQWBTPF0WKbjdtKSPAmeczJ
QuiCfnw1cE93kH3GRhBEboe0xXjfwd2D1Vjk7vseFsikNUh2FQElyDTZHEDpTCg1O5AuOuWyMcXY
JDtNmlJG6+GF1+o3X70kxNGN3u/R0lUKNYVoPI5kyKXTnWXsaWnkcrisWhY2sF84p4DJ013QZhgh
DKB+z8zg0kYak18+Hn6FuXLqw6VA/s+mzF1g9PagbzXIP6T1NmCQxhKb7mtaHmI2dLa7cg4Tc5mx
MMMudejwbXO9TjnjNgSeVqgAxM3wPz0eE1sqC74/OZgLpOx18HI5iQxCPFj3kaUHMxyT/9bBSNvy
43gNH4/n27Iy7Vhy6SQX5/L+3yleVp0XEwSaQUPatfqUOg6Eb6E6Kig27VK2YuDtV8n6SPETXUCj
m4xZuPGYHBlXreCfKiaK73OhpaoaE/HySEfsDAWqd8dO3YpnNPMlnB4/7MkvMcfqZUALlz03/auQ
xu30P1I6RxDy/sZks8oHzp4sst9Ph2b2R7gBueeAJCruokYklp7R2B5NdSOQET/jCIfyzvzZvwj6
DBKBun4lSKLmIAIp6Ccobp5dfgUMMqQju4C6/bPaqgrFCRYVhpjZGCxscS9wcUJci+Eg3XKfa5uD
1aVmv9K/68vqR+COxN+xABWvIV2WfIUsB7Dlo1TG0eqYLrIWkpzeMpMzIjlCUMwTwhHoVawP+pJ/
cQ4DmQokkTZkmIY4VaJ7pgKAUfzyBri+S043trQHTvhhG9+/+j3XZNbXq166/GKqLCRr+ELogiiJ
DVg0A/li5s4ilFcS9YbKTBRuuQ6hC3LE6+DOzQ607Qsc2bhUJU1pM7mDrcVwYpE0u//SmRVFShP7
+RnDD188nbc3JZ00NKW6v1uAaeCmFjLkdLhwTGAiZghHgCsNmV8FLPr3LeOux6wKz5oPAL1DqY/v
djsI6qWlmHy360wT/NHwjpDH5i417dlA8xnHargjGFp/Cv8TySUNnsm/iHq3dQf2GqN3+VurBrBH
v2BYJ/dQ9wCbEGNAlBVGBCISVUJYr/dh+TrDtlkuqLlVq9Z9DgkO2z1FaV4iVp7AoVrzFXxAvZK4
GiUq2XhFlbQHarpAhiX3C3fYZs1kYATz3S+V14QGS5PBOCafKS7WfKYm5u+oFyjmC5gfn5LCI2nS
VcrpzvRr/0ZV8Cu6cWxJp03ZaP+laEluG5nISzPMYcjPkGzvlNc00hZ/5VWOSOAPyRxn4R5FCFnO
4bU7lsDOS49x2dhS5V7VBi7E+k57vWRRtF6pzJ9Z0jao0PcZ3cunjqhkAe/9ao7zPmXfQRX9OMQW
nYyCp921L0IIbUzmsGTZRhAxhSmeCJR7/vhgOWe4RFU02YblwCL7+LtafORqQlvmIPsBVpu8v2hW
bZK9Agu/vCafNXLzDOHEt6X92ZBKoaumT8NkrS1KyIbQrH4lQpBdnFR9IpvgVVgGvZSQ+qE0IDvz
wEZCXRLXU5jJHWuCaW9hO5st8aJQwJAfO7UtA8qXr2cxdOO3zCSwoEsCUXm/Z91oy432vF0dB4vj
S4q69EXecpO8LBgMpHK419U39qzhsFGVB244m6Op3bt6jqlb/OoifcrtO6GNChl7dV1e4/zM316x
V8a+9X+7yaNEQPYdYEYpzymTvTreoVjnYGA1QCwFX4I84gNbkhjuYYnEG5i1l+iSv5hFqB4kyz6e
28IqaYF7fqwNNbHOtfI8PMv0v4nf/Uc95A/qg9b7fHEgz6S5yKFQB/QH4xa/00MeMo66TF1R4wgK
6nO5xsAJkAARq/mYzKzgnduobwmXVqFFEkFcr3siOigoiwrBEBojHntPzTw/7tPszd++3lzZESUl
VLgGyXUzmcirb93bd2+9IyXDGBxuyOImXN7xMzPtEAr6xDH6ViJD6t7RGO0+AzNUYRJsf4rs9p8d
6HGxsm9ePIWF5z1C0t3CcuNJSorTKyn7ocr1s0FZCEG7eysxL2vYQqYmG68jMCx3CwoNYfcU2BGX
otPm4wxPoJ50NkLEc7gaJbdtJZD5teViE4/Z1AWJNB6zb8nekC2FYap7MFjjEQppuAvJelpkvJWj
3Aw3CL8k/iV0CLBc4MmAoojllfaDQ30W8fSWqZLPz43rofxMg377v+iNG0CKatFF6nS3vQnUlARX
LbDSLU5GwWEYoXrp07AaDeL4ndUuhI6Wu0mdr0Ik56lWwdvFhNUtxBzVKzA262VHGjpMbAq2ZzNx
0qpONm/0Oqtq/hyrlw4FwOgrd8dYevag8JXiFKzPOJX4QCAvWqCU42WPC25Uma9z0z01RWyMR+Go
eI0YuIID1csCMk5mbUfmmBLI/ozfaaf23gbTfHLNprBDytYDkkzqOD8fYGLx0rG87lXJzXKIcBBt
xXU5GIATMv/To9sumT+IlBw+JbAftlf3T4yhsDe80UMmsDnFpy9DItFsGJBckpeemzaWWDeNIQYs
Y0os3EiYTNIcAuIsiFWbvByxvIDzFHr3e9zkV3cQo1lf5cwNAtchtZ/auO1Q1MNHSq5cDa/ahCpa
hQOCnl1BeyUFv9YTN9zsPWXmyva0NGY8Z4QdqOwN9lSy0oD2ThXkzGVobCOcWsNX1i1pTuX0ZEbb
FV4LBI9USkDYR182KYD9S+aSZn1Iiwhg67Ge414c9yuFKzkRNHKmMJmHSlK0JCzvczefzSh+E7uY
eqvsZaUHs1ELR1E+fe3td4b+7CPk99LU89DIWxitJTOrzfUQRcypcUgy929sguoVDBG6QLWOjD7n
e7q2BJO86ZO55wD1VdPO3GtpR/8ScK6v8WMqJ8Iz1HEANDGjmHnwpAdDfukJ6Q4vppuMN0y26MgU
A6rMASpGqyUzpr7FKjx+nqnh7O/7tgWKDw6ebprQz505q+55ygCmHnSmivp3BoprNcTgWMUBpsND
aCd5jgI1bSVG4wCLDbhmhNFQBI6UzE3nppgdSShzCdnMc4xrRiFdR+bAvQcYn51dnoCvGWnjfVhu
zefDyKOLw4DSw/HXiSpdCS6YddSLQdm1VLwOfiBUSgyN5xsTQ0XwSWWLynPqTAvYbKzFMWxBA+54
9K8Oapc5O3z/oVypZLKBXXerSTUwcmxFI5sTx28+u2Cxm89i380OESVxVp13HPgQI63HZkB62NYZ
Sy/LpUuxI3sbn77dbX1Z1F+j9ZMfOpO/Ppnaf+BAkH+O/84y3TPTnXgEUNzrWvxo/PuYLD2lZWUe
AkU1kJYCFlQnoTlREABbCeCqhT13UHPWDjo7/MNDEVWmAhWmmn6+7LpzrkB4+rmz1O29C94OD2em
wK4+hRq8boqdXPkl1zkTUmGK+t4DzSrXjeHxwo1MwpN2HvTjaInSuMPRwiTetSHpfiTjuMELA3xv
AZQn7XAuqGLXlCCw/6PwXQvHMYqD/2ffbrqUWnLdOh0ljY8t+GF0dtGG9koc/e5YmkSI5/qoFiiU
objWwGNTo2LzyPjiToit6xjC0XU3H3lIpklSRzfTHefM23PX/wKEy9BsT8yzxtEIUG3rYne7wwu7
tAVB82hHMCY4k3geJaleN4a3x2P+Ag1zmhTMWH1wBp+pLP5u3kLJWS9BTOglMAvkEh/CCRYQi3/U
qWLuok6tQT0/agTGynHlwI9UxMs/KV6uuYanOkkEZpGxrUMnteaF9MrUFqAeBAGUam3+ElUvkkIG
ECGmlzqLEo85fNtgYX85YUBiQlp+EpeT30RUl2rlKy7JbGr/C+Duu1gJh0aExkRENDct9BsTeUcx
AzxPWV/W6CDpPATboVNAT0aGVFd4MNJPVBlqaakHG0j7hkB+BtM7tGu7efVy7b8SiBcWvD/w0ZhC
ULdWWDSO3b/6I0I8jElbaRuhsbf33TuJWqNMJlEkOrGRPuDSVeTVo3PVLpemUQEzCLEtVr8Ecto4
5RoIGl9HiHDnPVwlhoemrsJxtSAZ6KhoUR0ZdU+JSYeE4gMdLyJJVelLEjDToOyUbbfgKDAHPaCt
IuGFPXSjF3ObAHTWKTUye7RBtJWdAcPQ91H8OmBF6U67jy8tHXdx8weukQ3xzQZ2MtmaotEelihQ
U2583nD5zIgcDHvE4kaTGTMuwaRwfgTIhcBcGGSmhWRC60j7YQZTR5eAoF+S41OnGX80nDa7wkS7
ZRCW3Uz+5mGosn3yatXobKs4YwXeQAUol0krNVpoWJH86aWRW27eew8xQqtM0IDVs00W9bY5SIsL
Tz9oMf77MBXSuMw9wrPZ/qpliX/Eu/HzKfl4HYR1esqQaQAiKdX2LXQD3DYIFsARajUcDoZ2X0o3
IAOZqCOU3NDo/jGaNG5RJB6NN5YkdIQpoUd1QpsC/Clkz9gTYJHLUkQ01E2ZR+Df4YVhpHo8q0OG
1WL7WLfX8vfUxH0gg3HYQ0gDFczJkzAxG2gRvzI1IOu5EdxP2qQyBMv+U7D6VJoNkF4WDz03LpVI
AL1t0Ab7nHu+P8sd7/06edEtF37d7EBRnwYgvfPivVce4RxSU6uOT5Y62nNCGiNPQZgXLeg7wVXK
h1vxcILTxJjG6LXdFG1mtMRqwZR1MjxPFB8/iHESQTb//AQAMVnOVmZWyy+7ryjZ92+GCowAJsIK
Afxw+rcjZF3eLY7vVkwD9fqiBzqHRIGXwxwG3nVshl/GY0+sUNkQhQqpRHTIGGYcIGkxjGGCCjUn
Vl7se7MuRxfaMBXkdIsuluOELwlGnBo3ZWC4LB5DaEozllAnInXApD2+3Xfyd0JHj/ge56FWZp9r
7uDw9xp682ozNTZ75e86iQJYj/GudfaQ0/LD21nJX3xzGYy7/mdV/DNxovQaLHBQSIh3GcBdHflf
EpvlRHR0i+eT/a4wlepjAKU2VdAsJzTI3fshysxkqG6Q3RaxqeW65IrSL6KJZQCt4zU0vdgvmOeS
IkZczuRdIqwAF0CnBApBbWIFqVBhZZ/kx23mAXuzPOT+LnZEkGoS/U75Czxy86g9zqjReMP/Mvxv
7H3pag8asOc1q/M7UHs/BphYw+08YMV/q1/88hILVG0Fg39N0Rm1lLnQXeTUwMlFJk9zDhCnmZTn
e5XWWmepzIA4W/m8+ETvidiIMHcb/Gcll6uxsxLlSHZOdji3ZNkj82g+jAa/il93y/KZywfua7MY
QKHFC+Y+s/CuddTRGzQNxw0b6a7zPu681CG29s5KOvbbAfdQj3ju0e1bsCFywd4RNSpKgLcCBPsN
PeBcdFd0qvASnix2DYLTWRJ6+SBDWtJ0jMEtCSq4PZ9Mhltbfgjc4/X7R5W2YDc1VsZJAT6ci9EO
gNKZtKrJihWC1b+lWP3HdPggKp09O52PKWAn8eFVKpaDyjtAbx9z+TmIIC+vd2zej9jLFfsIMri3
y6JQ9o6ur8Jt/BHJniZfX8m5Oi3f+/KD8jiZibJZvHjwgyowC7D8gvWjJNkljjBDPl67pqB8Vq24
MwBoNtwF1IrtLwUPKg3a4yYK8fCetxvrG6HZx/bMCDcqmgvCkUzYLhzpNUeALbexsWBGhOaAy4c4
ONLDUALNVQtwcDQEzb9uS0J2pmsVhzkHkpM/si2D5Ye13/UOwlJthaMx5BTU3bGF/pNjpdhJo8sk
0Bv3RUVAMzw0sjpKycGoN/p2X+85mOVprevT1ZH3a447OADSPh0cmHs0hby2hCpTTigt147KMz5d
9h12mWxOvMZBvCLp3z/XFcnIrPKzd5MMQz5AW40KH26kItBFXI7XXmPcWrY0auGIBllwJsVyS5D9
17t4Qnuy/hGyQwbc12xmctafK1wZqHIGKngrlRJFHGMijMtnMwJ86BLmEHro36Adc+gVqD2Z8gDO
6u5ALxw57lXIGIreVPUMofBraHvozD0+DO/MiqglQR5aev5jeK2n9dEUSQUtfuoKM9Iu5KQIlp1r
wffh3DPnEDTfz+rXx3QdsYaIrwaOVcLg/VpdNZktfW+oQ747bPFL1YEKt7Wllrl7X1xhZStqeJ7e
FxU0lz3uxC6juyA7vf6INPKrFekNbPcaQZ4cD2lZ4dIE5VhuXCJc3NaBowxgQwqJGth56Tc/Z6vZ
va+Fq5xsYZgQs+BakHYZAQZR8W+Kp2f3R3MaOhlumKpwFMvWMsqartSkYOqHMA2Dom8D7bofdcIa
Ej4HSHrA6K8O0nFG3ak/7AQvF2YMgo4p57HmfNT2HYDqyF83Us/FvN2HleeSC1OjtexVKTX+rzpX
Bzc4A38gj4dpGb6XSwS+ypYTFrEvf4seud0KFmnDTRXjtqH4QMyRVBEy7/qPK8e0HKyi//RciX8H
0G0PuXNzjDlcQHYXF9281Nc2w0TcFtlgiKWby6OQxjvOstZ+145Ta8w//x68gFsfYcfrzVKSyq5T
MMvhNc+LxQBCfAJGU0lM29WT+fXcKT+8MJg4qC+jrriosv4fFTqGX53rnStlgbOsPQGuHNhv7MYP
8IrcV44rDJDoRrwVYsN6v1j+k6ZbccVq3CQYitdFMqTDwYhJJ7wb8dKsQO+xNORawSfgUnoy7dhl
QRhfumPaq7YzjBzUkWFHj/jdqV2A1VxDtSYdVDZ7KLfU6ia4wmd4N6lsmttfXUEDEEn5TrvYShT3
z978AfKQObr420bBkqWeS8+3X5id4k7iAWxW8OBdQK54nZkbU5FJi/ZcYX9x3lMJeRe0qI0QMVea
dwCeRkQpYnDfW48+bWZmLmZ9jkBN4z1QgctC4YuHY47z5dqHVsXSneooKD7VBsk72JpcBXkCmA+3
o1ddM7tkdsKcReqp0l0a5z4SMxsr2vO3v3VhJbnjtDgQwhlxRXx7eLd/8ihryeFb7wbckZumpNI0
XXgHkDELtvAN2Tr3DCGq4pg5G4djbUX5lZ2zM6KrHamg4u8Z6/K3TTyfU4TlVnMXgiWBeMSCEWB5
4iAsvvIj90OszIVmFJRg+2vUcRgqglVaFg1bu3kP0V1Q4N64jZHBRanBgT4Hk49jYbweuUgVOD9K
xzGsPrxybb3zmQJ3eq80UPJgoHJFW5XoAT+eNjYPhBNhqPUHDaSaCk3joc8MI+Lz+d5DTbo5qqv1
nIxQhLwO+5Nbmj7L6QyYyPBs3GDtXmmlC8iJZ0mH5b967IIhsbmYVMyW0dQguzWfKwmTeGaTBlS1
ILaTl2vRUcZ3BtqzB0LQBCmqfGAT/Vdc8gr11uONf0awRWhiT+aHTtm3S8UyDqyjXVfeMfmEKU38
CROu9HVQQQPAv7aWiWol8BrCiKjtwT73RZ1+ZZxHVvOKSxo0gTGBn1iY+8Z/+NVmqru46NsgcNqH
Km+exobVs6RWfKkqmMGODfmsNOCYdRB55CwBFX6yNI6UQjzaGYgvq/Q02wwKM7/8oNwlz9AUoRUo
/VVuNJ2oaaniUZ3W68oQJsvgyljiqAjh56dJwR15xwEFYeE+hjpVNXNpeD1LgZVUvPbmi2drCSB6
o9K5mrYTgWHA50bK6i1GUr88No7aMRP42m3FicDOrkQfkz0/kuzN4Lrr0dtpPBy4wi2TMOxUo3X+
Qwtd7dnoWuQx8eN5EabrcEBKics2ckLZSTGlcXhcwuRUlBLzEoqMqmBwU5ZeCQ6hqa545vItEa1C
zcxM+00Nk0hrYfVmt/i2rRcrHpPgWc/iUTg7Cba3OtxKXQdiK59GmAKaEAY1BMfXfRPbzf1euxc5
3Mj2RkQlwpz0V+RuNG+GUDCl0RElHMpAnO4eIEk8jMX8VkXQ4TzxOrhXmnte8Wbux3kKPbRmpuv2
TZIrAOrvZPAl5Tpfd6BzKSgvR9rV1mDiEhfCGoj5HZUqiGiC4noSMhL3QUkMJDSb/qZEhUka8r6k
9QtblyTLIScm/CB6gpeMhjddHb2rwqUUgtT1Ytsvrnw2bmK+9IZR4PRBxg+eqTQG2wZCcZy2UMUz
O01TSPRk0zrdtlWIPcwuKS0MJB8eTPdY9PI7n8FWSEeQ7k/Y3tTJJ+zat72K1HqQ7KEUISn4iv82
mI6pa1fu5i0kCMs6orDM/wCV5QQWo3HBYdGdGP7NgBinsFKdPuNg6XEjwhRbbLroZyVcAjrGAJrs
0JFcCWlsGVsO8+hK0/KKXrPA1DHogVCxE3fapRJGKj5wVNJUvMpED/4Sph3IZLFUA5s1g/7Q91+/
xJq72iyQV7Ti6bMdVG4ywDXYyEnx03uUPjOjZNQ3nOT5fGo8Jwch3VlBvFrj4RvhsekjN6HNv2F4
/pLSKBcjFosbbe8FUdoBrjppoZIjqZXsmzlOL5dGoDfkQO+xDvFay3gZelT7mLD30JOpRam9rF4S
QJ9WXTFt0Yqy1QipHkhLGx6WmIaiV/Z1yEk5C5FSNq+A3PSg4ibEqdtYZzbc3oTtR8awz8sy5Wy5
50J2hdNdaIiBofeUVmrJP+34kbI+V2FgewMDNKR6+QH6s+hxcgC3HvBOwOgQ3U7RXl9ZQ+Ymdyty
pzeDJWQRAlH18VvXNFu1qN/FLH3dqzHCxZZJVSc3CztXhfemw6yWW6OAKv3/bwU4ZL4AVHIFSncG
ivhefM4L6j3ql2Tm+ZEWBVNoenripZlOrtfzHxbw+aBJX7l4cE4hausdXFo5S6EvzfNz5V94Ctdk
vdXtQykRmJqTnX8VXjDTfWXTq4GtPdvw8ICxjck93+8GzNNbjL/g2VUOiImIUG/AYEOTHZrTUPpt
JyenF6CvgGCuenK7xAbUKDrpnK3+QTQ2fJdNfIAd8qRBwO4YtMzJ8QnOEe5g5LIWZ771IlCgi94w
Cqr+TTGzbrFiCYoTG+9KG+x83eQmYJv6dXehrNSnuYTYlhAR2VllqZ/auSdxOp/ZDpY8gx+SG6QS
iYV419F0enTuKu9CcTyDoXXYTV2/MfD7gfyz3jBqiiqjJRKgxddiHN17oHN2DRmyOg8Dmw6mVRPZ
3EbsvkgOyE21jtuUH7Vk0pEFhAVQSS3xEjIAiQFmJsP73RoPP2QGOL8Z/xBx9So9muInmynCJoyk
Z/zQUaPlUHbJQ6I9/wswIZ9o3lZ0+pqWa7LBEXq59vByNOfx+0NyTidfPjGxkcTiR/LoLmM/fR60
k3Dg8sQJWda9/iDbeltgR1+fCVErg5CXtxa4cd4SE+ixegtnOa40MO6Ez09nszjzcxXatT4VKvim
dye2deB5xiDclj7zS+y/ODTSvUInu5QaWRpTjtjwLtLcytC4YliSuCnHG3blONZDGgNFISc3+2zS
gRhNMW8BtzGh/r9DF0vsnIZDHVJ5q/fEhAiYwZuyZdM2CgAydXOmqUY2JA+cwfonO1Da2tcq/Chk
jMUh0EeFkzLjgUBDj7BF8jn/p1TMXI31SYI5Y1/3ovk0D/0x47DbLqXQikmFlN0gAdFLhp9w5Y6a
fsHP9pbHmegdfTr9Cpi3gOJ2u1bCgFvnwi2jTlnZJBqudmdoYdUK7OxeEn04tzK+3+wsHsk/FVhL
uU/SJFsE22K9CCJKEXfLYNd4TVm3tGwipGx/kIuRHnju+BGRHAypObJX3m8Q3el7Cl3JvW7Mt9vB
YS9TxJpZIKwmDQcJWPJcaLKcJBjL6wvuFs26cx4z/tl3KTY1+53H6POrRXqeCEQK3A8KDTbNJ+tE
4VmoXTXG5hxfMjRsWSPGVR1822cmqr8c6y8WKEQcppi+yO1Z6+XBYJFBkOWXAl6qfLoMNM9t+jPg
ASjKpvHkC6VOzDAmBfI+HxWoMrU0uTTp78IbQlK4y1mmMKHGF9jmYNQOGjDPJmTin4jAmJ695XT6
t1Ejt1JlITnmQd0GKOEDAcrEA6akloDP/CUPc/XXuLbxerG8D9Sn2LGfRui7E3j2u1PckyadAWdx
AXb1I8tf1sVvA4GnOtCJAJjSoEpQmbgH07y9OobGWZ6nv2EcxXtBUUkrUqLvD0+jMegdFoH5CQyC
qBd0mhRlIxw4kOZQMaN8jdn9PmOz4LwfflwWYX99RsP8y6/v5ya/O1feAJu3IEUCa5ksEDdFVRa+
qI9+Xl6CIO2UmzhpXMO1P6vCqLLFHTdGKTP0XFWnVvCU+Dp2Igla6MXhNebzpUhZ5LC0B4/qNgS8
F/0yYxTx9lV7SchylW8w2FMXwN7KuuuCJJLgVXRcnC7d6ZVMOPE4tEsmXG2YlbpJy0NBjhxzj1Js
w5c0N+EJXtXEyNw4tYWEkRtf9cjdyTobbkTDWcK4cmAjOWygML7Algx4WYu2At7xl+Rx6ho3EUoa
um9fIEKfFLvsS31VTNGSu+4cPa0+d0teGlDh0fIRiMYQaaZgJlMOoU1sGVtMwMy/GtNCW/eDHMXn
BAkvie5Q2Hc4Q2GlEzasZ3dUYKnnqd6hlkrFIDjvIoIH0GkYWqxdBGrPAKK2RNojEoV4bywisVuM
OJuZOKEBDq25/pf4ZchTeOm6MjWv+L320bu6MZwzFP4Uk8u0Wga+MnsVtois9VEEuOvmU0ynxPOy
gaQf5ixvpnUOHtktQgp38TKYAq1LOTEREYMfU0ZGaXng7pbc/kPx/tyrpyhPMDzH/vZAaw2gxrXu
k9go9MpJ0GXVaHLZDexvTSeDBYElE3ojGKNmak/Ga+vyNiN1RV8//c1ST+128zUIMVAllH7s7bJT
Po9jmu0UtLORtSY7VstRTFJOqgr4GJ3VvcNSRMJhT529/387Z2daG+fY0NW6uQz5n8BBiI0Osl5q
xWZ+JI5EM0nfZzvf7UVH7H/oGE3m157aRjji5TlNBzL4tkbeNlNgY3a/poyqZbXdxHCRuDighjuu
Emg0KIqDJdyuZGX5nrvXxmXpcGcBJLo3Q1mczFRONQBtqcWDF+cQavgL+6os7YptRbbDZkyvQ92C
psjk2toa1tdsQ/vdbVhzRd0+i/jyoTlTfM9LQ0gl66JvpOTH/a9zHyB8JFZwLByATipo6/jj155m
sCi8spy48EMCL9YjSjXqFrAD/eBiBf83JJDhiIerHuXNvq3GfmgpODW1xVnQt64KnTEjrkgaRb+p
4LoG5YhSggBDGDH6NoKE8QhzxmQTAtletOA8xVku3pUfG2uGHcYV6O/noE9jplxSTCiq4wIsYGNJ
acztIVrA+o9Jtiuox/7Lydckl2MI9W3f2BW8KfynOlLm0OPsN55+nqHF+Okx3bQw3Dmenxyn1g8Z
/IOO6c/KplBaee/OoumqUP/ODOmFeybrTX2V1CJTni2QLaVLZAWMRwONYdZQlld0vq3KuCjmxmQz
+KxXK6Vu12goFQKNtZdiH7c27kSf8B0rd5KUjXrcA54TddjmKLj0XncfOOxv8wO3zdxW45KVymRn
0tbpeaFvbDVtQE0+jj30G5IxSxldfczx0IxUXa4pm0t0GIuiRcE5ef8itO/WixXBR/78skJvJ+Eo
QDtnNWXOjuTA0gd4QhbakvRxwR0RWQjMe7WzxOUmfZvAZlrmB9A8gIGbuOGzv0Bv8O0av/rk7JOA
ydhPl99a2CB1MUZTBzzuWeTAGXVdBLVL9oL6DVy1Ax9s4MLJ/QjAyFBGO/mt+F+/fvgxPsdnk/Ui
vBs1ZuI3gm0wDHX0aoM4i1wt9PzfMQ9mvcUhPX9fMUkYNZOecthhhpjWWb/Li5hH/Q5Eg5xmkiZr
PrbchGRnjwxGQ0JZupitynaPMbnYVr90G698eKTrXtIZ1RQtoXorC/1YHoPy5MuWc+n+PW+9jNGS
mTE7tUaGYiSgWB2MRLr9MGMB/W/wUPLHsFrlM6O8o4ERz8EPyBjb96QmpKyxj1TuYmGQ0GvhjN1w
ycCvTgBGDD2+gvYGBs4kOlYw76S17Swmhy5RHyBnvU7kHHHmNSOcfXm0lwSZjel3k01/RvZ5uU9u
zZtvKsFwwN/tIKd3gRt0Udf9x8uYERcruk3K18TfCVXn44ZFQF+HMLnsxaV75LRiJMAPaZnIUd9k
hWJW/szO+Kab0l4B9Q4Ag2iYRyY3JiHUqwKV5otX4O+fgFH+MuGAdpAGns860x3I2cOY1K2iF6MF
qhNGZvIRMzM6HLh39wuvSDo/CfO7XCFmS2B7qc2yA//p2Scm1CPeDJ1zueeapSTYecBg7zvhqaAE
p+UnYf7vLHxDqe7ZYNNZgfvNN2wylMv3SQc+zKOyoQYqJLLKEmfz1vT/jXG2apF+nM5mL1yjHocA
wu5uioS2U8sl2139XzcgeSthlAzeB5kLs25tP2j6myASZLeuyRUTy5hnLK/uF8Gf+5uqnfJ4/lHe
UqIt3Y3Fi9/4oeicKURcdcRdRH2fzdFXVTsQdxP6FzK4QXcBPj5GK4rqBCipevER7turAIUgLVxD
6TFEcQfNEu8MuLlbYpPipPt6O99hGfcEI3HhLTgqIXOZnJKMYu5iH1efTNRh19GO2zHBTcO9cIS4
dBxAMZSPqgb+nno/LRmdDlzDlmuTHaJrYFInfTWkgdlUgzVQTdaCnhiqA63so/7gQGm0TylrsV1O
GZTTcx4R/CenpeFK9/69Jv9Fl5ypxWVrjh5V1RaESK0hNQSOyeGNEX+tiLmC/8bLuaXhiay7SKQp
xmDHHGkkXCQj0fWu3ky9ruX0m1E4rhKkYjsFQYqlBZCvwRWdplQK19jTmRhJbaJ3Q5LTCUt6DhvZ
XDBOwmSZ3qcAfjfMk7KcjA0EHtM4eA5ktbxoBH5GipxJGouux9QkOG8kDxmf/0JBr/xV42ZcGAMT
2PMjlMCoPQloJOftLjkd9OY0XLlIdgdXP4L+aJpTpkAfQDKvo8KLbow8BHQYgslMpwtEj3ddPh34
eci5YV6OmiCDKCH165Qu2BadNi061sT8UhDGoSH+ZCgniA705g6uFEyXgCZl/KD+dQXOCdqMUmSn
NMIRIwUK1CwRfaTRHGyUBw773VDVM+Az/FdpUFBTvHRoChnESE9WAcF2Mqxd7/q63o+2fuDDpa4W
t1lnEFFIEqdRfCc3tp5POc3LxaiasO71QrS9L4wDR7nI1AWhlj1hrPbb+kuBHFNjyyWGCgIvHtpM
PPZk3fOUe6LSfU+ecA21O4yyps0Cbf8AmKblRdi3PmzidQS09Fdbl4DYUAJHTgxAG3ow0PJ7wNs3
5+H+SFbdM4notq1q4Dv8fcDCKj2nRJDOgfpi6db4cNlL5BTKDFXI8LtvCKNGsDp+sTtdvtOXh5HC
nOOhQA6Kd8wIF1kuEIsdwKpw0dLDjwb81kXdIYB2nX8dwUk6Ua1+Yz5b+B0Fj/EFQCc1ZOgra8LF
BP2dK0CTfwkUJuU6wdgZzcU9QuT2ZgUwQ/i3OY56lt8DAYLhKFjLQ3lXFn/4VB3Z9ldyqRqfjggM
u10R59UAjxuNriklcsl1km9hYZXZQ4gq5QNp8ay4u4QVrW4r7OAidQda0vVRCXYZ8d51eZr8Nz/O
k8KqFOR8GrL7n5nXCZy4gmO85o5WU8ALUrStn5i/Tt37TwX230NFgjluxky6E8LkKfewWPQmxQYD
pf60+nTp+6f6OqaaTjNuIGug1T//mjbe7ajHaWt4YIfJGH3OZ6wteWwbCbCAndEtp0XmuzRL2jtZ
GTvdYaBiZ6nUuBpCup7Ov/J3xNU1ZMFdwGzhTGpB3DALayZjJvLmI7CL+8w/n8lahT6cJz016OU9
98z1I2VVwdxdC4C8aLFvIXb6DbofBGDBS5tQUZGlvxPFI9iD/QAoqZuTKEN8l8od5G2zLupwJGUh
hQDLyKbcZ06fX8dYrPtMa4KTzskgAqGsHbE231F4y1SYAvPnTbpf19hcY3wEQATmTDcKYVfLHfw3
DYajnn2++zJzpgEakDXalBW6bqi4/ef1/3H0fzNfBFKA1Kw81KveV6cpGJ06Z1CVP3diTqVZIUiI
KtpF3JscEimygWxn2v9wH9IBlFF94mO91oSpu8zMW6s6g6XqBbO7rRJ+lVS0vbqyMK5zD3jP7vkS
5yPmdfbwITUdiZPPTjkW/38i3lFBK2dffeL99S3aOczX2CKlsiV9UyT/SqmMcGmmkWoYhvFKQyik
ZbTAga8bQB7eZG632EllU9kFtSaGqITyhHF5TXoMEanhndACcj+W6ByFy2obIl3Tvp955oSs33Rw
LGd13jhikDhT6oZcAvBol+bG5o4QhkSsjOnZiwho38MLJxWLamfyIxVzrptB1VUeiAAIYQazbGGl
mhVH8H+G4yYYmMIyDNf3D6M8l11kWxPSPaVpPf5y9w80L8T51GaPXkuB5iaQycja+oYnoFOcvp4+
T+EcBHNX9CAOYrB0MpX6XEDDxYijJajAk1yHnCRf3W0veNlgw5kmU0HgvB2KS0JePnEmb4MMRwi0
2KsxYQla+8WrMdZL6MIC6V8+OmhWFsBx6TrXIfZu0eE27qlE1r/vkCZmi/6qrVG7GEogzSG/okTK
FbJFbFn9LS84TzRE3s4Jg5m1AiSgUTY7WhgHXs/d1NrIRVruyO2aMx/KgjQ2NeQ5p/FTpsJDW9i3
DWn5EbxbLd8tuNyK4DVsf8MX/qy3bcdeqgLL/eqfp1z0sjS5LOGtBtP0yc9beTRkbkdFeqEewPCo
jZTHLjyNYXKDiyROMmlaiLe2i4pW/a+tBrlcuEuvhuL/hlpHklf937zJZby1s7te1HrHEBpg0i+f
0gSiGSKM74y+Az0DDQZ/ODEvAnvTUNUTrRw7YBcNbj1JbWCp0s1VEC5vB6dYUqer76BKZz3dfzWe
euWho1zY7e68dWGolJ81BtPx9p+w6o45w4NhHz6zK3bkVvZtpRC1DUNx9nPPqwiBVUpn1jH+sEZz
WICxH3br3WwodyxEU0ARbnjc2HWTwL0BwG5pl4Khf+3wguvbNhjCiyCTKH43jF5GW/ltALLckyQV
6MFJVXpJzdyokMlg5xzxhM2vTcGhZ6nskh1ZsdO5HPFXVtV/ksBnm5NioDKsiU4a2oxLcC+K6nKz
GwODOr16fkawF0ibgKOWL7UPAwmdVcC7jgczy0PajvoA/r/5qQJtUELxfiTJk0qbWBcDg2YNO/xm
33DZe36AmucfPqpUXYfkcz3mYWFniK7AUacPa1HZkrUMOqaZP+Ia0stDTNNypY08tMV96Exrit1w
x19XnVOBbnJfhVg0Sl49MyjlMXVDKhLVb+MXWQPvJ4nTfcbzkoT6oO2p7TZgaH4Jhvx+J9Ra3MCQ
NJYtxidsUAIOr80Wo8DKVv/eNEsaxaPzYqlRtGUz0aW8ESVK6iA+alvQ1Mkwsr9S7jC2sPyBQU92
h6YR1TayeQKWRgek+mbcPnlEWkZOPdY8sUlENrc7BaAoRkJBELsJO3imVaXt3BEg9yAWmf56Gnzq
ECSSiCT56rD3+kuGHu6dCfPVW0X43Z4wbMxfNmAzjPNVwOzTskhVytgdHTs/P2c5R6R5P4QQ89bP
Btgv4m6iyMXPjEbjc88V4jLm3KH9d8wXe7dQ6/Bc6KEG36Aq3zEL4IHemUXfi0Lo5OXpEr+fs+gm
nL/oOHe5D2XszTQlSXzep95aeFtN5vjRPYg6hzuxsHH0C1rfuTODy6WBwN0ip0J3rP33IgVCSxT7
YZodrZQtMo+9l9eghy8nkybtDhrn0C7D+vliAMEaNA2z6aP7PkwAJJo42wu+ysQ5BJ6TqcfcRC/3
yEYSAN0oSp4ZHLN+7cBD6y+SJbvW8RWarR6tbPFUXQMmrDNLDD1mkyEKyPoQjJ7R1+x7Xk1wBDuA
TZkEA44CTRGgM29RxVR1dVl5Y0co9u9WDGXX5lAZoiIUczFlQMIdV5ZlbeM+mHVoXeT0f6pzQV8i
dgmIJwmwycp5SZLgUVfnqlD6hppi3aS6g6XX4BkeYrSx9UqctS4m6L9ipoJH9J8a80xPAO+6c4uH
PkJ7iBKhUHCIsgexJFaN45KuZYYsrisEo8na8/wTVCS8Rpr9FXTTuv62JOLM8e3OIFOEJkStoYgP
fhA9Ts7dJmEP4UcpzoqiUBUYiSRKHwx6nSQiMiXsIdX+gchxonxQU8XoGzHosg5orVqt9fzNbzi2
XJeiQtjmf126MMAws45r0zhQBEImtGji/uqZbFQBaF67y1wsvwLqdegOaEsLcukMwoKliSQxwv8k
o2f2xSTDKMtlz620vqmD9mKvUxJHHwJLXelfrrnSFow4heBDl7G8uDHEQsMWde/f3v8Bc+ba/ZTr
P1hch8Rp87AOTy2x3AQLwX7ziPtS+3Vik1Cz9Kju+gR55/Crna0sbt2s6+dW7N6dItWW4795WUqp
d9gwxBFspi7EBmiixZDYq+wf+gS/NFWig64mVZIbznZv2a4ZmeQ6u531LeDg43o/dMFSmNrQxax9
u1MzqRnN3bOuYQsgNnbnlXP1ZaxapB5kzRnw4GOhaKSna5+SZmhjOQ5jOUEUuUW55TevIEUdMnVY
F/KO7Wta7ubGX57ls6kOaMEeIRN4gM8U/GsLJA7iCMjmsBtl+I0SYJ+IGLkib/LseMGQv6Nm1feb
IqDIfvZbhi6etnK1dYErrNHPHtCHVQUorExXSsSEClNyBR5dg3+FN9pkNnemuxwbtEuKPzN6YLis
CwFYwO42KWJ/Jwc9LrghcHwpBRsrPr7OgmwbUtvYujr6z3YoG76HxPJr/rLNIfRPFOs9zd5bHb9+
6vMKgmw16qEnjSA+7kTmBx3/e7QMxGoZscUWttOSztUZxVndIWibOkfDH7CpHDfMk+2jivCEZ9QU
mVPXWdAHcvz436NIr71pZ9Jc+fx3xx4c4WOKsCgbPy+66eFxt1BZzY471iwssag9rIBh20t+8vEu
26Q3lMor5G94CRsXZRQo82+sOiepdUtw5CSiV58vghk0Wop3C70sciuPphf7rX9sumJ48vgQJrdq
0GpmLbaZGZ9PsuUrbZO6bReSZYT60wivFAz8eJsGG7au3k9caFzmBSuQN1Bxhx3dox4LMWtkuknS
Y83MK8xr7j4flPTK7D3yxRVqF+s5Z9PuFz/Lei0+02GLoawAIuT+55C7k845ouowh7z0hjSKJcUB
7jmsYCrA1clF4aatci5uAubDY55G67QKe9K2sOQV6fcrkzJv8OUqv9qsQEq2cDPODDqd1im/DRFu
YyMGKsYUMoWojDcpFMNKPdnmzEc28vBBqvmRJb8m2O5wU45SygM7WBgc1pOm4vsLZB5y+mPtAvnF
4C9KcQjsOU5d94oLYULf9AmVYoqXCYROTpc3Hwj1BIoFwOB2h59QdrBg3wm7O0QfunUxgUWXWHxa
OVPrIkuoiqmEO7iHTZ8Lx4Wst0k7i8ZT3qCIXkPaI2ZeZIMcYa0PK1e6gYtNOsF6cLzL15OfqzLq
uio7S8L/YWvXSz5wGJrI2MJD5SsPl5GneVEuqPRBmOvBs2hghwRm7YtE32Bo9kJO9APD6Ks3Q0sL
culpDI+obta+24GV5/cpF0mCfFanVatgdlMHpy91PGn+2JgGS3RUcrHdq31gY9y+1MTMraa+NfX9
HIbG+AkPplIMRCRLomXwek1byJTERWAZOgnvQehXVdTdM28SDT9XSGQvcHUet840PJbcP7ESgxhC
mDdP6ldNVOYBfzrH3ZLC1IO97XzrU+llhdsK7yAfPu6AM5b+xNPa9OfibGcA7dYBfXkLL84bndHX
fpcjOAx8yVN6LkMOBCpcPTiv+4GUTi0iRqquCHPHnIgB/jBjN8uUH/EEC70RNh9q3Mifqj6dtCNy
KFpzSOmU8efTwND5gwCprgbej29KUWkNjaeaX3+9sme7vmZK0770P0gtkyW64SWTwhQ2jbc0d5NW
axkz0RLK7DAkFDsyphxO5U7DMc+4R5FNUEtHUzOJJP3U84Mu7g1gy3ujK5w+aP/2RsvJNPphbOtd
09TzdLVfoolqG4PCy+vwXuO3SOFitDd5e8g+2EKK0lVo0F9rRZJXrWiwAbgSEgmZ0SKupT6XEC42
M9AIRVIaM6r7K+YEuFdtwJeYP4opZFdI+WB3bogtlVDpChEXBSs11D/GhSnyllSJpRCpwHWdruWu
0k14Lz+IsSXy7PZ3SZyDKQPyx5h/85YN57aGRxp6Y7Nuz+tAnfZeV4UrMoHs9jtHpWrCs7rPIVg8
O5cWsKnQRavtkUkCSWXHqMg/pzVaBz7LIx+MLHcBfuZ62Xil+TZkdfXxvvFnwZQTF1b8YIwV5aR9
4tqUdD7Eq5Y8ION1QfW22vArzaNKZxhBlfQ02nIDnPzcKhWUrlhWltWK758wgBZ+6Yxa2vkd7XNC
yeH4YuGBX8Q/aq7miPsOw6o0oC0JK1rf8xu7fDDRmB2ap2x+xP2ZtuVPdbqNSD/VTOOOatT1U3Wg
HcYrl0+B3amJ26mGVPKTvMMJKvvyABnUgullb6KX5px4uATnq9KN05oGjE8iW15R5ztbqfoHSIHD
il92eNDzb7X4qJLpAIxkri+ouXInsOLexTTBF+kaJC2/69RGKzcoBAp4W7UK1/rN5sXOQZ72lJnY
i+pK9/aIDoTPyox1guYuxM7GcDOa3jA6Uw0qS/OwKPUfu/Wt5Euj20PmTEwi8Y0fvVtgjFvTgGEy
WicPYZIC7/VR+nebpr9NiuZtt3zl7yaj+FswRYBnVvjEa3XtO/53m0vjr/rhm01CMZVNOqejSgAQ
chW/HIgiXWYr7j1SSpE9cKf2gkXDixmVpdlYyo+ssz797KymZEMjWYtcjf9vX99/l9mNGIN/5DL2
ju8ZP9O0Fg4ol96lNNo5yXO0YTx1HvI76mJoNw8ELjCViKgyAohQIJBVu5qxnO4vGvJDRUrIDSD2
cQmbtKiItNrmpUp2mGEzY+6TYNVdY0dJTGvKoNTY5K02H/Eu4TUFH3VvcTPjoZfQgxpgA1SDqhrV
H5Ww0Dy35y5JJr5KtALwyWXOOkKnBanCxFs64qAQlGowpgOd+k9PxJHYpJhq3aWbpmPpBSHOQFjz
Y8NcxBf1eFoAb14LNy+xtsPF2zV0Hfy9SaOinss46CV28KwSN82G4vHF79yqiMGlvGIGgfndnZyS
orVeKIDRKi5d0Yl8X5GH7drvdGJDLA6+maKge9wu2gLqxsrFbsnvGtTwnplEwluegOiCevDNmRTM
ZdYAF/Srr3Hb4ThtRnm1TKMq3ptr6hEyAzd1NUbPwwykDrRFfzoEbCzAeFbJXd/o5s2nJlzbHMqQ
6MuLhHYbNZWZ1+Brs7N+IHwsl3jCHnfc2mBxuqGRAcVyY64UA1m7QzDZkba7vKPzboA3BYsohMjH
2Ked3uE6ZJ5+EVlhb0e7nJDs3m3w74X96fl8IQ2zzPGrx8reCYhZtxJPvg4CORKGCKAjNxaKy7Kh
k9h1R/RRKMZf8Ah55K3lhZhYwy1eS+Q+++oI/GLzj/ZJgZMKlp2wee49uwqUYN2s0DSrPU5q4mOK
E5WQF5QErQPY9ZzqZO5dtpgtWXTy7menkDwK4OjFeOwKVQOgh4oDepZosSaJkdDBc/3bPlhA/t9Y
RLFsh30nvWR5D/cB1PTvTrkUkci9Oo7TsNnaMN+eSWL1Mvtq2y7kTpPIQA4SGLYnPwOfHm9Dy8ND
xTPnP7MnyUiO6uATpwlqAsiCHOs6sGgNf4s0Y+1XuI93HQkU9WuveHRq1yVFFvqelV8n/uwu581l
P5nUJjMOw8QCppCK/Kkz5pmyCrx7t61WULWGjDLtM5RXKpG9FH4nfCeCQ/LxMqpuvn135Vs77V34
I70BXOmR3toGfVVefg4vQhMTMsEGiW5c8w823dDPazaU71sVYciORM409c44R4UQKs8KcGZvzm4S
8gdpfwddXAd4fPSxk8/KGtwoR3Ts/rDCy0EBqTbyJfMfdEaBPWuIiK+zFJwZhiVKyCO0yBYADrrj
Kf0YVMb8c9rYjWnLLANAHICGT1RONAwNQX8fY7wKGaE9rGolDej4hThSMsR/j+X0J73gXiSSrCCX
WxrM30c/fBFo5z6cihPFIot4ofj2rylcm4CCtuzFOGsf01tpOJxGKVdowdbEaX8ExeiBocI9zTyf
HMjltk1blAT+fr9GD18pvZ51sZ34XWDVZi1RN2MiM3md0Rn590LleRDn9wCFEEy1VeFzzCSpBJh0
fevIR0+Up/KPZWwDS0CUc5D5qCGByoRMD/ifUFeCIF8Mue58wiONGj5BPtUJRnMi1mDCT+pOlRyb
NglXsWhjVfRHsa98c0voh9WNV+X/ZAY0iT/D1i5/+YfmVRCelw7hguutl+iQsjjdmV6kPf7LS4HY
fY4yjJ+i5o2YkrVUmu5aEzNTfzxYAC6n1E6xZlHJZbTYmVBrbudzWZTtx6N0A+zV3a1Fo6Iqd3KN
6gsx5tcBixMfMkNxG8FK7erbSor43X/BRUeJhn7Fd0k/4sPuN6U5tJw6XQ5c8rUPM/Nt1Vyfrs25
o5zygWUHevHRMI1HSINpk4a42cnQ3zJHSvIphiNmi6qqTa/zN6tgDAa0cmQtbuFY49WI7UlgFr41
rD4RZdJsVl83/x20OxdqruCKnU/VvPKedxq61xNxntcyPsyEWrUhq64CV6M791E3nlTS47/nNSpu
OXZDiOYtGE+OIXgUC/VQRjzIg6ntj+MiSnDVhZCGx0rIr88nqvzOtzCLWC+dCFPJ7ZTskRS0Ph+i
A/3qMakKC7TRp4+zR7twUDs13bKpuDOUA1k5gOXv41oSzc3BoFWnYRsmcAC7ipfLpvANUM0cOcI9
10GZ3j8lkaJXbiq9VmSphQG3UtUh4ic8LdMfHzqhVarZHZthzG6GQebo39ei3hskPRNsogQqk8Tc
YlUw6ZrBknkqWdz8TBi8t3XWiPfaPCG6KeAUCOTiIsgthkBMzR/ToyB1RIiPiR+R/rwvAtM01dJC
zVjoRHQro5aZ7DO5mRSMCxxKQxUlRun7w1uB6GT5dMGT4y9DG4SuKl8HGv0WOOlrbaefR9I9FrV1
E8C2EOuu/YLM6luz2bJ2eV/LTJ9aDM0VYJO2T5bT49g9qIWk8jD7oskneEMOvN6EajxtGZb+BZYJ
r9n9FnrxuYcrV1c9umU+Y6pbrHGCQBis322D0Kiwds45zGARhfIQVOh7x4ctDDzFr1hz8P8zZHuP
m9isUgeqnTjGjxCqBG3Q+jKwPjdluLOmh9Zans79ZOCBuBLsBFDOKaRukvn2HWlrlYicfObz+Soe
ct7sMVjOHTPddyZcGb7py5AqTwDh7dsu9QcPj711IhRPJqXyOlhvbUbE7GJ7IJ8SYCvVzRvmk63e
kBukcwR/N2kXn9kCunmygOpSBWravsOJvPXao/3U51J8ABjo3s9iG2N1TcbG+OEGNLecnJH8OL1f
1v7vbMXxwGDisY+nfwzNBkeJD+6R8wVQsJDO45Xvo88MzrNfdxoHEatUkyFx+8vPg/+SCrukytDG
/RQUD9GMgsvbp2/sCqwmn1Dz+ajck6J4p8r/e8jTzqcRLGls55NzMw3Ka/e4KwUHGg2s5Gt63qkC
31vjutmsoRt92dHCT+u1smkMSvqRfnoLEYKmDQO2etKTaB/oWNGRf4nKBLsilErRGqf10NHCo8QA
K6E0Q7/HrIUj1J7MWeGmUP7D8ZHRVFVg3K0LaOklk33+y0Ut/CC9xTN1XFJIvz8JQi44pMmvUuIl
U+kshBh95oHMVh+Jvi/UnwSLh6AaxgnJZdKxnWOEcyP7HziPJosUwUFSDTkC6QigZJCN5POFocYR
nzOBaMJI/0xws4SQtPIg/2fxBf0BjLmT9m9gSHW7qjTGKeO0vwzE1L2mv7b3PyJzP5ndbXAZbKWo
yqn/uSRy/31pAxGDGvqxYuVFQy1WAO6bMe46tnvqUldFqIuxarEase7Img5VshWi9OL+Qeyoncp7
ezCWMe5jLuyFsCpoK58qUnKl1O55ydwEoyy8/ATCdHM+36Ygm1YPrF8NMvA7LWluf0JD2l4vZepo
xjIqI0578/dfzEjHY+zICjk6MCDvv9DENW4H8LrbWBirqI6yy/vUadKsaaVkVle/RVtNhkY3AOXf
m+besLngtfFA7dG+eFZfUZIIoyrT0Z/f3Jk87QM1nssiP4a5pE8FD5FJUZlLazAhT/FQHI2wmWVZ
IYm2jalFTJFxFo0ZC0L0+XOCJ/3ht9XQDT+OePIJ/+tEH3W32ASF4fobZ56LRdIu+Amd+GKFwAJv
bO0ULm/a87/NS94MO6/FlRGam7+55WkA1ujWnv7Dl68irBe7NucKH+yEIWw67e6rYkLdrTnZqKMV
IfxTkSqt7ktCNagnbGLPSnYMxepEJ+SPL5iq6+8zkgjRXtGIkS3+0zjmMatYj9pq0b3UUNLOlKxD
FpdI7lGc/3MN0AaKWmtiY+YECAzsSxjfPfQ2+HS93tqy02l3rEIfjnradjobxpo2dNqeEJpEkuMY
P/dcbjmPWvnKo+Xuo/MPNf7zg2rs7AIGfsxu/hWeYltJ51ZjpSygpzccawaWnMH0VIPH2DmECxXp
btXNCG4/xxloNmhohZpFhsB18pc21jIIAOBIQDTAr/DhmiL3hTTE030mELo8khy655CTaxw0XzVe
pGKTUCJ016JTyb4JkZA2sEx6ocBU0vYVuuLxNhzJW5tbODsaC0xM0OXgH3Rz39nV+U7ExIkUZ61e
BfDWrJoEE2XJhyqFluVNFoM9qu8GNQwOSOC+dlsv20kv6dFMzxZZhjzcnq7bBkBiw5nBxCyJq+z5
tZJfb/S5lKvmibuy/EeGfGVb1fxZYOuOxxQLWflrNxHiP60LNq6d3F21YKIL1UiyObJUfcEs38be
Wno9+JBZ/H12OxnbVu2kRqIHFHQOO9ivTJH5stKG32V5mzFRRk2YWOIYH8Jlj2bUm3fccyhlgVGv
kPlU44Y7kOL2jm9KDOeP7p8TlfESiGFbRpBkVuknLNDuGMHgOu4snsir72GSEcjsObOpj0z1s+si
l3cZ/UZUhL+Mjl8RA14WFOcdzLr6i0tOwxev6lnEUz1dysZpeRd1VByx+dOmeFO+99n6cXeFezxf
yvrBDH7kgo1XJ34dxCGX8rsN19RCRaC2CDAtUeMEwbXuxkVr3dZWZyq/17FS0hsTVGfEza01y5dd
BHeD0tXxGc7L27iMibbLkrUf0vC/D1VqXyrWF20CjtHAwgUK01oMXybhBgK4dZ2bhUD4FJ5FktH3
PdiOLnMl21vuKLgs7DUN9HN1Bz5hodwfVNqCsuWNIdWQvh+Z8kg2T81Yx8Wh8Qhu09rGLH53w+Un
9o+DypCN5iJ+k5Oy5spDKFqjqh6HurwGY7iY+3z6/wNZWqnuBbXGR4SaUx/Fk1oPWaGUTGy7F/da
swepX7Aob86PJDJLdeEEPk16DRZ9+etNPJ/+0Kg78VxQavr8XMZJXwCvH3HQmCIH3m0im7Rg2IlB
6eEBorREBUg50To6rx3vO/HDix+plSd93NTR8WTnfHc2eJNRYrIInpqdlfzy0CUU7pTR2qOsNil3
jz4xOA1d2KTgNZz1EFvZWlLLrofq3QOp1X3AeEziHqa3Rdo0V7RRP26oD7du/pL6/Ry+76zwb6ed
/o0Kvl8sj0b1b01nCdfS6l8bBltaW+O34p2xe30+ZRIdxBoYTN6umVarMVUHULhqDdC6ZJnPIqCP
Z4u2vI1TzDAHpBDGKuSqnLINxTHCUFTX+GDSRgKJxDY6MzNS7MkMxwZZtmpseHMihqipW1yM1sSb
fMxJzt9KWjx9L/PkUu7rIz0auP8MeYEBXRY0N6B/KQMifMxKIcgBRRm61oHxa76Ok8L3OydkZbcm
lamPOtyyNW3iJ+DFtIEmtJAoB3BM+z8xYtWch8b8qJ6Kgkt39pj19lrQEY2KcMWQRk3z7DEt5mA9
gsJn1wyAAX2hFwtLXa0ctMC9lRuLwg58ajD3WugXK0YcBwBG9EslPON+r8FIY0Br119QO5YIdjmp
fBp3k/eQIsBiYJXKifeqkXpwWGl/iw2JEOC7m3tmtPJ2fbDa5UvfBNLUl23FMldyAcIsQQadk6UZ
F/nk28Zs8eavHf7zaIZGNyQmrlr+rgaQi7Zj5/fsUVkbPgWD2tz75IsDqWTIxRXptbf0HFl9a/LM
z4uLE6HhVW+sGI/ZDdymTQwLR+ByUSlfM3jiEvs1MLKzE1JdEPDOZBVitaGkEp6LPScLtADFbkkt
BmZLq/DbFENkDTkbEOMCROgq800AeCFRlrVD/dJI2eC5OJBZGC6282NDE5cm0ADcThwUeTGHFVUD
3rmY2l252Lh/Q2hVB2woMd5ZJTnDZl7ZDBu5rCpskVKic53Soq7FSI3RL3rQOzE7S3YGydy3e70A
lAIdvejxIn/hMakFeEvRkGbeS4Q1dsHN0BKqjJwrUTrUp9op1gdbiYZTRh6Sjx2EyJXBW5qcSimj
1YFIV2Hlu1Zy6DPZ1G5ambOF61d2/ohB5blntEDbKGS8Wxc4ClllXpmrqXfcXa+1zYuwwt2e2wrN
uFkgUPHzssaUbS72IDghxkzA4hkp60XjTCFaTGG37j8ZaqiWScNG0qrIutkik6sgfV8qwFCjKrLT
AVO9cDj1NNQdzgm85zckvd3VjinvVitxRI3XLo8mTmwY3n0O91FBm9EM2/Xp/GF1oCRW0D0rR8ay
sIX2k+bGe8kozyShMx1z5RIe2mfeq6ddhN8f//Wydk7RbpexUDCVGxIhaoAGiP0Kr4vKWkokaMst
molBNxA5Z/SF4HKGoP9hHRnf3PNPher4W700RPOG/PMBcBu+TF5Wwv9bEnzoljHljrEchetz23s7
zcI3+teiU1fwbAPhttEvdZl2X5HGAjPsIjzpnIKvOLfm0ZDZLOngPC6A80vRqqkzUYs5e1HWMMyu
H1aFHkigHDv8oQN7blHOiPhsqC8MML86EIOJRXwrgGNiVwNsKtPcn0H/7IbJpew+AC8SYQMLUIa2
b4DpCuM3qGeTIVEc6wKEkB6LQarAna8PciWWRuXlcLqX/8yz4PoETtbqpjgDQPSQ7JzjbBQdTzwl
BwTS78uxIeUlo+xoZR0QGmAT75QQSwQbThkpiaG6BQRA+AbIEgVCiq8L9AdwoqS7qyyXBzzpHcuy
VYNrzZ+EGiFlNeSsYe+lZ/DVVg/PAVKt9L35OQit98tztgGmaJjAvIqnvg0/ul9q5cjIt/vwOGZy
ili7M3hFefRk10dnSK32KlEUXQJxp1ut3n9wdRw0uZOZe1zi8ypALu4Upd6Yng5zVvyIoNSiuIeq
Pr/XeHgm/YU2cnHPzdj6rY+ebBIdvcuexTdAyUOwABYi2nWiLqJn+Og9WIuWk3IfDTlWqrPSAB6I
Lt7rBcBY1siKgQBWhdyQNetE3qMw1RIw8JrhWnS/m8SiZYxj4rsdV2x54uBo/yyfL/y+O0cLG8zX
bgmqs3sISPMXhEuI4FI9mHCLd5GKtIDXWc428YghzL3vQ80Yvm/MuaWAS9CgV2bwPL4wTV0Jw+6l
tnqxQnDT6INs95wym7r1ZoFmwEevlhDkbN2C6D5MBUvMystTY9Mp8Y1zdqWgr3r899QfHFcKtxgy
birbPiB1qLMlzubyYP9U78oxkoUjiBIodyXlFLkZL9HYzj2dUCX0jRKLJAnVteQhy7RNepwKGesr
T+UhsyQ+HcBFvHwD+voxtFJcNE+YaWUZ5llNloGQDAwFERInd9OgfS56zfNOjHfgXT/7rwMy6sSO
5Tzr3BhO+Pcy3A3h/TV112lfPtA5BMYm5XAnT7aFJaHpKN+eMm2FKiqBQC+mJniR7wWEHL8AzfOa
SjyAl3pCdZ+Yp2UUVOo+6ppT2bkgGyohzCrZRPvFkrLSuhhqSbV0ydx4I3NJPuoWdRwGd1SoojyQ
TX1OkfXKDKabXk9RcjwyldONBk21L4ErCGYP3KH3Mc65Hjti6WvaiQPNL5L5LFaNbux8ILrzK2cI
NfXsIXMQqzvfC4mHULuldRykUn3YpqhACeNocRu/FKZNYT17YaT2660wbOVFvVYzwX9SJlGgDgOJ
cmvBTunWofldJwTYArGXJgk7UxoEJ2oWlpwNSFZu8OpSNl71s7lM+JT+ol0GskwRlFVpNqX79JRN
GZ7nVZM3H+y9bSD3s6jnyRUKuUE6WNtcqCQt5jzaXzMPFZZu9FMZLaqWPhmOwcLo8b6Qs0hH8rVI
iXRMnTrDcBoOjuutUTbsvuWwmxArVYBharf+HTCFdfGKkjvyroy+NhCNNRiaRtVGNqR/5uyYt1nm
F9UW/4D/JARoPWyhjr5I+awsYzR5NIx5p1trbgwAvx/FyQq6RlWAp3pZ+rYcEZj4oqWlOG54crGN
pbbL6gLdQWAvchbld+zQUubnoqf7/Z+D4cDwobBG7DEa45xFJq4O8ZD5CEzcQclXulgZWSraHYgA
y5TLzcdWZ9AlldHLcARa4/i0Z/lQlpcWVPcmMVloX7vaffWnvI3Rf/RCj9KAFNETL8i7lKFo7cUe
mNWVbLlBg8iLw9298oSdYl+hTQAJEQE704wEYITjxx8c000eyC1laxAR02UHiCf6iJOJbSaSaVTH
XiXF2sUa0N15P8xuAwjkBWL3LE1VbLUPDgdmgyYRdlLkc6/jPAw1jXV8Zpbk5n1Rgq/Y+qX6B2IL
qHUrKyte5zPMkMlVCBcLKWA+slReDToEkj8wUlWM4wJ31ac7phierReDd0SG3xHNoejanJhzrpd/
VgVvqlkTl12OUsFhrM/UyOb/tSNkfigyVwmjm+keAV7+PK0W+ifdHUQ/8kf1g0eDSNYf6S00xofw
gUUluI5M6C2/DeFgmdzuGoYdQrn1xdvJZx/71YC9rihP00ucQuUt66UeUFaSDpLUqDo8C2DpDfyK
wr+sXSXC22xMqZMd6nJqwvT2fBs1yXZSr5m4X9dh6TGAIw7r4xj7Ehcu+gcIwViHnbGfchaKlfTE
lpvgyGKRHjpeZIe+YeRmQ/+lnyw3NW61BrLxD/jD2pneyxxaHEhRIDhxGSShkizxDttDvmqxVZtO
4AQMAQCR3hqwbdeG0/P3++J4n5L6cf+ljcbVwlhy3/vCVGqkweXUc9s3OBNP8FQZaAaHmVIIYVN/
RTHI0J5TetxSeS60Y/du5niSg1WxIZwbujJnDHrttjnfCDGX+dDqQgmuTpF9kMbUgj9qLeEw3Git
4UKDgZ6fGQPnfwZCPVip4rAFAmz/UU59ICqjzTTxTewa8wyZea4HEojyMQdmZgZo6FkKDD5zNxVm
aRZligL5EZL2RXXii1Biq+nfpKSZGN7BQG6W50pspIuY8XPwSYVwlNfok6URedF0MVfSrJJ0EASy
Fsp8293WXzWaeIoPHaRrludy5rhXoWQ15Rp9q9RbHSGnptF9cN4Eb6yqq2M6EpTKDGQ/hj77E7ov
yfkpXqF0LMGrmhTLy/EbCY2lG6q04tBwyqEwZaMBPktmrWMS6TwUDAjiRORldG3G3Sx7RY0P5fUK
fNTY+wVz6GNhza53NN3UC8CegHfhfAOIr3MzVhiicbbng5AvBHx3lis1gXe1NhGeCMCDiuRWBQew
7gTXsNGr1tdIioOyOmev4VgjZ9ZrCQobIlnQ057/oEWyZJxdEY+AJ8vR993k2arj32r3nmsoMWNw
THb17BrJUDRwYytq4h6ch/kz6ld5Qit4csnYBAgKI+ENQYxR70ZS+fOqyPlDjXvP6wFRRbInUQCb
7s/h9X8ocsfJc7awv8NzjfDGmLTuO9+GNb4yVzR//BjFOoe/0TGuVtkpcvnpjhgl1bzw8WNaJP2v
XpgdJNYzMVg3Mm4aRLlzlbLPioMXQV0kRdZ9FyKVzZue1qsN1xSoGa4ZgT7A1PmEBkLvjU5Unkju
cn/VN+dU/zK+801m0rfZ6DT/f+DJsOcNJ0mGk2YMW05xI+DDKKSrLw/VF3dBgPifHPdICusbBNtT
jxFsq0wrIuGHh8oDhFCC3w51tKdfZeVH7jnz7la90tGro6SS6VzJo7L3lgcvODl05Q+N+CaCO1f1
wPqPVS9BLl95UsZxpHzv653J1kJa17eRtrLJ5rMFT+6FoATjKr0UZdy7smDpMDEurjG31btoQfQZ
4XyBFhbOPR876EBBJH3i4Ia8J3/3puVqzEUf0Bz+Q3d6EgTpx8bHFXvQBgDgyXrm1G1aIYVEtIQO
IlqMZP4w8RhaYezGcZFHrqQG+MuYbrQNVoleWwieTEKce1PKKNatxYWHhguz1SaIdFWgC6MhqFrq
q2TFr9CBFb4jc9tst2WBBwODVf0tQ2+ybSEl6npuyF/aTktSlkIs0TU3W41bicQd+PjyZYgl8CXs
OEyoK1hMtlAK8UGxgFdmd7BVWijRTcJT5EpcndhfxE6ETyD31XQTeWT0v1J4Oxl7GlYLEg/vad1d
b9zl/H/u4nrSoxzypo1cxfxBADfyTp3tKRKf3RH0j2SbMBMXJQDG/P0Ounswcpp8634TS7d0nPc6
PBJS/uHwTYmKplZny7KqRcfDydvtOIcz3+6jHdVXNQTgWQ2pJX3kWH1YRtTKqxv8TOUsxYEbub9Q
oBJ/g0DgajWfCWudFGEnUkiDSTubCBykFriHbU93Xvx8hPY4JELMqU9yC1zJ3lA2ppXeDFU2CBzp
rqinXE5Ze0LvJ4NRJIkd4ApX/WFeGBhhqwtDzo02zWtDWCFMTgkqgFYzopaOnFiplk4PAJvx7eoA
NayRncgwmlAI7H/jtW+kDVXtw/DiU9FT5FKLsxT3g8wzltCXOFT8BWycFS10tT0Knt5+ks1uNY3D
+ZEhHVyZZKlLEcnfIy1W4kEM4R6HyzrQXi+LZoiD0s9WwWWbfHRZmtFohqd6A18g8vIxcpO1oxmx
iFeda18TJeB4vbBOD4kxHhPaA18W9Ju6kb5WUW1YD7JpBSyF2+dxuawV2E2CGnPA1Wflv/PXQXAP
Ldw5ESbSOXWjuSWCm4O+v6uAcVDLoxqItq6EAvLLQaIUUknA1uNHfDRVm7ZX7ML4n0HaO9Fm/d/m
mn2zv1+E/RRgTubmD0bozvHopsl5FaTRRjsn43/9CxJtf6jCE/dVCZtJJgp2XZakEF41lgCeCJzC
Z2gK4TYnfrwP2J4gpveR0uW16G9c+uDcCwIk44M/kFT0Tq6kHX9rGKy+butUhvDsX5+sz/vyggrD
XnxbcInRa+8pe4RnRxi1XiZd4YAid4Tly5vABNY4aAYwMKiIAfvFaQOP609EB/n7rndloaiVx7NF
85xLJuWUkt6wSfMT5qh4MzMKNSw53uMypoQBNQeEpLrlCz7KFuDrCP5A+h7bbpsL9rOO1o9PzeNi
S91W0asgf82EQQr7b86skt9qslp6XF/gaKJGsQytryXBG6tRi6BX25UZXc66QtpKkXC/LjMhYGOu
TcbRq8wh0xJEw8nmgX4b7COOsF/2PPWXRLtHOrmh1aHifUCC8salNPPGK9cKEEOyWcKL8PN8wRrz
lherU9xQw6ynY1BK4QXykXeH8KJaRUneWHrHEnhtGtfj1m5CBRPYVfRjQTOsHQjKiNpWDXAxN4Wm
JUFEiJaGtiZkLGnjfYI519f7GLKUgruCg5YZoipzmEjAjnTMLIsuwiidKCOCSqbQIDImHqCNcCR4
aSjs/MhYEfy0ASFyfwY3K2doANN9h44l/6gWaZq6vjgPDbU0+0OPr1vf06bp1TnDOq7zC384HNru
MWa7E2A6T8VtJ184bZsP4PBO2s9H0iKdQuQPTd/HEkfo4q9H7tHMigUZg/vzZ2vTGfPgxOsXeVx6
r20v836/U8QqGMqMNmz0sXLGDt78QioOsaUg7tN8YwBrwReuG8ryZuQFo4DnE9ZMs3wy/bZLlyXq
jlPTU7/ycqgTCg9vEzBsDuXLgM7Dv93fUEEdmkHjzZHIBRqpF5WpIO3P1OBqp2RIb/rgRegHqxgj
TuNzFym1d4vKQJ7E5xo5zZY9OJFoNGcKz8Ifkmdw22Tp+dgMRi2hGKhnytMBfWU/C6Ef6wHz4f5I
ZkglctSHOcAT03THq+XtCwhEOs4Q7fOwvruAVZWNYzMS0eg28AXvBHug7U20ddSJ0YfhUc0DJ1hk
t32j428KGquSV6IT+aTmzm/0gOZWcFgruneJJ9DY44JfVgTZ/cKQwMbycrDc5AQk2ZDB8+5Rriy4
MJX0lNjhko5+RoD/8Bng8Cp0oINdK5vF/h5CWTyhGjQG22V1LNq6KsUvw6zsQEB/kCWgYhDvo/JU
1T4bZz8Q7OjSt0g8eBt9e6CuYInfxawLRc0QiRbw1uymHzbLKceA2RqRjQTqNppXDcKwDaGAPkUl
rWQzdp6zQSNLOTxyHz7Vhz8t4l8zfnbdMdhyG/zqvpr/rXO1nXaApvtNvpBTtujYyOP3beuEvupX
qxap40MgoDwlPrfZ6QNCW4PMn0o4QpAjEJ5otTBEYjc/F4daxl31jf/sLDWikojQdDnuvuLXe1y+
C25ULI5qSOFFIOEOoL+GZPVNHrOCfj2dudCDZEcDVX6IfJTV69AMOCaV/B0AYtwOExPSqR6QbDYF
CDAjUFm2z0fl3bjcRcgGoWA5DEjk46CNrZS2XynSB9tLAzp4AdOm2+ivQP5b/ReXOOKdf0INwAqd
aA55yT3lvEhJoumwZPXNow0bXwKmsVr0CD3TsQyyH7C79k72qy4+HKbZPCxWZEiZDfv0YVU2Nfdl
HYk1XoDoLxI3lYaBd9BuzS1QaW5epNQz6GgSP4v/TKAszsKFYzZFd0QautanN71NTGAJK8xQBSKK
DdH0Iu5ngUm6L1gzm1YgbicAxa8W8KdMCh8A3djxXoFZH5UywR8Xj9Ybf/CcfO33V9Veec5O3bgt
JudqrDNo/OTVW8FM0bnPq6XIMEaBN/G4h4UbVVfeENiIu8HLWpvfv5KkfHNwrjaznwb6MRmWWgRF
jfa8MqDXQvIbOc82eCkqcR4tjVz88ABnZYUzyD9FAymcCsgZUg4aFMTYZXdklcJe/iCl7ZC7BEYy
7mRXqEKSnF1U+pQWKmHLw5DKJcNfm4RVyonYh5zohatrFvJR/zqW6vggyJ44XS8sdPO1fQLx2bXi
tRmPE0SqjVHKiV/y2wdtuyCBm55/fvnROvp2dmDac1VktkF+j+CW/FTkpWkDBBUChnFjWym0VnZL
6IKqUhtWGZH2cEWcuViB/xaRmUVpPbwAm6xYZoxs5lcxWHtOisq+2UEWITG97MMAQUO3i/awU3q8
dUWWEQgLLWWHlg2wnN3IibBqvB+AK0bZRvAkcKyjLiT32jCwYqd4kgHlEbNKZnTBd//mGNhYs2G0
aj5uIM8dgbpg7AhS+KfR6PH1DcFxI7FpmLoeVj3gUAmKPWtw+Dbel8HMmd4AfLdbFeE0iiFekXAG
8GWEVNzv2qkDBKkG2/AwJdBue0Tnq3LdvAz2HBdO3P5suQ11BnDORaAwFcAsnIM23AQo0lhp+Hdo
/+bMoY3iy7bRIDJppXepiNXgmzM6cQgMOTWOjQPZ4qSFlRd1sqhE4odUOs86jq8yhPu7IDPtszqp
OHalpO3ww0sTju0sg7fhPCDsfQsbPCrbzLPUIICCGV1VrxxFMshZ/nsCpJWBJKHrUKyKZLhfS7NP
bxL0U3p3+jW5GZGygRUYc2BAA7qqfdnCTnjlcQHhrm4quNiqHAQg1r1/WzOAiTTGFP1Byou+mkwY
IKWOLEDMc112VrbXoVMwDWhsH4lnht2yILk8uf27+deBKK4Fa1knVex/yJYn0A7tjSLiF7PDg1y9
M3Jy/0nsvejg/9F9xSj5keV4Tr9SBAOW+vfMrOhUbfBCHnZWThg9fmQl3r3GwBAEA0/MFdwPXf+O
vJANhgW+tCBxtJ+cFNVglAOHFxIHXLFAjp8Ei+OKUbiiSGKm9Y0dOz3mrp02Cc5zFtzz+yGLHGaM
uBIibicAmvSL5+0F+vkjNfJBas8vOLzEUzCKmET2fwXfCIwkDLwQXcPkbaogdFBLDGPULJ86io/l
k+HYu4neKwBqJPpRE3fU/mzQft81Nav+2KLX2/RJoZMmG2/6y71CQxjO9V9HN3LJW2GXOySLMJuM
O05d10C3ylFVEp+f+pCXTkSAxcns1jtn7mASAQqLv0Oc/1+ADUbLYikrhXgESWlEle+nbYZTy5Q+
wW7iUAQk95sEvbEpx+RNvKcb8PV3491QqWu0DCuTlYYsus+mWb2gbOB2v6CnMqqnWjImUUeHJcwx
XkqHWqblNSxAwgKXYfd/bL2gBdHMGba/VbDZl/87iEUElvU7qeTVLqW5sdP0uXq2pmGUAnw8u2Bp
Boz9N/ok7W8RiR5WrnUdL3zH4vxT+wBlDVm9eFa7Lrudgcn/oC9t6Zyq5vhm2Qq4LZWai0RLPLPy
UOgSViEKrrz23kj+povmhxgqxDEbUGZztpz7AplzQg3UvXGMCYh9pZYBF6tBpjFmEB9QDTtHofRw
ixycBsXWur0A+ydI7Xu+ja+n0fq9ru5fVR+IZB3RXAG2/14qBC0Geu39fMFBW9EL3sSHJYxglIBu
dBNeRxQGoi2wJu5vTqzzaaJIbRlyTgFMhUcJlFPJiwqa03CpK1UFyZ3N2DPqqMNyNlQL7lj0jfEP
DysZZJx+58+7jsF48cLIf7kBRTfZ/US4v6kAxBXyR15i8aQZhzsWXJY7BeQDabs9ibiVRZm0GGur
fFfm6tC+NL/3PpbzUpD8P8+r5wyv7ikUu9Q+JKAKCa8ZXFI6+JcqKrBu4Sbwm926jRU3d8F4eh37
Chzz5X1rtSveba1qUWQyow2Lp5XFUflRpucTsEIr1xgu2f403vgiB41f62EWpALGjdAhPYsiQbf8
qT1b8esMHAQNtwdFc959R4yVMw/ezW523L/o0w4YsULRuRHeHxX9B8FsMrM9GkwJnrAKb0SNpksU
Ay7ZDVOklHnLtom8mrplTlIEghnvFb41UglFQyx8Fxhkd0GKJWWWJ+nMFek0n9IOM3zONN5QldUA
O2RASSchkUopHCJ+81tzrZTSntGrzL2eki+173uh1e4pacb/DOdaKwXGB3Z5REUocwSlVeUAStju
b26PrBolZAv+3T/CSQQzcn2hBlPGY+rUjUR1p7PX//OH7kuv4mZjz/JOLWxG+XO4kl8LExx+J16P
ODSpdO/Gt2vxB/lh7PjKhD87UmCtYI0P7gntrBvu6WE6+xElg8HsK8e66BoG+ALJ0WkiIRzJBdtz
NV7SOhr0p7BTsLTUEbUdk81Im1y2pAZLr2j3YlO07KFJBkjpXBaAeE/R6i/gcYECMASCn5Mp7Jsm
87D06LRWOzUQ+q/HoOLIOyf0DnNw3qWmR/5pTC6Xo//EM1RUMO9oRPNJIrpBm0g12E4Es2CiGjuh
681g18FeisRPFbTvN+19rJcpnt/atbYt3HCpoFS/G1RlQX4O9zjYpi+8VoyqoQ+MiZq0feD8KtCF
ufM2LcxOwS2n/dEzHh0zHDkJ7ZZpcAl8Kac7vnVyuPg88CFQm2QqhII7mmWCYV3yhSVbPPB+wz3A
j1qKQuRZFZo0GmnZEo1tihAUHUYoO5jzPvfPAf2xZhPW3BW+Ub54P+v7p8s5fiz+dIlbjs9Pet9K
obcLXUeBnmWSLph0babSzjKNLoVA7dn60VZxHxh2q+0AwnzaNAa972VtSzMzgvw3P4fChKL8zntj
V3e5wEs8oovUrARrrn9NO9B/Tbn4ak3PwTkdwP9PLYb3+K9hl4QgyNEnVspwPlXNX4LaFUSHJKH2
qrbJdSik5o+yflDW8GZPOtJZ2CRHCRPJfNEd//AoSgTsaE9PNNvIpmmvlvjTG2xX5mCIS+nw56jq
aARZMJOawvsvMd/uC9pGyIkXdo4bWqs3hYNZijWQ3V0FYDsbIrjNSkls4r0rpPoq9cjOxKkZhB/j
vnAfKD7BdhqCrw6tU+/DHgiAG26u2qKskGNy//vs68MKEcqRHDQRl6Ib2bXxzLDFRvpjPscYISUw
c6tl/j8z9+o+L4ylNWpJCwX2VaUuWoH+PvdX6KwtY/ZG1HkEL33qLs6tEDOMdN59UmKKtxUL9AkA
orv9HI44030eilP20M7hL7I0Im8bMeYsp/Q0JReEiRhJRQz+btKnYhffBOPJYcNWIYmW5Yzcef/q
OlTjxmqbn/jlR8gQKGXBr55Q0Y/tYG7cDUdJG98zuhiMgISimFvRr6WdVKaWFpOrdNuL36f6PG5S
e57dPWopF467CFn2IFZXMybOpRObAinI9IiGfuHAs3GYQmST6NAGnz24G6uNFbC1IyF7RvtsjKy3
jKj6p5VMdh/xHp6E0/kcA0DGwe9tr0ecmvnvACLs7HLK8FMGrhk8gmgha3TgrEsIAoVsoAL2ju7r
18tLgsPXbYSXFkyIXo6MLskVfCTY0jou81c8bI+cFzM40Nrq8w35ZmdU6zX4NfXcVTS7ayq5Q+JG
+SUFU5qZIIFIZ785FUw318582dYbU9Laaby7x5eD2xk3t0dUecq66H+o7cA8dVEHNIAcgrJ0g7Dc
n7hzbfLNAaTPk3TOF9mLkeuhXciUY6Aw3xB/IUiAZ9XvoBAjlvi3NcYLEgYtkuyhVnY3rK2/SMRs
OL5RPpViHn95OuUDWCrmCi97ciUgWhkUl2kw6EJM2ttSYikrUfn49060ZCsl7yDLPqUsItgDZW17
0XPPGj+Es0ZaKNw/BvDHlkFJM0zsbiXNj1YwLaXowfb0sOH9RjExN1P8TfZEYJxg4d9M1ni/Bz0y
lFuluWBjRguAuxv9CXVJ7y23UEAYydf6pQAhrG/X1Z/pBZgOuMlL/t3C0kgdW9MPuFi7RmvKvKgD
c3zGjBxJGMmSqrUQlxNaP2AF15I53ItPcgvnDZKcKc2LDCCL4POxcyPppE2yLgAfY0CS6olzZ2d/
X/xkarA0R6Tp9/3gQmsX9K6dMRsE5HxXq+pR1rNprO4QBSpugCxW6k+pwWs2KfgYfiLiR6m4djXc
b6GZGm3P2T5iIpGnyYDJFyvwZnHU8d3ZMgkwQRbzf3bKgdztDzcolHo3vaJS2yZq/HWrIQfBWVmU
j7F+RSS9dQuc/H0l4VRln02PQ2H2H8bHVv2fy+51IrPxuPEQDONCks1fMjCX6vj4gWdz+3i10J6s
yOjZM+0CM6veltzGMmBJ5ZQqa7T0yzYwOq0AcHu2KtypDTGhPUuNhh+efqPOOyEzmV8MXd178PfM
tPiI3lXBcOAnjaPuY1O7urmlpmt33HWUXnwmMX1YxBNpfZ4cMCvuZ9cnQnOQlXEhtCY2lmU1PPUb
Cm7B4GONdRUUDrb0+Rg6WmKGuze4YOeFCGdm0imAwp1Qtzfpd6X5dWLbD5oZ7eUqNDwiwHwvdnvi
5AAudgi42Cl8PWTn7vqTyUHbjqUuj7WmjovScREnjmoQEj1/AkGTm53zPvtZ7Fa9cWGscKilc8xw
AqPyrCM01+rYFljpUUXu6JOss/C0wSgJEZDsy2/qPKHrL8d1dENF5A5CWiBtgnCtLal+PBtT1zVy
eK6xlkVUv7L44IMjekqeAmZ1kXLn+9rtqLoGankufZZPmmZkNRs1aNv9VXOeesXStGP3cjTaqwPD
2ALeCbLMm8+2El0sSjRBx3s7mGD4uIGYXJ4zaQpbetEEOmok/rJLLlyqblZ5sYHTDCeVoD59uU05
l4yzmHkEd1jFelFdZcCJlW0jAOXDx0TFckN/fT4Qa5kgj36ef2D6QwET/d6OL+mFKtBxbcx14icB
3CV4L2c33Z5BDsQZoRZuBTc6ah90vP0ju6bwOia43kChxRlnt9tVHTK0akOLdL30jNomA8cLj0ey
VX2Ldz71QdjcSXZtB7ahCRupArXxZhJqniGSHrSx/BJ4vjVsqecRLjQXaBGeH+zPKKS/OK1GlbY3
/mdiJ4ZodHa7zPBWbuMV7CGM5RwEdphfqVwM4U3Ox6xXTZv98JqyxZzrwJc832C9LsAAeQnhW5QA
yt401ix6uod2y5KgGYswvdK07S/LJ0cijAcQPEBwnEOyA85FlVmMznc22sTOu7iEkhm3rp4KAFEp
Fn3mMoJVTtQWop8a//CI+evsOGFJxY71rxtxuAbXLiB+rI1iWinJBu9dmA19LLDEAqKqszLDysK1
5uQl5cBR1Y0YEGR19uFc3Tng/goTlSMqZiMRvavDhYxWG8YfYRuhISmqMnS/xin7ug9WOSOfoMqE
8mB0sKi+k7ZSEUEbDWjms/G/TPqAulo9WX/3kD/fNHl1Hkso278t8FXoIzWRNg6kP+QYVtMaeIot
2zzuxjk8665EkOJYUEgf1QNBe0F6z68Nwbyw3ysyUV/tBBLGzZOhAnmeDCocfquyTQQo2TrXGtvJ
ip7gRd20OQTTkiKvQrrZJMA5LySWBLliyESL152GU2brJXjDRjUOopVziNtL3ovqghjfC5Z54mgC
3w0J9K1UrrmvKxbO875HCfG/ugb6rZe7YkZdHZ8OUg7kmpfsrgSdiAcnQ893o7i6OjPK39EsYcra
VqiKA0QTeg+qA2kvrvgE0t7ucEe9p9UkOGt2OtNIwNOgAPlO06fxkWPLbnKHvgvDKeTdzaWbh2KD
r9VWulN+60mx42ksmfpaUajC8/c6a6euUw5AbT06BVo/Zb0ZoEy1YHeKHmE0PTmhTXxR2o/vIQCH
cu6q6QGKFCaVCHVwt9VI98M+mTJeI8nVjIBkM0yGXw49CgfRfbxuZfnE3vS39Pj5P2bNJ2eozewh
ThntNSWBaL1yWHHcVbaMPJ1GK0xZc6NUuOTkLtHxs/i4+X4zxmWIB6ECdXnsB5NY8xd56NbWqUAT
atC0mHz/4A9Te8QQC8FFoo7bEBLXDllNthvpjycxSK2F6d1dcU0+xvFdNoeV2gYUhHTSNTxcrYvZ
MKKQFwjaRQlqbel8PZycZefsbjOAVTGHfOe4VkTRQPVEHugt4yVc7dJNxrlo+F4QBvA+31RSTmbK
pDQNaPgRgeJNwPk9s4t2Geza0tVNQqmfHXvEf2kHggL2wf4h5qz3hA3kn5T0aKOEQZ0bfAapKk2v
v6347r//nxWA3zEZY7NgMDohD5Lc3yI0Jh7F2PNEnX3CW8zpLlC96lctmN2jbvIybP5ME1LEpAm+
JMV8VfrOfXSEHrHqHS3En7vJsgB/5UoXi8lCW6WQvQYVsjDpfayhkjoYKX+0dAROtL63fTVQSjqv
pBJnELCWm944r3JW7Jer8RUtdcQb41aivIXJGhrXFidUc6DfnnfQnO8+u3eAwRFdXiL6GKaTq3lu
PxR+SH8PVVlTNZyHotFuxr5fyIBL2WWx5tS/afj3kO5HOdkPxNmEhT9JaUYhHa9OJA73xhT1PTwG
8XI2OH+coEWYNAT9wyCubsXXj9zsU90dc8gTdY6QJC0B3tmWuaMTO554tsgRZWJk8BYeB0pjtXrH
3ytFLkdzUI68l9L2LY7QjMxbJV5ItosAXMt4RrI3my4dQeLlZGF3ObRP4a/Foh07t4Q6LRpgEbCD
QYXgSPBYsikebr2xeEHrUxUXVmMQ6ubf5p4Clx2vSiSEuUuGA4k3Gw10Lobf5lyerb2bQ58JMQxO
VJwhQNXWghnBjt3S5hqZKYE0ZHlFOwkwwupJPtckOLaDNSx6TxEKnqy+QB0xkV7nsTiyTRI1w6OQ
Tz7abdZtNa3TwY+g5kv86IrZyJm40U0c2/SCmtLJTBp4Bdt90TwBCxO1ZgG7iBw1kPpdINrMKXoz
ptnoL9GnsdBgPLteFf5cJ1jBMJi2o2vLdzRflPnonecpEe6Qg57qaGMDMAldksB2z6NrkjYnHLd8
cqjigQfMog4puCu06MdTdKtaklWAkNdxFHpstMjwl75Nc4xf32tdYV7yQpmfW+w2gMpQhz9S7c5D
BgxJuoffem/qhkUkn5dAA0EFSBM2mc2uXViQRegvz8QRRX8vG/ZJaOmTxj/0RtHR79ovPfHRECsn
ngb9sakWw+Rv83TGN4w3dKwbTeD6nbWbN44MfeJkECft7OJCC311OnjWR2B9gLBgh277egLxnfsY
cJT4tZLyxQGmnbett1xadzourUEek1lUVCitk7omd7nOYLzZwT/nxCK/WKHIFIauhSQ+kGSMEDaj
qaGjVQMgnouz6XZE07wP+rtBApa09B9FJEtUrFU0ZVU6xdKkYaQ5ITUeYZCG2sBZQrO8xpWnlZLN
/lC036ktw07+46c/Tg4EeplCrslHZOJNDIoyK0y3Zg4wfcsKyHzf5MFjDl2ufkXGWFsBjfo06VgJ
J5SuaLdMIZsCsl1R98zvDBpuJTjjCmvs7fUjg7LfxJz4pYqdQljqNTiBv3Udd2UxEgUQRn3FwWqu
vwlqBkh5oB3BZtm/4Yjnye5HhVqeLMW0LxtZobLQxcqGNYaeZPkVbHTWSw03oIuKop4gtWMkqt0T
777W20W8Qm2YH/fN/VhcX/sOI94PIehYlvzL6a+RtYIh6ijcwquRNg/Kj5x49f3IVaB1kSLCLudY
b4Zwb6Z1PvIZtM8grINalX/2IEmiUWhkhddvuwRFc2AJcdNTdumKpArRxdPMvfuwVtQBPM+2cv89
WyZfsi+8NzMZIdJ+gY9u9i4wics9XEi1bRpYU3UBcP9igYIMeEdKrqqKpHNWAQQi4/bBzhRHMO6E
Hn2LGPmt3Mn9SRswDCXO82Nj3lxZlPCWvY+NiOS/THV78Z4wpJUiQeh706KtpbaFXa9l2lCavJdn
8TSO/Am5HbFCNZaCpPmOTYVHj5Sh4U950JnhDjdvNkRZxkYG39eWiLuFcOgtnwBCvEpcDl6hHBfX
bcolHlHj0OdFb7ZLb853Tyg5LkE5E4J+dsoayozUpeq+3v0vn3+yVbnpE5b1GcOqBL00gQMawdjW
vjW9pVO+0W8Qx7ikQ2NTkWczFgIU74cNQjxvUoxzaZpBoRcYrOmQ0HSyGEkmHJKFr2j2bdgDcoTH
tmiWxK0HRELzDm9jaAkOurDGGI1CEuZ9LWYggijEb7cqXtXrk2qWe2pUOmxwK9rHtai1hgo5Ld+e
fjccWWkz8fHsKybJUWXQOxgKl8qHTSfbFs2+e0z5IpCrvV6cT4kKkTaPyA6xAy6zqxDH6TuIlkZP
fkYHWE33J94LOo8djnxaW45cX3HtFbJKMS/NCZF7CtVI/aNIRFDkDQP8MPEt38B4Fz8FAnEODC5f
q1G3PRIXMtvSbb7dhCky36yb0oc8UUSBqnBALiyH/+bpIOsPdPAeqLcAzGfWFvbFoTQ/ayas2orR
U2997UlbYBu6M7zlMe0nLrBIkec7cBY7Kg6iiqTN+2fBeZ4eNFmwuqnRcIDLXtrcQD0Q7IWPaKy3
ww5SK5kLQxD7apvklmT+G2kDYlGoMyP+3fhCvTEaVm6ao/hZomcm7a/nl85679Wj5Na70hNKt8oQ
WWy1gNRtxNtlWNZo1CnYuyHMwyiXKnNL7NN8RvaMSpDHA8YXmOfB3oWuF8nm+7QuWnwRW1oL+yF4
ncELWakVrXxW/ZsVSmNThH7mL4cLg/SLkKCj7VUFQk0p8IBTeXqJsYU/TpM/ETOVBC6HMZ8EV3DL
leFe0VWJOenMRurh1nFmpiUli6Q47o1KEfSiY4jX4NY1ki16KTch+5X5mr3MbdrM9Q7hmG461142
2lrA+QH0gEsuUI4JQi7b+XUE8dsljjFYf61pLj3wli0b6vttV7tVd5nH2UNtDWgVRVqff9mc62Vz
aM+KvS4u5BGi8seFrtkikPx9isXhTCZHrDPxlcJMlB0DISKq5sDIFfF/Cf0ZzX8B2LG9ut1KYwhC
soRvAs9YysB/AZ8C5rgURe6Lg8TLACRFySwpCzFiQlBa44Pq/B2M0IHUD0Ti0nWxFNkIjmRMobS1
04NXxymDoq9n+b3mynCqRLtqByo360rhDYnC18Gw+ObTFmIg8rc/kmx48GHlpq5/hnHS7anpPCwp
XVbWxdJS6UyeWU1fjGn5sUgcetXu5K6KspK3k+sM+VXBUr1W97tvPw6DpssrBMD4HvuM6u0i9Aqx
cj30Oc6W3YAkjDfaDkOCVbf/dr3EWWbuk69bYrRYVfGOVDwmZnvD24yRWzxP1Jw8jgtK/rH1O1xX
QNeslOmxdb33A5MkajgsvJ1aVIcyi0GUJnuenF5QBenKZbO1mUKtfNyNZhJ92C6XsSRJIlvU9ksh
FokqsqQY7ftsV0/Sd+6WnerIcEqctMHZThABL6XIPVeyOVMd6ptpZV/OdDL8BuO0mbAiVn1oCJ0z
1/eGW9IvzljNq8szV99qOyPBM0EGxkZfdn3UdsV0ZjCSqlNViPtTB5zyLaS/1DdC3wxTbpSda+nm
Rtp5Mw814zdX6Odj/2Th0ETZeFJMibyJ95zAPUhwt4T4X5zn+vlYAEBN474dGeMalCAZcE9w8Qm7
9rIxq6yJ3xqsYyeQPQdfyraVKT9gPb63hZCCKWw+lfFAluEOzPqozqxAEyhOjUe4akcZ8Sybcc43
6KKOe89LmfM5ShTMs327zttQoVTujHUv+LEV6Qu4/xLvtAJlb/9o40COFe58eGV23nBTiqlyyR3h
+c1BOivGmbO82VWgZex3BL+oI38XICukpBnM0fpSG8SmpnOupBR4MQy7tMdFXBGit1SKaadFEBy4
bWfttS+PrT/Rjr7CSMb6Ys+lu+eQGGAIrUSrBRxtX0MnAG99VRY6azzxht5IO2Txsu9vfQzbnLfK
bfoRXJ77EQndaHtAQAi8ah77sk9kxDTxgncXOnN83jBxziGPs2YdyFn677rT3Y6QaWCr+pUCIG+i
bMGXuZPc8tczvp9x4JOohXTsf1Nt2owD9nnCaL9gHOcskoutNv3QTBSlLN5+aEXoLN4an4wAFjWv
iaaZIgXl7HwhE/bs49NNQ0NSaE6bsiF19tHjB99Wx+ihbAUyLzzCsrHMaBvaBsMPLOsKztBoodh9
u7eYHWvOEIydcWC0rQGj1gwcaQw6U47lpZP4xY++3obXVFi3vETzS+WvXXkh/uY8n2pkHaRQx5Zh
+VN10E78SZ5bzCKLH8gUjfsJsziIr7dGNhBcb3g592RBZCJD2t1FU4kZcp1tbHw0MQY1XqM++ZH6
bGAOqgj8mmi8rj6I6XYFoA8RVMC3EzXlHncFTR6ASR8VY+A9MKIfQZL3EGcKZ/rQdoucwnXzASlc
FXlIaZO1MgUi5buQhOgu3/pPdCatR+en93jFeVZ3q0gorV9HkoDnglcpFbxnxvN/xw8F7AZMnjpV
ztIpJZnBhBHQv1EyPn04Xpr/l+cbZ+oKzpDzhEEpTh4qqTMi//FPQ7IZEkcdZgAvu0/Alk2IGMXm
nBgsSqDg4Iwh8EECLFzeYbVcF+82ChSbJ20aTHZJg8/mV011Fnp3UsvXhxRXTJEMb0jUDAQMvFjN
vUbty9atgdYcGvpU4QW9NHUwkU3Js7SOTKz+QxZAepyS/8AoiddGMvJh+/byfGCHhDfuY9xAszYA
A1ubm3xrlsdJJwA7YDJU178DV2r6MFzuSSgnG7vf3/Bw1zfkN7sdvio4Ur086fPqh5bvJGhXu5e0
KCnrYQ10E6KC87aGgW4qFSuWcRtbVfUTpUiWcJ2ciQyYuJQa10012ev+CWQpjlW9Qw9Iugfm+1c+
Ygmz57+Y8a0567CD7CTfIqRejt949YeAE1FS5E1Blxwa4o+1QEEvplIa6M32k2MfEV+h1b71SoKe
Y4s3AR8+ADHOurQ6uSZTkN8hdehARd4HBHUMc5jiW4UJ0SleAw9ERMhyea2uxkdixwJDpWNtmDJD
HPTibWVJVO8fGAJyY6PeTdncf21D3/RWDOwRp3gWWAixrY9xF2BzE4JlePhwLCyHochcQw75LdKV
uvQRBfB0nKwTtu7xYQ5kHq9RFEf1pzxgi4xCWRVzYkaLgY7mt8v2Q7+DGuBMmZ4e0UImDRc3EHEL
EPp7BKwhjzQLSIFQaL8Hdd7aSFmsGrTttITCFCZtzfIwNgSnfjQ5XKYsBhrN9jCkrI+PdtX2Xab9
2hkvuFvClBuWxx+PBEruVFEM6jnnUBayfWcOmPiWR3tO2tzpwtx4riz9iCwGbbLGNtmZb/indcTx
02w8e4TsmQTzGsDJ3Nk24nss9BeD0KqkCwQfHDaMF/XSoJO4RCvFWxS3A7uRSSg7bW+YeaVsqXeA
nQPVIT5xzWnQQxuUlFhIXvD8eg7QmTB/GIGD4MRSftoFJNja+Xsu/yxde58qzIts6N89M26aJcLt
8xXR/Cwayk46I/IMILli4NpxIsCRR3PQvh3GCARmqPU6SlGc04/+bE2HpIbnNCV7VeTZrCWZD7YB
YYP6xO9l8kiCjqg9mWOAQ4SagdzQdSLru6i3Lh3fYvn9LY0ZPC2QAcbIhQdjHFrX6R+ED0SlIdJd
DtIHbD9NGdp+xxPKHhwrH/YMlQfyTcjz4R29gD+LvFRxPgYRIqq0ph1KFAp+hnq4s9HzfnLRFE1d
6uWI59mnWYy9kKE/QvWbTXaZji/ixpGSLyS4NlySDxnLdZJxWG+oD9NHaWZtNerg1Zb7kQZcLYfh
ey0Rigk0Q2qhdyq9sgX8Uumf0TTkhooPslpS0JlSa+j1T5S5nKTDhsz+IlfpNR/0TDyrp2zKrHoY
JOhnz2WC1ZE7Ob3wg65GGPm8vOUJ73Ldn5TFKorAWPRoAJC9X47FX3Jo8SnbLIviLXXa/2PMeoio
rxIkkrlVgrZ/S7khJYesDQ5jgRZXVuXVWPLct+76wCuWmZzx6Tp4Zhx01l8HWc++t8IXi97xmC5M
jQ3tSjZ/wL9enuv1wt58vbCt/n56ZYp0UP1XusbPefYs3ttOGZKXV3hs4W09aGwwAuV+FzBRRr/V
Rc329P78GdtFWo4M+Tk3f5dTt7PNp5COO3DJ9W8GMyi74y9W7cI5UmB7vm7HkAYMVhWcUilCpQP8
WieJ7HSKqnq+JuS/4Hm5weKKv1/Lp972nOfPVR+HR5sqFiWZB+SnRFUzbRrOa08tGFt/e9RoMxcP
bMKKx3NLQClzhqAJySAs8hkPHl4yDAbzmRAwkc6Y1t5qZVLCqVUYYe6/KQGX371MgVjOU0MzTaVg
EXVRFdpxb8q9ZHRnLcrzXTo1nW6h6DNYtI2HqzpptfOhNCtolrpMOEyMPlX0GbmmSZqEKS0ixprW
d6U5i6ifz/uJ+EcHiG/qUDQmhG6j8guWXhLQMJ5uD7QFSttqXxcGMhhv/XvJa5j0HST4ZAJ4DpNU
gFZ2HSfzSDOWgfVojRuJSRMaBLgeHxTRWCkrIbKLEZwDK3f4vAXInwKTkUQU4Qcmrwt6g6FeCTbH
52ALUJLKjuXmMpKf7voz1lO9L7u05NfHkcqj1mEp0RKYlQ8VCx34czrXBOfZUZZGQIM+zLYjCb/D
llJzDRyWTaZRWohSXAbqaMv1oz12kALDxYE34WqtoezO6914xQl84nbfk3hd3ubh2EUqisOMkeW6
3mzSiGx7yqeQrYejHwaHmVev26co//iog5U59whTeMKQ57pV3cEhMO5hoQ58wDrM577c3lJj0o3Z
T1zQ3zZ5BFBqVjvs3WPF1+FCCFQfNkQunfQKGGw4hy+H2RnWESpC2EovhALRVqoDHGje1wBJ1JKS
olnyfZYdg/fjwxKhfx+Oq4JvxbBgDae+dbshBMyY9chatTeM9tsUdR3teT9qfX/Ze25k9gDBV0Oz
MOXhBn+1g4mx2sbb2+AGhRwuyHq4BbPZtr2KEj+vyKdb0zssAahKvMeB54+UOuedhHpYvpL+r/Ef
GHIH/wTOomtGAAwTWa3+8YNX4VBUgCebDTq4C7zqzukmP+jHY5Zz2gSEWWVzrQsW0u/G2RpiX7OJ
ungzHtPS88t8UAkx2XE8tCxZgFxdm/AmMRGclKOzY/IduxDYCs+wDyobnAOCXlVxQTcNpKZWQSoL
DJCsd+9guTtgGQHJ97v9+mtAbKVTWqBXLOS6Lc054uVpwXEAIoVBegfoVr/30PsOS7eerF5Xm92E
r2CG3VMvifIrLM8lN3qPrhWt5gDTHYMM4Rov0bHOLQ+5SFwprjSk8LuPWy5NHdFtP3YwBJ1eOioQ
F9XaeLbDDX3bEEmpyh7mELtbU3FmMNm/bUgAezxbpf4pD9nmbGvqyv/WM0e+WsP9rLxGpK6HQBk3
BTnHn3aJQThcvQtZSzTHefiJ41AViTIOlFpuZ9jZ2VRq5nWPtMW18jOk4dHztrshfRZoMbRdPttW
5hwXkURQrdayi65FJmEB7fvnhcx+R9oa0bGTrb7gxB3QpWGbeTroLc17Ub7i1x4QlkemHT8+ENWC
Ok8x5UuOoOnaFm8lNV0Gtz5bcLlqBOaVHFNquFTTlROgWgfm7qAYVVhd9HRDJLqW5gZ4tXs7beS/
gwMV9WOkY8EuT7oifn5bPOhZwsMDYl8u2O/xlPxwx3rhuUJ69ASmTYnlLnaDuzIaYm5+nw3+W8vU
VY/OPKyloezZ5gEchgs6kmLove95J2yp6D4Y1dW2OY57SMqB3fqbcGLMhhKBw3VG2yLHe+DP3FZ2
yhdqrnnzJBD6zosxnlJ6TRTwSZGdllj+xtlfLlV3NSdB+sTjencPlMmbLLgXlcUemj8+mo25ZsuC
4Xnl7kaNMx9ktOqWCVLNnIv7UcfnlF/fkwiz3fZ+qYLTc/2w40My/Rs4b71ifAFu+E7NfhXYWIMs
J0B5wSgJc3tcwIJvPNi1HSGRCjN2GqToyk9cdnS4znqcFqMLg13UYgGudQeXb2Le6blhip/Zuf5v
nDi0dZxwqoa+BorrxMKc/BhJvMiaU8UUqw3PeQjJWRsZ/lYezCQJFRWnybuvXQ73132cl+B+apwU
AGsLXTnmgil3OQVWTMmxKE7ahfc7Cb6mNoiwbEtS0kXOwJDil87MvDyQM+vDrfntrbJEAMFDpHtG
ArhqsK7rzdT+1dNqWuw/aIfJZaaUINgPmehrMB265sjabh34DObg/YdWjbdFagF95sy5PtOJXxVH
qidOHmg4azHHSXRjV9gZ/Qq+VPKJB7ROQkFcN3z0FWFsBq6GUCMRe90h5q7TfLlLTGHmplT7r9NJ
7+J+agvKQxll9kxNeKnwDTNmX4S+3aKAu1hUG2JODoxknEMaRB4Qu3qf/DL9/9bRQrVx6MXahDDG
rPdX2djdYnaaW0YDAQiB5L+JXht+oh7br2j+YfyztUUEuYZ+tcrsDBg67wPQrWpGhHC3+tjdFCRF
Q/AYuTJqezyt5r+7wjGUVvfDcIhCUwNSONzAe0k5nHCSYdeqi6Vbi5aMrgFm1apq/uTk4Ax0UMry
DNHt9wFCjsBphzWD/r45kdhQZWos2VLcKF9cMj1RGhPSUl0J3UBg1Z1eXY5Xcj2clnvKzM8z1ID0
oYH8lp+MpKLUqb+66muoj2Iauahld/+qta+R/LufYfC8XcbS+zd2+3Yfl8JX4F5/brzg0pGT8FHY
Hr6RMiSGVOeuhkgMjDhhd+afP7LdcAoHl0JaYLE7pHFxA9fIeaU1Ycwe10IZ8lt+kLA/BUj+xRiI
dUoWrcEf96Q2Y8fD1kx3Dpi4zO89Jm5uFcjChGMRoSlNRlakzzsxSmpBHgkII/EFFYbDH79X1V8m
vLr+b6HDgr8753t1BeqaEQCrjMU14Jx1W4SJACDuD2NLkklLeJwOlOp0Z5PWX1isQ2xOobrcZKqO
5nBZkw0icDJxfJ04tV6wibxIUO3C4e/Ba1lKqlnchixIyr/xEPwpvG5/LUp1gEXXNtgWeAqCQwXx
3C6xorB//fKaoDRh6ZY6beuwwcmkrUDwlMCzBrOuWLPTGVCkte66kMHaDkX0tNAZBFEUBGqnkjXL
Z6Pt+bZfUKHKYPvN71QJKVONstdOqhja06paeHqpmnuxvulbtOUU4xNhJPpijEOK+d6dNwN4uIhL
+YTnQYrxqEOAMmelnKajf7btb0+iMwGQxcIr0gNQNFbJZkvXQoQwOfjBLFF44Is3mjBXUDGkmyDV
eXY0f4JOYH08pZ5c/IidG7x9AkKr1ZgOAG96iM+NDzf6xR9jjcQrBXSvYBYn8uYY7OPFbW5+RaLT
HrLTFc6Oc0UFYNCyer5TCKIy7jaBDFXOh6rDGc41OPMehA+io4m+KyR2Hp/jfUo4kZbRx0EWR+OZ
Ie4koWIIqEH3ZIAY5/6qsqdEdLyjxQJddTPZA981HLENdIfa0q8wZbbAkZwRVfU1zUudQVwxNeft
iy5uX3SUwc2d3s+0G9T1wUw7e8W61+YtrAm81XHfbN5Rc7S2mnUVRbTZ0V+0C2N2FSXt7Ory5LI9
N2L1ot8HjPaKDOsMF64jcemyj0+WuBrzoQnaLu0nBCEKtTHDEVJptMjSLdpGPa2HdlA4Mc7nw1S0
mzmLDVCOkRvkyM0UDd0/vZX29gBXFlCB8ZkTosSjOLoqPoQzEL2oQA0NWWQiLogxGs3glLB6htm5
PZ7AwvAJoxVxGbY4UaGhiK+CogDTIHsI/cAjJVrx7Z+u3r4z85WALmkbH+mArSnMacqS0xwhFur3
9PdWzvx3VN6ryu7m6dH9/vTZm6t4O2G1Ybsr22cZocYhtFatzKPcE6vbeWCTkxTHLElW7UrPN34j
MFBsmSRhIxMq45RXj9i0/deFoqsb1x4ROhdcuKI7fZKgmx9fblqVSDpqytHGlUe8jTje82CG5nR8
hDa4UrRj8oZD6ef60+FN/GlZaxDsba1Ts7NhL3czkt7VnKbxmMvAo8dKwK1MbVMmeSvLKuxqkoGO
DxQhHJNQZw1t6GC8tbYHJ2zeBMA/6Wa09megAx2kJMO0IwugTSCKg8HOJDp6TVEr7BJnD/v8f7p9
K4SGecYDbejMVcPH0IQr9SH2wzHLSrUOKV9Dl0w0n+U3l6qahumWfqACJfPvdC9goY4WS+cSBgxe
zxvT5MFuDt3s2H5TIRm1xwgIUv+DI1gzTKgfWq9elrk9dIwtUBTPo2fv8VI0QKk+2Mbhpq9bxobu
ZTg3HTxh5ElsGlmBZnVppiOWrNGvgthrA02/iogCKx9oQSRm0/QttCRt5AdBQG4+gNeuIQbiHM8P
fSI6Xgh9f410CDDzBYVVhtJJKgejpwYE2LNHV1w4xDVuHjFvZcktV1ncNfm35rK1aDsXyl/z5N/R
HlIHmBezD1m4vb3XAQwutAwvVk8yHbYfqHG7ZRp5HLhFUiu3PLaa4oqe+9Cjkg0BBlrfSNU39xmu
hvenDws/zRHR5sjNIGF8ZsZO6osnJpIdjW1Fj7fHms9jXhkq69FGH+fJ1XfEA30l/nGNSjW8mN6i
8rf4m4nuaLxHRe68q7HTBwZFxE26hvNAftHIzIvRnFihX8mltthfzT9Q51numySgU/rw7m59q6kb
PAGOhA7EL0Uzh3lTZeCQD6Jr2lXVUHP34FpxFNwq1dg3tK+NFTUdkfHb3v0f7roqw2c/Z6GB9vZU
lkR6Nja6/kAVWeL338NpbZ1ZmFOEyFCDXDu0oWUK/ougAgn6HUSf57UVTmkFn8Mr/zLVe0Ko5WNJ
eeFF//9rvZtGELJqmqibsADwd8SfJei315qSvWiZuTKtJr2fK9ityrgpSdQiVB4CMBEBQrQ4kjaB
uDHFKmO50HUNoA1WFJbZeQDlfnE82hTTm2R7QbsD8Otk8fUDJJ6VP/ry5GTFjfEiYSDD2OILtd4F
1pfc69qnU3OD2tGty4RZLSPkdAvH/kCmrxrXHKWEmUumfZ8NvjWT861iSjqMLWM9ilTNmp69y/xc
drhokzymlI3iLigKUr+53BIRlYUV6yiXO0nUhCzPQMZHUcG5fNwrGYzmR/3T6UlgOUQFClrwuUvl
svyMQy+zlErb34DTPeT7fzI/c4gKALqfn2LEzr6CxsgAU2DKCCz2wXqMxbo1UgmjCIx8DxKDnfhL
T2X0phhJbYwziXoUGQrkLxYmPSTKgShln4dQfa4qR66u1XnqFXfmpZoDq9muwC2FQr+sAXmf/3gY
qE4SO3JrPevW/gFhZ2eBuJViLRuQswwcILPN/TSSItlGlPDsIgvTeMHGmEc0c68MSauN7sW70U5f
d5IUnbXma1m7mkXSqw5MwZ9C7yDYcEQwawUplsTMVUTGHfu+CT3Y2KOM5EYq5cOaWapW9MnfGQ31
Lx5OHv3L95FAPmc+88bN9LvllYt4vO0MFfq/Z1vHCjPKBPB8MS56Kna4CF7A0wGYfG2igFp/km2U
DTd4t+JIvPQ0GncFVpM7N830pinN0vWlOuxsUIctOM6J6YhwBQnL6SSozEJOqoDIE5BN7Pd9WxYU
ldGq3qID8xPjvrElA/gMe5oWgmTychNryamcRnxhKR3SsJcQKMEnSfoTdzzqF19d5/kSfKWx7Wl4
IBnIjqEy+DDnw97Ni/TJlnDGCXmOx5e39cpq1/DdStgH2d/rpHWIhrjSFeQuCCqag5wwUJp6ekwX
ICGm2NMKfIfR4R2OtoPZX/9jU1AdSy5gpqIBoZo2RvOlwZA/wzT6z/M455bFJJYHRjJn+lzKKd1V
CMUYNOhnH7YH/JV/H9aIfoG1BKRjm84lW+opgK2CzgpW1qWY+3weVJSQygURKbZtbbQIA1PRbFsz
fu2kjOsEe1P+moo+8Uxb2Eo30FkX2Am1ztuYlo31/pSXDOA5rNlUCi8EKf/H8epuW6IcZp2U51iB
Qfy1eDgwwZsoNFXJ293yRUQEvzg9Pj2o5jv6ZfuLL2YJ2XrEEvfogxADHeeHEVoIww0Q2MtL+4TQ
kMhs4hWOwWXywjpryqpU4yhz44FNTkVfwOaTTW5QquNiVuGsrxxKdqipkMfG8W5MZwDdmeG///li
dvZLdEja3jfRl1/FYab8oinP9/Q7/sFs0nUPMZfWLFruO5xP7pILNDvAd42UGt1uA/a4zqM4JIdv
8Qbwj+jOAJxneUaEOh94BPMiSVU5pdTdjoGLBssrayUWEhc8G+D9Hsu6eXt/o7KMd5L1TT2Riodj
4r8sRxg10+LopNpuO05bXUUuGnHClryLPJCYT+J9zK8paiKSX8Bm6Lxgf+QIxoo8pez0lNdbGc9O
9Xp0TPsAkGs1ObuvmhTmYsj2FqtoGhK4UYsqI5nnIhf92xK47nMfx/kYQOkXXWmVHJO+acNTw29U
ATlv78abLjVftciw6NBSXC/OSWFwwAtxBQPg1ApNYvq4bi1sUi17wp+LRnEqNKQsdJUrZJluowbE
7SziFF/O++LXi7mHvItnj8XG/FIeXmNTrC+sM4PiBiwY7MxW/Lcdp0sDHCuKmNah0HSTFWrcRZSx
I6zvxIwnSgkwL/CA/69r2TPSpbwx/nBJXfaBGAbK1PWU+tVqdv8Z0gGK1vSqGIQ+HQDSrtXUkkL3
yRwQ/OpcDuVzB1aBWYMkvd8lxyIlgbhnrr6Tuj22obicTXCzSyfOhI4tm+r8i5L/i7Qwa3aOn2U2
wfsawY67l8GYXQwuO8g91FAoeasT0XnrO0NjTXJcn+EiVctTOq0yfkOv0BwJypyNCjNqNFDx4M6L
pQr6aImVZK3zqdYxq61UkllPxgtkiWyWGQ7qXjLjxx6RZPYmtUBspDMDYw/mgnlgOfPKx5zWa+As
lcIR6l+nL+1zV5/TFPSJOpQr4dTG2UgS90tx8MaMDgncAOUGmW2tRVDl6xGkJCy1uQgRgGFP1vlf
EWSXrzpOp5lVZnqqXgywR1Et1sRzTjgNqUeKhtm3VQ/nUxwr7lTB4d6OXpAO8YK/slElOhHD1sjd
LyOxy8OooP0C8BKG/dLWPBjr3Igqi58Xm8YVmZrD7lm2G80AX/MWkpXTylOLv6gbJl/WjrHnx6r2
HgKNW+jo4JCLjbext8/ohnmpgx5ZfGBrwTrH3tCTY5LeMd02K7jJRWR7IpKiRddbLm0HwTdCzZMX
9/U/PyuKxs2DFBPvtV7xKRkmraBPQlmpUmVdkr4ifo/7jR+KgY0S9dH9o6EHLzdwi2zQDeSKQuxk
RCpsIpu3RScpDsbGplNHm9BBCRvfgx3idJ9nukyZzdEl24+Q+KYKIqYmFchV2S60vTw+49w7gaeY
lNQ6sBGJz0AQiCz0FXyZgEbPCtFDwhdKK2/f4u01MUJP7A3XFHdeXW8vLowdoeHfqxN1XO7y1UDL
Tsm8GWwfDh+eDgY1rO/0utoBrJGiA4kY7G13/4J2ypnwjG+oSpL+9I20tVWw+HAB8ftLO3hgNzwO
PUhQ+H78Yv18dPUiTkXutySCTgMkzlPdz0f++FuFi0um6+vzyjjF5LE3FEscMPrU63XyYqBi8TaY
DBH0vLaXJKW9dIeSjIvQowaqKvYCutZOmMTJNEU9g/4eI4kxjat5LR3zcDoM+2MpiXUxS7MxXARp
89lMHfaAgymrMl8dFHXrZeHHqdnUQA7zvRc5Qol7MglOPyUILTw5M3l/amvkiSURDmPMC3/FcxbC
4pCCJNBaTEfBBqlVwKOL1A32n3wiMFrINCzt01hcbHda1wj2/EUdDAJOtOl/m+uQSpPEu4ZTdnhZ
JwhsYyYCmCcPfGdBuVZkxOi7ufF7Y58wLaQhnuBK2wtEDt4+Exb45iTR+vq5m+w/x6lAIxV+rTxf
fohSRJAKvyL3PsV9ZrpDoY7zpDEir9+TCxLrcFZ4OPoYacd+zzcLX2vaGyIRisfkw/dik4rNlcFH
oWKuFNbYgRd/oYBZKSuK
`protect end_protected
