-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
isLk9brM0eEjxEkjFK2hpVnzvaPuH/ncHa+rFDRtIUoCgFAIdkeKzEGWb7hWhZkm
6r0Ey6vaUpwbjoFBAwJxci8j9SF/RJUcTY5YwgM7uG8JkoOnE1gzy0dRPZuZoVvh
mDPMaQK2/NDqm4nF7Bf17Law3x1Ax/JI1n6DdupEpge7XilMjc2M4w==
--pragma protect end_key_block
--pragma protect digest_block
7/0mUf4c8qiXEPnFMVNeFR8NBxM=
--pragma protect end_digest_block
--pragma protect data_block
BqqZfgKxvwjgYipARPYtumo8Drt2WpiR8qxUMwITWFXYB5ykQYXv5cYdx4AH8hzl
sGdTHKccKkC97Ek8PyRwI4yX168HzsC0Y5/69PUn68wubT7o8tS2e2UEUOj4oYY0
dp13k6IT2GbYe0b9gLo+NKTYtuBz0X80M057eo1iRum4sGTu4O/T5fId1QS7dEvo
U8n4RV7cMa1rblXj0NZFP10UTGioFULSObZLp9uuNEQU0BhLDBzFgTLnCfHFuvBt
uM/i9+CJvfXL9fSil9pr95olByHMCdGoGmT6tTMahFbatN4lnUFXdSLUpXqy2UBe
oYjmZyA0B95UhY5hTu7Fo7hNpuau45AsEgaf3JGl790CWWttH9EIJ2r25u5nINoI
9IKJOmPWVII6xZ0XJnErHEhbUnYa5MHtzWvNf0Y/Q3XOkGTdyrs5OK+ELIMxaj5h
WowBBJn3FZJheqZew17QIj2qL7nuoEKvarEjxZdHSLXoN6cdKgfJc+b/1cv+Ivrr
x0y6JaOR+eGyC/MRvYyyvXYIsSImVREBBW2MpTcjAsKMu63LWTwyfbVHvSOZXwGP
7LqvnhMljuuusipM/LzNlm+7qSrRcVcJ+NHuVJe7XlJ0guCsWL1dDyFMJsVYk/2A
RA/zVfsqL6a3PhDblEmli2a2i7nHT3DxWUaBrHONnUdKgLat5gBsuadOzrakklHy
KQ9XAP/AZ5ZsuLlbd4tg/yTCCZzihrn0SgUygWAfxZ5qcmAk5cglr6ubjrCLZm3W
5GZFrnrqmyDI7Ja4wxDxy5wx+hi0vLw+QES4+9OW/o9T76XTbsnstNGiNHQYGwIe
2IDB5AgmvG7UBm89wZLxqOVC0JUTyq3FPz7tSflQY8OQRCrT7ksHifSchv58OBqO
RFkzObHCtI8M0b9OyKjXpOHfQKhQQRESXtNmPNGdh/WQl21SCN6WKYi3AtkMOqrp
JEMTQAhbkR/rzD3GIyjtgYHtIDUBfzQ4n6p64Z3lpq9KLwkptAzhxxc/zAz8BV7J
U4212FlNjuTBMlx11QZYH6YKozwbbmnx7PGICz54dy35f5ptf2Bx6IgWBycQOv/t
2cOfrZUmCBLEz+d2a7sxIa7GU7QdSzgbxXaUVc51efB/4Y1DXcnkhJx1pASa8u5R
HgEzDIa7tsQDd2F7RdFMnkFWg/jIV/vENbM6/3oglBL1Z+keaGoh44iYdYVMkpo2
OzXMVaxhFLQ93mwHlfz8Rqc0sCN4AUzCS5V0LhK4N/0i6wUQZTy/mpaJSM7uDuPO
Y7wmBlctdUAgUBDr2wZbFbD4IpBCRelghFxtUo+fOFQDa0hKO9ujQWuJlChubLXs
y8tFebH4G1Uo54WWQw1UJSiamDjF0BOaCD9GoR9QDw9CJI1PYkM7paG9tdN3tf/W
KteKLQmfDniz4QO6hU3WDAUSGSYjoCE4ldTwCFHoPXFt+/1IL0XjULtY4WldD1Mt
hfrEDhpJQWLYHxjFmuVb6suQhQ0ptMuBzmGMmMkwEO1hPO2pu7y2k8Zan4T1zoNm
/o6j+GTBKfczQmUmMKoolsF3Jpje/7f5j2chipq/sB4ufqwkxM7OhN80Gc9d4DKF
mw+HNgCsJhaelSCEDWB3rl/eCXscYlr+MjG9R1+9aPSRJpdWBn/sjpkt/ndyVUsr
orIWoiQE+mqHF4C2HLPHRhQsHUHuAXGOJeE2ss57HCrC9saOkuBuwx5yLtcdO/tx
FJMWsoPXiXnv1Iog77BJe4j6Q7xHBblrPSaJdOgkTob8RF2BQlvfsffIHfgdBDPe
hbbvY/KuSa5lYl82qI3n/dpeNRXQTLF9yfyuwMYssa/Lm2iCO0BXm92WpZZdJjrB
Ik3kZX464K2P6dERiONZ7npM7JUTnG1HXC6H5HgmNl8ZQca/G12DY5+3Gtru/nlG
6NdBRJW+gCGdCnZ2sfThZ/3nkXt9WogNCei12NOJaM94CF3B4z6MKPSpwaLeen1i
kV8wmTDcxq0kQdh4dNq1mxsP18HUSqb5TsanasVr6avIlAh5mPA08D00p8tC+/Sc
O/b2vTOziQ/QGbnsff5UvDzakQ2KMCWCNOo4bLJTrZ9BBwJmFBnHlQuQnmO5UhXG
dDXPtmaFdWOa8XmBtJgwIWYiXp+YAGU//etLIMpQ5G87Ra2QaZnOPPhDrfmN7CXr
hEAaMHqRiYs242YrugAVG0++dqvvb8qHcz3dQaLgCxKRbHG6UqW0YY03j5eZ8clj
L0c9ew1Z4k4YeLvlAewWtchkz33LjTQvC9hnmBQiZz4Gm3GdNADFsUy1BRUzzETv
d1ZsxtxTVf4i5ObMQNF5i0q+iICotEVQ4yzOJ050zflx/MPkSmaj2OtAuJ9YbR2i
56dDqZmP4VnlRGqG9sWEQmtuLKMZOTYm77x0Sy9WH6jTC9HqVsH/iER36CUB1kw/
MHTz/bQ3gKDwu4Mkvl+Pnk77d1ble6iqJHrC9uufdvnF0rUjIm9R6ittuz9V0r4z
h+qcIJr/hh2rAtM+yERFGyXZuhB5rqe3Jo+GljuF6A65IhZOq4kJmIVQHTTGmBzQ
JbbqcNNpJx7WC4AEgLdadZR3FRCK8QkalN3K7AP3Odu68BkpXHbnt6hP3UB62lIe
GtT8bwDLdyduDA/bE3zUzMWyp0g3OZ+r0DvWNWp/RbRQsdM8vuS97CKeQwSPSaaw
HrmR6+KaOHvr2WM72l9NUKgcyCKk293sdGQcJFPxP1pM4UYEd8qcOQhO63yT/4jL
x3GaxRzvdjQ+RA7YJZyloJ5ubKW20wE3Q11nW0kY9e3ug0lyWprZ7vD47VsrRb2A
mAGncYXxfSna0ZAqCul2ifF74QNZQ8aWC/x6+1ioKvd3NXRMKGc42S0bvDx5O/nD
TElcwI9Kj3vWXsw9xBX03FXPjSJ1MuPq1MrttSVZkPuxIa9O3bTKnMDdAUpVy4o/
tz4FpVcazQayM3hVltPI+SuF1W3lriiOMGKbw8m2Nc7Is3usgp13y83Aa5FhftNu
gzrDqCcA6DdgAttREQhFlKFJqEppwuzsaDq4fYiUdjgslhK5aSfXzCB9BYJttWrR
ZAAdsC9BqpH+tCKcqU9hCzMGY2AsnXLm2iPdNPwL1dGwkTKsMkztmrJCO+Dw1NXj
L0T7zisvIUyFcHjWZQdk8CHW1W1m2Q3oC8NDB1PGjJNrXJlVYaP0upgI2tevAs0D
zioDeyoB2OdixhcZbfg8rRWBVreMkZt+gK6LM3dEx4zafjz57QMoXiY7lcwwhxhg
GnIpJ28Nhf+05knc0IZD4Z5ErK+WAq1v+H/e47Oz32AnvHVj/9bAW5ESlZr5P/rU
A02KGEmd23FAT5soTyOLH1U4e7agZ+Aa7o86qvb1DGsWc/9SuWDn1MXI8H/t8y4U
kI4iOtnKSRRX7YC5HeUQZkRkiUvYdpfehEs2argUMDsPeFErR/F0VoTuVVy9BKZz
4AiU7DarGyZYOq4PsKyg5zXXZh+uvnLH7Jjb8x+SjoQMIemgaEW7TG1OmZ4x/HPE
MFdJ71Xxdxqd6LGgaliTr++rs4g26jevjVyi2e41jQ6HUVrxDtfBl9qHmegKRBdU
v4Q7WXOprgPoX3CRkk0mgdVd9NJcSoLUt2k1+9+9salXxjVaDsug6aycx2r0erZh
vn3yo2lBTl3VU6FMXrmWTLywznrGfFR1wzsTqCIKCFvf/czmUTNQvRioybVkAkpN
gSjQngWAKUHZNulkEmu1Jn+vXd2Rzk4l9hpG2DxI44KGlEgsilPxPdAWUS6IhLGu
h7HvXMVWhEX2vFy7efl8Rzozdq/gumnXtcE1k6r12eZlqO0BNbTxxOtAnkqxPslE
iN3IDKSxjgPLjBs9Sy4fbBM8P6ckkcKprFXWW3uxSy+o/h+lzljnhw+yedv65YeF
RkhaLiIljcUvUkpFpokxRGJ6gHIG48J+Lr+G3N3swAHF114O4feVsh06eK1xVoft
cIN+RoHB7NBFUaDNEArsht5WGYxvipI/0FXHA7ypq6ZvAExpRlg8aOMf+cWNqsjQ
6ezi0Tl3qxG9Y4Ap8Zp5KnzqLfB6d1zY54d0PUWof9R/Ck6oZzXe7zyzjbl4Xx6Q
L2+Boiynqg9NaHM7JvTYiaZK4gFtdfzUP2SRAckj5IhWeI3weEBqk3fD7ApqVjpb
upz2IiaV5/gr9NqDvlAkNmpr5TVPFtlc5TF8t+1v36rSMfioDDg5pX9S1hHBKwGJ
uaRxBXpkQWbogZCyIvekf8oby0hDoS91aZLInnaBH4UYpZP49nWc8SlOO7p8Kynz
JMQyHzczOY7ZnWdoG6mMYvUIe7n/q585F0ClIlVJNEgeYbcOzrLzfqeomEOcvB0S
gbTkKIdjUKYnD3XEhkh3M0q70MeGsXgBnFe+1U4n/zr8bbPKtadnp+0wzGQjg0eO
bFiu+htSMhH20lM7wn6cF8sEW5895Pqyi0ncRSUt0ypXP9r5YSP0gi/1R1WtVzbx
ddlDrtd6tLGxMN/vT0U+PqUexSboPfhBgce7l4l60PO2larcT0IQWe0Rr4iXeQaW
U36KcpShCHb7eRD69Yh3FV1ZKDw6hxMSA9C+VZ0pYoz2RVfU7hAvbTNGGRI/rQ2H
WcThQ+ob1FKqSVW6NJb0EzFdPsqf36uHjlUDQ5XnmdHyJMJ3uSW34teykW7BU6RY
K4s56kZyJ11KsWdNVkTubZ0hIoHlJfO0edw6d/EvEvf01T6m+8OnMTrmzqIplGrh
Y3tGh401ifG4p+1kidxKNeUFweg7GbuM9Fcw4DfZXYCNEm0t0Aq6rIkppY6rS1Bw
RUK5cDqTnHW/QElLHSjv5kvd6kA13SGeurMdctqkkgRf+EFvspVM7jBfyiZ0Tvt4
Mf1xG6J2u5QQAxe+5eOANFDeGAqpcBliflEWE7sS/fzf5vOgjqdDlAOIojaQlgpd
fHiUULPWCm5+FOSRfhLwkbCxPwj41v3jwFi4gpC2FOi3O/bX6yjvpV3u5w9+0ZYo
osM7nxSD1AqI5rSFpGyRV3YY/ZPkvswRjiwEcdGlcIMmrWpaccdHK0nE5w6W9BYr
gUTl9gJVYWMzc1qJ5EuxSeL4w5W2oN+mWTf05jeswGwRRCwzG/wVT2/yoSJtKmg7
mXiSP3MZEDgQVkNMgZlfxA5b5V1mvaz5I0u0kkzRLr+Ssg9o4UcxIu91qKdaL5lt
p4rERhgBCd9zq32zG0Uj2SWs2nsJXbJhB5QYsNKosS/DQ4qjzVNFr47mo+SVOfQk
vF/Xj9qImtj8wd/XGE3Xm1Bnm3fYsgawFjnocWYGHUUK41SqxcY/GBqJ9kL3Tegw
LcxwhL0+IE3sDRwKg1N3uSCUyPnzEzHzrICMyq040o/cVWF13sI4GxKblOzWcBwr
eEQP3aNhoGrk047OU/+LkFD33kJIsXeCRyACYAf2NqrdgxgEt5+vqBmdLO038VLY
eePkMSaTqHuRzVN+r3xzisamfgOmj8pdccDq1kwBG639g/EwlpLVhTl9Xa9vmONI
RY0A6Dwamsbl5j5n8p5/3EmqTGbCbe3AYNleB2shRPUIMB+C4fLPlpMkKl6D9QQh
WHWl7138wSlHJfO4C9SpprQNALqlQgsADQODk6ZLBW1KwrJ/MHKWcmq4PdN+AQ+F
fUwFtZnVB8L2WKWXHMwetINjTUZlk30OkGimqmsBBbvtM87pStqSmoYUdUfEFe13
tracxk1rqwMjmyItfnmPN3Ow2OfEBrivGPHdA0B0II6yp3WS9N7YpeQ61Yzrde5O
F2o0mY28CR/Q4IKxrTBxoRQuSJEMbMjlzLW7xHbw7omunyQ4eENpuMTNanbCbdAt
jicDwkkrCEjovRGkGEZgGQY54OgiSGEnDjp8vAZqlfq9qjWU7b0lD9/DG7LAM7QN
p+0Ym1l/w0tKIa6kjiY1m1R+tCMYalPH9xQ9kGEwXiKGtjyRIAhNJ5XDVaUMgX0c
0cP8vTrCiwrOxSjo3Ci0g4DxtHkH2FiY/1PyEbJXnY7sWzVzDQQlJRf8TG7UTDIz
Ks/fQ3RNYYMAnW59gP/gudBfITupLzk25ZKp1dyX75dyJJIpd3ZYjnZ4dzAAgjVx
2Omig8XVxXx0NInqixzde0b0lBxnvTzb4iYgIpI41Zx8uB7INrj5z1Tyk4Zz08fA
D0vB4U5lxR1+FgfjxnLhlo77RcCu41SLX9ES32MAgex7cvZYoVz2C7iNEBJUr1mo
WKhv0iLJUcxo1w2tVN7ZaUgkOFgbf+wZRGZeUFPYiT3OJYmresAIBtPbCI/UBCbM
noazpCwqGU2MMx1hkglbWP0SZc3hm5PZbdw7pkwkQLsO22tw8b6YnMVGpYla3jwY
2hcqxBWYu3AZ7EIRPgVAzXyGq+jWSpG8U3RdmxnxDhqCLOfH+MgMCKU+8PCLILlZ
gx0vaWuKujSREjganu22hBgrfMyPTvp77oGDdOv4pSc1lWayJ9As3RYRNMgSH/K7
lKMGbeXIeXs7BXoKuatOUwxPeXPIjV13PM/Hqbn4FLAnbWT1OThNEH+SrkQO8vcJ
K4eDnaakJWkRKCgBtOgefmeAMM9eBT7YDrPKGe6xBMWYQbO1/cOnlH04KH53oeH0
SPEMxsLMwnjtARLyY08LGgz8hM4RK5NKu/UBw9b8JTlY8+3GCVEfGOfbNSR4bBzu
gPi3Z7GVgnx25uKE9Mbtv95rpK5HOWMUywXxSxZxV1bTegwAluzZXMRDHDfvzLRz
NE5ExBjz/piR6GtDN7Y/AL2fgth/Sv45Ph0kmwclcxXPkJK4wUh2asVMqahmTb9R
msdoktybvPmYkkn8bGQBFXmmkKiW/Cc/sOVKC+D8zstTOtoGtZNZ20QXQ+3vk56S
PNw3dtPUjp8j9Ug2Es6iewVwpMiGRottrFxCx9cFdnvaGco1/78zl8vNk4ANche6
h7TDi0JKzOdX+JJipnNteTQUnIjGpu+nJvmvlgFPH3yNujzsmzT9hlL/sZm0LJQ0
nMBfL9EybzCtJBbGCfGA4Ca3/8mstY35RrVfKokKhKao19tzW7xjBJgIoUXSiYWN
eNIy1X5C+5dYPUTj4ocwrRturkZ8CVWsTyHt5sF1ZpEfjKopQXwa6ydvuAoKGwsz
gbHeWLhpcuSswp0/cb8m87gtDyKtzLyIqs+jLOWKPrcinYWJirZZkzszb50RwIUo
cNTpAQbsNO1v6Ksg0z0B4EwmTdMHqeiz5n+WuxeW7iZcXp23k5FlBZ351HuOJbG2
/IeKM+kTUdUMn5kmhvuSiKxxZkOzf/CG4TRKXyGOO2fV/vsnTzOuqxgiWCvXzJFu
BzBSCbX5/47tmOxzWWQKBnTk8JPRy5F5tNoDbl58JxfDgGjF0nDJrBaRkk0vi0iz
BwFo44M4Q1OfRlNZ7e0Hz7Z/g7SDsxajJMAapw+cMZSd01x9yA0YgkptEN0F/qQL
5R+DwZrgk6nGLqEcooxQhAVMzZo0XGsLaZSrPyldaB+lO9/qXwSoZJEZF7bdn1ew
YApa5rzQ6tXEbT9XSobJOxPV5bjtYI8TCS/VbBuj0uTyrmDOiZdh6mFFRZZu9lRs
ktlXkv9obHXgFwRLcR4sJrs74TOEVUPN67a67ByQP4McA+weRurDF1K62lse0MTm
Y3z11hswrGEVYJlvEahO3dOBZcfsY7OQeLz9hRCvis1Jz9EhAXqQMiKlAGP/iABC
8GQs6LebSESGvLXW6PFj8RI8/bRiZ3QyocIXuvOMI1YGJa0gNkQOLBglFPf8+LaT
rqLh5iQ7X/HB0MLz0B0gt6/dzV2pHvdTAJ2WIS2+4Ro++25qkuiNTpCdE+P5TLDY
5hnTANjP+8zOycKfStkRyOnuT/drp9Rx4N5gpepZ7H3LV/7kT1koJMXXTZD/AWM4
kQTY2+HDJc8or/AVq3fZQ9louHn0KhxxbOZ02F0sdF/lWjJjpWN7FJnOYv0xvJb/
wJUQSvOdlVZme41QJpHyG0LSrqy4w+OC3SWpIbxnwU7/CCJpN7APATCZwOofEO1i
V+BgHJThqsC4byGwV880V6Ux3BOZXbXCkxW553v60N6DxtH7FTFUtuuJhSnal9Vd
RBSP7+Cy6lJJkWPAJn3wb4VwhzBb8f2VYzFWW6eKA/YTVFhpoB0Xi23Sg+KUo/0Z
xWw3Xatv6VQYKwbPL7Xrp3mAh3YXU0z3064x1fz7ZutJ5n/kdH0oKUjNXG6GlzJI
eMItMLRfpIAu5rT0i/oc25NGmHqtp2yf6J1xNcrto924ibbbi+LXZDDmKP37x0I2
DlGafRYrwYXbfQwdajE3PURIG5mLnMhBcdshTZsCet6epgCFsnM6YxRNOmUcQQrZ
rHcnTzQw8WIhChIYrbJ1tSkvxTnQ7foatX91+Dd4TK3ajoFHYqXxEEG1sZ/2xKmr
XjJ81e/xvlaV1xSGwr5LfaqwjWSXWU404T0o4pEQMAbpqHTy3t4F4em7ENcRktJw
K2rKPUzBecImuVBrVR6c8wO5Sv2lGIQ36bOElBKYqDqzrjz233SXvYQzea2+XAnA
wmrnEDlHGCMpeq2JOOGmBWNge5u66hfw6Ak3ckeMorDbat3l3jKLV3uEPVg+/0fy
kCgJn1CKTS7rZJSItHz389tsFgfz6Rb3KZ8nRXGNuzBrNpfFjnBjxsd4FXSG5u9J
KYSDIsIvh4c4SKWB/3UD1BvJAj6bvNMbufnbbKkBE7aan1V/v4RFZUaWlPQurRDw
WGPEXQqCfPYbYEkQveys3ByYcxc4lehAL2I8d5HEzGokz7808u/AZEd91e4uMnfw
UaIesjQrpLFdYMLfzRX2pGbxgyBj3oqPR/CkhXCq20p1TmtTYjVkmOXctwEpAtcZ
Eei/s2f9vb0FmDjCt0B6LTSVxMHVpGpNyDntAHNBsjHUJu/kRrs1DC/qoVD1LAqF
M++kLE6om8Msm6jXToKVLwiHJ+l9mK7lCXI/nloWZ47EHCG/bBM64QgF/m3p4Yum
QijXPAzkwYzsRbPZEg4MIvq+aftxcQX0uWynFPmIfDRbSYEAPbn5XutNKA9E3HpG
ohCcWGXfFB+2rEcKYwQ8Tt2gHqGeGwUfzZu7phkds1/Vg7CwuVU6JvXOg0KEeGSW
ayB32LpkXC1OAzNLYs2Lfh35ACkVsm5OZ2PnYAE0dOVNleKx55REjVqEONDuw9N2
Owra/X8hUGdxSUS/qk0tbVicxWVuXUecplKQtMH6smiXL0coO2d7jp2CucCaABZC
8aJji+OkGBsGPSttHSWvD7iOsUe/Mvl5hsbeXI7PEYvWw7WD/SaI6ow4ZS8dh0Ne
HtaKIyCKIng2bGYaq9M44Ym6j7XnV3ZtXLTHdlXLvX9zL/wvszB6GDmERsXnz+JH
yiHhgwYq+Pj557dGzTwGdOS0Q18h9lasKKEw3vBh/HmfzCRA9TmN8hExx+j/+60B
feZo/fpRhn9PJBmEQQ5SuvsJdgMTaTWcE1Th1lBjiWttiTXAfpmd0y3rCq3HB1Ph
QYycZOCk680ope8SMM9U50Gk0mcJHrDKlMrPprjfD/lMeBYcwl3FJqpUN6WVsKyD
ytOlfY95i3SANyQV8AmMk3rVnqINFpVW9PZwhdofVtb7QlXW1SJyPouFejxIFtxu
O4uXBb2/qAS7inDUoNUKeuHUJoqZ2qAQ77FG8bZZTkTIR+q+LFpHYO/mhwV8rnwD
7lHDIxuyhRTn4Fr6TPSjftM03hZ+MCVxeH1MJUzew+6Y5HRkrr/80OiDhJTK5M+y
Co216C8+VPlDhdhUfrwXRqu0bNXA3vRLzeF/FA4e9VH/j+oExO0Z9Ev6DTAtCuWG
uOymvMB6BVWePD8TCy0wZH2UIc3jwZUD/vDM0vN1WzsHppQQIzRQNg9OjiC0ztim
AEyJMbrJ9zRDWJSV7/EvJ4cSjlxxGkjMAe3azASPEDTi+n1iK7N5TpY8i3m5nUvy
4M0RjkiBLbQCht5p/rhYOvzjY7AMkXh2LJbirBwK+/J+zStvGmwhv6L8ccvkED7u
hyPoX14wQJ4evWy96tAHpc1S2/DGdEyP8gsyfItGqTAIedHnJvrDm8G7vlXJWck8
Hl9653hPFc2s8t4BvKo5FNIJwxDyf1hKFt4B6XnXzT/rvMBiASR5n1n2f+H2VBf+
5K23bfIf9eBn0antfUS0S3C3Zbkqx/t/MqPgKwDUAbg4MqKM/eIKQoVXCuQwOHfn
LQPu6fMFil59+95WNuf2kwu/fbUXL5lm5LJWarfwxpKanm/Qx8eElDt24hGNmnTf
lecUnnPtk2dQ0N2TasoqNoytyC82GhFKQ3Bqmp9aVitRgGJzivPJXNU+TY6EMY/N
KMR44FFIQRAB7BbnjSS0h7+PXQLHu15kDHRwyJCSWlXGTc3D6qlNPNsa36iNbV5A
6EgPwvfHut/nnIFmfiQJwo6iz5I1IyLZNx0uIWLrv0earvP4Mu1sI0GvJz2rrYGe
5YrQonU699pvf5fgKwnGJyN0z3Mf4eCwV66xX+IltyadA4mUbHaXe6SEvnrX8Hvk
197wRts5ndlcQY1obFpngZ5O1t8M2wGbKav5gtu4JOrOWOYhbWlQHEQbacg/w8NQ
sVKrnkfeC4Xfizc7RhvbTNRmF65QH68zPv7jo5jvfcTmmQ3Rwn1MakDDPnM9u7FH
3eC34aFaqpiRrOiJ7S5ULvf2QPxys8vt5haxyhPvhjl2KDLyiMJ6/VB8rMkkNWnd
0UYGVtQRUbe2p7vF4bFUHGh5KcIUJpKGzi4tMDm08IJN/PY/BiVaCRNUAojiYBgP
W5Qt1s99lXZxyTexjGFACTdtxx23S9mvlNi79ZsWL+j4KolU42hoBy7+pU29zNM0
sIj8OFplciui9XlzOfK0ubcyb92fO9HP2W0UmP3z2KElrOEBGTYMX7OHHoHf5FKZ
11RK6FnarJu4tYO02Y4Sjw8N+oDSgwz8R8C+/qz5x+84lYywEhAWHROxx96Yyiim
Gz8oB1LfIfKz7Cz+P5eYqpJs0dBYEcN5w2LEXgutdY+niwMBuoRTCb4eoRoL6Uj/
5t9zuXXMC4b3SiaJNpmce4iPffrx51lSsYLMMpBgK/ieERbCowf1V/4bA9cPvnXb
8mBT5BYY0776WwlRQuoi53uYiyc+hSj8ujvrojZNG2jXlb08Io69njw9B7yv6k0R
/zBM+/vX6YqTU7xtUiLI2s2FeQcMDYHsNw7ldi/F/nTPG25HcEZDKP75wOMkztVg
+oNNDbC/5M9pmHS971p5MA1pnWVezi7aeriRtxDknQgtgocTDGEK0/wO/dcriSDC
k8gCeulFRb9yuLDaKPEC7uvZu15pEH9SoLE5kiLKA2OWVGXMNPqfYN8MAvd1aZJ/
9LiYkbYV0CL7cEMmq+BYg2VRAKwK9b7cMbekVXz1mknVEesAoSlEEDUaVrWa3boG
qReOg/i4gB8We3rmnmca0XHETd9fYqWA8k1sa/CwqB3eTmUvd+PmkQ3fqsGTf/8N
YcF+AMyZGh7K9B/t5YBEbafcw796CXI+Zr7nh7SssCj3YOyWpVcVxReVX2Fbsq+m
UdH7flxInRKQe2A8V5kWv+NcO3ec8qSDxLUcblJOFR+9w4IfCD2hPJpOMTl6oGr6
kOWRkFe017YS5nuNx5WiRgKCSQu3ykHG6qDhS9AOKgkt1gK/DA4fCdW9wHYNt4mw
hn57rp0YCwICspR9BrfLjeQRh8hguNxenD9IVnF6cG3hHgN0UEVu8iiFkAhnMNia
VZLyxMWMUXiutzqJn3AfuZjPk1b90EvB8jZvvyFIgo9/20O1HR43ZLTFZQFFQhfT
ZcC2dAnjgXj5finVf3sTYgy0BAMepGGTnsiPDDZky1esI0eEkgaAXqLEuvGki3ih
9uTYBUM5i2pdBL8ilfiXXc8qg/8tI4NKKBBuA77UD5VvbFgagzXGyQTYO4oc9Ywe
gzZV3f0E1YihOO37vEuFILFGm6CaoS2a/ues8NJ0n9ld+gBU5hC26zAiKePdVtjo
MfqRh1wL0SxkykWoP+dNorne7cesNvN8qXUY9yRqs8KOAQPjDXzF5XAhBooXmqHF
xAOrIOde5UUqq39QGQ0tXDgb6iRMfkGlDXIVZngxsFfTj1SggcZlBDA7bULDgKnQ
LkEW/T2tKMvPFr6iGc8aFo4EsHw4H0fKGxoRnWtbzsk+f1VYld8pFSJQ8TC/n6aX
GPFJUMXyNnnSp2ATp3lu7/qY4oalUSl4ok2rPZz279R2Tetk+EYVd7SEm+z9IiHh
AUYA4TdBVBE71Og7xvwwAFspecqxipc6IbpCu8/QPxBfRnfN8BUL9SeX5jsh5du9
H9Z2BHWl5TYl5m1IxD8OR/OAXLmrcki6re1XUUy/UqEsRehOxJuntA+UUeiMvS7T
YLylw+j6DbwOw/wY51ugF0wJNDTDWejFqURGfTbpvvtxY8ZtvjXVrrgcUPsp3eDi
kH7PH6tqvvfJMMK5ZlTdHkD5E/KwG7r6335saugNP079axK21+7kn6HQjXCgxIuc
Mzidub48zLbtF1g6YUu1ZGF2EUgH6ndeFNgJBqr5Ve8zsD0eWVzDT++QGSafHNM6
InM/ercX4Y0lh2gzqq26tYNws/JCsPMozXMTZIiy8VNgjHQqtQxuIcipWkJNBa1G
iXjFI05nFSpyaTcLCidBbhl4s2dwwvewGLcC1NPyQUPTYeuf65ejJEsSOBjtifnl
FMsfFClsmZbJ+x+HTuRnU9Wf0o/ZWAATOVkc6Y9j3W9tDih9hWBX61n+LEPlcQ1M
dfHnwws8TlJSROwoLwxpYkFo3BbHgAslhemJ+G5pWI0sr0lkkL5P+ofk0GfihYj7
qoKhz/8phGI50RonExJ25jOTtlLfMGUa7rqvhhsIj1zRH4GqGJEKs7vD7D9nzE+4
RaGwXCE0lC7dHK4O3fTq8utKzxLd3DfczA09Rkt4ff6o4oaw29eR5phN+EDsEd7K
giUSY0e7a5zx1wJPC0aO0H0xrvrELT3q933n4QR6EpPZ9REtlZELyoNbgC0UNffr
u2D2B/Zq8agXojq7EQ0r9IamFRxuQcQf7QYEicNZOg8gYtQCtnAXD3Ms0A8Fdkum
hYp7zAePSwPTrK4PyVYYjlzjA7swwr8lcqJhhiITaBIKSexmeAYZ8myODstssELI
QpEWZLSi03f3UC+0VkNhNNbhj1CkXV0d2TThFH92Wfeq58tXINMNcUHWiHcLFsxp
TtT1kyPIbmEFVPj83X3Unn6OD8lMQYWBV0x+xDvRry7/jAOGlD3RJCJHcNpYybHE
G2ZQQkPILtOQmhD+tp645OtHOe/8qRaxdWd7CHTOLwREPTnOpe2W1pUVQfi6ilru
QzJu5BYPgT8FrugzpKQtXEU5GHaiOzoGRCnfcPhPwcsPiCw3ozIitRIOR2yS+C0u
HXZipqYRAxJUxwe7+PeOTg60TtTwfyORgLaYCKQ5J644CGumSpisBlAaqP3CVjTb
Dpzk1hQysw+LDHElHGgra7v/GfKQSJWkMXiWTGMmkPIpPOz0Hme2B7OYn+bdK2KB
shEoEiOgjsKxHVL1zp2DGM41IEpWNPd64ODhuYGstPfAFg3DRSWU58PfYr6Hc2az
TrJfjVRrc1JPpXOyVBfGjRjr4d9xoMeEuHTGwdFU9zG7fwsOpvyPEXou1ZTVo1Ty
YIPSjYN6Qd74PF6ewDGbVPqYgVKjhSH2WjfZdvqsAIC+SHPEeTuZRG1P76AIRjy7
cHHHuUAi2oBw23gDoerDQDnVF1P/5JJLZ2zgwPqmiK5lo+5M18esUuvJQVMrj2OQ
k7Hbh/WguNNz4s8FI09M9zd2EFH+HHwgx8EPgf+dJ2oODHp54YMlwiA3q8oNsaj7
usKd6Uss8QDge5/P72gAwMNs0d1DRASfk61dQbXDXgr3/l88/rODYH1UYnFy33Sm
1TjI4ju3DPBG0mO4B7qMGQYAI7ln+Jz7rvSBjIR2LVC8JPU1ZQk9qhqdq+GXaLRw
LPn1iVi4JO1z9V1v4t/da0pEYFA2+hkQTHl1OJ6uZ1Inndcjo6AYLVT7Y24Xl1Br
oHtYDoYdm9+nuoGpsmu4E6HNhWw+7q1bnjk18MjlvubGxNzWYXiJPxkLrBX2axYD
nZ7lPqbizoBU5l9vmUNveRm1MX4HCTHkxdtA5ObCBKHaTBLC58raK/pU43rmDPwh
icDi/a6F3eMEXXgM9096rgPW4TDQaOaxPN17R83AGBp0EUjngIb6o8glsOcvwk05
FtuQhlrXLr2VzF2AcJpmCgYS40hwbOPBIHtKrjwQbWe7MwiSP+pk816dRHgLGvLO
2rq3T0uc9Apnnt2KrLRhESSSDIn0f31k9RLvtC34sxCgZ2twD8FDCd2JBiz8chAR
Mm1/tbe1TnYGYJXaXxkoLNCldTMTQS0rXAbrGPaSxE+dp9OdsZNT5JhpdNX6vmxx
FKubWsS23LlzpJPFiYtSwBESD3+wq23vKp3d0Mj9LgORuKXYJfxJQk8NCUiIxV1m
lYwPLie/ecUwllaArxwYiwVSrzJUghRN8J/DaulsKZg5VBZ2hXdPfAlImEld6fDK
N+bQJmZSybWaRDAIIyDHLTo+60CpfIB0mVaQD9HghAWw3rxnmot1b6VAh6l9vAih
Dpft1mq5xTuagihw7FA3oIJ2M90I3mSMmOzk3azKGP405A3hIY+XUN0isel7Zd3b
KrdJk21UduZCggnbk6XVV0CmpVRmFlgxwhhNgXs5TaoGII5JYxAOahGPS6MURFSp
+OThDA2ax57tSNM2YE0G5K648I7HCbS5WKn0Lt/r7Uw3tEcsp2nYg/5TAlp6KwiZ
q0JuQXcjUOtsvgRbWbHSY8it+dmUotij897wLHXLDWXmZydJUpHRBzr4m8lAOldb
f88QoKYivNV0sWmUSHzvKuhEnt4iafmPa+Vr5N0XH+Y7hJFLianBtbHdMqRwKjxA
0pkHn90AfFH9SejlYtxlRWCuug/7kVsRzdynp8causBdv+9Od6g08F4Hmk3H3ccA
2cU47dZbmmuejNNnPPbNj0ASqma4m1iKwmhiyCcrbqdDh15PQnVtFAfggtvCMFAN
Ha9gZoC7//zcMI6F4zsyogTqaPyCPAk+gloyuxsjnZvAsvv5PZjgbXqpyPVDH+Sd
V+zMhTtSnlzmM6NBzp/c3fmdSdzkN1EtIF4UKStEzDroIX3CQZYtUVHEXjk5NZXx
PjCJ0VM4aDjDEYqN0vocW4ob4J8UR0XIt5/bVVxjgyssb76zJb1Y88gRJTCQWU47
ZSdHapohxkWAD71/Pcf4I2kSYfFGu0+O7X5l90t55z7GLH4z1adC9+LAtfqsMBaj
PGmiIxB5Xt+5bcCz9TXruNTgSwqVFqS2m7TtKZRuGmpTcsbJyP44DPaP6wBzV92r
ccvove3UThzjXxKrwmfU3Km/2kwSI6OzxplbL4yuL6cud7z/W+uKaLgr8yaoqdgw
juqC9F0uiPhP4PjzI4c9rudvKK8Yx5hdqcTaYbWMumbz8qk7wBzn79/AN0Prz09w
3CEwIZX/j7crR96vuBBa3rYYZKadmljBmd0l8rZPGHvI6CL5Dzr9tBaCCoFpFoiV
huAdrUOx/lLdDJrYbVdtro1SYoZ699LfsI3pfnhExkoQ5n2HAsfS2g8nXvur/BXq
92GQBYdlylZV2w3kYedJcva9EbWMOREg6DBi5NjNkAhXtzMBBwjBJ87a1WM7TYse
LMylhXxqbJh+C18asQWToaanay6ykfBIpu+HrxzNYLCIxx7N/rBwv5r/zrHFtLE3
KTo1zbVXIXT7XGIYa0c3wSSURKvJGX/ISIJYk3TvLsG8oaizVvutCxCjgV4VVY9h
adioWc2Ob1KRT+FsBpzEzBpDuhHSK37Pr83oVNanigTV/Fv4indhlc5zW2zA8GzD
rY5f7fL/xe+vNWDgfv/g3aIRdI5mRrvZszWzqervBH0dbeTnJjdP1BjgEqUxNgWM
se3jehb2TFASFeIqADL7YE9QED0FPOfrFPUcl7zMaxaqaaybqtqWm9GjkMvFcmT1
MyjoGSeq98q0haBtxwFLU8Z0EZBY2tEZXTlofWpkMFq3yeXhYNiMhYogqwdFwicD
Lhasln9YS0p2GdFHIf06iJQkV2vt8x+xlfOOOjSz4M1r6faW+JKmuViIrktdDrLU
z0CnOEqtF6hCKGmpTdTEBCiYKWbrN+ObpaykHDVwByQqV/hKa9gsJ/7FyxfCRRGK
ELtKKWvf51blNDE7+3k9Dnr8oCZ2bbnQptOqfmiExi7Bn80Uki6Q/sCV2M6ywO5o
fLPvSBvo0myuKNdbrWu06ZhSFPoivJTQTIOs+n6YWNyK0wd7x6Qt+7Y8D3oH12dm
v0ujl4rSud61NjiwOz8SZHcRenkc64nQA2zfbKeN5dH79F2wppaxnYFhJc3lY1Ei
0oFyEf7d08qPQU30XuFTM1limh8ogR192wyh9M/oC3Ef+ma7hcsc1Q6/Ubtq41iA
+x2NmhmOp8Xe7QSZZRO8DtaSnwVwvA5xS1wguD0JyvsW8tfo7MX5j7CmJ4opryoY
0YfNU/ruFwybDKTVoLkI512idgqnbsR4ie9zyJ6IK5J4NwCnpq2+qyp+qdIx4aEh
opTtdDN/5IMboP1OdO6Xb/G1sVNeBoxrM09GZApwolVid4MiE1JZuYiYfBTQCa+l
JchYV/r4ixZNNosY6ayyN+2Yv553YkSIrkCXN1zVZQ8NbMDSAfmtaaUEkuzOyG+e
Dz7Q6wKjt09tK3uFFA5jjwldKznCTAH82B21n6IiAEQ21lrK4Uk0htKRLk0pAHFM
eXVTom1yEu/9IaXMPiwdfDhm5iwStvyDvDa5cQ8A6nHl1bxpSHEDuqiSb54PDruo
11vzEARNFSTCDjjBxTPvo82ZN8o4wAdIAkeDJF/4YlF7L7Z/UeAV2r3KtBWi+ZXF
7JprmRbpL48RjeBbpM4BM6BN04ZUy5o7iobgmKeorF8XTQ6SuluBek3kpflreGJD
7YoRwahxHW5sn5ltf1lE0nudWFnBHt/IOk6p9/C6DvajjjRU4kZvyT67YFhSKKzx
t3oZ4RQa/GzNWSovrtCuERLho2NqBqaVtg4FRQG9HdHmS4saC1maPvZ6r8G0Mk4T
6HwccIUN+7nSoeAVZiK5ztwsg+R4rIU6bO9lA5yloLr+DpRX3IAurme4s6+kd6FT
VU1m/4JgDTPNOSMesTFaCrSJxxsJQYx4ORLbRK54uYvqtrA23JqCix4TjilqWzb7
0kwjvQVJcx+MFKk9Xvvc0XZgSrH7/SdNNmO+n19wUjpVWylxxILv1Lyne2mGX1Jo
u/vUQju2mgrBdLhp+6rDK3wWIurIZpEaWriisYUjK7avOH2GQ34FBfGxM2Oujynh
DL+aBLWooyJZdBlnF4B14yDoLNNfNSqDtTSTqqZYnc9ZgbRAcnhhy+K/OGhhYnQa
WXABrEy0GO295PgnHgj8GzSmeGp/LjX4An8cTfWpEUQsyU8cL808FZ6qdjIJaSwT
BW0y43j2m3ANQdJ8FyK79zR6xyLy9xGrhigO1Uzumupk5R3o8yLy5GASjpNjujOT
NTk004AW4g+hbt+uBAjveF3mZn+0v6Yz/Xs+zA6qPzqo/YXoYkMB9PgI35QzsuDl
c3YKEqDeKWDsgGi1/EHqJeaBoNDR0hoJeHJ1X3RB4lHUAIvJyr7xl/8f4h+jN5t8
UAhMC7WBdKbit0U/DSgoY9zjVq1VwgGDHF53VqOhZWeMXAFPz4GKA8J7Z4Te0aft
7tjnOjK0AAqfNt5XKbJnhzv8GMICwj8GFt1O32iVO/tsVx4D4t2r9M0LMI+NOHXy
OZgB48lK9hbtzrJBMjxN/o+Z9UpHAMVSKse9AopFDaGmHMb5+B28/Vldp3A0C78I
S1fmF2MCZk/8icjeeUoGQ186VMTqUN8BmfVUhu0gBDzM4rJ2dAxEqsAeNWQBBakP
9wZKBiWHiV5TxXomKL8ZX59/nlPSQl9ymwhtY08fQtEdZ5p1PZrGuqn3n/ZZxUsB
Q0dlV676FbnBqPRRymFt3ghz1mHfq3om6sgN9pvjTLBGYi3t6Whvjj+kCRWdyaD+
yaXYLjdt4e9fnMmdIVFO7EVayHVsi+05GWyNK1vNU0ecP/xSkJyhUy/L8VXJB12B
mR8G9b5xp51gBBpMJj50yz2dDgSGwjDON6Ql1E76WsITosiwXrB6U8rQqXQakNjq
ODAP3xeqM6VhcmDMCBh9kp+I6Wq0wxsfAZR0TEl3L5Frln0IZcBruXX0Wcaqghv9
X3NQJnYuJ3oQLkxnBSGcAKX2h89vqGRdgfGkrYPgnZxrJAz9Gq1C32WdWEQu5fYg
xdAoFKZg9fc9WZU0iFwRW38O5hI8V0SuuTVSPJNsUrbhz8j5YAA+R1pZiHLBes38
iKy8M67e8uwyWsBqh6Eg/uo2PbwHGwbYsPrt9ql6eEyFFTl37+aNv39eJqXD5tv/
TL4i/r2C6F8Rq7JU15b2ltoEz6uYWzoqAWQRNgr9HBclMTfq9wwJgQN0rXvIUkIy
K+uLZENZF+DSvKCjwtJoa9zE2hrwa2yGLDJwxZQg1rnTsmQxheMo7iKxo8atLmBI
J4uvMtQN2peuqXZ9VcRlqbNBtfX/Tu2c4BBwGTkU9Kx6XucN5HcIsX2ii4l/+McS
2Xaws+uZXvqwKafwCtCujJ5O8+6Svq3G9jcQoYbytCXX3A45xSgGqABRmoAmFuij
gBMuqK4VOTzNrlqfI03ghASuYy0FFcqrVMPVCYcUsemn0a990x/OnGUd6rnd+OtG
C0C3ec5aeWru4PhIfkC8RAjTqCtTIED5PymKlOp52ZwjAm1PoV4mlG5VItxLSujz
M40tDI0D9k1Ne7jFg7ytek4SQOHpCiVyGgub0OTsdMu2FojvFh2sOgLNxzkap1VK
zRNKIdy3n57D2aH/yhvHbCt39rVEKTDlTFaxUExbgzSa6IUz2CZ2/YRqCFKgf8AX
fi1BWnzvysa/3IFiMYAK2/yjJZ/kRaSEBf96UNdZzLm9vF9n+23wVDXEjO53TlbJ
jb7o9n0mLC5KVaCUQBg8kE2Y4bzYGB0H5IywbpujSC+EGA8jGcoThQrbM1DLhuLO
DxTa/FQfTstyUgxP9KWdy1UzB4elv2uyRkKPGK5yuo0RRahmsrjvR7QlapGqGst9
eJ9DY5snX0uCqEiabGnTX8V1EsvQAg/ueRNp06VoQJ80YT9Xu8Jlg7S5BTd47Qf/
EPAgo83nZC2owJ74sFRafbq/0dR7hShTcOctszVBMIUFIIEp/xCY60ohPwrt0083
anY/N+kaRVOffoG0dhUVJNf3Kas5HqlDS26rlAkkgh6UfmD3npGO/x0xRFk2GqAb
hfqCAohks2WklONzksdNqLtfNVUeIx1pXaZkKIOwNt8eEVUbaelmk2hC+ZMfETwP
K63NHEO9HqRAzGTIIw2qkXiy38jh7KrMuMK9KENzjRXO3Rac5R2bHf5b0739z3kl
CGPWwciTHXy0OSgs/Rj4GVu89jzywRRe1qFTRarwiwJPtzHi6K1CGjxin3kt4z3r
zZvD7W4QN2ji0oiKua99t9wwvuzOf49CbXj7wCt07llwE8LkmbghlPZaIKK8Xslq
1aUTmNMIJxBk1TqsbL+BdzIi7WGiDbAwiaqCxPz3n1VimXmiU1VTP4BwfZAGhMNX
3eT0wef9kVhvzcrqw65DBJ8twbnlrKo0KzwPkg0FOpeQf6X2/5sg+ykmoEEew5A7
KpwRaEyKK6NUZryQ3lb87+GYL7g9EozjyeCem8bT/2a1uAue5xJzBZIylw/HobeG
JS9Rb9n+dhQK9/0XVUFQOkUb9diPiusbM1gL1FTL7g0ADTYJ2Gw2ORAxiCz0PGX0
XOPKMrXid96pogf8kHwz1oScoBr2Mp6VF4uex1T2dD7iGFTnbmC9bBlgHuZQdrxC
IFIwh/rzDAllmMhHAEg4viBrdHgj/SSwoLLG3Z+WSi3EuqoZWYAYB5LCJphWzMzR
uYO2mNQuNMOGlq34NonGwiTkCGcaTL8GSR9YtcKAblaEpvtKdM1b5hA1ZLo/9myU
weX3SLtMgYGvaKQnkFpozWgfREmj3vrZq8lwG+vxznhUQmIa4ZSzVXFGNZocLBTR
tZveu5p4V+Q+pQXlPDECWqBY+IYuQt+rCRtxdKve/npLYsXBeHUFC6CYVOVwCc0g
89xHLKwPPdq44rKUw8LFmiOsP3XPvsng8rwo0190VeOM/MQo7JBQM7cArYRLNJjs
gmv+nl5KfqL7zC24Ba3Hq0NNJNS973jb+zIpuTeMJ5GQxM93CLMPOWOFYxUAB6Oa
56YsKbrs+f752uuSy6fktWbIMDBiAWrNFsHe79jMpBZ0sp6DIZAuBNkcppUpsZf4
fMm41tERPKmv/R5GlMUoO6JKjyZimyCVRvRrTmOIHRntED6XCI7mxJjZ15nrs8vo
J6t7IPn0CACCFVGQy0orWBCCxUL1CBJwWQw7HQ/4ZFB3ROSCm5h7Q9RbG0vq7w8D
OMFXyOSYm+/9kHL/gelFFXJqjQlTYVQewNtvHsUdoE9L9m2mXhtcejAectfLYwY5
UfbkOH8fdANHhZVjXV7y3K57OxQ4I9utVcrI/xpOr8SiWjp4zeeObtbzAtfwMOoH
IpRLGbb1T7aij2bSdqbKkybbtCffqxMXDWn1Tr0CIbzNTnJCwdmDvDnxKok2bGWI
1VUChwyzNEh5qnQUY/ndsS3wxgEiZHb9kxao+m3LGJLiaCGxZx9HRhYdu5vi5NDY
845zgVuvvI21FzxwVQwaPjImu4DFsVcxJBxT5S9q6YwerMUXos0D0P1gORE93DSM
HEZoNEwwEibYg7DH69uOFU402zI3IEj1r1hqd1VSOG7mAVCXxr5vQLLXiPbGUDsi
C57D9INeSEV9/uE709EGF5ISMAZZw5cp8jwtNjBC5uof85kWewWo77v9fJO98+Sy
5xV8wBdR5NE+2Cws5nuFyT92REqbEpWZCu5bR2zvFnfZYlXqgr7olgSoWvjjc91l
ESndwDqBL53ICm5kBgSoU5B2Cxdf4zXULw7dd1YqpckcrtrerI5xNqIGGIPhUhsV
FIft4AlJ0wYUONaFRY8rNAV/a/PGlupdcAlDIGZYTy48ZpQluGuX6cWo46IZrfnW
yVYO6jnuS6ZAZL4JirF+K6djkc1+VsExrEjYgBDtnfVXFnBvakFtZnxGNolZA5rd
q7G0UJcorr393mMLCytmRH9Rb5x0k2b8LGnQWwVLVfx2pOdFnX13NREneLTWSJ9h
MB7IUf0zm+p53RgOOop99TQQH4mkwdQ6/WzfY7oY5JuQ2NFvcG/B1lzmEWX9wJcE
W0X7anq0FuIO5X47QG70qVjuyk8VT2D6FPsUuda7bVzf+nvTJ3UCOBE6jBNqFth8
pr/b3SufLJVPAQo8prDA93kuyU5PYT0kkheN2HBVKr7ohA+TqeowJpyN5luQZYQh
+OSFov6M0ksDjo1mMhuRa3sB1OFkSry2tmqYoynmmf0Yqu+kjqz1OkdwqQcKICEv
5Gle/9EvTw23IAE+ujUMlRp2U1w8sMhCimnT7nHj/XX1NR5LAJNQvCxtjJJKWKlj
OY9mAGkc3LZJCDwTCKM/t1nTRXcyT/kGkgqG56Zp6eB1hOFuj8tlyyyvuFVCTz7C
k2NMHTeD4pdoOjJi9Zg+h5hyJJN9qelk9jjIYffPpNYcjaVyU5lU18mFf5rARSjM
IcM25eAIYBe9d4S8SGBx5WHOTrC3buQVlDhrAYySYXUH1S31LDG3RSNh+kOj5/gW
g8lCdhf1qhBQ9EkhJaiAMaj0aup8f2/ZLyl8GR3KVabrBIxUrvg9WGGQjQAUfR01
FpfcvUkmzNyhfdLmJwqSU45/jafzAkmWmILyJ712ZDIzHcyjBDil/tnBYNZ/vxpD
HfJGmFtGD6+3N5ouBnNPaMABjbiXOnOofhTZw6jkvEqnrMMgeDI/lazzCtk3cw0C
plnxIIkDAO9uUMjqTPfcyPaXjYxDB+kx9LxfBt+jF30cP6AYgLfhXsVo104em82S
sCyjO53b8CO89z5YYkzHUZQwTSBwUg24dau/8QvKj3gOGz476MepslWlRnHgROzE
tMwA9KSoCPSVY9kGWP7FWG15fc/yMgyd6zU60Do/wjXYnKffpyAd1Xxz16r0jSwK
0tV5+WVZPyrB15kRZhWMzsvyxVIuqgZy/zIZ200CQnOhX9p56HJU5tGantz9aZpd
mawSyr1tNgAubKiJtuAOLtRBodmyxz1qeZhHdv4jUAuOcCmQXxzEEC4Qo16g6b8s
g3fSWjJkUnT403GcoUQ46LenaFommdjKk1pva+OTP5oiwVQiRkf0Aa6EJzfMl8Wj
VYnnmcglGhL0IPLTtxDpVkuyHMBC9z1P42ygmdchaJoVdq6gYX2FZkF/wxPiXwAp
bJxQdaws+1DIvefH62WuSHwV80+e5zsxBIJ7nEufzIJ1LO31YX2GUhffPy2kami2
nc3YrsMUVQKYwyi8BXKeMyUgYs8SiPOTLBgW+XtX8BkotN+YZISun7IVEYCjlft1
JJ8DdAUWEge8zAoHf+Anz2qb5bzlk0CK4jZY04zSR1fVqCp7jn0HI72m8UjArio+
tV6vroL+a0GyCUL3me/XS5yDFfdWx0Az4zKLPqtPY7deVWpWCMlyhP7iHgavE2A2
cu8p/fK2X76hayiXwyeGmjXnlEIOgCuVf3kV4SCrLEQMbZj0x3oTcod+ndPLeZkZ
zaYvN7LeUeOQTu6l4sTpXLRj1iomlA+dArtcqdyKJLvUqbYOTEv3qlP6/kl+uAJN
WUb9LgeKncaFgS6luiIGI45K/LJ+yn03QyHBEfzuZrO36mlAp6AuWz1xWWmsQDBE
F2QJbpU5iNTAiwNIy7TGJVi0iV+Jw1WpgdkxBtHNBoOEdr7sSCM1C6Xyz4wot3n/
/CGTcrszoR0v+fUwDjg+Jb4Dslc+OOlKvTFykWfgMBSh/2FLq4n8doTX4BsAEi/Z
NYsbg6ds66eMQc3r6ahfR0u+d0AHFZHp+y53DBBfaTrkPWPM2bTQOVUrAMdwqnme
C4q8pPcoYLTf0TgZfO6rqPTXo0bLT/xFOJBVMzNGeGV2RSOe12PY1dLf0GF4ZTH1
u4ZsdnkF9635WbHVPsSTdqbl1BqOZfd49MmHZxcmYNwH/SXLRqG6jXD9F2cnpZtl
5j/acRVkHNcnG7U2Vl1MX42ZYsGeXn2ELzzibFifQyhYB/kKsk6zhO3MGUJnPFl8
B4J+o17S3BJCr1YN6lO23qP6LythXANu6cdkY2Wi1Cl7U7b8EV2rhweglqFH4Xr5
UdbGxnQCn5O3kPe0nqwNFRBUtZVubpOFB7AH/6hHSqzIppt9cRJZJRM3w5KI1Mfc
D2eCTB4CWH62gUflE9CQ/VdfMYvMEpGZoFsyV2LorFgXRVHzuweKXVLXl4tEEw1S
gwLKy2nU9TSPz4vjTkjQNw11clU4VhyBC3bHv+RW8ycy8dy3vcwbmUCUgPOonrMb
CfaDENquOMwPhUo6tb2dBROiAXqgLZL+JaIy8PVE3z0wRt8c0Mmhex2XHEfDegx9
gghD204GIigFYsMwIPHL1A9cY5hST4Zv/0Z83VOA1P7+2HB8KW7u7fKk+0BBSXHR
5m7WkQF9sUt+tJ7FrGS4rZCrfnl/mG56VqvAZx6gJNr4gUsgVEW4xKhiVy7pEPi1
6jeQHQYCPJrRDNQZ1kgoADaSI80AFnuH/CrPe3unbZGoWAOIQBaX/+SESCyTquL9
27ReWpVjat9b7EkGofw1sdlOvrSQSBPC6AFbRxW+CqJuEG0eyekGRCkXuIaZ9tAx
sgVmKiPksAysjSojOXfhiDFl6Gt4Lsn7O4JghA8lCElo2zgaBk+8B52pJXdWPUxJ
nyTuHzWPfGEUMokUir8l+WbG83hvoKsP13GfLCfWQ7Wnhzd64aErfo6ZW5GT5brD
AV9F4kkwmCfBtYpNz38gDa0KkRP1gBT2UcFsjQvOzA9NWfHVmgOAxhGWae+ScrOF
WgXWwgRRt90i+BlSejt5zWUG4K3gpYFs7x8nJNqgJjcMwTxWxK2d7lDF1iwu0Rrv
XT0XtLt0DCYrJ4jg5PSEKSXAgFlPxuW32b4Os3SHRWQu61D90OINAquA3LHlLRvz
RMaUD4oVfRBcbMpk6w3Yml31I3c4ukLtM9HzbI8oJx41B7qD5iTIGe0olychphBk
XlaAnNlZGkHpyNhW7W/AFaidBVtkOb+HS7jntkcsJ9PKVPUYKnpIk9AQsYW4x3Kg
bsdLrM4g92TI261NmiYbHYriauV7GEsbSX/ZLvkOdEZwCxUrTfi/i6Sq4rOuG+TN
cDKiaDJLewnO59UJ/jTZgdutamfTmftOF8ug9lClEPGRA01U4QOpsgrCyNx8bO51
59KE438eV08f9l2IfHLZtevW5SgDgaM5BIYSoQ6FBXbbDLe/o8mRYPByt9CBY/Ip
PnCdpz+WQGkHjkQagoi0qSuBjNP+2i/t21UiplKSpoVMDOlb1N24z57uAfW4KxRc
SpSlSeBhCltlTf+OxMX+FWgdjBOY5G6URNIsvHiFvoP0fXvlJpzRVLPGcGzFl+Yz
gMKAkRhL3yKTGAHEoAYVzDmkN6OxZsHFL7VNXoGKjlikj4sdDcDmp3enUKyfBaMd
chxW1q3ojzgEzcfXKOAQYLzqQMh9NbwQ+v6/FYfjqgDMDJvA883ZONEuHlmM630t
T4za83E+GIg8PbA1Jl3eM16lJxL5X41cZSC3vgO+Pw8YMiBMfykWOpq6dydoDNB/
72o6nGcB1hk94m0O83KBEkDvGQGJbIik3Hqbqoe8GGtjw7aZnbLp+PT1u+3XJ5hq
HRJv61kto4zulrRtkf7xykkCgjqk8VZhhbjGjbgsjqjkqvMPGZYBVZiZHIDn2aR6
H6ssByDWB8mq1Xs9vpRCJ0NWBKle6mFcLrzHhGKQOrgTxWUSpguqGFSw06lOK+yL
bF+1C3NPIHJZpzQTQ1HRYogdlUNI339/3cp78H8Vs2Ag/LOuaWWLE6daF1Kx2Vz5
aaCTqa/MGpGpPD2yos3SA26pWcQzJpa4X0tTya0/vUs32dQIdZz8qPuiHfsHtoPS
UnSUf9X6+5xTu7QYqluoo2awSCue0txhsnnAVHirlBkt50a1jxVm/p9okQw+gTmC
oxtmPS9b2wod/HydNNbEM08ID7wBYBKnd86012KZaeCOxVFzulnLd8BiIU4qjD0e
ffLMcX3ITZEHFGO7yajCJwiCdM1ntW8BJV1qVvO/DnihE4G4POfww7O8peCINvhw
AhWCmRqVSf45wXxFyaMcVBMMvXXUeb66AM4AKQgxcXm6sEp2jNQgUnMEJ1JweYtB
kh7mIleIExFYzp7oMv/RqCshFV7vmK13SM6Jm9QHPcquKfTtxVWge/M/wwypGUqe
j0dYELJrgqsj11LIlxDf4yTry7lv1ikJG5VtxlX8mAe9D92rWTKKn+DbFEJNFImq
luPDWi2LgLwtjfeJg7nJaIT54vR6vZHflCB53vbnjinBgkOCn/NWzGFnXpMVn1Hl
vQNFd7QQFg+X4qr4YdVuJS5SMNduoFmnH5dECFxtwv0yIywEK1lSKUm4CYD1QLDP
AjxWZOQPSLcgFcO2iDmJ/SUV1/QQjWxvLhTSgk/axVQgLzkZdPX4CuqkcXWV35r+
Y3+Ag5VRSpAoTHwbIUrNP0AtBgwUBzySFP6fiymYsXnxFcC09ALYgmHGAnidGb/T
JUo11//iIuK+r1rSd71eAZKGjRq669QnojZghp8xktknPmeJWk53kPq1fCreJk6c
H2vOXyHeNVxhcfNTyoKhUU44sxB4uyi1ibYzmtN4m0HKAPrZSniv75JVl6X4Xnct
Yigcv7RvOZsA9JWF3tTa58ly85l+3GByybV9dPEdY4jW06hrMvbsYqvJ64hN3bVY
4/89RtVY/Zbxy0r8D2ByBcOp6srx3EcHXxZm+AMYpBENVSRRu2QvkvCkfAdpyvZz
eKu3WAiI7FJtIVVWKG4ypTztr2Jcp3kA2tZdQpJ7JM3zbTmWAPMXyfo/lzAMOkY/
ngxwOIvz+tQvb3ss/ZF3oQwbyQVUHuKZoGGoxgU/5AHdIwaT2bQOglzcRGr14WEE
FoVe+kELkdpuT7IdRuxoWP66xevIN0mCjmoJiw4cvQDmKEAkKgGv9SaDyuq0FucU
HQ+sXvjvROrUhhyjKCJxczvwDkq1SHVobBYdH1px3vbNYbHup+vEsJlRVImwg/tt
eM7dqKFHDAcojNgs//xh4Zb4TnpDZV28GnjYtko9veJ1A1LNa6U4WUCkHtmRc6LI
fgk9Dk/S68jr3J8Bs1a89kuSHOdBY7AG3VjtG7VabHdqvh0+ruNe07nGWe60Ka4L
72QlVzJcN0Da5hzjPS2n2VO2/57pOvF3H5q4bY3dGblC2MZ1elDjem7vJthq2yAz
SAID0Fgp2s0Hyce7JaBDAKEmcmtjnD4W+cwodYM/OA14R9l1Fk7RX0vI9eJvNq+8
OFr7v0zRYntyju+7zSitwv4XScHukACwXndMRomBOxcu+5+46izd2c5AVyXhxmoE
x9awwqSA1Ai9Q607zVv86BVUoCSTV4+PFXE5liTvH356RflSnn/2UKt79G5TyXxU
2LLZSL5B+mRt2wI0c0TEwwl7AVKYVEBjr8QG8zefWQbenSfX5AhK5MI+zmVMZCgn
U8IJOe5g8jXKmk1WVrcDKEdakp1ICdVHIuWpzbkuPPGUsBcnIPeh1P7dA+DmMJQa
YASeJ2jb0qePdupHLKyFMyve/r408wwX/eV9wGEw0snctDmFRBNSZDH7WtoJ3AIC
4dmhv72PVGZ6t6NWs1gJAxLaMpORSytu0UjcsuGPBU6TIT9fgf7J9WrS+NJh3jUW
4JwkGZHa4QGYK/jD/gUb+ToVqHU6W/zM9Q7v6FpXM/duqEkbGBIR7zG+Uo7f7mz5
BMWOyC1RuL+7rSGZccdR+wAvJlB1Q9wNj3IUKIRexO9dLr6CAyLlGMJaZEJCANmy
mTVVYA//2+m0LsqhtKh5q+NEracm9Oxwq2c+jnWupLC6snaN2sqsz5Bp/q4c0Rzf
ZT+a8dsmY8AElciduK+kMov0wAVoSa/59aamTpBYRrNjGDY35xFjn2py9K11nPC1
u4GVGTpKelVhniKKO8wgzmAPRN01EDV4U7L0xcgowQAFOXVf99+ROMK5lHfNhlJs
TdPgafkY6PNYkPz/bveJt0D8txJ3PaWo+RHqkDB42KMeKXE72sQzwxU388ldCI1D
f8s2SN1kjI2uL6UD6CeInaZlywZMww58ISu5soyCo5kDxn0VPpF3eux2s76YAlEb
9qyPl7IjYK1UYS4YI53fV0+kq1B2IZELErSlWebwLyoy3zrWLGuQOTRr/PdKSe3i
L5dO2kXCL65Cm5HkOvINV008LP1lIANgteKB8OkR1qO22t01o7dTI1mSgdu7VnUP
gBq0d4JBQzMyIU+OoMyLMLYcVJcUh70Yebs6LO3wATTocoDKKyCFTtWnTOuSNBKz
ef7VYhUWv1TFizc4XSEI2U5du6JW4c6dB4X/tndyuIX44HoGhn260dZfQ5gtRpeP
RWCcQs18w/R7ghyCC/nIhYUuHDncGqOeoIGuY82/gcBuAGyFzLOu5FH/js5y+KtA
j2aUWBDYzD/FQCNs+BnJMq08nqjO3VbnCXfZCa3fYfhtqEMj2pCRbXjejoLwmDcY
ON5me+qcKzllFyLaUn2nMWIHgewVs+9Vvx7KxMOLmJkgLsWYkA1YPg9dnyFQvxuA
NShDRYdQdu1WcYIZlCsn/F5nHv2zbM8/BZ/+WAjgjHptJ8JaHRsMk5IrjFqFey3g
fevjquLgdkr5lEspJ+AMX79cDDXJxtEX8zO7P3hoobxWS4tjsTUZK2v1BnH/0DCF
4RtBBVLEI9cSxVGmYHHGa3gaJhgoutAJV6AbLnnCZjIlO2VHf4TT+lmQg0TIJU0c
L6/uC6Kr1bwCecG4O/8hW1dpy2q9BDV+p55WpB9036Rpgw4tSmmzYOMNExfe+hRU
k5BLCvUGSGRatHT/D16rf8Vhnph6H7e9DAx9cG2Fzpf4Vqfaejx/KlSy4lmeH45p
Yo7kr9Vfp0JLgDtaDRt0zbZLVZqWSxwH1DW1qlA/iXkosxmZRh4NL20PSbjSu9fz
Vvp91JpOJBC7JwsEzoUXjTzLO0HRirCUlnsO9DRkTlyuEooa/vlZ4b/gDmhTKVT4
di7YyobrI7Hp11Ji5isjWqE7oOkHR+lI79CVhnMTNf+X9H7ovSwoz8/YCurWwbR2
9KscQGCAj7JGg6FQCc8SXIBYfVePaAr5/nJW+mxoR8vPVAhPycPcog3Np78ak7ZM
E9/HUg1gnFg45UFA2PG1+WtdRPXVVTU6nxZFEpK7g1lx0JD/ZgLl+zkR8+Yy3Rnu
7uqmF07THTo/5iobCxPK9AnKst57+g+hvkpIEasYGqB+WKnctuShUrC8PRMX4ly6
nlXx+U3Vf3f1/YOM2PpnEntzZ7japSyN9HtDzu/CyWytUKMpoMy0jDOb+5V317uL
+bZPcPtlM7ZNtI8rzggO1yd1iB4VXOOeyA+OErWPEgIUF6j6jgkpJVZ5o2Ap96Lf
QsT0keIzSGW9eHRu2TJpJVMD+emlijMREkcTUhOrFEm4NA1pJW3uTg57uvfYv7FS
CqzgeEuzuJI78aEfWEPAjARNXDAsJAU8fdZkXB0zKPVchpEsBWXX24rByi4lE+Fc
2EybJnQpT/rJ9CDMF7gQYPdiccBdYwfNjxVdNa6I4aZJVjPy18tgBLZ63YUNdRfD
yiu+y2xXCxnrv3hoYws9uRqvgxdm1o84RBcVJ/c8LAmcLTZ/rcdRn1O8MMK3aUpm
UV0TBruPEzN6p3NeGps5TNJO5MN5R4x/KpTSD+JukZdBbZf2DtEjEmakEE0aCnph
GIZgnDeuuU2+sJDfci6FU7YH8DqOCpjr0IM2anwPSWTygJcAJBmo+wXF5hd9PKqH
cmlwv+9pVhiTVkQuuTP0nNwtn1/8xkA09Kll4WWlxm5WFG/ZGqFoaCGqPnESVfQ0
CtPezOkAaIBCGXe8+ApPIXa1BDZBiOrurAfVeyLmLp5hV8aIeJLI8yYsfRtpEqNh
zkspJwypoy5OlW4KyGHnGPWrUfEA57USIreFEZ6kwdrLDmtfKis+D0lZekD6BrQB
Ts55HnZV62Cub+cEdpzqmQwobS91TDzyjFa39lqezBJvnU7Ph3fW/qI6kw2ff1YV
WB2FukDWV5RPnvfEJLxu+H2/CMg722Vl7XTLLZQjE7CbAmSetkrlK0KsnARZWdIn
ZhRADikBpjTzO4jXDlWUlv/Ef3nOyKQh8JWHESLdkfY/X/730QPvugwvxrdn/2xW
gLCrmZcIoKBqVCScZFeRA7TeLDFickQKTw8rD6LvGUy3AZHxTgFTvL3gPA5LUgJy
1foTs70MRC12cRN23wfkw5rlJ6cjFJv8+Pnvp97Yj3q47VSn8Tsy5/Od6Kk5/gzD
p/FjKMbJM/NKsDNM0ZO4HcEiuqGW+/0Fbe4NTV+Ststo5nA36Fk+J/OzSaognXGG
Rh0cjuR18RtMTX32OHzrsOUfOoLInedn7KwA+hl4XPzNUNjLjrERHMm1S2TjQnSF
nzz6/hst39n0WiSfDWenztopWIM5IHL7HkII4weljRoZ5HynErknipwMB3oFpt9m
xHc1CuyJwL1AedLIRj6YhRrUyxmqmNiuP3a+lQ/zktz7y1DhHpljrcMZWGyS8/s2
Tm1Djkh25GzXYRJYoXR5/szlxG3z2Q0VxDm9I+qCHZzkt7eyRnJamzXG33UVJQw3
shVsed5N+BLepr99aR86Uolpz+7sqoIHIh1VySr86XjWg6RydTBalTXLfaXKhkWf
4ITW6Km3Bv4OmxUv/R/ZBW9dYRff8q8wxm9G407cCvmyZSpx2lgHjP4QvFafmPzv
dDG6QwtzTSyaijoHLETTQT7owxk5lnaowCOccLrNoxJoIuuPNgJt7wmAmYxE10JC
/e53BJbAnltyyyPw0wXxVYLGls2sL0pn8x8kbwO5914WmogBb4PPDa3YkmSztiVd
sVYHHaeQJ1uOW3iolEmDrZ/YXxxWSWwSmQ2iV6u1KxVAlGhwrpdtEM/ITE9mzSW2
5GYUwTueuvLv8StL/kG76H3JhT0FQYJ3AjcRzRu2DzknhLaVkEwXhFwv4LAlkw30
i/43EaIxnLCeEuuJflFGmqgqRixdMz8t1FzecRAsHyVnwrrZm9d/CHx+MdD3CxXh
xlv2z5eFgvqQznJ0fyJc+fD8wMpKy1w79MvTRkOn+Rq/kaIsRldTv0kE9xs7h2hf
2PWunB6Sl6rbahTg4humAxUjY7imgnNBqNkTSBAxPyr1HgZ+Ig0bvAjRkKeKGTHb
gP8+YANsPX9vFrl1fj5ronbc7JqJOtq5u1vbazysY2rmrsGtx6BnCoqUptE39t+l
2JtImGfHU1WV+dt7IkE8c3WKuSQBBZrtjkINbRgIUvfpYSqzVzlUM00l1CfDVPi3
Lvy0WerzDQIRzbQ4nwzXczPcT2buMtckIXVDH8JEAiEeaT1SiwP7vl72b03jnHeC
SDqLdx868btZ8v++h6mlbZddbKVRjtNuE/c/DGoHzK2cJIqPItVq50J3nXZul5nw
uEwnK8FdAcIJBgUwOQRcRbzo3XSxlEO5CJmIKgbk20HaaXDwIlBcopQuNgyRRmRe
6SSfW02jzyYYe07X7vwSfmwxLJ+6ByJvjpFTl/TadrYqCd6nYqbYzqYZpkzloAua
sU8lfsg4a6xFqF6EuDmymamS5SJ1MFn9QyNgpQzN82+rdBk19TibfoCdwc09trpz
a9+esRO+oBw8KI/1K9rkiSBg6xijUsALs1N9wtv8n2dJNJVVTqW8eGxF0fy/EpBb
jgRHtS4W5LVFZkUXAG9TR3Fy2I7RhlWlpRvvu2+NXgRkT5yXo/8fgsUEV9jSJAgX
obJPoKFzA+pnXJ+PzgYYGUAS143JN2Ax+j8ReJekBxE9mQ5Cen2LC59MKiX2wvLo
xUN5KrP8GD37wNG88mn8CNIUUwQpJqj90XXWYr1kNBrXN192xbqXhwo2dMTqhiIt
xHB2Ttz0o+Gr2aiOyCgA3Y73RnCcqBGleyWlotj8eav4BtKEJQxQv3eQP5FpWQ/k
pPoGGj1OoaReqVpVp3Lkw0REdNe/EZ7RmsKC6fh1juFHiXI8biohZtAT77U/lBPC
Q6voayUJe5XV8PIB1/Sz+MZaMxpGhJAVYslynm12eGcEGfy/Uw0z/OmU2tMLMV5D
4u1rk+Ilw6X/PdHrn6mP36ehIiMwPH4Cj6UHuYMgcUkvaIPeJfD4fGkmr5+7h7nN
U0tQA5ySIoVCwEyKUgmWIKZhwwp82XJfNvuYhMhZCRFaEn2RaUMbxWv/ZVrX1yF0
ifpwWt2X2Mfal6110uN4gVrOAe0A/OkQUGiVdLF4829xrup1AjYEcq5hEwi7ZPs+
v216QBvXe1Fld2bdpYgbS1UMKBKOTitsEe+RSssoYgKt+ARAJAPOHv0X+58m8MaN
J4aysx4YG1EfVBIPOM+bXceqPjszFLur9/d+8E0Kdqbjdsw7xz+8weNPL2SCoIdS
qrrih6N71OEbzcpOt7PRI+Ox8nbd0Qj5JpV/yNGzHpUd+Oo38pyTQNYhUyM2R2F2
Tx/hQ8MsITQs+p87cmqOiUlB76WeLcDP5BjmDvpjMoEPNoWqPgtaYVp7OR7cNOT/
DZc+rDScRLy3lZn9wJuK3ElHznilA7ym9YdEiVwzOWFaD9s3lc4QGGH1lgRfzNKS
RvC9HeFLYeIktcwza9+IcqbZ3eT/FaUYHdGAUSmbkg3/+8RGyp/ykQ1hPfc+TWNF
MZ7zisDliNI9PgiMEdmSDTiJ3oszzdp5/TD96dXFg21PRQRMJwNDDKoQeX1GZ/zf
rYPudKkqydMKgrsUVszofXMuL3J31e2JuE19zgafVLugsCV9HvbOkj8G+TwYgm2q
Pk3/spU9Go6P2lQvZb6iZZ+/fyRVynCueXZ/kt6PHSU4MwNXQuqOaAkw53Cb1u79
Pk3FEqUEqIjJF+v7VX8dntpJgglZzkdx0GEjFogjxEBGNMdWhPjy+1W3HqSWukB0
iXEpgXJ6bmObUGsEKtptvxGJ/3ygCV+t09baNHmuHUB0K+9Tn85yvu5LuTpru1aY
BHNlBdrEMkDR+xtXfub5Awb41nM85kY0AJAwdjC96aW9R4h9OzKmLS7eLcrcRplr
ol5gp9alS5XygIzn2eeoa1u09rAeSFRAuOraWa3WKAk5bK3AN3AcDW1Eeo4WUoLZ
78SaT1Po92CTQ/DKJ41IPFWd2mZBnPSButOj7RlDMcFNoEbah10npXLPC6S4zIsR
ifKmAw2bDqGKODdziDJEWpmIRgQmZIIfjbb5adaTB3z7bNn9k/hcfaCRvi6Dfwyd
f5ZFgjtIPLZzR0iBCtV8BRvKodvLv92EHpynfqUpOXUefJVqANNAl3rXtjW+9XcO
lPJUR7fVr3YJLKbRhRSoR05I8J5kMBIvX515BGmLEaPw2rT9Kl2hJilFQKHF4O5w
sB7gjbxT2gVsZ2VMfKApK/XpT3hh/ZFb+GkU3sh0IYYH+wK05hhX2jlkEPqcR0g4
24UUrNY0OjUM4VCS6cGVCCDtJw94RA7f3g99xCCrupORiBpvOmfp1mqpoFgA4aag
7Do3Ply8OiZR+tIlanwTSPevvTI0gXfYEXvbqINqaKqkf5h+y2++XUSEMI5yol6C
I67UZdsJMxNhvogesoot+kDHZ4FZSipNO/JNX40D1Uqun1bODxXfH9xE6GitFRzd

--pragma protect end_data_block
--pragma protect digest_block
mmrzWwC9ro7fet/HncB5wjZ5pXE=
--pragma protect end_digest_block
--pragma protect end_protected
