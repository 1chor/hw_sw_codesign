-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JOUx96nGSt3ZavYR1kHMCxcJ6BgTIXOz0L1QfEqgH3PSg3AE/GOxqNEasmZZ2C0klq/iE90Xnhmw
7WeW5JmDTpPL1J4mefYH//ypJjtg1M1nTxXmtbZ0t/QJ37vq6fbIw+283mxFNULMjSh75KtGAeiF
6+v88sISMnMu2HT3//TXzY9ehsUouEaH2e74cGKwVPHTAoydKMR05/Igv1bKcsCZFcp6ZSQZTD71
0oEEsenbAi1JqRxK8aFZNlH8ItFO8VvIj8uVFX9mxa8lk5l9SuoL+UYpz7ajLvNxj8T5pLWEX7VX
EH5qhXLm6/wzLF8LGHjgUeGJbZI9GGnGxi01Fg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5632)
`protect data_block
aJBluVMyGLFxdrVQpK6ecOT+/hI1xIB96KjNYka8hDks32yrT7HQI3NEIiBfjUr6hqTdP42hjrnZ
XFK+XahPTidbziQRUs6u7RIpH7AuCwN+u2UYY0jz9d6P9+6eFWlv7RfHWyh44C2MxqUerDGF4+O8
HlEqrFEEfbIhV2g0pWJAVbyMCTFX9X1mx5lBzATi6VQ+P0BO2/Z4DIEA8qL7wV5v3wwdI1zuRwaa
Nk+qoeCfNBJmhtsB5xlz1jHvAcWiSSdeF/jsrMjS4s5BbJOhpvt5KlL1VgYK2xFy0NoNhjkVdFFZ
7TxtAj61DbMTa52cwqcyfe9/F7FjSgLOLyrZ6RPO4N09rnXj3DG4gGhEJMo39q2ZzutFGvBA5CK5
Hdshj+6LBgZVwFR38Rhqnk6SXr6PxF1GxWxHc/Hk6fKxqfejj94tsbjfnDrhHk0YekUUSBkZvKka
m34Fq68OxMvsoWJ+V1FwW9SPL08vtVkfV8pwhtqZqt8CklVj1nfJUhfqymGFeBSHOsRD5dN0Zo3t
hUOV9/hikoqKgdacBgyd6ZB5YLcIeRCxSxHjIDuo1AdZJaVkLrubh5KbTN+86fcQXob4PQEXFMBU
H7ZDyjEGSnYbkf9iYMVsxAJUhZqa+bNzmsu1ZUWqgvFurZy+jbAfCMBF3ccDZqnMkUTmDUNVBp+V
uYIQ3mUWYXKRYFI1P/mi3XYjTCiiLlBc3ilvFqFLvw0LdsmC3voX1a9HCVlNfsyxrjfJ8beH5Xtv
KFOZ963qarL5F0X6OLwTLWUPemuo4sxJiiNrow0InmtueFRxf1Puc8KnQrQqzEcBgzZvOGqZfO7K
7aYlZxZ2OHnlChX675FK3If7Xsy30IXxfmKeZeu/ty2Frz84HAXSg0pK1gGYRoFg/8a0AAiIt6c2
Nu8cKAIow+54HrVD5Xay0Y05oiq3cYr1LN2aJtlL8EpGTI79+8nvjjqRbPt2lDnOSg0gU1gPEmom
Gwax4gvVX7AOP50lAMw7uQ45ycA28t5gEgU3vJNj69ooVHuHBmiQXK6/maSGEo35UWjYT3YmdLpE
0gnUGOuf5pvI5/NL+Ler31WIeXmI37fRNacmxz4KXJOcL4J1nCFoA8BV/2KKRU/G/0W1Oh6FKcxA
+UyEqyChKt9neVT6Dg7YnfPJ/x4ReNJg9Ye65Jquiynleo799ZffHNSmuKCckPJKe8y+A2ibfRwv
wrGsS9koAmqRyc+83KJ62wYNpsFYuObuKlaAsioyRtCT3T3SGGS8Jld4BFI5e6+nT9qRZKsmSQhI
e61LXxcpQ4u30u3bVct2KLkzT2+1JCwVR9v+1aeq42aC52hZY/WOe7ks8q867HNI1afgz3gCvm8u
FivVHJNXnjB3H37qzGiLO2h+QWb9lnVFYk/wcU9U9R9BKbac65u2OAKpx7QN/nf7bgvWehFAO5F/
+K4PKK+i/rNGcaPJeK3Za3NhaOamXYYN15wKHra/JZiVf/WXcAiKJOHdBY0rtUp9pv60Ea6UF9kb
ANYwbTGYysY/9nYuo7b9zPxaCuMNJ1oF1aAWlnyAAhxAqjmFh7NnWMZMAFtkPEKzMa4l1B5SJm/i
jDKkb2zyrNxclqRIxSaa5zCo6WcGlxxfkl3GUBJXYbGz8wTXqSnx5EDjGjVGFb57iaTyMvmtU7E2
bKdtKJMF1XtCaLM4x//lig/jjEUGwNH5W6hcF79TNDmcd9WJehb12bmiR4ahtXzWqdy9WHJgVRqW
BC2g+euamg96Q7luF7JIFNqZQQaa/vvBjBOuquIz8b5DCnshdXlJjhq1R2KCA8Os28FopKEacEsm
qdGFg+oGJ9bPi0WgLC8JcaZyJF9Z1Csl26GkRsSVKn/8DNQu5uvg9+spgxiNIuOkK/rsVjFBzf/S
zBsxD3ty+1a2D7OHrSuTd/MCEkCIAK+PcWOPtQGZpWamBU1JDZWXP39HV14P/XK73xzKO5OyLzBp
eeZEGWkIuXdnlAi8g5SUrNpyzY/7UauX2YYUlu7mWrEfw4IvMr1capVA4hs8cIgUouRo2KTetbeV
4pF3asPwPepRN9aIGyuVm9xCb02eVrqStj03mOoR/OjFllESYA2EkVaMRHkc3nnf0oQtD0k8Kyiz
xIGZlDOiF+jAysZewC7PkSrd390+o56njb5dZU89YeeHzMXihbAMpVj0Ct2wUuW3l0zc36FfcRFW
5J48GNUo1cpWS+CZ+XObx4b49GLeJp2cEBtspbCj1ru8leAZFB0FFBAqZ3MY1sEVn0G1QwQMVZh/
DaFkLSd/4HAsXnQS2/OA0QYSCAAqZZ7ghrvg/7J7EXnObvrnzR4bUKaRVV2/rgJAx0Zwo/6gtBa5
1NHoBXvFwQ/sR2wdTlDT5sU3gPNA4qO55CTzRWdbTi8NL42h+kRTuSRYXNn8lqafANyI+HCoSLdY
LvvCFmbTt7cm0BugzFz9oqyOLxaM2MBQvg89YHLax4pxIyWjCKjm9bgGKUU5MET/9JD/FRh7a4DP
s/KjlOl1uRNaIK7F2WlG6cnqmq2K6Gjqv2beIl/8xmzgyPVg4gdOk3KZE54RCgP6Gj5brkKezB2b
VI+hlhUxg9WrqdkAmjui8X2pWMPzhNLAzNzZFLZVFjS6iCKAne+kuBRz3XcDDLfwSH1gPf9CN13R
FysuZ+AjiH0XVg0ThhHY4+mmsbsdw8xmq/+0mQ13OwGytEvZpomldWrvjhVd4CTS5NRc4xEPHy11
c1ZaqhQOwI/Qko2yx9Mn5vnsEJqRSA7UWJQHncg14ITvkWUXbQcV4D2b/5Z7vqOmcQo2u46wOLcH
Ogxr36cav85I/Vbqa3Xe0OMCRy/RtV5E0S3xvdzeGKG6dKU039nxCmMOG7WutV7dZupYeM9q4xCd
rKxecVqGf3v8sSwt+BegAdCBM2M7aUPoyeBgnFzhn1SqHW3Wzhc0j622jPyTCAVuwyyD6CnPZFMB
Lpz2CUW3Co6JZ6I950KS6/sK1cep9AbLZ5ml+4FLaJe1OJmexQ12QomalhKD2Daz4NyidvoaW3E+
5bzhsL8gmap+iNwkBC7MT1LHv5iUPFVAi0ZvwIEiaI1RGj79xHzjFCAlJ1lBDwyAuqLuGSZ8MBX4
u1iqI+YkWvs78U/cFKH5lZMu3NmoT0hz0teKQ9oZv9ezfvMYxT8zV9gSvglDqHSQ+JEdgxEMalNm
qlPNxYvTfSW4TH9zHl7J04CB+jSLA+6meLvc3zZr+94oUTtI09s2iQzxHzWqO4pktSeG9cisefyb
78XLAgXL8+1JUhjJYmXUS5zPw5M5SqX1+UkwLjbgUXsPgX1fcDBcgCupISGD13u7LrMzNdGZ6H1w
CGuUQFy0pH31USt9gYQnxI4VhL0OsQzSvcynbfCvlJIXvY8mEWGSDT9Wj0uZSXovlkk7+qOeT/pa
EyWl3+OBWZSADYjodZsHwewoR5W+8nbtw2MYPNqJhUECrlIm5Dd+egZwRPFry899FAYYSVnQAxJV
tymTar5udamY8TJUzRiz8Oi74hsiE8VsWYtKezqT94LEw4RTsQGHHxdFDvvGPIUqlHxEFguQOd83
zyKvWf7etJFLd2W8das7Oy2HEujc/cvprnNuI77GeSlqGKA0i6XqaI2A2yqKov7XKD7XI/7rtSYD
nZGfx7kpNJd9P0699vYtBAnAqSGPOgulLkY2gUYPixT0J07Bl9l4OP75jjwXutZ1D5LJedId3gK3
tkYJtOzMusDt36y0ANoPj4DaSBLiRQJyX2EBTESx0ykk/vuRDhnqA+b68RZuop/fd6EXZplih6yb
XA8pgYKYzKP4nBa10P+fYtEGTk6KWxaK5aiPH2UAgkuTw4g46ZSv91K1s/8wmTYPfX2ETiiOjEzs
1Q3LHfMRm1PEvzlG+qIZIRqObC0x5hQNz8Iu080WYxhqLY1UqxC5oRU2kcgiP9iJIowp4oScaNu5
vakR/hkqPIDI2KEOQ3qaX16PqtZVkaDXBecB4jBnD4yi3e0b9RK1jJuMgEE+oBZxfW32bnoy7yxG
RbxyuONXD1cgKKAIxxKF6VHuartp3s0fIRozuH3E2MgbxOX6tQwtos0/dSZx1aukwcXsDEkx8Zrx
iBxSPv3KXKspIIsPTBSNdJbDIx6ncTC7o7SEypNowC7e+jJ3xM5ltoRTr9p5ejF5eAwJeclkm5fx
6/E1ozCrb90wJCSsJHGcBCTyCMNEPoTGT56JUtsnPVgXA951MeU1uRiMcBWLOw02/ETS7q+eYxq+
dsKRLABOVQaQO5cfhtbpA0Vg3QxPxtAL4pGsvYAiHXfxr2zuB1qMpK3pw+kN7F8kWwRhh0aqWs2E
QMALhGlQwGN9XGKZFG93nS0rChZXO7Ij0bHApcYqbKvAReq7UDISvUoR8f4NTlR2zqeWzISbxRTZ
a/5yzhxc8NXd7aJXMz0htCmaOcfP4WxLkFPsun6m15DiFUNjkjeQM1rE1GARGh/dn2NkjynZkhJx
2PPMBZ9OpJ/OhbGiiBL/FGj/qdu9Fd16E3M4KgBcg5pQHo74P6vqLJOOXvWC/zmNe8gHy+3BkAy1
8tOMItaNzrA45kmO5l08xrp/Z8Sv3DM4a340WNtYvxCGto8WLukQ05aWdR70/x23GNuehhamQnmv
Zicb2pNhddQ3mobZH1lqUCtpBgn3hEop8T0LwGqVTlj+9rQIoF9yzCj0H/9TXaQmBkiY63SoA1os
6Ab5OdDO978x5kW+/MBCb2QcFjL1tG58TSixcC0r51JZj4YblDTLIrBtg5nxdJmZ9t1sgUIPinEI
gvpFikzMI15VzNzzc/siakvJQt56RRSCV9koxvdgHIhyzbabRL8fCUq0gpgT6dcmUpnJePpAd0gb
PXgP9keqcqpskMRZ08PCeOI2LBKjup7R12/w+y4GFYSl/JCgAUvFxXDk+S2k6hiqUHVpqk2TpgXb
Pd8aQxAhjhwKtBlJ5tA+UnfFih/KoXPUhKbOOeNJH8sHotNY9Heb3urpVQOwTE+TIvNScBxZIJcC
jdJUy3CpKxGqFt4pLLR8wtQUREOpwb+dGd7tUNJYG39CJW0GHcte2gFItBIbMNpJhNeczDLYfKOA
T1RDCG8NOnYlPieC/FinQV+7LbOLUrK+H5nP2mTFvwD0wcCLNR16YSr/qjUho4eoZKHzKsNw+cNa
lcJhV80TMK2F9Xp8jLrQgeWW9ORpVXx0xI+CPrGkocRvdsV0bJRwAEZ/Iyx4tNglm7GTeyoXIuWs
X+srafAA1n9aQQoJs2CzMwiPBzfvDk8FBksumbzSokQq7/uxWAfEV4+ZXVjx7DK6sHFICZTK0J9I
GI07LyrmU1Rss4rbMC1gMlVdgBTzCyULR3wq3TqwjjrakOfDQCKy8CyMELUPifx+Qpswlri/2Ijf
R19BRnSkFDnbY9/iGU/8/BC+bPpXKYaFYxRtOE1+BOx6MsiGzi3DodLm5oujy7f9i++pCHYlTG+m
m3W0mQ+vIbQ91c6p0SaCvU1kZ4TzQclaj9oGoh3AE7ymMSIjSzsDon0GEMYjeK9C0sGYXXDSDZok
kk2UEt9HKpIsbbYIe3+3aQwcn+sIhSLV54upOtvE1T9TTuElZcHLzQFaZ/tTfPL9HiGklmSlNnH7
3eHtuWqyzIHBr9ZtkkHlrQh1sAkCpGxbTE0ol8ygHZyQTyMzprW6CUFZGFLVYBXB+0FnCuKMfxpo
X2EdoLOvK0LTStOHgxWszzSN6e7Slw3ytBh+iHtHLqyZCZtHiaQqIncB6vKbHEJlWg2nC5ZdSQIU
zSGdzpWj+dqVVue/nMF3Q4GE9OKfSyfEvC98WgxKqILLPD/chP3Y7OOKG1XX7Xet9UQ+GTYqfUkp
Jif5RiI+sqEoISS6mIQTZCyP7Yox8KA12A8Sab6ruOr/4WMgDt3N+8wsil9cCp/nzqWux77/iPaT
B08RrSGqCp3sm81IQHmQqlUzMPn4gEUBSN2/lHc/bG6BQq08S4Dz9WX6SxBB/8p1HkEqIrsLQmFv
UaR+Oy6J/wI8prhWh6u5ydft88p5rMQU3TESWWQb00oSKN70VbsTpuR2PCCVOMXSOD8SFzJRdvyo
14Z8ss/KJClQbMwRkYy93y/Jziki880jHpppvwYm7XpnlfqncXNYa03rDZyJjHWx3Nnjh/ycjCD4
CUddE7sKb+FkIw69nIiFNpN3XhTDJ5XZY//OVSBGYcN7YMsBpDc/gW6h0uo5bAQ+999IR6x/x3pU
gCq5tgk7eq12Epoftj6K24cshF9epJuxwLAYSJw+JqL8rFnme7rW7Hys7E5p4LbuNDYx1Cqu6VVU
6GHpbl5xZl9rw6L7RLOcZCUcmVcZ8ClpT2b0SXQ5HQAKOTy8FO7UiJruMMUpFa8/KD0o+qCucIVt
FCjwKxmhBRhzRyMNtX8mv6kEXwjQMDR7SygUgbHhs2aAdYepikaUcEw0dGgz02jmWOAByQ4ZrBY5
Sqt3fGncx33B0Cozq0dGuGfOPyTlVl8lVOadmxpaCqQlfVX5RBKR/za88JK8aso71Sm8sf7qk2/r
SvIOtl3BXbleYQhBbMvEm6cPNxOi7eUJ+S2BDK++wFUDdVo9fQiz2qao0v1YnPLJdnAHKH7icQxh
IaLB5xpQUQEPd/KtbW9TKEWG+QEHnkPCbFnL7lmMExQBcKyJqi5L1oTa9l7Sm+p1ZZF836firgEj
bRaIB3JDrWkuZbSulFTgLgbgu88LWSJUKEn0SqiiqvDhTHg5E5RXd/W8+I7QsyFhBhI6zUh8RHR6
MkOJ5brOLFrMTseCTpN5PFZN8jQj3r2NH/4zQUKfE087q3nH5NbbW+LwFqnvsp4wow7jWa8Xo8Tu
/JYCe4hr788uXxXBL27hIMJPHFXzkxfNRCsetzn6k/yKaV/mKRouW2kEJ3ZbomVxNLrWoah5QIuB
1yftVKIXxn7ZeO3LjD6sX44VjHgurzwK/AIKm2hk/7gPjtrVcE30fP2Xs1Gk3NQ6tGXWrBEgq3oq
gbFD7QNtDPYlrI4Ih/HAl/NwjTA2QCPLrf1W5/iSEzlbsW93bu1Tm1eNtF9NVV4tFrg59WjGLwPG
t5meQEu9xML/p+cr7fcZ/u4VpA+nB103yzanQ6dMjHed18verlrliwGjyT/mbTZAi0p5IP1X1set
iwnslKn9RyCS+IHPMOwmjvoG66ksrSRZutL6W1npyaE1OeqdjBP9CkHLv7zIfslQY+9rTX/ThuWz
f0z2bePf5sDw1C0WCOLTqnSTPcsJrHpE3vwRbXVvdAbv9jbeXanVOAFqgyahyCbt5HAMF6TLublu
PcEK9PuKJrCkut6prT8XlHm09dDFxp8IuYvq5cDPtHqraBRNOzEUoviWUh7fAeIDRrTnJq7nEZPQ
Hx4LwqI/7KoAVIb/zxDad4VXhzrEbVl/OaQE6MmZDZdGIHRInSJ8e1eRwdjULQATuI/c0qUzJdo3
VaXj8bOla3DaHmHt7Ax42APggkgFyB6IQK21wu5kvkdz+T3q1K29XTP9kzJ5Xg==
`protect end_protected
