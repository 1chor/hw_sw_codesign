-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
C9cdtnCP3yHsgrRinW6qPeuhZ2jWLICYsdfA7N+3glGjvD4IGvgT6zHqJ89SyIvo
a7ct2RKISk3V+jqXJ98g0gMYlSwNg7BzTIt9yyEyYhm/zQB4fuU4B8qhXh2zVYHM
1APYc9dFIxRQdQKAbOB1RoB2zPh/e2BxF3om7/DXjmo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8324)

`protect DATA_BLOCK
9XSQdUFqLwLLkz02d7P0Al116IqojKETZGBKAhPlA3afqjA7lU+h7LmH6abYIJrl
8+Bqp+vKMo9Zt5TF+J8rWY5d4hAWY01k56szxyixjxwI6TretnpHTm1yijucOxDd
/6i8dYsV7D27/Z7OsqpV8aGndKIkH/Nf+GvEuglP3VheiSmLnzxHQueNfm0iEwU/
fxpVw2Cb1k39tHXNboSg2Av22H/rBnRtu1SmrxMjaOlfh/DKk/Av8QrQimgL7yn6
IM48tqjKmIxQhiCLifOrh4SdWjIA2Nt8B0yHp0uUxM2WBYmLpQ7jbpS+NBfbQDVx
3m4dqOxiBRixc+TbfrFVqWm1LV8W9DwohVR7bJcZOKL5TaukZvZe50LDAR2de9M8
6gI0MPz4zg/HfQlNvZ45O4TXRYTiTT58IiV3X/W4mMwIHk5NRsbe/Zkc6xHONX/N
UyOiuxhRhCtUwIc2gYbJaNW+jfgYWtasEKs+2XsnSeSeitl+nPofwwmNsDmUWuk9
ydAjdnPFlLOIJcgk5kMut1YvAtg6xTjkD6bz6U72UzsBttg9MGbAtwF0it1g6RyN
xH5CpKr7Q41YIW0E2ghptfhJ1Gys+dTVsj1aRlHXsM4x7aqGxlQ7eEO+b/UGzswj
Ih6EaMVHQaoBhjHpUghpmx3iGX7qIjHKo2wheqby13lZX2LCunzvPOPVM5vhKUcc
kX3dc6ciAp2dD5oLtSD3+NRmGK/PuFj7z0oo9DJSv6+w2fbSWC74z1g6Klfr4mde
5+JsjUmzwsi54+GAi4pfMsaHVjyjOUKYtT8SBoZtKAl/l2XPuN9aBK7QXd5pYAta
eXnxpA6dZNLsZJxlEkt+rtaR1P0lkMgiEYmkbYbprq1+ULlXy2SXmVNYIqlpOiFd
jpqlZX/Af2V5+f5SIQRmZSO2uJNaC2xG3CXjSDigYCtRlN22Hec4traLuj58taTQ
+eM5itleGcmK6TmjNMePZJfTuEpFSEdRa6jKONCJQ7y6btxaxvXKxn0rKGvhxVhN
YXZrxcNGqGIEK9DufPmfwaq0ruJjF9MAdNEZrNtMk6yseJC+XXevwus9yNSvcLSW
Ur1VJuHfQIgithTP6N1Ah7MCMYWO/7t66b4OJe8jOziF8VX6rVILJ6cQCm4J6+Dz
2Ic6e4pHEDLMYnOZA5cEqUeqM55HGVx/SGofL0eubSkXpdvxWmZd8EvjwMoP+lDq
zLKJEVgAJTGagHYzSAwENHjsazznNhOCiqf7Fvsg23h9s5rMA/BACzLj3sKUeHYP
FgDlLPgrvabtkqNHTGnaCzkLgs5yE00uW+/6RkztZ2MKtbJtOdi+o6Hy3FrIs0BQ
uw6Y6M06zDistzbhL7jMrCGMKG3ayMDtx05gps1Y4cXkcffX8qERDo+tqUFVWy0x
CT+jRpmmSmYTDKXgZTRNCDm3M460mvSX5oD5FdrqGVGG+YNkIfVvhkJAkopZMTdx
ThRiS0lbgTMTRPvwnyTlrddkXZBBms3Az47Y8GnAG7LmT69D8DcYUJGLedkM2Bfw
i5juve2WOJHGmvCncoqx0wlWsZwWAhPJZspUSasBuuH1EWk2nBhJuxXvGmbrIqWZ
ixNcrgQ3R1ic3Y3m510CftVVzisAWsOGxqv+tzu+oZi+T0zIO8YSsJavBxRI60WS
TX7iqcXqrtzDjbMXTNYRzwReUw9ajJngceHUe23yN1Kc55TRhXWmJT5GbYVbgVTw
lIfHuv6YqqTCHSOzyCN4ochBfaJD9zPQlYgiTGZ4RAJ2z7yyVo1vlHaOBc76ebx9
8GvtqBWejlJjfr5bPEpbhm290XggiqnkLP0xXWJsznJKgbo6od3X4hmphxmqzhkv
g4+R7aTU0FRmv2b4mrcVd0GYkQWFK97hcB2yRdWJUb+EO+0KLdieFQfIvQ0aD/Qx
Aoo/SltEr/+CfWc29hmjzp3O8sybA/vFPSpRGqnMJo+3S16QBjHdcZa29T2EfN4M
sU5VGMx8Cji6r+xY+x+iOZnAcV3UaP2HzvPPxVRVzpn2toODH0RzHC6DNfat+h1e
5e1XQS0NHt0xjCbPHF1Y0RGQHBpdXGq00Zcq2CH+hPg820lX92OPZFzt79G8NWHk
VPJILDiSSZDyhuL7BIvVwBEQDKkqNuoftw31AQo/KITQSOL2MxBk254vlRzRLFL8
IyDWWlis1dZcGNO2Pg+RY1Zp73SfmR+HF7ojnHrMWGQ11sGD6z+xRlgvfacKwJNb
jaWuFa35399ESH1YkU9MC6i2dVpoC94EiWhKhX2ayZrHyuMbdDIyd0zIw+ZzTLwV
F4XkgjFxuDwgnlKF1BiY6hkzxBeZPXDnGjkR6LrD/TuDsgSYohjIXlhJ9163GytN
HWVRgimGHkZwGvV47i6GvI4sSJPCJiPZ6nVk9+46pd98OfBElLKOc86BHohIPf6b
KDWh6vYrlauNFOQx7wCBHcXqRIh0w+gT7fwlDWFHjBkr04l8fm+31we2UEx6exCG
r4JjuZZBHcc9RDh8ZbLv9rqti7/bMMC9L2Ag2934KzY3IOgy97LE37PKrjfjfv/K
FLf2gRfk/ov0XjIC+Mxej+Dw7CvWmfxaZ7zqd+hKCeNSwceTOvXNkRGOMWfHeed5
/U3aaQ5L/hXFba/4mher4LvrsklRw92Yg604k2i6vMmqWzMQJ+xBc5FDLWJzNaYk
DHnt7kwt2DYuaAWIdU+lUG1wJyUu/W0TXqznAG00duOgTnfr3NQA4B48YKJT6O27
z82+w9/EgxzVRLEaX6BC9hAqTg8LkYbmHhyUBLLY2JC1ZDJnoYEq4uguF3y4tLyE
oQsNJXQg7GPLKTnA88sV9/5xgQxhEUcIBx/bmcwD1VLX/yD/opaf8ICJPndCmJqd
CV6g2eOo4oN4AYT4ryX5+oauLcoctg39gSTIq0ciHHi1QKbDLCC4z+VB5BLkuVmz
VBMYU1Ohrn8D2UbsDLQd028b/v4kqNV62dBkzUItpO/tSIuyT3m7Ndng4XrIiBYc
5e353w5Ms1xAi5KDejZLV8lq6nnrQQsg2B1EJtDawAJkii89VNDXhB1xS1J3XuUD
niYmrwDxxItlPHl4UpINEopoC/E/KnFj/NQ4YAPsTTEk0nrL0TPAIIoR6/ue3TCS
PaVvXhLULnwVfHgmRLwh/Q16qkX4GEPjnZeeR4KuyAp7iHC7GLxs4NED8DHOsd1h
bmKovuYFvXpYb2uXUILIEE7H7Ordjcr2D98H77L3CFkNmehJaLkNU79fACf86n7K
Oy1ks/AcpOQtERZe2jjnkmKlcQjgqTTbWhbho6U9QZuladr8YEe8Qqy6iNO/NKKA
20hhTmopgJH+nq4H3m+aXD0puILLkbHyzv1vuHPjCl8XfDmEURy7X4YlPKckMthi
5ROfPDo4d+fEE+5ahfjqGbEzMAKz0SmFX8u4MqJGQxND3GUpMJ+C8o/HWOO6sAOX
b3f/KyPlyQ4MWJ75XqH8pkZeIj5moIeluqhqL+tTAaAGh/1KYQKHt/JEVWGrhjPm
k/f7j+EtHj4Mzx7Ca5V4ao2NsGOqqO8eBwPtUOFs1rGTdXnFgW4hNw5e4T525xkG
vOTYrHMMVAU2WOLi0KeZbvGW6tnz8A7nffkwqKVA9wdUTF8F9rtkbXPIVj2whV0f
97x+3mKxgQxpj6bM+CK0YkuvCym/lBTlzl0QFEX6qLccJogPyPopqnHe+0zVNNLm
JNHJu6jT7gGw6yKUq4Cy1tYDQXFMoYmuekrjQ8zX80gxrV5G9IZ7Zmmzg5TcD2Jf
AztWvJLcMMESliiaVzXQz+CviJyNhM0BpUWZpNTKtVf2sNzxPe19zS5eDVy+in6t
CpLR6rIi+nCdbHkpkGLfStz/kOo8vIpTPkYksYtWr9D/4n/045lxn436kH5PhEA4
rqtI8yHvKdba0nPbsYaL+kIIF5uvhU/q94v18IqEWQVr+4TOHFjfFrL8NBEnArpF
MdVmWnY6jsrEgPcVBHrv+94jDv57F3F6T7u3VKn+KPs9FpR6uGanffB+P2NLXxmr
bzkP46Rd8nE1vKulq7Bbu0JKM4kDRO3veaQJlQH0OqrBFos3B2pPSAqqee4rJKe7
xLXavvf7tGLI5u/YocBfYBAtdRmtsMl6BJoNoGLtFGTBgLislcI902w4OZg8jd6d
Q1JINwt6SIgCn7rVKnTmIo4kepmFKBoPBVdAQkWzesdt6bns1D68eeHu/1w8haYF
BamFFZ2JEpWURfBcuBXD3/5uMxegqXhHesdxwt6vqsHVgvONIWeZRxo7pAPPfP84
qhVXF+tAhGfv7HW6DEF/rkQVCI/2BRPUzHCX5fYtft6TaTZx2w4q3e3tRzR/Gbgu
XGd21wNwI17DZtU1K7a28K4qva3GY8BB5XyEFrxKbDpLJMdot8K7GtjeiowyB41U
/fGTTfj5bT9sNybm99cSNVZIicb1Dt9crBuehDu3BAVYuFpAy+noH9nAD6UsGUGt
Fu521HmjO0NCgM5/c7K2ve10iqHdpyGvSjIYLnutFBiExW4pZ1tPVaSaNjaYKptT
AIo9Hm/mNI0aSv5FtYqT0P5Kvwud1QQAlUBQciB4UzdbIurCTggqfGi8WpYGkw6U
vYOopnW3DaNFqcuQuiSy9J3JPLzMcND3MJLyH7RdRAqFZxj2NhW2qUTW5N4GQy4V
LjzJFEX8J/GafOEvIzBcNh7CPlIIq4bJdoT7Z/tSRVRgoAMkrVmqiVM7ajCXeFG8
HbOfHAnDJ4iKF1iQpfEB4iI9KtT4J/Jj3WmSq2Vbp8m31Lc5a0gla445f5QHtit0
frXdEFn/p6A6Y/ulDcIg80DIiAMGLfz8C9r+BgBi+gWDU9d6grt4Gt5Fp18mAyHW
FAPVb3rPJEeYubnlDo0ILphUghauRuZHLupLJXC0GqK082Hq20PvCc9GM+86asq/
pCutpusV3KfWMujth3S0u0dp8RVXoHvmo4Io4WByB9AkRhbeDbSieC33oVJJq5BA
Yjr3L2n9r5rjWqMqYAbHYhznLSC0oSP/gK+T21scCw7qT/Po00FnxwEwp5qZC7lu
M8Yj8I0j9KiPtFpnW14ayBZ8G+pBN0neQj0FjczPmz46QMjyizOWIq6/docvwvbG
5cTSvnU0EL31lNUFDZONuOyCj2rZAjSaRCY/E1S5HrR+CBfh3RrQGEyXxzRhIpr0
JU7aVrSd7WcLItAeG03Mt44H+u2IkpcU6/OyIkcPiKE/QbMeQusvXUKUstgI0p5G
bnIxEettZUXqc0w6Run72HWKMW4G0pksS7w4AMXp70vE9RIat8T4Dcm7VYZBMUdh
zVqabHSRuyvj0HDc9vB9VNTJEpfay9hdlrk9aMFzFAQ+mJzDwZo/z0945rvdFRbS
qy+NUiQGzSdinbUJPCQ36Msg24ARxZA9sOWIrWaJDxTc8IpjYWWEVZJaPVP6fpya
5ecZbT7ZAiqSpnd3enjZ33qg2XmYwz83RZkdjH1KNRuF8gGjKvrwJlgbOFOl2LkV
Kx3/C3mXYvcQvz06IRnB5JgEmkCZAYjcBp8NwPbLLdipnpxQcUW77GVq/wSSXihL
GOodCaKg9DhHY7CurqzaC4fp6oj6lAjoxr4unROOGdM8dfpvJ1/O9hVDgus2ik9e
B/uRGUhPCjRH6YFj0u2cRFn8VMS7NAIp4c5z2EWS9i0dNZQB3IP2lB/iVpKYA0fe
4+aPzL9fjAZyJ3vZ/USqMrjT/c6MmN+wcz+yP2weGw5MHATa4MHX5/QjFa5OSzbu
+WpmgSWfsSWfBjrUAv2oSBHnR/rOVdoRUvywZh59QgeH1+sk7+IQbWPHfBBcp85x
Z4A79vuSsVS1ekiCYbpey8kGFRRUYbPdHzqe3/jnPaZXhjr+a3vkRcTZgfY8OqE5
p2s6uCEBP68Loyz85oazTA5B2gX1JoP2E+tsqmjyDAM15VdoTLtzCiBtVKXsvqoM
6/xOAMiHn/5vf6R3Eo8Z2vAgAmynVwZ9JoGwLOVrM/kROejeHV5Hqth2I5dSIRQZ
t/D74vBkCi3m8AeGlLXeP6+3O6U3XhH63hpQMwgl5rTGUpNqDJbQ7i18DZoxNAUp
+2ypzvZB6vAk3cLrfeebVun8F8ziMTbjoZQLY4jIBbn9VEwYKukzNcet7pH/YqO9
Bm1nVwFRHJBuqSgBwpYN9LvkXDII3y3Q/ZAYnEdm4oJgCCS/x6Il+sn0mGe6hWH5
IudXkXhyUYJBSTSELOwaodqGjKQJlnFzbMGsaI958o4X6Opzbl35tY5QfpMXU2yI
7K2ltdc2F8D7f8gNkS3dhziNsSAhzwQWOvuZ/ZDg3AF5h9eBFgJflhjEHyOsrEwk
tvI8XJ9F42IjginHGqBGMg6MteGptjcE6Q4FtwHXHuyjTbS3M10OrLNXAmbwz9is
IVkLKeVEBUUYWGPVp3Wj6GN7WPqdkMCQxpQdRyi4n4OssH5LJzjJCZc82iVKr36k
pShsl0jbS6KcSVlYyJT5O7039pbJQQ+Qzgr/BRRsSnXWOrCAsyUIpaitnO2J/3/V
WGVIFPl7mIZANGvHyWxXEdt51BJ9nC1szyvj+5rsNSWkmxTQBwAYuITD8Jlf6GBo
Re9C04nY9QZbDly4vb+QqcOM5/o26IlgyaBxbpJebBQ+4hoj8huDDg9qEMbiGP40
veSOIgPTwjmUSw8x+hJWon68uryTI3H6iVaupno/B5wlYjhBsJ1WRtVoIO+AbDku
h3v+vtpBNjYTOhlw6dLsspg85Dr6Ag4r6BtUFaMsAObWuMF5tPM1ynB4QCWkAf3o
2Dxv9jS76gH/+iw1oDR+s95t3qW4aJjSOq6Y4JTBN7FlFJFzhYtE5kc9MDw9SPu2
INSBFghV64KMx9PV2Cu5Dn5LSallexdIYLyFPUQv8tZreE2U28HEK1hOhM9X/fiS
Kdw7n1oCN4TXMR4te8QitmA39Sc5ZphtnlkLuC5mdD/QDejoSIdbwVXVIbg66hYx
twbBm6Ni8FB1cAaKAXurd57MBDEbyi8thIQM2G3oWdAfrPDFlNo47T0LlOehUOHY
ZoyJGMvidM/f7HpJhEhPZueaEcN8zhVxJa0b210ZBfuzVTdL8J4JwDaA054Cnzua
DK2TX7AdOWYJD5EhnXM8o3N2ekFerF+c3ChSX/hQX20wBQTPo7hi7yvuUXlrE6Mh
RZVh0r9EDnSmkye21t7WX+sCdYNA7mNeH5QRUQuYDQtrOP/TmjAXywN2tu+8QgMY
D2rVvbuVzn4SRKe1eExbrgxgKiq7CYs39E41VDuneNG9Dj3qhZZUxnLovrO3t2U9
UeHGc3Dyvm1HuOZuM/9aPG9Map4EFEVDNyYlYr2NM4Avpx83hjarv60ugL5jByWv
KlZwdhq3cDvYb7WXCJMtprBOheB7uJFusgR/Z71be7leBX8uud6MC7TkDOIBOxcz
S47Wz3AaC7CeaS/2VYkZYLXSnH0R+JfDJPB7rbdZFl4QinUuAZC4foWubt61UkOh
dIZ50DMYlwaaIdYEeELqPs0+Tx31pr9aQ/0SfD3dYsCx6P1A5snkZ74kZGZFQAQl
HqYBjjLspT7O+zbLb1FmLBJ/hfxydtNDveUB/WFzPveeBBQT5aT1gdAT6TE6GWmi
0zLoUvUaQa+boyncQHkCazehyyZk2xEfMBlFSqBlcRgq/iKM/hhJEEjAomUB9GCf
65oBTmJ+UUTWTxi4FV1c8cmdZLf5GyXrYca1sGGM8kdOU/LjwaEUtAOnrxNeDT0u
IgEmsoXx0l842eE1konWwqDt9qQkzOtW4oAc97BRCQHOXD8MndNfX0OzWlXxhY2Z
BnT77RjDwGU9ALENiCCpeVsyu3R3eqXREbr+GBHA/IqCsWjGlHj9qUgflKGowwv9
Qp2nJ4xPwSgSWtecSdui0oIUqXAFWEl6OyGi13FVygOdei3HFS6UBp0+tgTJiVX4
3+f4GTnhOJzRN5ApT1h9QhlGFBdwBNm34cFz0XoBkA3+hSK/S76xDKmClbyBbP5J
YYihJlS+A6nbM6Px95HyFP0LCbIXoRoalm9yCydSeW1wFqU/KdUbzpHcI6qCH3Tv
bMfyW2XUMeKisuSnDj4BXsW0/cNwybcgJFQQa+1j448+WTd+yYGHau+dTrlseUrK
LhHV/lKUjtU0djUW6pNyZJQOAlrltRuNwhW9SyDFAwlN80ACkNDWPbJIA5KOfXll
ZgtMOtCIpjVMNoU/RdL7jkYruBvYwFCORqOodmByoR8S229s6ZT1vO0j/97VIIcG
cGOHgbhfyTYgHkMwUuqmDWWznk32pZ4WBnmyhDABoNWyS68ZjEHcOHlQOp6yqsPZ
pNv6aL2XX4cKayK0wWsUWo1KeRlfAnnlRX2bEDflZP3ZqraUqqQaZA8HzmtLI3gQ
05n80W7+NTOhyvlFmzqJxZPQGjcpxS8QOBjoLkxX9TPV8sA58P3m/PODyifji9as
8y2Pb62/jDLfduh43FaqSsRLZbhj86EGMEtl/3vx30B0EfV9ZgUQfPwjYNOHOpQV
ID9FhfPLNsR64mP+qRGutK2/J/FjnAoOlD/cH6dni6jY2jvMaa9hBs/NkVwJXBlk
WVC6cOp7W1kio13S4+k5Upy5liXIwHRFtR920XC3S+h1zlSeSqBePRB54Co4dtvy
5bDbhGj6q2yAnKXoU8YrU78E3+Xj7ogFn9rGWe2JrBE+eAQ0A5lA6kb779mzpllo
jsJdUBPiUm/DjrwxpkViRKnOVN5OUReuUw7ziNKokSaxfr8hji1N1dIPJPx0rywU
WY/5JoWMmJucjv9YFoghO+74JvYYn425TrSjfzlJYwyzIWB/cT+ZJgsQAFMRgoTX
o2UESmsGYBQeKxoQ9YxtZ+YY0tLCvL6tWvYoTYDlFM+ahm+T5qVRVeHSQkBoAmmy
Qhxyx+30Qwh6k0LX9bsIFDxO7rOzKHMk6NlRRdZnpHa83pNPwCtFJqwYqN/XPhzH
3GzdiqD76Z0DTZM00GhDMdppwv0jHVTczv2YueN26a9+N4HUTp514Cg5GLM87pf3
/Nu17JIeX4XEsBarf86Bf6WnkyTJAml+vD9Srj3rMMZ9SwioWJUW9tLNAU3aEELJ
AU1pWIsnhVQo/6UkZ8gPwi7/UG3Nnyq3nYwMvmH9OpAJlTTk5hMO7im7jIwEvQtf
uk4xC+No9wlw9RCu5M5zCnlLVwKjXRm4PcQF5zgiw0ll/QLIk+naNDtEKijsF7IC
fYSuuWKtyxmG8IsZTTMkN/fpGm5jCPQQaUDqjSXhTEK7czPpsjFEm6TB+sLj2KIz
gUm0HbHYjKsUMJpzIXzLleNRnljnyproSo0xVDw5M9nlG0d2cbSOaRbOXgHjAL0Y
Pu4hAVOPwT0uE6hJIh3X/blGWQmllYeleCPxMKaAODsIqVCArzHkQrlnZpO2arMZ
NBn2pFHRseQmW0ey8lRzUiUdheTnGGfXFhaEZNlesOd2kip3pRBeaRZkDwPznman
5NEDfK+fVPkjJ4fdO9iWPK3J7pWUesxnm4oXL5bQ+8QDUtl3E6yp+q9u+hdsRQd2
kIrt66cuZ0ZJ1HApSQafchR3aCWX1jPxFZ4r5XuppSfkVYSN5bLC8QCPKgWW/Oe7
Hr/jSFfxS9UF8vWLETGcTIdWIw0bt7uq/VO/SJFl/X7sf5yWRKoV2sjsztwAKmuW
I+awVYaM72KRXtGOhNf1kJ7UwDdiDBCkz6IV/99CiYj5ROuFwCi1Hlb0XFkyDTjP
p1r1qEsVFLlbZ4Aj+Gf4VIHkW7eu3ITA3bql6ZLk/zYKYeob2bZY+7wSWn1ZeKdo
ks10/bB2wSdIahkWc4FkWI/hEwSoUMTcqlLYI3JI8kf986Ok7OuTUNP6YflydCoT
THJT+htmrJZ4nLq3jDQyW8d6Q/QP+3Fvq4YFJciRiFb3VlZPB5pZukRhPSmKSIW4
LOIAlJatBxvMFm9481VF4sFovvo/9Lo3tRyy0U88L5CbuOnjPoG8gV0mCnkx1RO3
Yz73yknyZ+LQLOhaRwz5xotdCZvMEY622jUZo9P3AKCvOLCYoH/OH2nwWPrhIojE
vSAl5wbd0Z4pV/TnnvkTe7z1um6x5oMeKmV56hzfWm4DP4rzoxWwiyO5njQni0/4
bqJ0lDcYMq+5J+7XUweT/hDoYTcXcZWFFLE64Dx18Q0QkM1gLWTkrX8NSTsaRbps
ehQTiEH7kgQP1euqB8lxkuj/BEaJgHHVnsf+GO5DMAoqJmlpHs3OY93X24yiTHYX
YpAcSzHt9Dxe2/XADXNoP2h5mss2iG4v7yi9c2/p+gDd4yYhcWRtASnF8JxMFuv4
971mC1ImUag+Y5RI/7h1ElIWqMAiukej18mWQgTijTaTYhaw9YuadBxQ/IcGhJ9o
H44M3Cq+8s2STQM9jYRQiiP+8oDtRZaaQD+VjzQ4Yb2YqqhcQiMKM4kamyqAhEYh
3o3j+VDbq8TXh+QSuD5AJ48wOHPr7FysqhLa4ghHRAFj0dKqVje1NAcF5S9DhxqL
ivxRLZpjVUZ6m+037H/TSArwZ6mTjOF6eJXhLq75cgOL9TOti+7fgrEXscNNx5I2
64gzd0bRwBE9FN4UgUEb0kkgCShSHBRNyFODUt179lKrfrZ4z69YAmECmVhgczqy
NfLHZrwzXpV+PASbDUCo3mtrBRthpkT3eRoLZKzyfJyXN4xQU0QO9EedSVvH5AzP
oxUvk5E6xQjynOmHXSTo+Fe+GJMo/YIGQnhebxwE/iCgI2yPJE+Rm2kmEPWQArQn
uaVx5OM2vJHSk40J7tYsqTBAiHGFGvWkNgH9hqYVZ142BadjCDb6yDe0wX/XirJj
Uecz+aWu7wQHpmOVoQWuwo8W2DAGEeczR4uA/oi/z9qG390y1S6X1MybVgKb2G1t
g1AZRmROI4x9+B5rEUbmt89icHj2j8Iga3hF5vFXPs+Tr0y4o+wmtJigPWzXbZ23
6MT9PTYwhvciVXHMZ3x2LSmlbVUKyOvYcqxCYg3PPVO75csdavFX7J+ooqGiDAvS
hgY81lW/Crpl5CSA0sbnnWF2G0vVs/svvEDYaRI1qFXe7pBr2HJw7Le5GZtiO9ud
KrxO9ViC2hmGmZZmTXsUtmhGaCsJclfgrleUUbRRDmj10VqLckrhiugk6IpDFr98
`protect END_PROTECTED