-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
pZ/a6y2zMk+zJ2SWTKZZblFLA5UJTBjLZIR5l8yCt8AhlDK/pAJLEUVndbzEdNCM
Gl7pUNr1wrW3xqfo0zAUed8SEpInH+Wdl21XaKV8prnwBwCr/E/NH5h+6LMhPW47
q3E/rx87CsWLjDtlK98O9HiTcXFtkxKF6xNcPAzeY00=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13001)

`protect DATA_BLOCK
zPT7PXGUVMrY60D+h1I/TI+sStUVv05zkmVDBqXw/SKmDRjvd/K48VdhTl5QTFUo
VQXXUQPZGEKOO6xTB8vSGeCyzAq1qoD9VahruW0A13e/DKCKq9Ng3uPST/Vy6rzJ
YDtPCFwRqaO4XC4Kp9N8iQnsbex0o2MV0eIbThXc7hNbbztvptLWxMSRjGB+y6wB
5tRu5rHOB8NKWy8HDz4Cy+Cwada5OWP6PXVKd7z4rQPbRGGxUPyQbMkFZGdG0GOJ
gJTHwsFZJyhZeRz7w9j1PknYPh3gjNpedQGtSitlYbZhnVcf20P+hvS5eNbSslnp
IVOFw2FfqoEyP/eBtd43GhpJ8l9K2fDajM545s2jzKQpSYAuhBUEo0uwqK7d9cZZ
sbFLI+f8abEdJz/aHEY+FuHEYoq35LFJ04czD9NnzsDISU48LEAEMFwUb4pGdERe
WerO63lKFKeg6sYeUVyYIl7nR6aovXoE18hM4eIvgv+B0f/8OJVM0fO3S+9/CEpA
YkoIS95Y3V3ALYosZIhmL4lGcX5bOMFQ1dBtXqSDkujXOwLvABaCTfuKL6HjGrFr
P3r4dqQry7mEcpSY5fRI/BJtFjpA5uJXl1zTi699z7CaOCedhjejnJz1RwZnFFNw
VFpTyN6NFx5LAK2eSgS6sSQyy2jCE04WjFigXVbsYw2Vi9qWGIzRr3cpMkNrt00k
ZUDVLjNZN35DhaA13Egqdfy6kRqCm16mc15PArDCpChpx8ixzRKpENQc5ZS5AA8s
t5Sx2+yUlKfS4tlE25Yo+vbchMQPwoIKvcZ2XULbwqVObphxM3sgXmB7C1XAdlD+
Gr8YcziA32YUJmMvLUcEp/kuCrnBrMt1kJo3bZ5dBNx+liU0PMFWWCHOquWRB7/X
kCu+3Ona4wQqlHfIHV5SHA5zKlqdBO7vjjKKGdWq5PVU4fZoaqH0wYeZVxsVA4HI
+qIwPXZ57AK9a8XiQmZx10I6NV5jtLzt+CDvberNeghsB657UJBHO/PwbMmrr7YY
kJc51WDNy4UrPzq58QACqBntFGOfaydhalUznF/xQD14QI41czrsgM7245s0WTH4
kI3F6hGri+HWuK7yaJM0+D52meXlVd3u+JFMA7JqZhZSuiH8RPTTY20FR88/vnF1
Tehes8rCq9tguvHJdB9cM6KS3LUkB5RuMlGcRt1AndQd0GjVjq1eLGlwvjmn3LcZ
+ihu0zYngxUZpK1JJRKRU3ZSFxJTUcEH3fHdprD9UeKCFKwvMZL55+pAAiJ5VhOm
04JrW8k1TSsz/2FzwSQA8csMTIIysIX8A8vkR+xNcmIFf07e18W7OTc1uP7vnBYZ
3XrniZiIEDdcrAhruCaftgNMz75QJy9qyYWTQzXe08Iw/yix+zm5Nq6+FZuESMYX
mfMpw5Q/kof0qofFnK3XTlbLFOtH5SWA5j1PXy83cJ2QZrK8lyRPYPe853DiiLsO
P+EoIs36s//TMDpPhtUn7QcEe0AjO0nkgFYObmPrLPgTrcO7qD6e4vxJ1lv/1Lja
yUNzl+iyEfVmIkf+pyUoLqMnJtyApwdzakefnPc9AoWFDibkgMz9P72Ro8fnlKi7
tszta9gbpwxyGbPdbRFB4/SJyR9ZSn38auHIu7AWPnWXVsMMKz4EIQrTptmSiJTR
3qxOuEJRZZZvMi/6DzAa+pUF91ftlCWhOOlCOW/aVdHPa4gQ5MWfnhdRdr8QjVVg
KCUmKUnwkCAybFNc/pLaLcu6ioy+37qRQI22Xydo1+jPPfSdG0WVj40Rn0hAOl4B
FIuL0Gw9xIpzdYXCNhTtRxfgAIiaVOoye9/XBlRKGMQaeOlm2FKoeptTXnrkrzt7
jP9siGwrKYnu/9GMkThkJ0hJGQRw1IgcsU+TO1EdmsI/ql0OvyK1IsNIbTKwnMov
marsYVvXBIU23OcF8Oa6/Ndo3j42qiY1r9DGAA5s64QzKjS08DQFRi/Lk1Qm0Wmr
AfNX5iD0DjaoBHUDYTcQMWLA6/y8jmDCpAurPa1/GTJi6CXnpcPBnhLHXohnYAZF
FFyiQmjkqCTMTJMnxoXXtKDhxpFRbw53tXzX6deWJ0+HSCRP6gS4E+3DNusWEThX
MJ3rCvDCwk0vRIDcQZmx485NWqutd89RSSfgJVIyM67CZe6OlmfoCNZAjYoB4qeV
YtzvmXPftgSh+/hI+AZu5e22s2Y73AU3BCie6diP8biXhZNAcPRjUcMjsZNw5y1k
jtJ9RBNwr18qEWmRpYTKSd8db/90nByIXW6kOnMXq7Z5jnxP40vslhh1DycKOTj6
ETKk1XZYLBF3Zy3u9cUCUZP3wPEmLLcbGCVfvSu4Vd7aXLO2uskW8u4KSU0LggkD
5DvqGN/86768LdEqVMXUm3gcRnmYPowRqzSqyYJoSHTJsrnMx1LJym15ePctccTz
Y118DeHBWbMNy6ZfaOApkDKrkDf4RrdhC0T2zpPXQ8L7Y9WdarBySAVij6di7BoF
8Chb/JCd3Fnpqx7IEOeNAUs75knzb6UdoRPwPelU3NOIyT708PtdHmkuO15JnGwF
HAFzAaZ9fo6xl7TxummqKTV2LB+RYid/1TsnKlpKlXmB0WGZHzi9CBzGe8vcO8fY
fiXvUFczqsgyWZ1XLdye8KM35y59DeaPU7jiaauQuL+MhgbKTFIAbNeJxyOlm1Nn
7f+dhk4j46iB+tldLXMKfKwQ5uN5YBweaFt5Eh7axQ+rGSjkX3S/31hOfehXSbxD
yePXG3+S3Sjh6eG2vqgr+uce5caU+4cx4+tpcUjR53jseg5W1LHT8evE3Ah6lBTU
MbpuxD2muxRqxgg5a3Cr8aY3aqcMGe3oPntqTS5y7IFZn4qearAjjGn4DJzaf6ev
vIgBKc0PUAFPJeP0Ymsu81mp4HVe55sXVlKy3y6MWSVc1zTSUtr5d+kKV+/h+onp
cZvmfq5yHF92qVT3RqmTx4UMefHe9atritphEoy8z/UjApAch4X9C0UJ8L4T0lXk
1lJ4jG6wnNLRj0fZNOwVlcv19v7/15aiSCmPAlmaLi+FL9iepqKn6hWiMyPtUfMk
lCSHD1XgqBUk4lZH1sE0wAOFdOh8r3cGB9e9SDUS1u9IqVjunnnAOsqr7+BaxIYM
sOS7gPKj/ZJ3i4HqtkYLh4DntNkb7nq1SQcR4fvaV2rPFhrVZSthvk8Ogi5J6fdF
ghReWStEJxhbqW3GSHlQTBzppal0Ljv/IXYRdqV6Y7eh18LLvohUJW2nn+glseTO
ARbz3e+q9ZhAt977HX/x64mtm4UobgMsMRKJERDpoc/DnggE+Nph7AhPeWLqTIfR
gGgr4TksT+58lAf2tCzbwYprrOj6yfiWk4Pn1d7fIgagowrvq2dbIwKn6H3J4xuK
L5qShm0IIw43xB/9mEnSrxkzAzqvL12kiUfvWmqZ/6+HByuuFsnZODT2T0Y69pBz
JL3CI01Ap2BJSgR+dPTTrKsa8lbBlu8a0Syd+VGanklqadcPZdgnX7FF1w5yHryO
X35KLzSq+9sq8cG7hZkEzeQeuMFuBl9gskvwrYO3XDbXh/5dogb9nMyFxq1/7/wz
EgT6KtzjhKzUlF7IyMl5kCplZoj1amqYDY8PobiuYY8f8qyu0zscbdf8/ZQTghU9
CIIKkDs35WqE7VvlFdzLn19LPuig05IdHXbv+tsTAQ4qq4Cit7wnLU5ZwoHUQOWv
phcGK62x2GpfDNs8tQdagxtMGfmftTJ+D3Aws0blNF73qBEMHd/HX87R9JC91hVC
6KkPRnMNPii6UiVc7GKCmRAEXDUMvU4j5t+/jJmp6b/+cCSw4IT64bnOhEnu7354
6q0s7tZsaqFO/0MbkHVrBT6/TyZWHjwScFUwzhUNFrI5xS6QcoTru6dW5Xi+QvD7
ZhCszzgv45dWx+4dhGiTSu2LTe70sm4RWOTGvjeZErI7aBxXMLQyimhhGBN4GueA
YDuNkxvB4mQm86iTv8zqr8VzgRCXw4a4w3BzGma4bJMC4bUWLajgLHPTEJWkaTbr
3qAB7cY5A4yym2AZWmDd4bIhY8Y1mWoYtNAy6FLIvx5z26vp4KegU84I5JhpSLyw
TJl2htMbX3KACH3zaRTsvN9H9rbRv40ZW2GvcO+T4QxzRxxATsT2v2yFTxm42jhX
LwzZ5J0+kxO0VV6dhOxiP1W/VKAnm9Pmo00IfzQJVL1fwGoKXB5pD1k5RHkBUAWm
73H8M/zbyoQCYnPMa+2aN0MsiWdNVLdPKODi99EHyJTstHiNa829oI8xZFEx0sKC
VewtaGkqD4qnqcBxQVvR4biEE6wskHlwfz4D3DUBUUGuCgucvDYl5eM1UHaI1M0S
RwIM79yYQNpiuMfH133Wo3/UT1pARqS0ROC8a3Pqf3MoHtO75yQiNCiO1KlSLRs8
TpUliXeid8mRuyb9ntiSCdCRi09ljNZ1ExR9DpdmguncGHSSZ9HrS5YR2J8il3aw
sTOiAjApeT4NgGVolpRmTDYw7X96x2K3FDbqdPZu+JyxqKIoZXqHPTMIbWE6kNjN
RYTOgbvUW8lpY5kRUKy/N/G1H1VXf1H8XwjoeU1h/k8KktApboSJty9vee3vlek9
aFEdkWIgWrVnee7TUTHuAYKxUWx/exYrWvBNx95MffEc41aNi4PCEsCYCkJLaOe4
O1yBYGrPEzf1709+wM1lIWA9Qd1lYEm6RHRxadPxY+FMGjMJHEVrZaNo6ofFX4E1
Aq9DESc0or+ARI9yNFdXyv3s4n0ynudC6t1NQLsCTeD38u+QZAlX8uljRL04nB/m
XZyomlUlbhzK1L6uNbuqZeAEJuamOqIt9LHp/eH3mGTBnzNKHDaAuydyD22XrUew
/ciDw+Zg+QQdi8t5b6oN3Y7jLQ/cFE7GI4fgoN6PBHqJ/YPb1U4Y4UnAZRYIaJLL
wyEzwQYRtw3X+0/Tw+xVXOCKIrjaM6QU5exzmOQkRl+cKl64/EC8l1yYU6783Xl5
Ydn2l+w+SwVb+yWTicREaICHr/OqrHz0tXu5HayKA35WFa4/L/js7F2Nj8YO6KSC
hCdycOnuUkL6ACizk1+699H72XvazQF9kHQw24nwsOCrlfgySHL1nHK9G+1wZEG+
7wuvfCrfrV5K6OkJghfYrLMS7IgwuuiZV8xxtFT5UH8/tw0R2cMFKj18ljOBHJ49
Yjwl85SYtC+toVeFys1pvFdrsERT2LQRZEKyZIfo+b5Ef+6xT53PQL8ofvxViJWi
xT4RfTzK7nmpXTZpZor6eH5MpkczyMgTlj8S9xxthdL0YF0Jf0wQfnWUeCj8iJuh
j6+aPBiqY71XvTK5LtyhYmTmgihdn2d+a4uGAskQ7YzzPNqrq5MrGfudc8hpusHd
ElojQYXQ9PXBt2ZvcLadSkxxHBRPjzRBJvaMR7wbVxvzKrOz0aNAcRvzHzmOeGfl
chFWMOmObc9UfFcOa0ylRIn5moyTjnuuTS6YDiGbjzwWt2lDAmeS3pyjV/md/qaK
vB0fmZq+xSNU5VsJOG4wt/nUSwkMmohhpbyDO1GHiL/QOfYAsluBqiGCWOaexq1t
q3vxch4IsWg2HUww+knnc8x4BejmUU+vxstvxEzWTsbceWP7nhf+XrL5lO1U6Duw
6zerNhQR6YCivJFgjSNFqVXHdMHEnXR3MaF9zUB4PYl/ZHTpQUkkYGe0WTOFI7xU
zqsgpewLWp0VfOQjE/dbIsD4Rh7puwaCfeQ5u3RCQ1UB1drziRU7U+aG4qJmBMpK
SOkyfbM3ntHiz0D1I5gyU3ktA2rENnFsSVcDmUulQJRzMmg3wCx3ztSug4ADq0JX
NvJvWE57ywfec2yH+e79227z1dn69hewws433LOAJOfLOlMHqPM7p1BMShRWC9So
7EPW0XMrYuNSfZtKHwM6o8tu0pOrq3Da8JKXJR7I7vp5Q/mPWBAGFXPRCA7n+gjL
1kwhZtu3ZwdYWPy8Js0tI91i/EsE/F79X3wmD206oORll3HjAyoraK/4UGi3/NaW
w3jFFHN/rI1mTHD9Xxl/pzGGLQIOGjhaY+7EO8odAz90jb3dSaCnnX2YiKTqVEQZ
qUYkn95qwZVOVfhu3N94bTE4XfFVSaMD2NHukH5+uXQEfcX7egJGivsVApE36HXf
gdL9fK9ZuYgDbNer+HECt1pgFtx6D31vKDg1O0/ZECurxXBbbzLmRj3TNlYPJ1j9
6BnxTTZ0cLRRI4qROUXKIMOtk3X9T97jIgmuhKCn7spIsjvqL/CB6q1+DxWU49JT
Z2zObPC9S/GJ1kv980NJSKQtD7rSeMPq5Jl4mDN2RPQiImfjYD8YjHGbfIetKgqh
V0Z03vvGUP2tm8DDcXpHtlk9YXL44YQNraro8hAh2xkt8c9MsORMw0tIRWOLHvcl
ct63P2RKXLvIKVSSoDNP1dkK0nowQK0M/i3opPVY6JyO8DV/zp3vseOI9Knj8My7
DdceyZG3U5MKB+B22FzmkB0cdqbdp5BW5ivg2z6ZezKnhJduxPPB3bJ7xlmGC3JH
92SHreBXr0k5XlWMjuTwadtPzb1HVsfkpeFNhfu/2dTVgqUypfdEj6Cd8Cln371c
MsmG1I+4hpg1X2/iwclQFWev9T0LWvmlD/dy8SQJTx/vf5uKFiBdruQxVP327WOA
hs/s6TRJJvyMu5kvEg1HBewQZnOFE6qH/nlRLLP19CgJA35t+vKxpU8qkXuEO2Dt
ouF84KmeDl+P7+sM/L/N1F0neCgIN78yIzGsv9DH6aQj/n++xhJJ0VvFF128/eBP
c/DQRZ4jj8lCsL5vbt2GcJ3pP8zE0ffm6GbgM6OqPfTqS6ucZ0mTFft1/ZK/7Cmw
Be4DsaZ8M+QkfBu1SAcfRF+6Tpj3Ei6m0QbDRYCHc2AjWTAIBtk4DM+LRsGfVSXP
ev+ZrG/RkF3UqdvRxfZSqPI0kMZX0MWZrYXyVBi1CNWQLSH49pI5quS19BHEzmlw
EcT2JYI4aGfdC54qmKCLdXUN9MEiv4OyPdqz368i25zMmJ3mXOn0Wip4znpgfYmh
k1zdeMApg987vlZC7wuiZUxQOGbLsiW7GrmrNTB9xZ6yFOJ450LvsrDcRuqC0iKQ
Av/HD+S4Y4XFQl+Bu5ka7sxjPy1fm1yJFSC6rpn71CuK1wlnVt1yJDfc9Y/9MUxO
Id9U/V+aWBg8LjdeEz1+DnJwkVkrKTOSfEUTakcY47Iu9egm7deqECmB7oM7arFy
WIAu9cqvqJKOqLQ9iDlYkMKetjqgNQPFRZVH1Napu9/n3ljSMiTj4JTQp6QqkxB+
KP3CG/xvmBfu/erQPumB+S/Ft4tWd9SnYBNmxfmO9IrAJ+mgiIATl5VrA/lPz5my
B26ZFqIOoXBoRsf4ptRyJplSdOnM2qGVk43jC0XAEDPuLe2+iAatviSh6jHPKAAZ
0BrHi+8scuzq0GDlu58SmJeD0/G7uLxheKq1DaF3flh1jnNHAH8aaCIoN/HKB88H
vLNE8rGXk1tCYc/XNFC+CaqvBfWORjP+uQBcFVCFTJMH5IROx7YArPOolYE2oSxz
zCqO/SGUZOeiEsuvdw1QkTgxQMJW7CrnaCuKJMNpGnUH+FMH3KZEordoGl//6m+W
QAeJxK1MOwMyUcHydf0VTFT706LZWtcnqbhDeuFJe6th3nT5XHOVmG/NxFdjqiWW
ilyNrvxXji5q5WTPn+hu1TFDpFOtnwLzzf+aCEpWzOk1vb1SgC6FCGs2IjJqJK1c
e5EbexB4qrw+u3LgrSKaBkg3Q0Ai42TnMuN8O0VVfq+WpCT67WMS9bOUwypDzRb1
1sBQzviGaITDaR9pUe+KOWMv3+8R7/Vs0OIAB8h30QvBpslRl0z4vDqbxAMb/djj
gKApxLgSwQG0AffF5230j6G9lo5h7EH/vTvUGzTlGQn1vix709hBCibJV9CiXc7m
4gUx9WRfm4tCDHBFWqpgC77rd7qa3Y2LYyn7mwo8z0Vh6eIBWbGA1JFYKwzRhKTI
W8JzE6B1Si5xw6KihQFckBCcyuAiT7Wzdex5oaxIJUJPvVCJaJmkrNKj8Sq8jiq6
SNjV4uIbhcFLZeLXmvemizJVVN2qFGGVkqE91JdI33KLxf55p/wAQPPo4VYkToyV
szALOBT9K2Qp0Kba7Flp3CXionO/cYeDT5MZtUhF+Yd3di5HezAv8tnGzm57SQd/
ehQOaCo1xS81lfgXk+0btTrMEy+jv+IF2cpgusoVXroyoLxcvepviqVK8dB4a/Wo
KqbptE7p3QVc3PKSMh7+M4TfArXG9FMURnIGPyiuk4Cf2hVuB/AhRvbcd1xGZDDb
4aw8QEnyTDDg//V12tnUVv7ruHqa9GSVs0BcldAEaEUqRes+cEQUFE4cN2U0QGZy
2FhMBf7UMwrzJTmujdQSvSctHrS56CAPeLxHCCIVH1cjYiw5yLZ3W7I5LPtUOyx6
u4OYYbgOOEFfC+4jstcS3QVCrRga3WYOnlW8xDNEd2FMrp/q949uk2/ahQwIkw8C
9UVDXtDNHGK16iKFRKAf+81ErPX/KGgBuPQ6koisECLKTcgkQzZYA/MvPMyxDO3W
QIAfX1BObufwl2pan7vXTuyeMx+nYMN6OIs50LXk6xT3BMDW5+hWeKkFt/XW7xBb
avcP7056LzCVqVDHn+1SzjNpcY+/FXOE3TL/gQfEAvEdbpbUZamCSgPnBsyqROxQ
TAXvjULrB/Wp9KTtmCknWFDNFNsyraTCdJWOcAU16qUJcR+qxiLoD/NodJyvvCKj
RStRvYHSp7PwL3IOebviIVIFLVENKnSj1zrY4z8oysOPDTK0iBZtB8+42JhQ27LE
6MyyxHt+q1VN0k6kEZsmkDTTMzRwNACCTvAqNecWSwGkRWZJrSRnKA5JKClam3Yc
TtJGVRHNgkKuZeo+j9haJMyrk9hMQWz9A32IA+9MnugJrx/AqTlYht6z1nx7t3s+
/wx/wpaQ3tz+27CJfRLZIFzIcYU6WZkbSxvScNkD+AIpyOtb2AsV/rRNgJyRcpZc
PyEszttdzJhSeBJ0eqv6B+plCeYYQ0zts613LDxAL16e/PawyVxO4ZMAKtpDjLl9
GfcU7nkztKL08wX6imOL5R2hLmKJnSv5thHuAFR9nABQphs3M0rLGVQYT+723y2r
oGMINVMxq5xogfOsbQuaB9r1yKnZVO1pZj/nYTipfkssqLdU2hlwzJQenIjpDU/m
pYgVWxegFPOeRS1ap4QMeveTmmc0MWytN9ryDUgcE5IQG30es1OBHNpfdnuUZExe
qoiy/dvrfrR3ka+9LjBo0+tKY1s2L6wcDvRndvw1vxvYxDNE6irwKzwFRZIORNDf
aoUW6jtzlBN7SdGB/mCvtRW7mXIVBZ0AiyjeT688P4SeWYUvZ68JqNC8FoOwscJw
1JWMYsjfYCukKEAtoGrn3OAHIfbfOpmhLq+b/WN/bW7uESbEiqlSMG66qqYmYb5g
bSJs/XCv/QcRYQFHpLAd5nFmfa2QU/4dm9hAqPJRWfKx2IU8ByTsyEbaVLtBSKnY
K1T4LECL/7DbVLBAn+nEJ9+6yNTsHetKdKdU7HVhs/EfSoXhIndgXeyD4yIiubyy
6W3Uu/6pcpWFCcUh3cVqQiYxLf1lNqkN2MNYeF3FxDrdD0YwOvIULai8FPfK0bGc
qnrPyZ8d58qZUSDKRae8euT2R76xvHBItX1B95YnpsurPQkbnrjkaDNaosv4J7cq
SN6NxkebUiqLcLr5cMlEn5vUU+Z2pWqUaRdz7BPuSDtv6Z+cjO9a+ZFwhTgjZFZv
b4n9NiaJPkilCsr7qNVAlYFmp7xDw5/KzMDZAUokCGQdu3YqLAjnNa+1CQLZcTYu
BjkiQAQKIefZaVRkeG1HMjDp93b8ato0Nk9qrnYEk5PzmZSzVEgf/bimA40wzbOa
JkExR3V5ATrI8fv2Gv98tyBgTnhgCjIJjGnLh8UrLzvkpJG6E0MQk7k8DaVRJR5C
5hipaQ4/SjPYjJy4mcVLQz8JUbYoSy1AKI0HUS2R4schEFm0ifpMLi0PhpQMqTOZ
6kpLHXosrvc6VJs0CalHYk28MDLdUHtwJtjWE13gYEx0179weIivQug+YhLIqfB1
rK+8Z+5KPYHTjcmAOehY1Yery+c+mGryYXvX+hMvAcv7UZHsQ98pjGf745jJllJR
+ijukJj8TUVTgsMjZ3o8sergLV8K7wo5ehpUSr+QFbklPhQP+Clva9D3m55Wewyo
1Vd2ZbyES3y3iOZzDjR1L+6VJyK/tkamcfTDqPQ3K609lFGOOp0ofGzr303W+Emy
2ToXuQO+XQKHPI51eWvd2FJ4vKziB8bGi8StX3z1DwihqgTfkMXxh9JrNwS5qSY7
TDEJa9EvgFztZ+J8MieFdk7R+qgl5d4nsWgq76XZ3A5VhXPytzuSX6rx29PsQXfA
vizd+4Sn3r0eYnUMdmNmFZxY8s32nNgtmA8ydarzoj7iAUK/RXoQQP5Xw1d4I0Gg
0vDcqOu0uQuYOOcqICCvMAU2XL0Abs0G4I8CyPWi0rXmnyOq6xKHK8/xh6TcAFF3
RyQwfv6kd/TqQYQ9hFcWNi0XCfUnwiO0n1uWqBQQZViCUjYkB9zOGSeE6uWB8Ef9
RhWTxTMkQKq/mg+KLdHUOPVVMUtd3xBVI0wtS4Aw3FS+KKaSX/mx7y2ukTb3Oacs
ohqcFlTIb1ZBhvPCpQdrZxvSIkEFxZjLNbIPAKeAtksNOFfiNE/4KIEeaAdJ2JR0
Aq5XEKtoAUiCMkYnHRqQoFXdMyhUm1P3Tr3vkwDcfsX4ZOsUWonuSx9o/w0PMv2/
gDO2UD979WDnE5EWvL/OioXY0yv0DlJSEJK3KD7QxuRZCAbgA7X8sz/+XJFYH984
7/j09XsE2QxmOhP6BCpP5Kp/OAHgvJh+x+raNnd0Z3CpZ2SfTMp+XZBf02DjKaDr
8JH1YFbtLiA9sNn94oqZ/R+lYaAKLQW07utRoK7/af3PwP1n95GV7iuY1QPbByTl
EholdJx5zqKp4dEuKkEk4s48GxezVIAYUTUqkiqpVm7g5JC5Ue4l7uO/uaaz5oCV
Qc3vhyjoQyMZbfxw3I5KVrAbf6qijj30KqgJi99NsipLI/JgksI8uJNIEsZtOog3
y8U9yByzinEHEDXh7H6o+EGOLCDRv9o81gsEamwCafR4T+Geg5PrEjSOMlvCEvDD
0gCcPR3sAzAmvIvNxtbVLh+6rESi/0285lnp87igL6WjwdAeDy0wtLlHTV2E+9ZG
ZPBBLk8UDg+b5Hm4+zoHClG4E3d91Cv/yQxxs7AKS8S0GX9nBwUk5AZ1U2mEBqml
hzGruKQLW3qPFJxJKtAb1DfNEm5Vjlry/gZcS+T/hfhHwl3RPbCHXF0IS+eq0swQ
Re02OtlBhb4OyDyoDNUJGk/jaIfUky1VEI1hMy5M4KgXJS/nheNbgNpeu3rD5TjY
1IByYjQBKiowKMDhep7hlyHmHb3mXrmKNFpX6dhDJzp6MsdSwfkwYUoiECw2zAn5
Gw03VkezI8asc6gag3dUzLDfOurBJHQ0umGZ/gJDE8Hipuxf036cQ9jSQGXkW05u
0YLRzkSqOAVDvRWqY3U8nBncoLqr8BUIUC/K+6S9725w0yf/rGGFDTLgM8cE4r2p
KsepXReNoAkTe1ip+Ab/OY9SM4aJi/rul877dJzQHOTrlxj6wEx4DsgAHLeUy9cW
IhsQEXTGbsoTXzOkjxhpKi6MbLpJ53rbgTqdh07B9zspUnH13fyPL4qQi1zQrKZc
mKe0+2gNnhUgqI+PQafMqVufcc9q/NHSEunMmN9VZMeq3Zh/SCqwvLbWxhwNW+fC
qpsRYTdTmfxJAj+X3fCqCWXn1i85/2T2XsQEgnaPcQ57wx5v/Wvtd8vKPT0sQJc2
/881/HxH4AnPCjczBArNhSQZxX9OuTq7Yt5wO/wneU9gFeKDaS5wlsFvrBP8VT56
SPQd8GaU2FiqLzzKQjz0wp/QzjEqyBEOujwA2BNQaGBAbvjIgvv8EU7SCnPZ2gF4
7mlOSgNchG1GUCLIJlLuuJJNXfcXF2zOuQEbDCOOC92Icmpm+NoOzGqt0pI0Lz0c
BH/0hktbtBumdkd7ysuSvRteEaqJ1OnkSvny3X1mxdu6yw93Ar7kMSrzbnr6xQT/
S4E08xr4JLWmGYnU4t/T+u154lQh6vDBmnHrL2blj6fx5/dWf5fn3AI8cUgTIfQt
wJYm4rjW7RLNH78Y3Br3NJ+MTncx2tXTdX+f7tT8wDZqp8NGWXal/XSTcHfuHuis
ISTQR6DJFyHR1bJss6s+c/AeO06bRZIGHW9yyr/AfxrCtPBPhzNXLZQqBgH1IbtN
UEIQJ0RGwFIf36NZf47Lh88hyt1SFEk9ac4FmxAf30UgpgZ0/dUEnCs26AfDVjLs
hr6tN7RwuDuCI3lyZ6tQIPoIyRWfudeI+cgRkn2X1s8d9RupiMPqXgDk7/eM7jtm
A7fN/Uc3AQPxmshTf8TJVFq0kQW8+0hAI59NsG74qeDS9r5EqxyDPJS4cYSSMhWf
WQyeaslz5tnugM4l7JUuoozrCj07tCSpDain+kCbmA1eAjp3r9ek6/z/j9ol370G
P23NoY5ZIic+xZ76vpIWP+GSxNfwzW6HmHfYPH9FhS/bLUPTFsvdgjMNKmQ5mUlz
rtKYck+WuiQiSK9siUFhChsBgFoc+YfedQRBAtxv+F0E0ccoy87wrvA6AuMOb35L
eGrhgsfcGIWXxDFUt/ZRNe45avDOubjBSg2NV6jvi08OFH6UiIp+OnBq7kHT7Dsw
dXzaHT8PyTAOhSwMlWlB30pywyyWFBHw7PIkiFbpKm44qZU9F1ZCpXGWsVfjKvaF
b9WDUI4aF0ud5zSC1aZLuZSdv9DZdOLgpw6q/WxtGIQR6mTk3IhzFGv6zKHQHt1P
MHB8Z2A0o97WOJ75hPROmwJnJ/7fmAjV1r6xKGpzzC1MIR6D7k8mEY+C33aPuIX2
VG0hzMIq8OtBfaLgTWhSWPh6+1hVYPK1vrBlFgyNUUQ5Mh2m6rx0xd81ZNNBJxAv
tzas3TjhyowkE3atOzIs0KMqt+Pgv1DBMxhDYRHGSNprjymBkD3aIDXNmxotxAHK
zAVOcbtj1ziemc9VPwz8IxVXQrKKT/WWRQUO9zavSJwcRfy3riNyGe6wYl+mOe7D
UFBwVtEcReljhNrCqrSe4M83SIQrQOtG9t5/3pWjHqRX2MqwE4/rqMUKSJwel+QF
hARCnv5jdCzX/eCQmzlCDu3XByK7cApOoOn4/8NwqtJYYz8CbtbaJ5w90UiVreth
38/yVn9maKMTaemCO7PTEkdZFaSBdZa94ytWUKOAxODEoMRX7UVMD9aM1rSb7pOM
CrgLA8IX4+ZawnS7ZD46u1MsD+66cPoLrI2a1haqXe+q41TDQfYTZP1t+RFove1O
tR/o9jxTmrBzAlOakbEkDadWUl8LSwzUkRiiYzM7FK7/bNjvjpyJ05oVhsZSF16i
j8GqNNtoxd08bHduebOsEzMPdypM5KIcqfo9tjZHD/Vmq1O1v1ASi5RjHUS2oX2E
Wt51sMMv94ntlhz0/ORepQa6dipGwUubiLJXQv2GGwqDhS5vKL+4sOVMzKiZS8v5
C7QG0WIfl1F9+PCM06LAAgVQ9dHu5LSgFLUy4TyTLVe3GQj5IzIe3Ja3artgvVWF
5T1OaPLEwbeJOihbAMF1t8v4Z5qSGCjkB5ifROXZcbByYqD3BpoywmJUUEjt6T8y
K15DGTGqnmV97I2iVSll1Fu9xngmqPScPUMYYe8iq3AZpHYUmH01UYJL0VVCJ9wN
TFGdOed6NQ6mQKxAIr4FybgeZCKPXcPRvgZZ+9OgBkZqZjG/aTAHrgc0ExvU0Ol7
CepjuFKwGcg9ARyZvuHZJhl0o7EvQfg6NHdvsjqExCg2UUiV8ZZ0RzGF469e7vV2
HzXOkiUeEgAcR+tlt/rx4ltGWd3m7xJmEbWfcce6Yo4Tf0LDIQkobBdz5wfSPutB
X6JSP7RZHy0nxAjIenk79XQaC6ThQdiKoOq0kUnSh4iSB5wLozkc01ahlPDoT0lA
Z3CiSNEBhbADkO4yuo9Xc+S0mNxibHNQ6AawOs7NA9rjFuMoh6GhN73YH/XBenOv
3WxInOsLYfa0wMFRim7sqsD72kt1HJYZcsiXayHrNFcaBUo410MQzYrwN1b0CiXg
UfpnuhRg6GDasKupZ8CK61w8+c7NDltOGRBLojAszGJdABO45wwHPUEq3ng9x2fb
JkINUOtjMiAfabzMqH+0RTMLBssLXnbmjA+T186zddWkIoIR1DWI/3c3XR6h7qj6
sNhPpHm68XzWEdl0vp1s1jismWxl/kuXxLN2miXKrxdQ9B6CoU21uu6358lJuY3i
9NTRj0hACzb92WlJMl0TmrdzDmQ12KIccOydRru1jYHAEDzBuaX2kYDgyr1o+uVQ
enA5qoBXd9qrlwJDSsNya4LNOrBmVccpNSdTiWqon9tw7JSC95UDb6dNgvoSHsqX
qfehm9o2x932kMXl1bNlafUv+KthZ8FdcByvV/atV59xPCsr6G1Aqv1k+heky1MI
JaFaqQI0CpjIOQ3HCeU9qTDgXVMERb+vG38JzC8J5kIKG5Rl6guhtbgHZIoC+fc5
JO7KDzZUZcn6PetKLhjrvQUy1uw8z+LoqyUOh8s8eBCkKmJIJL7lKJ/Shr6B/vAM
EgCqeVTfEVnRPeL/d+hbCcg2ISCybMSHk9u/RRKFjMIdCyRpVOJmh1KZlx/tB/7C
Tl9DEXgvSK1hA7qWo5Mnc8Ym13lLVUrZI/cicLUTnzqqBKWJo4KeKcIKaDetHyIH
vV3DFpVj0EDrAr7jobK1ch85SACv+CZWUOEXBKSCKtco4fIiOt7PELc/BRB26RH4
c5vdIXJaLTyJhwYJOCUdCX31JHBGMCMbDhPLjE/18ZYRLdkPB2Bv645rqlEcj4NI
jaL9X35AszkagrTlF6MZqRvsC1oQ4Qst3Xefr3PVFjPxcTvnTT3zvJkLiFSZRKhY
AWhqg2HDtRVN6kx/76AYQPXh5UD0aqSl/T8mZwR/bYtfYguZDyNp4V/6OQeh477/
/+hwgy67k4Xp366BSwVr/MyYB92W0KZ9cmfOA2X97cxJcqSMTHbI01krQQ5lN4VC
/D+Hw2SG57512nuLtf51ovQssEVlAyxcTUm3uSSZSkZ7K9wfEzBWbaZEsK8IliwB
p2VfTQVYFI9YPd3dprNHKjBP40KkpG/QpP+XBgv1TY9M4I48zlqnnhwfeVjGj6NJ
iB047rsqeWyYDlaeZOFxei5HRbnOrkutPF6QRczvSRRj8ST4ZXoCi+vWx8NJAmVi
fJnTMXoQ7TA4k0q59FYhNo2FB4Y33T0LAzD/np+rN6i1shpd9IamVtfHq/vRrA/A
EZh1CfRCURNj0c7GCsElEZC+eYufNINij3kR6d5MfA6HBop98K2Ye5qR2rx/Q4+F
5Y9yNVbC9WoPLvv+lDE4thAODmLWQBV+6SkAcrNR2RjUmpPQdf4wW/63U1DPJhQ6
FMGsfwU0msig05q4wW58+TRE48QO9bAOhaYCjtr650dXdKftBeOmVvuvljDuXLdY
po7GD4USZ7QwI78QIR9k33tK0i/xErqP2qdrTJVBT/2SdVndnOyQv7QuzPS6HkNu
GCjGQ5kXI4E/Znpj84Lj/QIC7tY4uv9NS1j2soOE0pHBmYYcySVlkdqYUm10MIN3
rm3IFBwDQ5kKkxxH0jllJV21c6TGlKvbirvI1bz090XJtQYrdPxisJ4hwn3CHVJg
2nv7nZqy0NT1iyFtcM5vu+53GNxCNx5oSUulN1rNqkOEQeb+dLSKC7BxS7VJAp92
MN8W2oP5vR+hiMO32tuOFxf8HJuexk203ApCYKwT6gfSRt6DXLWvs/di6MYNPwM0
kYQNHGrGYrsWDxM8F6trgyjDepwIHNvYqGVWajJtvAu3vWD9AZ0cYQFNas/lm+j0
Rg13QRJBZEmg6h8NCsYg29xijePkpYbT7nYiEtDQn7V/ejtnNg/tmbPMgMnBGz7F
u7OSUqV9hNDPnPqwqUFfpXnOcWknIyPklQKZq5oj/8fn1E2Lcd1ejHqNgnkyHQ9y
s3REygji66HPoJknxyZSTKJLIx8/jzXPs5pxyXWPD5RDtERdJV96TM/i9AmKzv+a
XxpUFmbSzT7hyWOoE64zEPaj4vGoJ2lplI56i8qw5ZCffwcl+ifiZMsdFZdWljcQ
jXtZtE6Fwvdpp53WZ+95RpAcCpTfGzBFVYcx8nfmdW47Vvhg4ouZh/OwN5gJqc6i
v7xnj7nRT4030x9KzBkPAoJ5l1ibCAgwZGdM8Wz3iTPQSWalKQyd0GpBvS8l+Cn2
9JmePH8R48xj/lKk866V9/scJ7VAomcJ2QmYJm+ogFuXV6me3ss2tWBgZPGw2VE2
y9y4p87jC4WE2c+xPLfSi5Zt338+slujL1w2sawKmKu2FAcD8D3RyR/NDZAYJ6FP
hICqIRGJkfqMKMD/NLoNBY2H+xPS6zM/LU0faUY62t1KlWYkC2vvHH5eN9nfv0No
jqygUmFFiOLVWzUZqEnhkiuHatpU92xIN6OtnIoF53sWwvcmiRN82AAS2tD0hwvq
fbanppmv/iqO1c1XPNlSkJyB5Brg5w5reetyiFXjI73sZhAs+Rku/eJl6M7eYysM
CNPZ4vdWXUvbBUx9Qr0knaBRL7uPfPmw+l/tN2QuCwAb42L9JHHO6maT9njdSUH3
Wmvrc9Yr8fSTanZ0jF/XAuF7PqQ4kHd8EQUX1LHNBEWHvoR5fYkZUoY2Zqa+reXZ
e9MG/Ho25DIxj2JkBZITm30gjLPcV+Lis3LDvKWOp51uCNPUKrAkTJn3fWc2kbCo
ou1n8wG+OeGNogk6D3RcNZ9uhbNxzdAGiuGOm4I5Ej88ZRuUGv64WT3Ib1fDoudW
j6BqTh/D/dgpPs3CorAdnXvLv6HgP7sSHsTDyY60xCrEJhP9I1t+Zv3of0ize01c
6/hIgSiXq23sBtpyAHc+UplfhsnpjDVnt7FMVlCjCyisU8RrSgV55P5XCBpiMsCt
zNah+Sa9LtGDWCLHqkeeqgHMTeVw8nul2YaVCGe1rjfAdgit9WWHsMTfc7O7oVpx
8H+G41WB7eq+VyfWF90h2ComSCLQ5nFOuQ0earH3SBfIs5kiuQOks4h2tOdJ8un4
pPuW8xvDhd/UoTjd+CFt7DMSsFLj8BDC/osbdus+OWAH1FtTifTQSEJDxsBkQSZ1
nit6npOM7N88rBawyU8NO2EMLIJu+otmRY1Y2oewiDGapJQ8NZlo8pFacYlv70GY
tByINMhglsuyfmRFoMdgEA==
`protect END_PROTECTED