-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
W0/dQz+1I7TVUn3UxG6BHXHcNqu0qHXPKstSIt0niexxl+gUuKAfvGvsSw0E270c
lf5KDQRZNC0IXm8aEMw3KY5Chg+3WhQ54wHVRyC8xYPrp7DTHzecrswQ9fttU5TR
Esq2Enn4FhhwNODYzu6IyAQVjuH/hcYYmdb+P5uBBMc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6601)

`protect DATA_BLOCK
PABjdNuF05buHVbwEfA6q5XsNO4lHKR1NKscNdZxcasT4RNCe3V20XLR104+sinf
J39TqTGze63ktnOQTEmLNwcN3g8F9M6LgUeaB4rsagW11TnR/jHV/rkJm3wJtfuL
MK/MGCJzMjjTZho63kqtGx2JkFHiUuA4C/PyXgBaXl3nX0FBJGVJkggg4+8Ifmvu
zeGUmBXpA46ubmLM4HEbCOWsZ35YyWW6gGPvsHp8KtxLcxrGtgXd0hkCOgVQRkra
u1DgGGULDg/To2NK1VZJwD/dqJdxlKL4TdP1Icbyr4iW3KJmgdWLMS7lQBSPNHtr
8cYFfudZn0XqujNXgOK/lBs9IQaRv8I5fR+Jo9a1T7JV8+H5vrpRakcike2WFl/D
aiYSZ5qCzEJwflHa/FtCJR8vAiBkVx5KK520oa0sVSeNaEPH7xN51H2mlc5c8Nn7
OcpxITOWlPM9G47cP4n12Kg6jJMktB5Wm816+ZejeTS8kwGg97g30D02jr3JZZhg
OoSyBoehDYqAv1XYftXU+MI8pOhEIYn7D0VhS6PnN8L0qw6B2pkdu9zLNxq6W7Sm
hEazAzZbj34UN19tdwrioy7xorFN1sSf18Qt9JBFIRsBRsUo1H9QaZanBA6dnOEl
fyEHbbzk6T/wx+TYNvBwy5GdK6PM+OihH8/kyCYoj4okNGJ4Hdkm0OuoIBD41in9
PMYeglv+5W7VUd0XwQS4a36U+4m9JiJIrZJYeS4A3umlxiYTd9DMp9lrEmQP/+2h
eUQwF5OnW1hQalhj0GiR4nYNR1pIg7bWffMS1aHuYmNvIpZDN8nygq2xHaiGNjIo
NrZhPcstuQn0qq1qLD1kBYdpzR/7ZO56Xp2tQbWS6gJ4hYEgDlaPmwPvNr+pv96u
FI1LXHUvV1m4lXPCCyK5VXBkeOGX3W66Fc+ayBx0HqBDrbk5FRfgTsqxoggSpWTN
xub6KOEa7pdDWUcmC3Y/60F4CJWCux94kbbtSWrdtmkALIZX607HqVofTZIt5Z1d
lfYhd6X4ATmXMewxYU6d4bVxv3qhwUl9moWTvNlGA5DXp81anGphHE40pxuQ3PZe
0IRr2nr7Dv40NnTvSswdYKO7Skb/Qnge/PTh32SfsmQDsmRG8xi7fOsaqVVPTqKT
aHb5GYDkL2WFti22r07e3Gv/rl1giR0E99L53sohvv6fxjvmvNJfPUuZSasVSvJi
b7dUMPbtwXGz485nquBWU76G+I9CqeOT0l2KnsBredz5spopSJ9e+MJKjZJCdWUh
cICgYoQ3+krdHy9Woq3CWBDV7jItN2US+qrjypgMGOhxDoHRw2IvYfZQ+JY2Sj8E
t2buvsNi4uJNPHRxO8JY6FhcxTQFwwREwMll8GDfs+P1MonwmYXcwh9N/9GPGVFr
hzZxVcGKXzA3iZh63rSpSSB+Gpj8gczNMeGnDSOTmF9+ETvKpGbUCh7RMsVUedfn
uiBA8234RbKAUSQif7eKemjP4wjmIMPvRHrTmVeH54te2RpNDDdKRFjqvNzzUder
4Ga0O12is94hYn29sXtdBWhzzc5Gy9BLCbGNuVdbavf1rPrbToj82dJVfNqe781v
1Y5WkbrjPfxpp7g4x/YK6g9u3sjiXSbBhdUdXn1QjVa2hyISRhMheKpuLPMfpgZl
oYlY9J5uMw21BKtH4CdDqTOslTU4PyXGnHkIsV+05gNK/Ci1x7n5pTe8zRCBKctS
xbGOloSJ9zM23Kfp5ZeQ3dCnEfirClvUAgg0GMhGvUhlJ5jlgY9wzJh+iPbd4G7J
US2C5S62N5T9autYEmIcjeMiT9Bht3Zwa8nunjayCXd9fwlCmnJsLjsfbb8mhRdY
olumqaC7dieP18hO3vFVZGDPUQCJFaX2Hmtt6xIZ73Wm7UB1A0LinY2wrRUMGkBE
HygA8VjnZi3jOdc1Ycq96N2n4aWacVkAyDTz0BAZALriYevlK+vIDO+HOdVKjvrt
ki1AvT37dC4/xctCCi2pMxdmuv02FVoxmk4OvtiK7350QD2tMdpqhYmD5zu9Cv5r
M0S2mY1XV1qI6hDMOfc1pEVYneMIN9UQNxXrsDS+cctpkzr/CF5IqFUxnaZxn290
vTMGpvtB2iteW9+gFLOBNaRtWjWL2iBh8vXmpQt6MGI6aDTBfHAA3OVG6fXP+SMs
Vyj/SG40u1GmQZbynV8CDCqb7gzIuhpXZKPOz5/SCC1d6joXoJs1ZZqnjmu+cqy/
iAMt2sSzJhDnpEIQInjlNXwXTE4QjEy5EN0s0KqRfTwwlzuqh0rhVz3rTgGXlid+
LP1pOuCd5e3g10/pblMgE0nzZkVwccS0ZUlwqMjyRe2Pn+NsfZ4Ho4p0MtKe/9XD
O3n06dVOBbcAAxQpd+QiraT/LGCdYzsxazGNxn8YkBXdmVfaIbSe0FjhYq5dIFVK
16Mz/sBxxYlZfSXcLahRaUwL5R9VsSfC8KawRS/g3tQ66ezsWyb/R+cbo07tgYSr
ieeLHFH4uwzCWBJ5bQpOQc29Lo4WetgcMBPbV/B/NQn37oRBAba/cvQzoDGJc73Y
s2wOdPGrXHNNZmPZFPe9Tp5iEATq+C65Y/H8pMr24poKoBr+vMRja1Pcrj5GLSut
M4MJWa1kLNkKwKqFiFpJZ/0Ve7cwcscP07oT4DU+Nphxd8RU0pb1Gz6uooudjDqo
HBPfEwXUWJCvQia4JHP5wmog/4hD1ca4Q+PiCg6/LcxFSbhfpSWHm6ltYkSNR2re
tLwU5ajfPntI501ABG0njAkAUf6F5UQ8REdgmv7b2LnOhlAHhPWtximDGaXDevBB
4x+fKMoZajTf/V0uLsSXckZ4es0E8+xYZbLR8A8X4MDBjH7XEaBNgtteljuoJo5v
AprSmW/U/ADg+zPyf3bumoKY4uXZIiencEVHw3kwVgldwbVQX7uxAheFXlz6kjyU
XfmcK5rHiJCiG/G6JoZou2AEWYFwNTScizYtCU6Cbp5giSRO38X6ldFcy2LnoJRp
gZ9+Us3A5CG6RyslQNdq7mo0V8CN70jYJGk2TF1wtCY7UQf9Zyht5fDYR8eIfcHZ
putkxY7Cn7Uo4ZezKcxbXjgjYqZRcYi9MwMD+K3VpqSHn1NG5eXG21Cg6a/8um36
FfpvtHFX5hrKUx991Ti75aN9FPB6K8wlJUzX8h286PHQIDpVWys1CQ0TFEur1noP
7XWi0CccZzkFO2vd+J4DLkj0PDlplfBbxH0jSnwYESIHVbEc6nLyzkHua2D/Aoub
g407bNj7kgUvY7HjS4uzqfXp2yemGg/n1xZ6nHyFH5gCtedGyubcdTN8/wSanRaV
68pNlMhbNcIU+ZfB30u4mtmpjzz39swI6HGwDgJm32lpfcaYRlvNvZyOwbNNFf4y
rQb69EZJpN1vzaECtqWnBiqjZTdIJsVUjgF4oZmdPwxrqgCZnT11r5vcpw+YuL+y
IpEd+O2l5sWvliS0FQp6qC368o8108QAd9CpYGU7wN81+RSkLpWuWoGFWJrZF47U
MzA6xb6gu+9IuLJMbDTKTLjUWvSMPxBFGrXdildWE7hjqiMSeuk0MLbBNbDWY+6H
l9byckcYti3SbcmvHLl5FSF6pWJYIxI82HxI59mjbPWDbzYC3wjEs5SCn9bm8T32
wyjqhzCoW1LPhzztw/e7sh7L+NsM9rNK1QgkEPBH3eB428E9otc2oYJE4N01WQ0M
9bR7EsfWxg3+O+c1l43Xsgjpkh4srCs9vIvcqTGa418LbCmQBkVGKTdphXYaQR3Y
PHODwxs/tMW2vL8vz6CsHRF8XgAa6LfYUa9Ttk4OvqNWtcHmnz1MSoNf1vRtlcJ8
4VZfhCGT6Y9pwsD/QdXxs0DjgOxLrefnbfsH2NAR6u1RHCUIWLgglFShVvBONOKn
/YGyHZtnGZQ1/Dj0PsI3/jkf4aZprBThlQfN1osgkGxN85Zh4Nudx5+vyK1k+OVD
IY2Fd9gBl5vzPjkTJNWJFQ55JO84SQTW5NUlCEEOHsI3R/pDXTPCU8vwOgLPbRjV
/S097ms/ZRQyPz3htGoyp3mZ26FJTlF4SK5iJWUp8Vtkpf1cEmeDOKJQ7gr7q76S
yMmBDH1r0OONechUWTvNXScITm2vBGw5pkD9Zq7+77iDqD0bgA2DMO9Pz+znSMfo
a7HckSa4W2Cq3F36P5o6GVoEIr/aZ53zhiUzcxlsaf8htd2q2cWieQ/XHELF1VBs
3TW5ZZlwV9SdvH9xVzzNbzgq3jDCA/CQtvkUkP1skBM+Ji2AIcQlt0qmeLYrNY2B
fIgNN9Jlx3Abx7bsXFPMKq3b436+3ern7kTwGrgJZLue6ltbzaIkJ+YSy2Rz+WdB
g3LS1i5nXMjrAfrRMBAM9NN/AUZ0WAjlqX+6nmpqeIIqUpxLpsRLAOzN1wzDi/P4
UTSp1sajDvYlBUsRSBmsa14RlwIFT2IyPnQy0RPmSokMCZhL5bekJOkyII7uSnQp
iurnnWoxkCbMX4PxdehipttNrtf4OWN7JQhv5M2H0R6tkcIASSiKM2skNop1Hh2H
STuJA/epDHgKdTP+XGf3Cvq1EqAwtDHG7+PN1JHtIWbWbvoA9JFa28wgPm14+WVj
wXbjk8i6Rx/hilLNpUKWVrYfnLBvXwryzNWYqyzyYpCzSyFmf7lhcdE8C0zBW9y0
RWQitZC+sRyCLfPG+d2LxXpVN1uyNyHLmRnrHV7EVg9Py3MmMi5otZTiVIs3/wqF
qgayXoYtV5/R6K0m5nvcmZi+BlQOYmfQjpBlEhHW4zDfmJuY2Be6VTRthwhZxqVM
Wi3xNOT4DQ4dDCdGbJo5UIBvEsjz36dUuiL0QmU/E6KbM53aztzcSBrhIW0zJmUX
PTZXPG62UWjSRb5wZWgNPnnDbSbjhD/q9FqkYLfISAC7CGZ0c57CreTqkJc2JqI8
h4NFtgNPD8xec+dH8NT6tDU64yzwyLvOOX2JqZzGJDGWph8vYHyiYiJ+Q5xP+PHQ
/WwdFKgInHrMdc2ebMRiSEVlyXqbDM9nFiO8A3WgdPBbSOXKk7r+9tYlFKxWyDAq
2G4UzOWXrQ2zz1u1uh7SZ23gwcHdM+vRjLD4n4Ea/KVm8Uf6sAf2SyNwRTJW5u6z
znhNn5q3Rn557J9WRYZo6j0sQ5pLjlpgO2J5w3DOOnclpzfHWaYrjj3trHbrohuG
SZEvmsky0esBYoGG94319NtGPYjAYIRJDIFTKjAr5IdigLFeT/oJqvFZW9nfYjsn
3tJ1w3LZCybbektArWfQw7/mpxEmbdDrbpjJsfTqvjvTq7VNdTfe8q2JvBnLjvQ/
SdwrbAizyUVMpmDv1emkG8cGqOo+wEfP9e2Dd63FF4cJhMLNDX6TEapKI4sxineB
dTiJux8SfrCYMQy1FLksdFy61CM5p3gY00//7dg8HKgz3rA8kEWxC5UcxJ6O7j3H
Y2XFA8e3ZqxzSN8R+PNJ1EofbQvo7FA3OTprGZXa0VYNN0H7Nnn8BoF3V4+R6+bY
rzL2EDvbQOCcK0Zy/pJx6RRtHfStVzmWKPlUii3IDVsXENQW3RsiG6+FonanO8WA
hs4Ad+ns8y6G9+Rro6oTh6RDBd6qtM3NGCToMyDn6Z/s9ofecvup9JtfOqFcAaBU
busW8XdpNh7F1M40XKQoAc9cWVZPvzvqQ2GP+AGW8yHx8n1cxm+4gYj2l10YDBt0
qOJk6gqdIJ1Cq0tBOEs7qOn0UVvg3C7w0TM1+8WKq+tbfXDnor7D0UgUvHXf68z+
fKKBF4SHlh1K51fY78rBsITWiI4qjzwedEMCO86DVmJbujegRIQyKo7d8HspNWLz
Dq01fkNgtXpHYZulQfNIqyuHmWBUop1cY6zzpTgPsdPZT2dh9Pe3DODOS2XN772T
txUKmULBZMLahVv/KbjR0nyugLoHIAhjLOBOrnO4asuzQZpYc75ZrS8esjUEGJFY
BdgqrqfCVHtwLv4LKyuo/vLJI05CL8fauDEJfZGbgJDV7gU7WFCqz9NgXdZ7EE/G
ifvmWov2IBvEqflbr06MEXmeNkUZW4SYs1SXpOEcoqryEdxZcPSguxyli3LewV7d
waHipgkL7gfQSPvzLASb2IPxBChelCe4S2/Lfjvuhn9ZOiYwvZZBoFIhe/vp5q+x
8BSx24EmSdM8J4+3FTCfVtvSCwJTEKl8b4VYbLKCtNVmCuTBAG3c7sjoY+kGfEIU
RbzgeQ6jPfAKNhpqBJn3YjvtsgAU/igzNcOsJ0XqsFrNuWKkoC6xJoBWt3W+/kPs
hBNIp4EJEv5W3CmTMLJekdAx4eZ03p4bvZZIh5KcABtXT4VJNFEkAtYyqaVrD8WN
pHbFBUMavAA38xA+4lcUC1KAlF9Ngle25M/pfRnSmVP3Apob7IEAxz0fMdv0wKUm
z4PPFAqAnnbF47F4uDFXSpLAcoDgavSB72jzfwfd5b7pCQQraBS0a3FVBXqHTB4l
WgREUC78pkpJZ8K3XhIp7AuLWpNeA8nwNON8cVHJl/rHqGYT85o/5T57DMXNZP8g
uFMZ3paTDvbxTJ8c1hz43Y07mtoYZ/52UWaUnXgrudpeK6ofziWQ7iKz1uhADl4n
ycfH+EBJbNv0Bku9t1MUvKqtlO26VZiIfMpJum778qKbFBG9yd2PqIQ1sp+g8CiU
JIsKE/F7bq+BbhP5wxxAwn0ruBmuern9zwD6C77dLX7v6FbEFNVF9uQkMIpGdQZA
WrDBJN0Bq2wiO1WNwsHMf2Iutmm5IxYD8AiIHNH+yRUqyBFLE0wc+c65AL2hIUko
CGNc7JYCP4NaxshOXSz+xIxCND4WuDqc4fOtdV3ZcwhLcLVD3WtSJp91EpIJz2/r
PqIuiJ031TcGLnLD8dDhwx1gEAr/+HpFWghnbq+YfHj91y4J15c2qmxeJqHswS2n
5yuw+1lZs3zlZ6dV5yKmUgxaERQq9WYeAf1uROXI1P8aL6KP6O+0F5IAWpdKD6lP
/EEfkEi+m0ocAiaAIuS6fM6ad5I5VM9bbEWNN+zAiOhS9NyP0B6hBp9Gndwifm4a
Hn+48e1FKaO26Ij0+hvOowFgBJyKD0jt4hBHWVMVqw8W1FpPkq48gstoZcoKFr/7
/bXmZj/6FBg9ON0VpBLbHggCzywY2E53z4lhAT+Uusvunxg2eriNKiLsmSjboznH
c8Vluv6lEWmNyOL4xmuBQR3B2OS9n+VzBYwvBITBsX6BiNq2fWgbwa9f0CrLwni2
Kq8zzjDS4OvCqNzakQHrxZOopbQrTcgL9iwU3FmWNB5zeTtT0vHAsKO0OilX+ZuR
/WZDd7e93CwG+vho0Hq0oxa03aEd0CwjMavI0rXm1VdVAIcj3zHsPkxGCga/BhWB
pe7nqmzdraCIjHUWb/N3yQVeVDzAjky1UgpCMKPn7osdsR34kRhDtu4Y35nzxgnO
3KZ8a4k6W//zNNM0bi7ahreM3XhZPpBoTFykgzLcZ5LVB95HuYB2cE94aclXmZNP
YL1R4uHbFebz5tNHQjHfobQRlWiSQF1A3wb17aKoeTsyK3HJao3FH4LZAYtOjVY1
NJEG27nW9+tIwduaGOWweENw31JTBO/C5uGkiOw77I998Vu6paTmG7HRCelfJoRl
s9oxJOZuZtlRZTa8qz9ykcJ2RJ3y1ez4xC056pcsL+j715cE8ki7oBv+VaV3fmE4
JdmwN//9wJwMN+677tHWmLVaz2lGdXstFcCt6fQsHCPdj/G+erHL5Bz+QqBYjPS6
e+JKYt1KUNN0PGS4CtAhbAauj6R39+X51RrTWzmNnE4FRizvtf6vUZ7GNcTExvlh
sf5sqVrj//r3lckj9kkXNPoLYN1WQMWDwIi1nw4oeU5O5OI+56jUJHeVJJE724gg
1jMbRCspx28zCmcJZWoMomTn6vn8F1550Mh3RbadgYn0PGz2fYxjXxPeUOws9qhP
LTPIiB1ojQWRPWDHJ/jRxEwGUJB7WEA6Ko2e2fzk7u7t2xp6BQ/rgCpa+5Gpi37N
Efu12uk8Mr+REiwCwVOrevJg1b41GEFa2Tl58Z5NbbCKhsAmq5/nQFnzBCDqUXzv
2OyP1bYM2bBn2MzFNKD+ZbmNQ5NsIVqOCePpKdUw0/QG+Z+7VjMhSw5O5kM0IIyY
RhMHU7IGV6nPSFypQOZhfzlj6gNANGtMZNsOUMRN77gjDujgwJN201gwzLvURB/o
zVwwMmmaGTzGJoI70M0B8/nWHhU/y2XDvzlvuWXTGw3MByQU0eGTZgqvZA4ZPN5F
COLRJ7dAy94hZ7PbssHiY6kB17T93h2IwnndUGGY5I/vhSsHtZSfvcKDKXL5R4sE
8+pI7UNA41ThHfkyroD8jkcvP4K+ifUGSztgJ4bhD010Lbl1v+C1d8a8TNKBvqDV
vZaUrWM/cTcVToOn/u8i4G/l72pde1CqKtkenPooIctHf1gyi0iV//jPEvg2Trn5
jnpUGwtQYhjRjDZ+Cq8iyfyp8wnSgdMFWZ5ZiNvJViTyDcmbmdjbMkLv62RyYycS
LSwFB2yZf0v8TF3Giq+va6N+NbAqRWyD/Z4lGREezmtviF6CiKh27p53RH/wxL6L
4buT6rEthwgsWvGw+7+Iupz6+P68fzZK84YEGBTCc60yBFgxzA7noO52gtD8vtOC
tIj645Yr2DyjkPQGvIYUKTrpRF+ZxXL23nShK2j3akMAnbyEHofdqVvtbeQCDwaL
BYuv1YQniYKX0Nhv4s43xK52jU3wCxX0FYmeAtErUZp0vLYjCSRYC2692Ilaa+fi
m5Xn0BZ3X9Q6hlpq3KP3fxvogggJIyZcXH4X0j8XfQI0NIgFMZFZeyr2sXP5rVm4
`protect END_PROTECTED