-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QnNaUSStXPvaRapAOtwEq8MU/ZhcCrGeXoWWqnWS9IXfJMBkSaDvSIKtX2vLM7xMMaoVN61v/qFT
cgmzaiBT2vpiZs//r/TRyUVJ8RM9Z5ZEGkjr1FHIcjzHLUZCdxkJcLSHhlEkvzMbsUZGixOkxwLH
khNq/xVbXrvd3D9pbh8UZRqR0fXMEp0mKkyY5TIyYCrM5vWg4m9L3dl0VySPHmwS3/jUSAQsR+IV
x5PGWWbKN2CZleqXWQAXEaE4YB6xHEi6GUYJnGhiN24XqKxfdrJ4vvbhvG97KN6cH6su3sCRp7Ef
0E/E2kwxBx6z/SxPiDHLnWdnDMBjSKWIxQdGwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 121968)
`protect data_block
4FDHn9daopFZ0L240I1HOj0v04i3BBpZuCic7Xidf3mGu/VsmlFyvLY0rNi+f9SujTxN/b4wvYax
yYmD7wfQPP/5YMx8dlIrCVrFX64e/X9I1OUyMjFCqfOXiNifYA/Z7GXDc/I3yojKhKEasDSGCfx3
EaLD4YPqN7OpXiOgc3kap5NLxNYSTUCgo9pSp/FiBR/+XEf9gQjzlJwEKc0gIN5XIEjfHfvuvblw
rcNq4mFuSHAxLQAhmIAT1QclzPvojX288C1nrwdrPwlnWcP61QAlBN1zPYxBFFRJbrOl5Cxk0560
lRCJSvrX3Ak6TZwjbgWwddCBMBA+164ZwskRX2MWGadnxe+iIspR4Yz698eelDkW5wZDN1rj5h+h
S3jdL78U6v58jDQOQYqEHmRsCErYob8evdtM0D97IxaEKv5q5JVRwYRpVQ4bwTTKxrgulRcaqCWx
dfIagEXr6jdvLiAGGIUEp1OsLQ/UJtEccj2rjxAl9N0jh1nz2tI8ChmD36y8jtwc6vXIGZ8ISz5R
xWcOrBYWvT7kssIFW1smlnv/BGht+TYJlN72kGBIj6XDWiTIauwvWc2gVHpbddJBW2JO2qS4oa62
pQKGj4tHPJc8KEoTGJA5+MWjoNm7bIWkPpEOHJUR86e1MCtV5cJ7h+ETi06yuaoHvhl+iBaIJtcS
MhL6K5Ak5xttJ7YVZprCzhFwMWnN5ge3iHbg/uBko1lKz0QYCAnLc20wf6pYE91dpBgLx3V/iP50
S+Mv1oSYCp+dAiiaToBDXDwJma7TV9flhYyrVKrLAytsZBDmgU6JI8nWlkAHcIoP0PD8Ar/sxV0n
OzDSjuyOibagcZ1vSwKoAbnG+Y29JMc+qP9/Es/XGn/1F+qM8FZUAAkQYYSFpQzsx6VFY9PEY9FN
9COZD1HZ9YkSzyrHE4Tp5cIpF4+b+AP1xnlvdSR9BYeVSzjJK7CTvRvvMEKDf4In4wGqB1hI7r7M
hiUUlKUq+ShYeNmWOv6qH7u2/EV+VwtBqZ5pKRjeqZasu7pD4SOeIn6dOK/3HBjMnei7ub+6tyUD
+1q/dJ0fp6vI1pb1VZH5B0ia0Yufx9b9ylqwAbzAPUeOkGACwRx2d3BH6tMgx7LfF4zb4oCiRctk
3RCjfxrL3fuTBjUWTPxr63YjNgoMg+NSBQeJpVP1Ph/ov/wDgm8ghxliOrrF/U2Q991mFJQzMVRX
6JhPzfBNX/4oWBBa19ZriSqpsTl1RQtFQu/3CArU+S2vfy6/CSxBX4eMfYCAzv6rKsICnoMOmHeR
S+nsHooHaikaLHTXVSGNNL3+6iNLcDB37XjKHbfIq0E3XCSf6afBhwxbZP4vpuPrhoaKILacGK5N
5bLeZDGJSgzdF9kPw61uddRI6ibCFLwYSMgm2GpmMo0h3w9vPfxTzUAkTA4go0IaNIOS7p+PxFIh
HvCcAIPBmmQ/iIdOpCIYAp7bGVjFEDc/6RcXshy7RQcplIzoockOc3ACBS+S9Cu1ScEH69i0VvEv
+XmrKDP34QhO2RHm37XhZCUDL9Pwi8uaxyUpXrsa9uSUqlRMFHA9MeLJ69t0J/LpeHng8Khpqgvj
4/ZrGr3j3+oGssirM0y8hZIcFT2RofoJXMg0JXPIUHJabA+sfIj73y9QdUGYBV5DIJZV7WVhk+1t
brrOIpkewJu2QAiVA9JB2NQj1t/74mQHDto/aphATQPmZOkRbckxjUEZqfmhP2bLb7u/R6ou+I/n
C+xri5vXZxf9USlMMqJDqv4rLhKqZUO34Ga9lYYAG2GE7/kkPdYayFOvem5dxNK33ou4q2MF7PqA
GudCPdRu68sE7+Sf4JY+yqhYftwhIQymi+7WSiB3jwfbihb/r2Fyao6ZJjkBhk6EswquT13M39Qm
mZiCNrcbr2VqPDhGY80YK5RDC68rIYYeG6H9IcwNx6Dv1r0IrMNkZjkRKGJivmUXSTsRQSyYoRME
sokl943DAsb0TAO2ApoAD2X93z4qDjgzeMqVH9wB3sx8Pp1Yj3QDt369f1jImVEibGjtss3+5f1E
zXTc2zjuAqoCa60s6fglqVH+eFxB0Xhi+OIAv7MNgiakmGSqYn0OHOo663dTyuOChqEtRZMMXaSe
MGCTsagAdChQnqtCBDCq0M8gqeS3sEHY6S6iQuBDBtaPXoRIqC5ubDPeqkVrEsyebHSgqFzmPUe3
kVvAyQ2PiDzrs++yxU/rc9AUHz7xJhc+2X4hL8OJiGjTuQmUWYcTHP52OGjiTpWFFBS9/JjE56pf
j3lY3Z8QJnzREW37dsGYggydAg4o0UKy/qyH6UpR9feW5DJG1+J99pLpscpFGNjjCwJZ9+4bTpH3
3CCATrXoM1Eyy6FHZhoyFNR/7utpmxy19M+n0nRK/zpniHbMIuLgtJpCp5DD8t65uRNgVfAZAKPh
Xugnz6iP1JyS95QPtr2MHVJhELjcqBV9Tvx93GtqD26dLienBCuUdmktqx7FCiqFXuIEQ+Yrimg2
o3qEAhtWgZX4whVRSrvUN47nhRIsb5MaPpG/DytIavc0Y6oQbkFv8ph0duH8uHFhabY2JqWy4oXo
0A7hBboS0JGHGPdL9Iuy0l/r672k8+tWkcrAmGdV37R8TdqOoRRTzTuuyEsWeOV7chHVdjaAdDUp
Rdpmx5ozthsNcWwt4QzcNyJ5k4dzBdO/nlwlaAVjvQLAZRwGP6wJaoFEr82yOAEbfLqZh9wVkl0F
atOoa+wbzePBcg5HBx+vbP/Oar3OdNHdpPrhH3HNQKy/p8psFuxzdqL01R8azfVE9DAPKzBKNNsn
3l3IIP0n7oBdUp17QSydrwSTC0tCrXGZjNnwQ8Y6X7QBfBYONrg0qcIZya9PQd0g9oI6gNKWror+
HBcwIcSVV8ox1JMJ/HdG8PNZyHz+HMrmmDK1AegAVUK1XsVi8fwmSOTDfVTPqZmWA6JxxxvzWvMS
6A5PNICbI2fm8WVpHekSLw5FbQtaATiDyWrmrWvWfuf8Sq5K82BH4JeIRIJc7Z5SH/yk4PVEZUH1
hf9kzJLz6lyNxlx0z6THPfaskuQetCjYR9YNKALzo/8Tcf0GDxXjK28/SO4VnK1+rk1338yhqVEu
yU+cz0Ih8uvCfTb26g1qe9zmBxoreZOHe2b6KxN/yg8wB/6/P1ov/g/c9uF5gnhdVqVTAPTsEWHa
03UMu3elW85Lg7yu7nTKn6vWk9ryaq1GmKDLgUwFrzNHwhqjn6dN0FzB1GzS1vKM35SPTqZk6dxp
22RVXBbh/yhGu01qTySrV2/1A+2baRI8REH8xNIR2FGF3OCtQ1l3nBacLSY+lt+z8cyJer5U/kuC
hm0AilKRFCGNvBh0U66ocxeMwBkIVyYlJNOJNMR0wFVf4Q2XdOaSIPTe+t6dfUxYyInrQ6xR6Hsp
Ua3UQJgJ3rbvofeHh+OHD/vyVwGLmQnP4t05+p9TCL48c7Eq78kHJYRKea8Y4+Oho/gbaEYiVKH1
5wg//oh2qWAK6s2Hcq80fKUIpFsOra3n4D25+O0vRsI1FuiBj9yGMJCH+x4Zt2F61XFQajO9tgYl
zmKfE4oNmnx/isuWhrNmmEJYnSTBqXuvHRhSYfZhRFsyroBoaJQpNoQ6mCtT4CVZUnmL7B8EdTNj
R6VLir8iVfaFnqZWPYzTwvDvry3xNcUnJWOKDQJKHGQqGh3Qx8wnWxR30tcg6g2boIpOiE6rqfx2
FVoCnYxSCULPQPFZKQvGxhBpqo06yMJ3dJ3Om/SuK0VW4AQzKtT91lAXSEIvSJjuytEv5t0+cJUb
TbPPqnYiSOHHxvGRdD0Bv6u8I5Y4nu5AN+AyDVTCqRddXfEF/iz2l6VgXL4yvN7MQLAWK54zZHB+
k6CDqOD/HX3oOtt20+ms9i3PSIcgFI3StmX/EEj1TIJxfnWbcmoWsjRFRmvVLqCCYQncOuzUGV9i
rSTZZqjDEptb5d70sQbMUKLtAJMkgMnMZRVMSEbRlV5Se9/QbJSiZy+fhNZNRwoNEPvNkGCuX4ur
RN7Z7Xjtv91aowKVUHQcpeNgLQQLHIRQ+vLCUxAZ6apsQkFXf1qLr7FRfYpqXKjAzkD+WpTVcToh
OXjLv2+inTpyfJvTJTN5HUp/I0pRmyYA1lh9AZ+FaiOBE2Bxr+YcsgoSzH3Bm6AJpva2z9TB9Ex3
4SBLlsksJlh/uL8K9AKg+cpItp2LVpHWWPYStPwfy7BU8fVNzjYQJYAkzbGIjxyulSIPVwtOPipG
5VwStQnmnVYrvZyMsfyBo5sUS9gnTC5819g3+kf+RM+w6JAMsw4IeXJQnLomriKJKGsHMa+Te+xU
M0+5OQH1DFQ/lxqrhZe7McRCsG5UAdmplb5S4AkbQZ78IG3btBMPDV5kwWeSc1FouLxJmr8etVKS
IdtGBxm+FvdsUMalHKvMjKEYI2zeT57ujyPKOhHtMC7U+pbvSHTLhiVpDQGwrxzqsGxg1p50qSY7
tlMlIdpVNAnjDZNB2jrKgtEMvGygCDGuVmCtPkBMpgYxPY1suTRNJmPq4BQb9nfF5fUvsJwrJgmu
/JluAjzfTUGz7q6p+h9RUZELoIUB4k2neMeYZ1nKoVN798YGGEgRre7ytVnVUgGVHq6wC5yFQIkE
SBxohnebOH9WTRY6zkn3LSMxgwEn1DD9Ei57guHct++wGjmRjKvWGlMWiKiwdpBXceqQCM1qV0sn
PsUtr1Iv3UA2icfHps+h4dpyNjFHNkH3aezuAB05txX+/icoFUc/NQ1ccbt9/Z57tZekSpso9hHa
QIs5i64IkiWLa+Tc5VFr4nOs/0DGCkQZqMCE+i9LS5ZgBhaaIID2qON2Cd3oQZfd2KC0o/QvA/4e
X3rCWrr0HnYagt4MeYCHQIIF6QrRIotMIk2Jfkrsp0XTkb0f/3YJHheqCNmv3gikv22PCdJYlf2U
dyVGan1BOUZch9QyjSx0LDWiEHRjLFgjtcoKJlAQvqVHYQZLEts1U5PTzCgNop9DeTEZSfPWavr7
0DYUJ/Zv8Qz9+ywMd0bqLgIio7Jogb/1x+qukeWAaAWxjVZbFRnkkBRlTc86TiR4+W6SzA11mE0Y
OmJkFeeYO3KD19wKKyqdMKw5+4wYsqDA5wmfha6vTe/IOspW4xWbNiZ6PgEv3T9hkEZ6N2fssokd
3aXvNGxbU1yPQi+4m/tH1MrYdi7rV7Qq3VF7NusKZZO+FUNIOUwhm2jF/mrzVRYDfyZVQBz/goHR
7uVOcD4KtictGJTrpp1X7Q+TRsgm6pKQlumu32okiaj728zAkrxqIDbf4ndyh21Qayqch5Uc6ZOq
ci0bnskGZiBA75SUNtng4B8I9Gzmn8JOBfjm0K5YLy0fiipCymB5mSL7fe5C0AQOR8S9XVnlosd5
Xt5wgTRSDc5mVIdGToVcdgZLqUPkdbxXnBT7L1QVsKLNj/wu+A6dE9cTk0Tc43fXOSRlPEIYcIpO
nTIN4Jy7SeBUN8iEWd4kw6n7+gaqPWpnxXqaoi1LW4UHaTtOvKrulIw9of3dJP07gkwlhAJRp2PO
AMi3tnQXmYEEfdRUofUBwV6CtDfw/zcTR6Zda9BOosTOPi3a4zD451pmhSgqO3B2VTN4ypxjksGU
s+hn108hp9uYx5CXZfiqWzEREe76Qd+qCqwBPyDU8FFFYsQyeatDlrVUVErSZhgjpOK6ybigKyXa
mNH6kKoYGuDIPygVbVL/Sh/tahgmQZaoPSlibjVaiDFMpbNMaFBFe1sGSyyymGF1Y4HIUmvh1jZX
OaYVM1m7P1cFX3stcinESmcp+QnubjdxLvP6dDhXrqQobOCzowKha7vJdFQvK8aOsg/Ps2o6YKwG
WzA0N4YF55AWsYh7if9ZEYlC4HjrucNRhrBxo1xr5OKS1ACawjhY77USRa9rwAlNbhcPV3+9NPl+
p8KopP8R6qwpIVgTrIrAdEMeO+Pqwhb4g1F7Db/vAvWMG7c2b5/ZRJrGxyww6Yo4gNLN0KoX9gF6
lTp9I3gSj7/8mD7lWgAcXQPfXpqjPfASkYHQ0tESEwajQ2YHjoEJ0hPhdYhGGfBQfdp8jUt5BWXZ
mwOL85PJkPrQ9ajalTDox0GC1QfJHKk46DijCnk44V/fSQ7NrKYAg4saWO9W1ri5DTeaxp9HX3i+
C2n1InikUO/cG67yHK34kjLS3JuaWwPgRo8fq2KbxqI+W3TxVormz1RQTLA1+xAFZNCNPlTYAfqp
CsqG0l8a6334h3d3UQg1u8LhjJb2jgOBF2GhiPm97lcR5vJT7Uzs2De1TLxEAhtKjrKMae9fe2s1
YgdbUGp77he3U7deYMLqCe5EFSJsmlphXeE3HEAkoROhG1wRnMmZynRQJpp6F9JyLrPrMsBjV3w3
jFaOuUEJumwRJeXNvaIa6yAdHzp65HQmBrNY0zRoQqMmnBQM98CAbUq2PGXD5MVl9WcPIFq6hWcl
ZnVRJNyGF5bbiWQAWWfqI2YBq42kIX+oFxuINBH8OMtuwtHEwkeSA5DCf0uEciGyAkBwt+cdLzM8
++8gsvJKLB1lxCPFqDflyVvxCYKBmu/jAOdHd43UBmyXa4zqXGhm3cCs6pUMqDuAaI8nO7gw3TEV
Jee4CfusglhWvZrNT6fMQzGapayvZIDkM24l7IkGLwjNjnjtqrKjQYrQ1kw57v33AxYjNxJEgxqE
UjcggnU7+3HvPt+r/crQ5mqhq3DoqKAErKyXmrUp5dXEnneXEl/OzJyhaQeGRMwbEB/OCrmE6q4g
liifwbSH4PZBy3ltJS1jfd9E4FgaNmW0VNLBl4d7+GYD9mWR7mB8UGwOUfXC/Yx042PTRH7xZ33O
dKhQwvpCW5ycUHVHQEertvY9a1aEN9yfa38Wg5kHFscatjifWQRCrdQ1/lIz4qVixik6H+qur5bh
F7aBEfFcWXcipmbWsr/J9bnLVjzmvnuxHivmJtpVI5r8WpPPGCtg2//qk6ZubvdkXU0XUiuTmm27
SOeuZaa1dCehV1Y8+YRJhyeN2BqGT8RwkSFJumXjyyLQnnM5SrsCs573foxzT7yLyfuyxgDLskBb
jej5LTJJOFUpBtuu4inW0yx8bSPj3kYrBy6M+EIxBQHrt0K9ml/9ufQeqvGRfWik+mAcWgBqPv7+
Yu5wChUbjvtOnk4jqVMbtjre3wqCzdlTnJzhvH24gp3o2AtZMtjT7TQ/+sFsfgeySsvNUoJOlfsR
z7fJrzlbaJf7E6oQtZkjH3rRwrClp2NPMy47kB34bLSYnADU+I4G21pjQMun54W1dST+NFqtBKaN
Es//QzkKNKJY8P+mBuNfns6sIr/xpVBZf2SALBte6gRSsVbr9OD4jsKHyLFD4hpE5AvtGMH8Cb9J
OD8LzilorUfJHDl85I4LfMf+LZ56Oqj/q55JumDRodYQirZr3IYARRlfmf/cF+xfySP7ikJdyExQ
yulyHSIofJpvfkIup0ZjsZS8ffyzp+SztgT4LKFsFpEltzEFzcMvx3TWn8YKe2zZu8yYwKc1oXrL
k+QY2JsA5lCREvrKT1XkQp5+JB/RltXn1bWjY39CQoW17R270saDLx0tGvw2xx3Ho2kBcUYMhSjL
FCRu363AR6uyQTWZYq4NDfAU3h+nz1rHxCVtGyaUzFx/De+djjySsIrKX/gXg0mpvs0PreMG8zV7
tZopq3tN6dBB3cxOdELnpKrqtsTzVhiPBKINS3W7RmpsQwtaFRUjluk23ylEUPBHesHfhhd3uohl
QUc1R6WjF11vb33kIO8yhrmA3LBjgLGFaHUVyEqBC0C0XVrQLy2HPjeYhhoHwdm9Nij66wZzy1TY
ChJy1M/2jFmCWOcigy1itS9/e9DsGHN6P4G3FaZ5EPSseFNpSXe6CR3S5LTLtK+ApFI2ex0wnQdG
u+AMF+YMmcOzB2djSLt5i89jfGIeRg81XuIXXPAExK5YQA3Qd02N0MdUXSMAQz00nD2kiFiroZTt
UB0bc4gcwcW4ZBlELKQWYF4d35XpivKtOOhsbKrerycoqUTNokYHe/OjOQDjt0MxohVAK5x16tDW
Lv20f1UETpLgL1WC/hg3b6tjNp5vioFdgn+AKhwb++j2PnGWJs6uQ8ReJ1yIoGp8NSbs4SiZgLJm
CEzKwGifIiDvZLgLhRKOiP3USnkzveHzGTpXA7n9hOoa45tFgIv2ui+OMpFoLPPfeakBQL8c6zNi
dSxyP0i/teTGnATXT4iz/lGw6v+EEIoavdOB//VBwT5ZjHtwyGDPDS/icUaWLVnVVKtchB6ARm6I
+vaF0IBSRB3QWPom5+oIT+ruhmxm9uhsPGRcgBh2v0ma1Y85kbDvOe++ZNKm5vCWcIt/H7eq8/4c
QUJMFXzUDpIx3gch9f7iUjYOUXgq3AW9h68RPdHWK7S1mqxZb3U2/M/dR1NkOeBmVvx+4N78BO67
XhVUWB2ep0C8KNie+DG7k5K0W1SrRf0FKkmty4HtFSoc5uPm5pZTYUNRn+dN/KDpglulelmGTT7F
s3GD8VMmxAkA1ldzJFeCiMBDRY7g3APvD2vsXjUBYqnV1Q4oLp6F/xRsUJOK/djsotQlsufPTl8k
J3oBsWtjpMywNSwrLt3QupEjEOrz+8hH59pmNrM7Fv5Fk7CwgbnhoHbFEjX3u2kLyiJUjLc0Wrrn
iQ9l2Y+iJmZmTBie37CBoSt4SmFdPuShgzTLV5gwKRhMVdkusLkw5eKhImS1f/iRGgvus/gzUVXi
g59sZkhgur1YZjCfMlnBMJ91CmN2CG/evL4IkaKpS8Gn2LoZHYIvPlIg/yllxoErcsIDOoYfUHQ/
2g1jQdq+dX716iI7RDrFfOE/zmQstQIxyKAleleStnCksmAVki5CWoqr2KslIvM8ZTlcyRh/POx9
LPAYiPZNuhGuXQPmgBDz4FkkgKTavjRgWnGWWJJIuS+BcuZzaTX43nfE7RjKmiPmFdtnMmFqeMEF
uShymZ1iVEk2RPbN2UiPTOnNEjRM+M9dWL5Uzs/IEwVUZK8II55CHIe45oeFfUBBw35tgulPj41m
CPwjDb5unzQLHSd3a/2tTt/eojXiSi60disd+J+fdehLPR7JODLFn6E0ODmyMTw1wct4JJV1W/PF
L1GSmuGSutRblLA8Ub1fqp8A0MnwxqqwXJUDg5DfZcvphkH1X99ZRxx3FVikQQURhJI7+xgIaCGY
+vvzp34YRHKAo5Y+wuCp0v230PLx3zoM2ZmeeLDDD1vCrK/+bHFz+TarihwnOccpGVZiqLnsTeh/
crIUrFD8fqOMQc4Kmhr295ZMzpspdWkSiX1nwsGoYAZB6Ru4uUtuIXUrB72b5v9RBrEpMbjJh6Uq
11d63ekx4idq9SaUuIBYxxqwNUvs2uqHRrff8ldfc2Ra4XD623V6QYJwE0eCMpbTxJp/JXmPpbhR
clsHGrYl/afw238htwMXrbw0jeBs7AB4Sy7NYHcrA7bs+XAP4gJYjCck5jEKuSWbwg3GNPhlRWva
HPsUKnBf1SG31FWVPVz2uqEGuJD7irdbD28bJUihR87dlt4IQs6bdaxtkWx81T+N1GvDvNRAv/Fo
cNWwPu81sEoVrR3AFpNvbd8EOaKR9d4mIjHzM7vY1jA9bip9ZthhcsOGvosLRbB6O/ePMNZinriB
y6pJ6qTyYpPNdurM04vHitwb1FPPrnZ2l2OP0iKHAwSmTJqz4F/cnGtOQSDcbuaYLuhRRAUXypwD
/eUsp8EQVoyHuyyr2dIfDDk1mDFLc9DSm/lM1K00VVGdNbr2KZob9rlKcGhA4b1sM8ic/IGQGvDQ
VYXbSwCVsAHYb54EgSpg0yS/0OWs4hazdcFUqz3U0+J7/fHzjiZqqibSVKns3EdDqOv09IcqA7RF
sOCR7GQAVr6Xsw0SXMmhulrVUAs1R6bAIJBS2ILqvR7k5evxcc8crCRDgHfii31Q9PDgD78w+o4C
wXStgJl9g3qnBaXWoY3N8QQorybryQeNylUyGwT3iKK1aXPuDbcq7FcDNfSl4jIr7eVdSU4H1j+p
UqWRIwuJIL534CgMS4vF6gGkZ9lCd5h1nJYLy2OJ1dF2i143WpzUwWmraxa7zzWiD+dTeekfgl9y
U4z3jMS2vQycqdkxbWLPeNnxQ3/lbvzjE/fYOlotqw2ADu+U7uwVSsoMF5YjnkpymwzHyy+/FAvW
9VSp2F09zA88ascBUGS+yT+cR4lVvmukIWVGw1crWU6ovGilV0XlReSzwfout08rTKG4vkaTiTSZ
xmZ8psIVQtTUxbpg4idwJsJiLosjQ6GXhgsxCO3psuGwDSVGooKVIG5dWuxjrs6UtaX9PunrKdiA
y1Lx8yVI50VQQ+4yW8bqCTNT+oySq1XtY13UJBQLxo0V1LV1v3tCYZuit6xlg2UddbbJd2n4DunE
IGSzN/iw+r1SRpSNCrsQvXMCLG4qIUxG0wJNC2UzF94pGEgH6fgKKevDZH2AvYUQf8rwGEDJuMj4
JRujU28miMm6xeWc002Yz1qhokqNwSQFCXTG6fOjsAU/XvXJUe34q9jzXjYXm05Vn6Q0nL54AYI0
Yu/6RNmjOK9FDOKr66v7qhSUgivDKxPnYV26YxBUl/FbwIAoQxuVt4Ap1LmCv2QlyH3u3CglNNqt
EVWLzcUW7QM9aPuYXe9Qa/Yh6sAyGHjHRfsQy9ls0Bp0+rvPtBMjErABJfVoUnIL4nBPjA2y09GH
CjwSVCXEviMfM+nCcRMFASRXFGe+jXYmxatuWAJc8E4XJPXB/LbT670pmsr1wxBZSdEP+Y2vuuzZ
WVMO7KE0qIBB0E75T6x2TUoePc/W59Jw6lvIuVrpt+WbmLczH82mM4yIdq03lafal3bZd2QOiBqt
l1cPwWOiuWIWfoWs4WGUYcK8xauKX8r8JV0x/rv2fltVzOSqUhe29zV8s11NMoleFRAKNbZnnIFn
uLnryDFC3z1EyPcOzlyQcg3xaDDSUswzFN6646XuTCf+cZJvRjUS4+cu3ltZ+McKQEkFg5PXoGOy
IAY+1mvrgX0PtT6vRpcpHitPiX42UgZq8BkBJPgPlJYspaH1vva2pspaJcC+Z0qgbBy5ia5K0zWi
d6CYIIP9HdvH7/5X0SR2hZ7q6yTX4sDT6lsWaAzM4WSU/z5jJ2bLMn9nH+djGwCLJNc7pPK+fr2k
JTh+8KXDY0hZTNSqkqC9Pgas1VzDnu5vGPBO4Gt2bjjuPaNg8Olu8PzWVOmZDXoqO5ln18fNfeUy
NgCrYGLWuRaTbTmAb73P/iWgMtIocS//X37pDTtaZPz6rPcSi5MVhGntYNZS4UP+N4wKCFJkJkgG
3iZXVlRlg+ar2Uv+/u9+lyUl6R2pglxbLXPkKjaLYlbsCm5SckyDZhsgvY3c74fE6Iin856WlNW9
bPhxJjCkwCILai9PsLezCZT1fyVciuoKLS/AdvowS8CU4RGN+sucYCb7eMFQ+D/8D2Jz4f4wY9xX
nBboXhP0F1gOw4SKbOknC8Jw7ovvUJwG9r/KH0B/sSbqyYo4TclNQ+UqbzEu2gKt0C66FupJ58b4
aBBHk1kVXaLocE69WnLWEUOvXf2jmbYc0bC7Uah4SwzEbCTqEI3/lN6Mf0OSAyxbYiyAIx6fyHgs
AKqZUSh4NaDS/pnQ/qXxQXhVk9ymEKI37ScFsKbE98kRqO1p8VwB85H8+n06epB8rrPAJBsM4Xkm
BH+1mgvAS2zq1XIx7hz1A1ke09ps/O5vb1bEPQrC62aU3QgIWLOKBRzbc1hmVJPbQijtFUhQOdid
fuNcQbdleHkSiIJ/A3QVcs0DEkEjl0RIDl5sd08FVliEfDRSCeBoDIJt5q5Epy6go0RwMNnJTf8K
EhZ61Iq6duipNTWWFC+6ERc4gL25enw7Jg/MerJoouQkEJIbc0CUM6XeqRJmnPcQ7QLBYJgob6GE
hxv5aPF97s0W0GZU30QY99Qkqgb44ykxQtxa3LDTCVym+Eek/TUansKyWEmEIHit/nRz3g7M9JZt
utQTQP4sN8EMhubwKTCgNN63W45gnogfGQ5O4//6f/Cu99pxIY33wHQZ216UHej1fkmgmGezSH75
tlWkDbsCKSS8dOMDbiL8IXShAeOXi6Dr3lDOq2bMFDm8V+fqYGAUFLEKERAPrNKKrKEqWwwT8Pkr
XfmWcHpssoesMD48ldcMja2qluOjzQX/AX7OEt3IPjYs48m/OY4lHChf9Ne4/IPEdiQcsemnhNbn
GwpNBZcXh96GNMAM1b74IniaOkcUg4kGkx4/I3ItD73O6ghmjV1yBmtad3etahrdRHpH4bmHSGdZ
DevEqYsR7vRPJylolTudsWgd59wkEx6yiLFaMLT71kB0cnAvjlS/cWeaKm6EQxNnL0HqaeOEIbOu
Gvnj8gxgUrCV9lCE59CoYiZkEqe8PclVK4hp7umkMvBwN38MHOj4T+2xsv5ATh/RyFVW05Wsc0hY
iJYYZgLIdJ3FghspaF2RLebMS9kaZmjxhH3c2OJgqBpZti+M+ftmPVuB2WJZc/J80ZCBzHYzhI+W
B1Te0dlriJCuB7GNyVLQXkRwuY/rZNFbiexwd/Fzaz8qHkLEeiXRBwQ6bk7JD2X0zOj5oiAbuEXK
4MsJgXsJtppVOgF08eHe8kpoXcGojYS/k0WHm3JbWoG7wkvWB8PVZ/hJ3kZXv705r8DDiacLKEOK
t1rUZVPZTOLiFPUbDOJ2lKEZIbCKfV9zjY7jj3/njXmGQDTyXUPtsiI0WD/r5vdX1bUHrWgofsmF
rh3G2dJmoNYmfcCDZ7XTVjaeg09wI1BfxCRkhgwIw7uPeH3Pt1sVjbsiHhE97oRWQ7KSl/WdiJKC
rozJ9LMTl6147mbOOm59qhRwineN27+Co4lARpny08ipaL4HaEEXwVPhUviK+4AR/wjOsFJV4jNH
v6Dkuyix0SoBIzxIvHfv/RujvBfaVSmCN+IVZkbeOdRbW+DKZuHM3T/LX4nSTMUstIKt+pQL9TvU
e/9Sm2CU87LkGLqRlu/AY2vl5WN4EmB/CRrIzOfpxiQVK44xuoffL0yAjqdrEarR5BKrWtRmom19
YtuQB7QRoO1BfGFMZzKb8KP2TeVWInL4DplpI5sHF1xR1y9SAekxaBF72ciHBwatPKbMxMXQM0Ek
F16zyun2gqwGl1SJSJfSuJTNC4GNlnO8tU7XbX6jJWEu8amFT+/FC54YnUV1VM3+DTGc1fbAzD5M
MtZdJ6qUen8CBO2JUU9o3jhgXqVsBYQ/empPGejIItWWuaKtbTHKwPOaj+nmuRqI9rlAsOFWJCw3
nP73kb680JUqiCQRhKfRwodxu9UX5gHi9eA1UXDTDD+wstpWgNl2UUFaPgO0T5gnweDIQqwDtNnE
EAfJxzRIVZX5vRP4risVwjIoC0YnkusERKsYstBJ3/S87a8EXugglUqcdkP9Egn8OTNiJbmsQuh0
fpI5jrB5YSE4LIcQdoFpcNgd2qkc7UQmWQyqSXLhddX09Xr7mXHAjq0NB1V82XPsbYOgky8n57iz
9JvTmtHN5hyAEvajkt/Ay4AU5XffCEEtNl5NsfvHRw0gbIGz8MKFmfqrNmwJbiLfV06PQYBY3Kcm
3xiw9k86NPobdtuNzwkSsHse55voFGCgYLOTeOt5wLpiiiSf2aXTN57/A9IgLJDpGies2AWu7OiW
a1g3BsbXJeAhe/ppJnbID3rbJEnkobzzHIA0ZUUhD/rf/uGHg2lbn+Fr3LjssQMPAlrDdDdsFRjb
TJ7M8YKKPYcvARMB8TnIwTWJXgzIUn5iNUivLOqyr93LQFTbhO30xW+O/4uOPkUMxU1d1D689nFq
Z1K88tqWOPVEW27lXXtLCFgvXHrAmtOcoLZAlzzaJd00RcfVAq8Fw28YEMQ1h2gId7cy6L5Pnx/o
jaNdFzn+OWNCqEpmIn4iTK2W8CyP9oxLP9tjgGXrZhTKJFMiSlGGKIuHh9dksnX7Y1rSgeXRrCUR
LQzYulLDcY4EKf1NX4Uqjmdj2tqnk1wp9Mc53HHEeCJl6SVyE8IjVszMLmALKa8xf52Q0u+uC9u2
FoSK1zIWkK/2w+LTn/L3Tm7pOsA9tMnRlCnyHrNV9hEA2NvC0xihkoQUEazFuHEadMHPjAOktt3L
pWsxCi+JgkDKQvIgrXcyjGGwoIkk92VGPtAHQVOaPnJakWzuoyCj41nECex0d5EXvS9a9S3YSOvL
iKEO6j2B/Ktwoe8DrdtQwTvuRERx7Q8o70gWTlxhLPjPZKGPqnCHXOIjL7z+hy52dbkz3NN1Lh7m
a9cUBz8heUuazwLQpJ/9UeqLVZlW/JLD6j39aq2voziP/EdiOgXCpqSxKjEExeJRQhbTd2S09Yvz
ZudCOsZGCp1LWSQrZLOwmOFlbKTo8tvRTr2An0xIkJ+0WdglObESoYNd6CtVSpgngc+6Lnylw6dW
kYmOIADA8R5XDkrxHOXA5ia9e54+ORT6eRU/6glFEt+vukq6gQ3JK+QDRX7PNgHMO3edh3qkCNu1
jSqq1E4ykl7WKppwckL3BWgv711bbXRZfOHVgpbTIIQ5p3TnsePJBr6B3lsT/XDnDbCN4e1KziGW
6Wp2ZnHPPaBXsI8ibQOxRmtcCnFeckf5HoAfIR/dnNm10oIwnq2s3amibywtCHerK9qelUJGQyXY
uOeP4TrUeVAEc7ixwO+rGbEcjYOqDw90Alcm1cvJEX4oQ+yMzHKi3YdKb9faM/8//NcjgVTMRbxr
uPQNANe7LBPvv8WWm53Mn2VLYPcC2exjh3WdmIJ7mKnH/QwBLoeG4OR4ziz6c1AoIlfWN7GvXxAi
pyY/dH8ZjVW8sdGkfgGGo7tNLWLUz0TRBkyLtZylYpv8cZhzzTndBuSw25m6Dg5LhJ47VZ34C/mr
P4Mx5lM0fjB++jBx0Mv8wtqeF2tv3Qc+gtdklC03dZTgZaE4ViezC7a21jkDMazor3rNtQFSISis
dxJpv2E/B3KJNa/Rb7Z3cb7nqOOHmlVQyb3mNh2uJlIvDGT3CBe66zXQPG8jVgfqRI57/BO7FTqK
H1o6j0Cqihs6OrqhqJwn/QlOYW0n4uUfYDpa5GQPFhJcnzrhgiZtO71mqQFztgmZhEBuM8iyZmvv
H3afQfqwkPnDenMt8LQlGBUhYJ++XQrs6/II5YpiXqTymxCXFFmhc8a9BRZqmb5dtEYaBTtzZX02
X6d+9lzsKCSTsQNWeocYFeVTaKsq2HE6lratWEKMY5upKQhKy7Ail9ghecR1vZdJXVFDDtAtfOJU
PAUEYIUHQzQ8eAuY7JwNyYvuhrSBriu/v78Kh+Deye1YWI07NaU1hH13n8Fx8IHZ04SueG3np0p+
oc1nEV58AZaKac2R/NONT94rzdBXclyuvnfbD5941oPD9rMTMsX91qwNPBO8q1BLm6ZiN3t6vO9y
FyhyOrY4/OzI+NUoEmp0f2gwcbQjtjBdWlFCy5Ye3SB8eHiNOwKQ+knOH814WhAorU+4eBmTNV9z
eX+4NdiYckt4F7KbU9t7koAB1cNLmYHzyDYogKC+aUFuWRi9UQAoBE1J7bCmap4Q8Rhxr11ukEgp
MN23ct7BLgK4gKTMR5vxaTpKy/s/wpJNxcSRNQyYGqdFONt+M0CmDjpxQqZ+q5XQep/qFP+dv80c
0liUajCN5A6912Ds5NF/S32bY5PfEV419WKU9MEnzpC+VL2V6+CXopccQNMC0gD/yR1B4E2MtiGa
QOxAXSMmd5/v+sgPr5b97HjJroi9GDQHMnwSknhdLZmntL3BF02XdzIKMGYS70i1PQXEKgsmD08Z
ozvF+MiXiG53g3GnxUWiGPQV7Hc6NW7lXFSkspZDZQ3sN+erz+kT0L7OkVi1b+jYRmBrdOryGtk5
Qp4uRWKcY6ji9xd2Yk7YygDMkwPQBunJpzcIFYbLlOa08SL8J0B9LTW0DfMVKBourOrXc6/+ZRbs
rCKcf9fwMJN+CvJSxgxa1s1mwF2ktOA/tyI7CQMoM8ZKr8MATBaMDS1+aa/uy/SxPHUgX5HFpkee
AVF8DgZ+n04pVpyTmC+jADUCb4esbN8XVYy23HqFh4al/TIcuYQfcx4/XDmcHCEZ/9BIJcJzxHyV
q2idPwUHOo3JHgl/6KF1bXGm8DOVtCd/7dROxBFaiH/Je07gr3j9MvXjnNBASPyprkmZuQZKlGbF
2xpQGzcc9xpxofGC0Z4uYWY6bXRKEgpvkuyb32/SOtOImu+9ULd88Sc0eYmzfkc+pU3J1HQJ5z23
SNYymjlryEql7tDeGAOUX4HTx1lE5NcajejL/XOsU6bBmtpcpxeAEDK4suqIXr5EZMA/XY7u5uGD
+MOMxF0e8ppNp9NDPhqbbm9J8j/APAjGon5ri+XlUzWatqEPY2jBFr2vpDEz8bEydFYx9u6lSTXb
WZCcZlfnUTjCvXQiN1EQ58fPEZd1BqqBh3BhBctFubWYxc7YV7degWgoE2JLKUoxjOrFgLNuN2H4
3Ikczl7XzGSalF1MA2f7jFCLVeDwgWjVexUytptrqY560ne65VmCtwg9Vc0etlptmpNpcLWlF2eW
P2d7A1aM5CfrUNRx6WiHwEV2+J/hMT7oUTdP9gWAxNgIhjGz4ESO3kTtVyQoLkW2xIA21jXPc/K+
CLs4t9c04zmvzCcJGIUKmTHYC0GRxc/qJqzVZj+QCPRKpWEpMOU89641OS+wIfuOlwKJh+cB9Q9g
EIA4DFyoXoUBS8fmci3WL3E3kiHP/alKGM/yb1lPVGA9eMxwgU+8SEdVSTpkDZosm7nCzeZLxpih
qSbkPBxrNuOBmhIedP9YwarKIcS0QsX3AcBtgsK5Hseq7d4GEkZo9y0h8EHnh48a0xseNKWX8PQa
6JW7cEr7VRtkQ90qBPwwQA2RMyjdF9Za/+H6GcJqa0y0wKlCs4KuioE2KgkI++Yzokmck7okMjKl
vaaAFM7+Ub2abrG2UdljRSb+xNFq41HXo6VS4bnSBRBPh0n5nhkl5ICSw7tEvomq6GF/jt6zf8rE
7vA1b4xwvgFWCIm69ixylHdPcTHnjtmYnkSRgWSbbQ8TRD6384vxvKtJA+zYqljSUQvhMC1gC67H
iUirZ2hxN4lfelAAFufAMENHiGnxL5r9tP4fMWQYXaORulKtjN2DspA15bY3oEsp7C/z+yRbGl+O
fvU5E3C+uCYSULVWHKmvWyU6b4CdD6T5mHbcSE/aiZi2zdhuq+/f3hxc91Wzpk5NPBNoUVDLTrK2
teBS14ptOfeucd9w/9rBDO6EhpjMT+0voQaDs4UwdgUi5DYeuTifwR/maNdlemC/YIqkLLsLUs/P
GdaDGLjpk7JHS3i7c62IGdibC2K64lZMsLadNwDxn5c7uwMM+Rbu58KRFdF/xt3D2G1KBfdbR8TR
ZeMd7XpYCrS7hrU6yh/l6+P3sB6ogwSFJdl7aLx2WsX9oAYk51TFSzqybSjeHhPnjIDAsHFufK9J
eI7cTBYMBZv/RxjHPIqTqmma0uj51tcGoAsUYmoRQ1YOPbl9NIYiMzgU7ULzXlgpaCl7/FH4nGaB
x/bk7EBoi/k5jLft3hTv9yqLP3CqCcATJyyPrhjri3Q+qodf0l/m0wBCmlgFXFQELYWdGzzUItul
WtjUrnL59ysCJPTM32gg8C7NRLOBXPtlCeTdHC9ea4m5kw3k/FfTDFi/mRyrqnD/jF+sfapjCMFB
ogdReW0PHMECVTRd2bdwkq7BZJspKiD4xPIL0Dq8Fof/gkS28XUitaAUyeZGA9BM9vaGd7S3c6Ry
fnQNddBefac5ykFL76ZjHHRQ6ITLr2o9zqr/pu80/NG1DkCN74QMvhMa5cp4yfiAsCguGE5lr+mS
Zw1m05NCUbtJUzRccbIhhpGnp2rIWmXajrAKLIZ/1sqhtR12MVHaSSVOcxlpC28vATN05aRXqaKU
82lLr6QQAYak5PzqY5YlzuZ9pn9GnmfOxAaieWy8rOch543zAsQI23fDqoxCjRNnPo472EuUslGz
res0PxC8yH1cxdC3B9o3vUz8vL1HeSfArNWySC5czVQHSAzYufhIcQA+tUdee49hmexR8bGtGkdv
vdac3HL9Rh+jlwxnVyKS+ylzJAZfxlHgq3lZY1zYtSRljv/BAJGrh09zofm3pHXXm98uPAzI0gnH
K2OlB49mgRgQ4hznc/Lwp2uAE9a/PelPIfID+WbR8GJqHEFXgiHSJlR1C9U1OQLCpcUNq7DL71ps
t51VAHPlhOLqziBGmGdE6dDYkwBm8KEh3VnLfDAaGBTU6tc647NvfjR2hHRyD90copY499/hP0AJ
h0LPPYMf370F8608EDAjO6QzkzjSdPjKsU1Fh/GG8NyfdKqrRF0OhPTiauji5bPacyLaUu17XBTi
vyLtAxSFPaYAw4pyMg49tS685baq5ilZHfHhNZ0Qve0TAEV8yQUB6pV0oVpb5VQk7xkjE2/niafA
k2dZUNkZgTHx/UZ9b4+6yUf81O4Wa0//jFNXEQl8AgkJd0QBG7dFgAQ+nLX8x9YdlOcWHbRVKxj9
GL+h3h8zab/VxGrMosvpl1pzNsm/ZKWMCgDuqmbXuuqQp+dfqJzdQkXmGSpZ7rnJt/5GXFCwQfiG
NWPT4wgJMRswzHmEl2MAnkm7NpFksZnaxYUIWAliKeZmFJ52SYIEiPmm9U5mezTmqkHk2fXQG3P+
C1gh5WkJvdrUvK2hbj+J2SJlg+Soihvp7DT8ZeGbcYGn49n29TvVLwNkj0/m5LViLUKapFcc7HYU
IZMe/O59c5g5dJQwFQkuBOnu3At/1qnuYC4pvH1i/0rV/tZlzT2U6syXjFNDQRs8WyfPPGdBKb5d
Na4FuCVpIu1L2x5veQCSsewZi5Eh1sFn86kskSYbW4AyG1kUuBAazHz0JqbSMmuhPVy8u1bHBBeJ
+oeupkPjD01zSeVmk2tp6DcU1+Zso8E55K37iFjarcL2wsN+hb2vZCa23aAT286/lQ7hBIkqmVLk
IwZrGMnxy1L9Xc8/SgZwWViRVlnkzhrPUmYhXSLZrjRLC3QU4ZBwMEZeU+zksnoX61A5JOllEgRG
bdv2nweQ5tDBVQP3RhRtyfL6xHg9HR0pyXmmjJpjRQMavR0r5I5V/ahj6e7hFtr93AeU3xtiznPT
Ju3ZA6cXen4o0gyb7pg6K4uOB4AVBmvMeCswQMibwuFmvHETjBy0kO/F0JXKWi1uY0npC01W1UDt
8AclHSPzb553/YdiQ/Klpcmc0+KU1Uo1sfowlLo0VOMjpYOtHvJp1HWieCVC6MgOarzy+IJ8CT5I
JGh7FNz2QmwiC7sKiFowtA7mQHtrzbPq4bzFBkLaC5aVnDvLedHoxiJbTdOUjI4X2C0sDpCPn/RF
LxzcvgDPjTTFv972ESufiPwPx4aJQFxc4gow1D+sOaj+34iZdg1HMfOJQtK1Zn5jlEGSme3AOMjv
k+flvtjWuPCyTD8oj5XCNjBGCRlBK39g9d1K72lOmPqe7T3w8t7oa+DhedtgAhP54yTgQ9K2axII
6+8Haiyh4OskJ92dt6BG7sS43MczxzyHoGk8UTS5jN036r+lQ4Ns6f9GirKsRmTRLzMoK6U+eU++
s0LpI6Jl1Kkw734cBqqYjv+8yWqFxm0ppT8BsEHKOXfEzwlIYxgxFbstaXl9iz1C81PmMLnU1loy
hcwv51A82d9SF07WGNZeBfeZ4FdaSi4XTF1s444YCP9bWa847CkikgAWVOSiho7hX8FTmqLNvc7E
0dF7IJJKYKbORsdZoW4PuDAupgZKxm67ttt0Ivrn+tSpwd9fmUejbu/FVX7qh4YAr+qK6WiuZLnQ
7z6KCdhXeKbBYCZGfqW6OUZWsl1t3ZEk7rI6PHfI9CIotkgU6xoL+g0DsYNXVY+vwOQayWmXe2LD
JUV3DxYiBvXGwkteKklM8+AM1aM0HpxqFIpMXwQbRr3dIxoHtMpFVBNKI5aeY+dF4fe+uE8zZUNb
vL/b3nsjSOJ5yKR1VmU2sahMKVGS01XU5iGNRf2drF4n4df70do2wrfKAIiYKAkIzUrOMVSx+t9P
Hrincdq6hf4J5tQbN3UmcRuM+kxXphDQZMlCwrc0B1VHS9uQxekVs1uJC61ZxjKB82fj2hzpTnCv
nuvRuojNBYlWHv9gTRrV8ceBd4dLlbZjy3L6UnBYL8FRUUDldWu9X6pvZO+ypNqcseSJgUi5g9A0
KaA4C/yl6O3daA9cg95RtwqHhiW05k2xprJe9aeHkRLAOUT/l3qIY/sa/TvL+TaKnMXLzh3Jjziz
8baVtml28go+YMAukYeDQDg4O/+U9PgOFU7HmFJRT1qscNFQRFo3aOrLhJtGsfB6F6zuEeaSWYXm
OnM5yU1NZjKK6TzFmgj30YMnhzY3D4erEVRllsDeDphLObH1mbsF0J6lvd8RAICxGsEEeGxB6Rwt
XaVl80w/+nTfmRk4NVM7OWRDp3+uPfMD5Sm9UNL/viGG3MhAY54Q73vfmoR6vvAcXQXpd4pn3zaV
1UpnKHeqwtzRsjNvogUx+5ZNf9SUxD4UzK+5j71ZqFHjYMtC23by/1uZzqTlRfguzMZzQjaugeu8
FOJBS06yowBwY3VjhyOPOucpoyG6MwgUjGak9wkn15Tu4rTg0RbDmhVHGCs7cHfB1xtSA6J4hlFB
hthmN8F38J1+KUWKwAf5W8XOUuMtKw6cz6s8xOzbtZucfD/hq25e8aDqyGer0ZI1vdIo8Cg2NzkC
w470OfhVuFo3KViSksSDeYFAP+tjFH/7VVNlat/LDimba7BQrdBkrClWQa3EDkEfrv/jZQVJ4oWP
3vlnkPuonC9Fd2JZ4QRokJNYuhFNOJmufYtjqpx+2pagt5kxRbeIPPSQw+ylLwnMGs+ZQcSOi8YG
VINZBduHS/w3xtdbkOOEGCDdlBg7sSf2WfynfH5udr7ZIn33renuXY8Ngyz/n8RM0D3KqkF8+hFN
UVaIn6CKpAe6rvb/Tqs9vxyajUJcy1ImkM0Ep3ImSJoGL9XXgNZWeQrZArOsQSm+rBRDWvWft+H7
ZRqBwsQYEYSu0KVgkRndyexQS94Z0Af6IA5pBQB3KIuYjkiWG2CPmy1qfURnd5XE6xKHSOwIvLmN
SFuSQn36ZcRKYLoNiRXHp3m5p+v+UN2N/M/5hJjTeuJACbPwvn5e6L0TmMWLAOyHHxAYNH6bdzUE
RDcJnn3ieajFG2A+NBhH9POOyqLGoEy3iQETxl7561Zv9viSCHAFilDVeqo/Emg3OfaNjeQi+HXB
m2xNFnPEJY+bqFNIwnhTl6pZXV/uExx26mHwY7P+tgGIxjjgE77wnFfbyAcZfpcAVqfc7audaYE+
1Dwz/ejfH/RwCtGc4bDq5xvT18MPBmktMBPlTEDCb2HTiukuPB5qW5E9lj6x7J0DKaxHZVklfUmZ
VrSrbnBAj1XXIyJsHjurTamKi25/koSEOj/qeDws1vacRwmztu5xVvg+A3fHKiqUMLVk6ElaY07a
qy1ddSgmTQLhAJTH0V6a2mYD+ADvuO5up2Sd9FjHbJHoj0JbCXh2VKTlbji5bdLZl08/bdMf/dHl
AGh3JgRUcaF3ty7YF6T7E1XcnwjUfKZJt7YFjJqBHdIkrH97nAQI5fBDt3wydhECDK1LofwCbgkn
xRZDo4zFpvjwsGwMYvXAIyNDfOgj5GkjBj3lfbRtxZY2H/ualFzi7i8/eikfK4sqWZUREFUZBdY0
1XArTqr26NvIOjoKNE24eKIrT6ERmaNF5LAKWudmYIQbD0AychYerQJM8ONDEb09DLf55PYlEVIm
nAK1eKlh+N6ZC/oqKTr2a4QHdeXcj8bvcGHl2gNLhTYLlY3Qd3SKffuvw7sKLZs9T+FjKcFBYeAU
pHXQg8vh0JjLA1bzsS9Xwk32ubcMzcpjWJ3O5JHuSCHrfdQavDBYlGU8KIVefjz9atZGFiU3rHqe
tfY6oGfeXUoF3dTe+cjavFsELitg6d5DeK+abZFkP6UVA3ssGnuynoOHBwgX1oQHEOWzwsydCMgI
fjb/1+DkaBcAqE9Cr/9+85aDCoGHOlol8XKNrRzHEJcZB/4+aS6kyejEuud1ib0EXyqiZxaXCj/w
3bDklxwbsFzU1cFyq0WObT6vJ5VpdHa4kbc4L9qEiKyt395LGSSgsaAx6WEBJj6CoDn5dgXru3Z8
2BC1mEbN86HmJMIgpLx5WuQWesvd2Nu5QCGapyiDyH58keLQbc2s8bCVDLVqr9c3LgNpEBOH5m1k
woMgGr97DNTqPEH7rx0g238+nDWfoBFuw8b4x/dziSFbAjO8CERkGg3hh8tS0d0sMkal4sVOFLCq
FOEdfSsz07zj4hXrXNJX+uyAzTJYZm2i1GLRVCLG5z0pIDqzHX1MOYdVhMQ7+vKLzTo3Gbk0Bq3J
yFYuPw6jgj1hL13is8Ks9ZNj2bC+p4co4/pxtPpzxjPzq5NqZeD2on935c2HVVyMDeVbVAh5GxW1
IfnhfSGf+hBaCNY9hzUGUIgg8B8zURo98nwrlkP8mwVHYb3zA7o4T8X58dc/l/zLOW0msJMyIIsB
Ba5W4q0USE5oEHnG7BCjYDJRl8sNXlghiNtIH/BmgWSzLr+E2Wj1o8TsoX4iJ+A/eCkrRETjhUpD
ZtBIMHdMUx4W8Zqq17ph9+4x/P1wJ8qkTrL7IMY8ZPq1iVPLvU6+Yg7wwYn0XZ4/S+fdv8SF88do
rN914crNvLfMprTlVHAqvyHkv0p3DhZZAV44QAPXEUyBGCApkhzfR9M6VCVf7P8mFzzQocKHbOP1
cUKPtqcgquV85byueEDYlPe/v1oxfJ7v2Y0cnN6olul2BsP500vDiZPbHFrvrfM1OuY9zrG2hk1j
Btp0tEbFK28Mu9r5dkuK6d8azzUNSzfDYzCjdgMtySqNISPAX3uOwkMb4tTKVKnCHhPF1o0XWP4w
10RLaL/c5mZXpNDxgkaFzgRSCWU7gi7cy2Iaidc0Zm89ZcKo5jcyRXF/0CDfnse6JSmFZNta0tA0
noj0NWfMF/qMSDUCC+ZNuiz02YKGe+UjvpfhxEDtMbK9tHmn69EnScIzmu1oFPYmfUz3LEkDxjRh
YT68kdKdn2XaE1nC3PVGig0caqvTt/Q/nq1BsNKVmuP49mgDOBzlXSO1ZJWE5yPSwfee1WiMGVQH
tcnX2IevGtNk6T3UOacyuWS2lqs6YrxBcAHvBI/G8DY3ddxi36P9K+y1mPNiGdUGR6jD08Xd4qoX
wdoQO6Al/HWQnZeedAWvEtZYzk1RoJCTVI/mVtURuK656wtWvDc1ECNF88m5p9SmwgLAiNpP++05
9WIrI8gaYr7nocWMBFvo+YjIDS4/C7jCzVqfu8TKrLrxXgCBK5XeZB4gZDe3KXTGZ9n/eJNn0oq1
Db5sq7vTUT1HQm7hVkhjG2TFZg8A3K82qR59UY+6krIrbC4E+XkkkRN2R1HWV7ftanZqL9lK2lEF
tcR13PT5tJn6fMhKi6FLOIIzf7AiewO+PjB5AsT9qWzkKoAi+YlcqzI5NJjEIriBvWe3ZZPisvCn
ncH/BNFD1ArfsC46HWiMcNKldgIroHQMeMHreD3/AyOfpgTRBRssGozwhPx+FsW0f7T1bWpnU4vx
a2o2JhINj5eSWt3fr0UFDRM9eB5UmHmxpltsE4k7+MoSVa0XsFKvQRxdKyFWrhWs+E8oeGnuSC8I
ISwQ7oSaWYumR1zVmbl26fTwXzMBn681JQ8NTvQHMP2Ec+/FXLXwzybrvgeB/53CRCFuQLn6Topw
hJNEFPt9kfOS3T3u4dKajN81d4uRZSuFCubRB13FsE3asNsuDZhJqds5ABK/3e+oYRavPFIklQf+
GFjWnuGoDatfMSfc+1GfPUyGiihzsBG2J0Hu1MuuErenEDR8p1RiHavDSHvhyt0QBIZ97pW6E62C
CUwtUnItwIdpdjPdTgZEupmfy+tXR02zP2WdMlNjK4xWBJi8CHzIXdbHNDqpp8aYAm4qheVkmANX
XYITVjWkhGAUuPXkFqysdoiltfwas2PkzU00C4RnR5LxUUQyDGPMTiiP9TKmBV/47AVY8e1i8LDA
YZkleYkslJYQHC/a0iquYBJTdUuEVgf4xmcUREfUdd+KbcOubiKG5AdZd0tgh6/I/fhjVdX2Wg1o
A5U5NpjoCPijkzu5JYF4VaiStBVHp4wpU+yOYKr/Su4z3+ouXcQNmo+zFlurc0cVb01enBsl5KiS
+MTYlBSOwuqvrgbsm1Zgs2LjpFxSadt/ukm52V8Y77Cb90ahrHUNjRJzbjUxKlswJhXCxJe/ZCcC
PVdhvln3m7dQV9hqinlaZth9xSZDLI4px4HL/d38Ozs3mMUvrYr58W0sVoojKotGHI8N2t2xMIiL
nlK2Q7gNIMhK8o26t0DvHx9I06LM9OAx0r28x0ExIV7Oo6s3iCqHw4lV73S+c62LoNB2N83xDUil
jtQqmZO7f/L3sk95NGhBhdsxRqYqEkEY+wZGFmlh0koivQwzGsrWMrwXc93C8hGHonxacjs0a4SK
FsTxW73NRgFYTVVUsPFX28xLlqjen73jYefFtJ64hQTUlaSR+d8QPh5tgqOz3D2KhgVR9xCuSftO
tvcDeTkI7XpVJH3TQ42si2+nZfbngLGxbzTwGA4NXM0jW6nr+Z705lAVvsCzIW5pRc8W/OIynrqe
ya8IQct1QOEwnkmMCTymd2Kv54CGOWlVf7mChY83TVMyyUzfRytXyEHK0mWalw2pfopXen0Ik1nh
esjqp9Fe8MAUn3ly5qXEF7EvC1hxqozQMdKukIbahOaP3YtigZU2zfF9xONSuh/h75FK7ULR4m14
iODti9ysYJU3T7C3R5PVd2zzVr1WpBe44CwA/QWn3agq3gDb9KkVYlBsZoxyfbV2VbncuKmFdSDS
QVrbOUmkBPjXRIYRx+wAZO1QIs9XqDA5A1lXZdFWwjhjObjDcT98Nmr9jzYSExdBs0Om+0W2y98h
D9+Q3WeL76h+GujtqB+55pdSFACOlTGt6dEzU6qwA4xjbr3vjpqy5s6Jmdg8eeN1Rfdx+Rkk4uD0
3TVw/xVrS+KZiu5+A7LWbL90JAj1jZUIXowzIZKX8K3UW2pQM7W/yjFaZh3c4WrRpNoZ1MaF0yXC
fprwxveH3iOVxvfMyzfwv4Uayb26kZokqCjjlP85u8CGadilZLSl1ZFceaDtNvI/msjvD40jHR06
D62KcQFdzwRtLghELGKi/P+wwW9hxMB4zun3rfQa6rXTvbqF4loH9DPe637bP+WLfD/cD7FM8fxC
WqGIECWrIPpT/S93zE0xQ6FSqs6LCRx8KXy1yXFCkczSd1Xt3Fh7K/wgdmteRQSdFLWpDk9I/wYO
IhRHp3yqCA35FkDzzQ1ixWTzgR6yKeSfuJYprzxJRHKsv1nXeo5QAguxx7Imx3W6yUEk/sveL7OF
TFpSLXY3gWZ5IycLlnyMQFFG3N9totElwlD+GBdmnNnGx6XtmKSSsxP2wgdC1dQdPE1xhHKv0dOx
GQU1t/KD7+FnW+bC1+CqaL10WM/u6Rt2yl/le96lHBdxm7BNBVb01jr03hCV7wxpFZVbPA57aBVu
YBHsl2gvp+Ir/5J0bBrINKy7WDfWkNoESGaZWKZONO284DInCX++5y346kd3tuhoo0YKFcqiO9ly
t7XUJIR2w3kwKNA9xJAfozAHeCYRWPtaSdFohDkPR8b9W1ijelsIGrCb62/6+kSeqcLwGrBRhUF+
cdhysYHur5qhniiAEcdtTSNKv+9tyPH28Gy1qAbBG4S11AvP01FSlno+4Rk4SgLjgUCk8dgaSjkI
nKFEQHEyrjLruDBqPJgeTmuA2nqADLACPGgDKQEjvzYLWJDyShY3Nr20pwhjja38s4Xz1n9cS2K2
5S2yCMT2YVarG1Ut3+g/hSDUFEY8n+b/aFvGScpE8fpIzuKi0SewDXgVO1aPUcxCdpN4vQaw9DG1
kfzae5tM5PoTaNeLq7rScpnVoLjz9Bq3YmX6Dos2VW+tAGDtgmKli9pHX84ITLPIAiWVmx9OGCQj
hsBU576MIl3Jq654wNQaRe3QR/jaWy+yVflMdDgMS3gWzFdEEeZVM0wVo71Im/6vX1Zj1WgB4uS1
le2v74NDeQNvSAc7KfkhVTV85zuFWYZavIxLHhtONXm5sOFzIQrtrYHFnxctoiUL7YmKZn3hmsGw
qd90E5+HO1JssXsvL8lbeRrERHMK/DiuKeIUzxtqK4MRc3VFma0k1iMzP/5QMoidESuOUN7VleXA
qMT/RwYb4M5lXWayAhzCs6xZxSEmhV5otIAsz3tseaqpYqwP8XuVyJdf1euXiodSeSrOXbc6bPZr
HuezpvFWN+u0u1pzHDEsAtualKH8LlMK//tmu1c7oW5XLJZ5V3iBLKVYAcnkKQe0QqRoDfB/ZRwi
fOIY4W0MrSl7gIpblSz6PXlXd8r0HkS6l+haWJRjoGN/vUboxZ+vK3eiBVHqPLOW4Lc3/gXus+Au
nqIckAj+BfCIW2WwTLK/qHaUfQgH5smdf/5cCo4QVFGl/nHNr2JaGlJrrVOcQApKMpkl0KuilQUV
6+yekzG8cvJmfAH7Xjs1kFBGXoE6meeZMQo7bbr65XC5Q4ClIJVcYd5VfWYu3II5Q0TNQ6UVkGWA
FW5epNnaL8XajbHm15Y21eI9A3WQ/4hvXtDy3orc5jYgfc5F0UUcF6+bz0dWAPLr51IdJP29pHu3
y0FQygAjsgqyGtJAwpjI2eZn+pnrmi8Uori6ZqdPdVaCVw6U0mmlGkbJrJ+PScERdOaI7G2YflIU
NMCu2CSp5TozUk+IoXO3UFqNKhb7+uG9Gu/Jy4IKil+91RfiyHZBQ/374SnsjzkYZ/ZuWiN2fNAl
pjykC8r5rbeNBmeztBXaOGcpcCCWYJSOcJWvZsD6YMJMDw//bkx/8TQRsUsedYaG8Kqj4imcCId2
qyrMyH01r/zj4X65zIqlpHdeIOzW1SO8WKvOI+YBdAlYRxvnv+Js0o+d4D3exrAL8nMvRRsRGQzj
Rpr61O+qS7fL1quoVTOiu0SYMrlyfAahdy/S8U3SsAmqPoh3Ad3Y8dhBHbghBNI5NX9laixKGO0V
KlqW3WYTdV8yv4CAYdqia+c9a6CkATtMbVsw3SK0sr0jwxALNufHLRGctlnbjcm2ua5Lcjk+q0Dm
7jTMZ4Ap9fwN5MbHy8WhS+6gIr//LHkAUI7sj+XikWymbG9UfOiI+PYipKC80QEazMv+m3av7tmZ
E8mWCDC99CBOvPDCBO4JjLaagLD0R+C4x/SWxz3AUyyQMEPws16wdhCHF0m047ahhBW72BaatIId
L+lvPkvYK7ivHw5b9KNQVz8rKsiTgLovrovsdcgFCvdR0jslyq6HVqMA2aaO+FQaVbSi4aD+4KOX
ZojERXdyhuUtecTTZSWEHyklVNoZaDTqsJELjSG+1GmR4JLMG7WYo50wC/DJ34gWVkgHiBhJ/Xl0
uhTHAJ4c/wpFnp22vksxed86f3CUF6vPl6ZWd8OotfMYx8vzyS6N5iYcbh/tkTiJo0DUH+SJAvYh
dHKSWcqZBBn8XeADXTI4x8cpnMiZtwjyoPWZwvbkAsGtmtjJ40vE5ffMoetcftEvNuGWDWZtxoGp
6XmoRJS6i4X/otv8w8PS7W6AwJuuFjWPC7NMd3aU8hMaGu/u9l4mtTavEe/j1z6UDyRjjoQ2HjIb
125dloW/w4kMzPiI1BNQ3AXRDVXkiQ1gP1lvfxnZCG7VbXT45An/X6bQyfj9fSQLSeNGUWg0cdUX
TPpEIhTB7gtTjHAqbU5nh0XRzpGO56B9Uodq+ZHqKvVYzgpm5+ZUi9rHyBvn9RkXjIExGqZtOVzN
1MfWfdjvvh10bewUA4Tkoi3WhcEoTnF2pu4BKC3n2lMymbWWkeMEsmmwmFF1h8oXpHzX55VIbDGV
eFR36Qht/AW6gAvStUvpizdExchOfGxmzltB8UCu5KydS80kOeuQ8VZoviEu64G14KtkYRfLne4R
aKMwjRt68ItNmW9LY5u21cpO5tBPbokfxcoq6O2w7oUhufXKfcYIvG8DRvby/W85rtEJN+bh9s/b
jmZDs2k+U00hFoM51ayuJvmtbShLfszQhBjyAYj7K5IP0Qz0ggMkSxiEIoF0KXCIvEY6emdCPj7h
3aXU4GGyI0HePEQCurM9oYAgJ6cBhm45kujtS+Yffh1vS/gl5uz87CRACIPFZFqne8b62alO2cbv
6bMvZqo4LsuJSQTNFQ68pxEGaX7/4rrP6SCNiTyKoyiAVp6cRZk+orRhQ4yAD7DAUopsRb8R7W2v
j4ox4PiLxJjGRAm0md85CVEQ1mJaeq5R+AdMSWcHMBSIJRgWLwC7GtNIgZtgfIjtjxj1+bi2aEc0
KGqt4a6xPMWQ5EbjN7DxmQqk9iDemlQu4EiA87MYp1Ll5Hp3lAL8dBxniGIHOXq7T6RTq3gq5ngB
98DvX2iRqCTynGRN98q6KOWgLbVcOdzyWX3Qc4LuJPieZGOQmCl8IKyefAIf5UuBpnj9Owu0leuW
/oR0FLT9UbGz3rwQizyNu2Lc2Xd/RAEPg+zya5gHfZEe6tO5W8y8eUWJVpIukpswXXS/qky6kEGR
/z/aCwmxI8vlY6H2An/QLyUWJOyiHIFbxG/rlu3kXi66hlqVoAGStMPR6+Ttl+El/lym06OMlugR
FwCgEMl6DV2FeYEKBbi4mbVFnSzRAwCtWZ8bydjreg8aiYlg/p/zU5xqCQKSmXvJp0WdPClWQx2k
fj7mWJlqhUjNIoDuM71kIGahdeICakY6XfeJcvH5s3QCOJU+kQHrGn1XAXB9OHkq1F+e4yvrT4Al
vuYWnSTQQ5ZuvLCCVVreyFe/Pv27iQAiYTRyPkh0AgqEHDZgxgYjpwsjf1QFheQNRHBTmKNJC78I
rFo4LrJ3QuR6BKbMq1d4vISLUQZaMMEFqgdDcTg/H9P5RaHxpUZIXlEaOChopxuABenPBGmS8qwW
OoQEo6q4xwMt+OBStQHQh3hIB7VpMwMxCLSLVM/S5azEgw/HWw4XXRiymv8inxf7HqAU4nVzBGyr
EoAhuIBLeh2UEzef4jozpCzxWvJ3MjE/7uJZAWJCVt6rMN7zmrVQy0PyoeaiIUfnFXoDSMS6AsF2
WGAU+HrdM5i1nwiIv3JHkWjmDOzoIYozFNwNjMV7HUPrRjWPcmijASOTPtzh6+/bUUJsvpoiOBEW
dqF5dnhGtfiu0pp6iPVbtI9zkpCRKdnGWjGMx5GahAlhZJEOKJXa2Y53jac7m3TyhYdzAxYkymqC
zYgbZLwguxQsMs5mzQTpix91h7DfZq3AVr3tHdtzOvS6H1eVRZfZSl8CWGeTAR336vbJiLui8s4x
LtdhyfljJ1L6I/ZE/OHvqrztJE6SJClJ1a14pd+GAuDOq3ViQHubuzUBzv5Y/lvnUzSS8C+p0Qci
sRjIQNfddj+/8QBo112G0x7E8LozA7VqN/blRkQ2Mx1cHvr0AfmY+ujHOj4xRHfxIFGTwlKAXU15
Sm85svCMxKpi4AFl8WLsrPxA9kop+r43nK7/1BCME5PlIUemIikuZxzifeAtVatxdP6UqymleWF2
oyktJplKN8NAYXET3NI2VkruPpLLIgLC4lOkg1e0J4nKe63gFaDyd+mpGzK8rG5krWfMoUgwXerl
aC4n4zChO7HRYz2tOwUCsCbxH9IAp/XKux7wRLTSgW+F35W1gKYd2QNsl7oDjU4vRUVWO90wLQi/
4qklpxVqa33seGGdypHJ7bIHY7EEPn4aDUDVXBxyUS09DPmzotFG68i67NcGHY2VwXPWkhhL79dS
Z1BF/SA9lAL1o6BhsWZibke2imOM0+b9pUqUzQS57+0betxucc7MhMQhGnOM7B+6o+hfl54NdHQC
dfS5MQRHwbYS2HrIDzS9XH3FyKyzvosSn/e3N1Mnpj7th6YPyPbJVx0OQa55A8ltqeoozd0euEVr
/rbgnfXVJ2Iz8UC1fZtIwdHYOII3uo5UwhZk3VKNenJ5655j/PN2Sx4GHM6M4Cw94l67L4NqO/bA
EqiFxaov3mPJ9hUs49Krds2j4kwppg8KjGifvRehFwJ2nKrOXJHgZyMvsXMnrKe1dwjmCrrPWtBV
x6bol2IC1VQaY+PklxopgTa4RIkWq0bVByf7OXKnBAS4nezJamqk6Vi8pc4dg8lLBfRBD2iUpf2l
KMko4RheHMCtXB1y4sKwQIFt6uXWbc/KFzy2PgftYb1uX0vZH530lUbA/U93p8XvvOS6nUlhErOo
XGjjOXF5wWXHdsuhiAXQRKs6abiXT1xeW0foGFiF+Cs9ZQHBESd0LP+z5RtsyXIieiSsjELTAWM4
7CTEM9x/aWP9IG+MEsD/t4Hg6K+250djwYHYO/ev3LgG+/818g9omiN5nKr2bJkui28Q8OTPNCIH
iKr2Dasp0gNd26C0IJg8536NFGPl3y/7juosFvFrPRToMdyjP9YhGviewyC4Njwa2LM2tREQ9aY8
SgOdXy0nn7TCbGryAJ4dSS8XUjzcsOH1KbUdNdCU7UZ+VsGbO/DGE6Qzqm/x8ioooAbGlgLYPvxy
O9hMEMh/Jd7LilNS6oz5Cx+7+lO2BjS/wW9yEMqhTTHcKa2l5bl2Y9EJtZ/IZ4Nf4NO4xETbycgS
jFOw19wDXUEoCQC3XqPDuV+bnHWI6u1sgtCEQitB042wAtXH0R7xp4Agi+ChIU/ErsFfIalS8ccd
WkIQL8jL7c+qQPbpA/CWSn1dBfMFNUAzoueIiM++NAjF5sy0orjwRwVwF40VNHF2ly3ECUUVe7zC
RKWDBaEJAg/WPOf6/ae4WFWeti8R8r/yX8A9h5FUKObz9wUoXF9aan56xyH+256ziZSWcgkFqcDg
0v12MfSVJNLSOME95jDndxfKIfG9MN5G0detg9PHR7NqiKwJM+JBjjnweLwE6p+pge1Y8s9iybBn
f1aUKhRHK/BhkklgZAKSPX/EVgM4a3J8uvU0j3uu+nVlW6uuZJM9l762V7mrlBk54dV8CKxP14Rh
430Hvv++LVmdLkac5P6hAM7jhhtxh/gj1NpJ3pVOt+E6xSwgpqSooHQK3trevFX/crn5DuQCkW48
4QxYbvzjSJvxPDPB1VlKnwDoodBLuLCSdvUUAC4zjOQ7uGL7+qzxNFQivQEUkD3o+fuyK1XsQ78i
aUDWoG00aW+wkhgwtwRBiNSSSetve4HmQ1iVZTD1Czdg3tI5B3R+E76pFO76u6Dk0bRaFjGW5vHb
G8ae8cHSptwl+Ll3p/DCwYyfUCHZPAhSQgEHIo74p9be9AiNQV8WMQ5qUWj81My9FRc2WZhP1YYf
zp2cUl5C3s+dAITxEOLAqBstEOX4TIOdw/Qpo1Xvoq4M2lxs3za3RG8VZF1IARXizVefQHW9yOfl
vSOaRKCw85SdR7z0Molj4RoZNGqrP14CJKXMKz6fwXIN7rTofyt/8zaHrkkygOkzMg9OVai5O6dw
ach2KldGYYvbUshq90i6R57drSf0PLAq+t1uIhRT6yoH8TiXC0+quKjA31bkMuL4IPCg4AmlMegk
6uxsk9hLbEQdF5xYY0Y0SpatTtYqw1oHBWH3KhKyPEKlnq6VUAYLZUEBKrQKDFsPyaremE8YuqA5
pZDaH+hHW8aBART4XQN3E1ayDzA+CG6jJFK7K1COu1K8SJRSiIpkonncHf1aIxq/2se4vztcUZxD
228p4DW7y7BOlcC7boTzBGrnGvmNp0+TlkNGUZmC6JxPytG1edo34saFvxP7SoZhG+iYlC5dnrn3
jcS7K4SpyTLzb1d1N+X8neuHiKqZl3Mi87HmAHqrO+ns7kjotcPra4Qc3tre8mRbjnYYqFiu+5LY
4p+MvVI0ERzwKe/6HIiYtmWAp+Hz7B3mVdknzZHrQVAcXhnvvg/lH33dv9jXCnRBrvTNC+wO022e
/0/q5o1QRv7q53DAzMPOnixn03ynpbx5DXSvzRnvec8CwLKHKHj/Ig0hz/UQEFf4RLh/jRAGO15C
mMLQE9U0rVf45qf0curxd3HCWBuNkQ5Ki44Nq6bMjuKZJ2sLi/HcdCUhOIzaEsiXaa7K4rFwZyUS
sSUyvqtBAAJGtw6+PFLxDWHn5bgA2q/H2TId1093OTGXked8I2nX4A+wlyJCIq4yGJQASsFJma5s
vu56YG7vqXrZ8pHQX3l6exB9c7HNPtAv6iL/UB+2jgqeGJJeCk3yUxejPJKtDodMBnAxHXBjIMpv
P6cszhKdP6mruBKzlm+BoML3pSFH9wk1kycauLcWU4Hjp/FLaXctLMNn2WurD0dCQRJI5++wDB/F
LoA2J2KsQrtq4m7JrvqdVHOJks74sqoFwx9NtvFrm/NGl82gk+KEYXj+RKl/Y26ZCm2w/Q/5H4Dp
X+xkL5Y5ABvz0AR5VpOOLi0OzfVCbDJDRQIoHgLPXJsIumxDiPdvLIyRzVqxMsgENHnFn5xS6zDY
7HX5qwGQ6Bk0AHegQNf1gxu6tosvoPqVbScG9iz5BO32M7J/Zq6EavPnRtXBCHFFeVWp2+rScl5e
pXahL+t9WGNkQT1gpOYl1/ie3kpWdSt+VAEbd6UsfK6EtxDHvRRyuRhHRV2DbBDkgjGCBuPiieDZ
t7re9JOxvk1n/qylQp1pOC+QfntxU6uyCqY5XxdXRgI+yZ8+i1qV1pwM9N0d+oZvmI5wjxWSwXDO
CFsmpzY9Xu2ILE1XxC0k7NzCGb+KI/0Hn5sD4B5TLS95BEbGMUxahmSY7ZPYl31YywZPcvyPkc2U
ZkZehFCQ3wzfJ39Mj51nrVjGt8by139EMZw5hg365PqA6kKiY3FbTQOfGhsIpm3A9fMKZgevBGIA
JcJpcuKY+s66lA+UyQgYAEt8UUpjPdHackRXQnkeNQCsq+CYwLjeBGTajlLL9t7bKvXK3KZtm4Iy
Bu4VGYJiIjxyqrY9C5lsA3fUj3gZhUskRvgAX3sjCp/zSD2tf5EJda+IalTjaf8jq9Y1Ua9USWSo
3ZGnNie8RNOUSmnTCQoyktiuEAcjyYFpqhWenMoD82MRufdNbmDA6LXZTaY7ch9dnTCddg3T5aFc
GbS7tDWFr+moFwJUWH0kDknBsbLJBlr5xV3KkkhnCovLvo+ByNWzfDnK6QOfmWciTm1Hpl+kL1Fb
rrrguooq5Qs1wGawv5AC15VoOdcVkpQO08GHfa4eEldCDo4BHppSRcCnLqRkkUtY0vk959zZHwgH
MCZofOwBUbq2kmm3K6XJA+QYihQ4gdBfEg1Sk2KmxY2JAJO5Nvm8zGfb/QxI7dx8NM7nEYMeKKy7
poSl/qp/ysG00eW7qIjQuumHJ3WoIK+8g80LyW0Pl0/sUu21msGdLQ6Kp6rifNzrkYe9+UiUe15/
rXBHGTNou5bq6bm2GbZ1LZCr37a5jQPIPcVCECWhwNkuSVRalAPeTHpuBJyGLrcS+36vlcZ3eiSV
vr83p4pGVkVypYM+3sNzVRUgfV6oR1GtzfrJCnGB7apdVlQJmAu6SZGsOf0BWlWCEnNus7oE99IR
GrShEBZhsPwcl8UXpOIwhWo1QBy9evacTHgsPtGt8q9FQpYLExDHV6hcXkmNWwY0yFzvVMVsvYEe
F5yM2BYfgIT1m6MuBbcMpR/9IvcajDbSH7lvF594dT+I65706gQwIxImQMwu83cRTBHyELNkCqEO
hX93puqBQNpXdh1KhTvWkUWsD82iPLLFjpJYn2YBr+MiqVMCq2hC9x6+EoRrbq9kD7nNfg6cK3Xg
rVnPtv8lKI0WxruS3caLDPgTNHM2SVh2VCdRQIjxV62nd+T+rOGhLz8iiQKqkg2bJOUgdiyFVkJi
JKPPJ3pXwzhAuTCzFzyfQR3kaHuzjR1uax7BppxdKFUzgTtJOto8jjq7iCuG2+8mNeHCkyAKc0Z0
BVWEzfWyILak13F0siR+n8CJi6PudKmrzCHdVR8PPtRs5mQkN2eyi/TTFs/z/X8wChbMMKtiqJBz
tn/1gqvoaAKeiqkD7p+kfbKKV3XpkxSp5ATnjdyQROpHXevUMbnnVb2d9IgRfw2BH+a1SheoSuOa
8MgmyUoqTmvqkIrq13jK+SwqBQ++3cmzbHICCBI7xptT7EJHpG+yU1x59J3Ktfw2Pkqiw49bUUYF
vqPO9wgYEfvKIWyWwhn0oxVD9XZ5RgLcimww4O9RRhiH09gbOcIrwfAZvRzq9Ypb7mePnIr4JjHo
18SlngUNCgrmdZvdId4k8b5IhvIxhoQ986bRspxGHvzU0eB7vlz7jm90m1EVW1kD5tSoGym6072/
A2TRh19swTB2VKboVW8qegvdZpw/7KeuDmB/eDnmZ42ONLtMeIKjEMlZ0ir+IL/EnAVR7fnyBBIC
gbpzVJqY09CH+QGLGtv5AJwGUZCbHxGR6jXzq6w04VNwmpgPxjOL34p3ZIqyvjEIjEQGMp0D/Kl/
80J40IuR60LtVvQRhFcGjE5Qy+L38eYeVcXhUEnbwwxzXFg7sqX2zzPkwB/GMqFw3VItQ1oWenpE
4S6kNPZdoD+cy+4D/GoJ0TsEqP9Vcf9S0f6YBnhbWNBWYH2Ri+WGcVmxEPjNXF+PZdxyBtI43YCs
1+SwOIMxbdjb5AiparYEgfJJ2HMp/eq9ygVysAD0iBF8pRNRsTtvTmwCZf9uYXSLu2P9JliUCWlI
+tK4cV6YJXFWr2mRGZANvFdNQquivigIQc9jpIhQxjFh6EVVH5VFJDAv9z6XxqdAZM4++3utN3ZD
8yAHE9bDI5vDEk+6IDPT4hBOLpqLy5cV+9r1i1SBbhnpkY+cFnAfaqrYTue6Q99bO1HdaNdsSbjN
94H8li8TU36UcL5Kwc0ODIzWsd0e3tvqk7fv2fvtQGx/4F3yepN4VEAjy0iFEJvJUmL8eZ7C9JRz
aZ+ozRDAe8Xk/kqE1wZsOEnkM2Hv28qQnsNn1wLi1or/OPsfALZdDfbVl8yDwejL266zxgzo9Rva
33Dd3j+QWmVDfPAX0j09dLRKPE/9eyjLmLth7C+UDDgDBYu0Mp+WHUcvUx7TJUAyKMBaOSnArfXF
mtYlZBbokeKl9nnwsoMCnORa3ivKv8xehK1OuWE089T8sqeEicVuV9YyFxolxa7lP/ZhUtCe0onN
u77LypxSKK9PhYBgn/oEhUJocBGM4TRhaPY3kE1sngEeKMBmugGSzxmt4xdKkS7QM6C0YamHIh8T
gV0GXKOkRFRbuz7v8TLfXpZHX8EUULbCi0WgC40wih3Rl7YdJhw6cXOVH8gKJuLcaVBjoMTmw3GZ
YI0U4gl8eg5BEn9kNj0vUpz669w2oswUshI766YAWxESIZkP2ZtxJPOtKQLQ5+p7NWBmB0k3vka1
ZZVi3RRwVFVWlT0Ukdj4dY3XDch1oiMWHKZ9Y+qTQ34A136TxWWmAigCn6YlXJ8VJ22H/weGg0tb
zo/1tbnDPpw6eUAoiqOI2b3Fi3Ifm/J59gu7lZ3gXH/f86kQaCnFiX/tj1/YppsI2piQmnYUP3RG
3sr0B7KiekmsdUKHHIKoezvx8Y5QAbN2jpyDUfaSjvALTUEyP6sxal2a7dCksRx7u2a/aTNMew6E
2/Gw1om6ju5s29W7miwEoVKCZjJINWq1+Bkk46nxypkACs5T4j+RNuQy95xnPB+kgLbVGQYyjn56
1Dh8TW9RRWrVmm0sCjOYV/CVjJS71kZjbXtmR7Z5QziFm8693CgqEuYzc3b1yS2N8EF0LQF5BTbD
8JgWsjysPq9FwPlL9N9qqzmu77L0hFWAurqHBAl/+LrSrYEw3EXUMCcH3UCoAPgc+V6cFv2J/BkM
s/ViWk6uXpkDSEPq2g6a2Y1IkRggHSZyKqO8uq+dF3hNbIid2lGFAecaQPudPe7ZGUDsAuqoce+Y
wmxpWJL83KevAOHM4nJihyeUK7d7z6NK/P5awtr7l6cjN5emZhTSRnnPVpjt78S6l14ca/GfJLY4
SOdLvsb/Ez32Aa8OU7JCTI1FyhkyDMpFoHlTFTFshWu7LEtIP2TBkbmBnPznsBW57pnIE+GFpmKZ
NEC4Hs+VisgLorn3lSscwmoWIPFxJTdhoThUg3fhemC9RulaEegwU4vvyFxKdUw6etZgFEH33ZiP
S46WaRq/et29aWbGy8cwhWolDNJKkLeKG/ZsJyP3+nXfOiOenDCob3WkliJq1i0pkJBXBKVV83oQ
UCmXvMU+GsbRpEDKtcUQdLpAXN7q8tyyPQvp/E+iVmWQafyQsOhG79jVnwwjTDPAR0t4iY6bEDe/
EqtcAy5L7hZL4U+TofJChGwFybRkr412Tc8xDHNj9c9JyDnTciRb4MSSGptjqZJN63yk+IWWT2fd
n6JGXR6jFUg+g4DgA9Z5F9Rt0jN3HG5+XOo1GmQLFxxY4EpUVG+D1e0h9+bk7edhXHcrnRYtZXrP
t5vSLKrKsmweJ7Ed8RYg3FO4bGN7IbRiFQmrmoXBDKAJZ/IKxSZW3iCiMADBPgiwEGulA6oo+IgW
T+XfQlXAykPyMLYsaDDUPvXr4l9scKxjwUk0QWiDNzBWhgQEZysy3efnJQa2UiaYx7XSV5ywI98m
kGHxd7EHR6PxOwmFzWijT3PZuY3VVODJki3m83XJ0651Iyytp1B5Vxxvo8TdqsDTdsB3odHQ4ybn
/vjl2wOBJJdFoKaArOCfH2kNGGf9KI9RTK75SGy0cBOB7l58g02dLTIuwaC1qtwHeGKMgO95Jqsp
JEo+jiYoripRbKpCm8/rtLgO9HHOEPXXMO/OlmXDkNcKQkmCYoDbjMGZlGbxNWD07dEMHUTHgN13
cwoZEMLzPwXMGo2wX1HyVTpRJ/aAy4k0/x7Gf6h4EpY8QCBgKT+zGpCEWZVNyrY+ogchhVnhLI/7
4cdpqt9QIV4SI75VUrukAehJQ4+iwab810nVlq+RiFyuNnCzzEjnK9gEfiVNEyyYb3KpZqxdd1If
iKThPMGl6id3ewU0oIYQE8mb5VK/UJCVB1yNnsme8A1DtO2UCR1LHXrUJwhBygWqY+DvyjoHZWVA
3Ahr/0vbY5O0Krw6vNXqBr1eABjliDJsN5/fcE1yOe7cPn4Iazf0byI+PIZWdogmEO7mS4nmX3pC
g34jjM0wXv+aDey+biLh+v2sYZweb2itZjbZaEMr8XT3/cTF89UYkPUmcV7iQevo7IGMwO9xMrZx
m9KUbRe2N58Hg5tZQodJfmwIeBcyXnFBHbH88d3VRigOvZqRGSR1mFJ2Unqftn2BU/71J8ln467V
NpIqx89a13gdYJfGUyhO4TZ+vYBKSoTU8kZqpbZ48myyFQWFS1OEA+OIImh7qcJ+HVydb0yeAu0+
RRrNz46a4U16M6TBFNQ0YMkSzgSnutNooZRxWURn4PNBYGHhlbvPdFEeuP3pY3VnyK3DtxtTh+4c
DTh42sIuNRYYg0irwW1YBxRxOdCgfGJoJ2diPFX9dP2+oV2y2fCAz+tBjO9LUvZj9ic+RvXS6BEv
591i01EGeIlzWupaqs4t5xFRS+bDdAsy9STv6j+5+YwZ94ROEOt57mK0cmdeSDEiZIJEnHuZhLoA
kni8hJoRydisFtpYYU+M0wM8Q/0QuXY6sK3T61zj6FJxo18JbMpcbhkfdjySXcYfWIRNmIgYIBiz
LihcIdFp9dQ8Wo8hgY5A2IY37OWPrgaq/VSXaHePnZ12V4YktftDmToITG1u+yMHMcWb8pn/57Tw
Ci5FJEKzRR3Q9EzxaVHDxcQl8c5z3i1VEpv/prAPUDbD0HJFPp/f96B/tXPKyyoNvDunc5vA2gm6
d4DrM3gZK9sIkDzDbW1UIUwCPhtYhnb/9Hm2juqjPYyRlXJA5xrnoCWpvW+swmT0FmcHZHwgxyi9
nbaEGgwWxTC6hR/G2WWT1Mol69+blCJHqTF/L6OjmEegTGt1W6LofIFbpCF5QLii2ZSMzg1aKFOg
D44FbG70bMmV2xUxYir7a2TyGnJaYyNdFf0F8jgtfQw4yKkEF2tX8pFI/4/66rU3ZuK0dsegtLQa
HhyefSxzRm4pmTnJFrIzBuDVj+Y+YhsjTM8hUdvBC18errpk6op0OoHTaOKnhYycOYgwnbW1PfaW
yus2UWF0y68xR8tqOTOydU6fNJD/0pK3xdAtJWexA6b90wKKNm6Drqfn/suy08eyFodd0bZwOpmR
gex/CajSsA090VFnnZC652mvkF+Yn4ybt7VvBgy0K7HNzOx1s4PxZlLEX5I3Nv52+jHHF2CswPdg
qog+P1frIujpS1dtw6Xi0hzNuKukeTsgY9VAwYHRhxUaQ9Xc1z3wtBRW++wtl9okb6Wd8lfQClLy
acVuF8zeuPZeHiRvgudjkn4VCEm2nwePw/EDgc2klvmaKhXvcuW3na6y28FF+255lhpWDswU6nTa
NajhS8vbaT6OeX0KxfJIo0EiTATD/zp1ZjPXsniugnLEVRWywG3tp7dS6AfKbFRU+6+3saWJYK1C
Whl4wQB0UmruNhP0AOXrB5VLxCIdxF7GC7DQ3gCcSwEI96zofAG+8cIEYazaJDhWBcYCAqKs0RLT
2GW4cuWepHYRKlWopjUD6z8J0Foz+fl2TMmI7kvW9B0v+LTZ61Yb0v7oZfEC3DXuL423Vc0IZgdi
GBS2dI71UOaBdbHPJNSj03z2joUT+4BIzFGAAhnTpkOgw5MbusqKcIlqy7RN2Kw50MwMrfqDMJsx
VgoOat1+9I7zNrjwUi0UDFN3lh++pc0Ku/hytYfanf2SsWIdYTu9sXQmHAyonQYwsLWP124rWOfL
IJZTMEGNdFWaXC82oq0vKEWVXXAfz/zHN27cXOgZrSLm+0zmEeNNP71Uym0TJAQXTrI+Nyz/mC7F
5tpvayf3bVhxzPuf25SfnmAYGIRUKUXkVUl/GFMBmLCQVpB/NvMH14QFn/jZXWXjvk5yQONDqtiU
Xg3bJWMnY8nvkeQFA2X2JCPBNPjusfw8cLCfGj+77ui1ULUuQd/cSGMllFQWSs0kD9oHco7zIp4U
Q7eNwMMZ8xWCbQ5gmNpAjpb9/39g80nI7ny+JrkDHEVM2L+oqWBsjNaheIJWSqLM0MTYStK0tB0v
iogsEzSuLpLPRL22nYQiPNlPWC0eEyBntT1dCa3qbvY3q1dusitfP+NQl1F7Ij2ZQGzZOAKDtIx0
rHYkYyBmHOq2idAO5LOo+s+FkbUP8GJzPvoCD/ZKWEtsUGF8TqtpNrkDmeskRcxfg/c2+PfwW3Rk
/h54CUXx8AAnEcC5u0S6huQieDGdvsFiYRs5K0lrMy6HduBffnLLSXY1YkctYMaD8DIAvHXtODGN
st/jCyTBXVbC3JbFWArZIJLdnuA4gPAs254Dy9E1JGyL8Kim1WZW5ueo5jzjcrzBZIqHDiS+E47H
f19atL1Ii9/6faxqSPQyqth6oXh+V8WGTco6F47M8iEyY1JESHeRGDI/Wjo4r4oA291sfRIhj0lt
CXr9lFcFpT0cfVO2l7TZ0y33nmuMdRwiD3HPLfDelsOpZx0hAKuHct9K/ZYmAgrUcBPErp4AcbUf
fZqsuwrMyYGSjGiiJgSo/i0w7OX/RWOtZh6tx+hgzIq8IUjlUdWCYlf+gUvhsqCS24QxAZ9URfEN
xhsRcUHlpKH0Jbk+vx8oD+ktPJnJFQ4yF+TXN7xmL1EuZep2D/gm9jyND+pMQvwc8nX2oDKRwniK
aUCTOtcARrkz56pcCU0Z75REA+rLICsLAnXHoauW2VPDpRvMP+DnLHDDKJElN71xHu2/A1nTn7ip
fywftMV1mYL4rK39yhVIcMF2b1b5RGJxiq4YiIopmHpVA9wrbpTMhL3u8/iEe6H47rEK8sGqhDYr
QDzW447XZIG2KVmSgKcBX9CfXNgVa+SSXaiCAfxkK7a46s4pwUCI89GadxVi8CXH08G8GKo6fm6S
DLqlVOaJhqSxQkBHLrUaE1eirbW4c1RhhNijqUEQTFQe0mHKPtX8hQ0VFaRjYGZJc2pDhV7ZnOJ/
+wpVePbbt6ZsegGNhLMnI/mjrbtUam2s9biKo0Gv02LnWUSfdQ7XVpjmUXfVOendJyvOjqD2KWpL
E1YVp9QrwB8PxnRfm/bU6HZMdxpuVB1uMQJHGkg/FvCOQU99Xx7AZ4krZIpF2UJ6V7vRMxDCuINc
Ot8qtADPMDs3z+I/8AMCejAD0ienOau0G33B5QBQbMiZ9Zyoe8twjNV2jrmHyzFYT2wp8a6ME6FC
Vyx3jG/6W4ygwvbH9wvP+fwBWb98wZ7n3bGAy8+JMHtNKwxxy3YjyvXda8+SWQRQC8ctMOMUxcUs
C0JV/4JMtzamdvMrEbr9dIIHjD+hixTpAGKrKTk8W6HeRyrRmalIBDLYPvRMERWFkbyFpRkmxsyq
Dn1yPwsrl5JCZgDlrZi8OGID0TQmFiE1xbn0lBFSPr6F+cAXYqhJa3lcyfslRz2uj2BTOpMBzY2L
o3/61+Fj18hKMxZzhX78f6U/79AVPTzD5Ccz/ONE+lgo7BDx+qMWkkZuGDRrh6AcNjsraDirP7It
XsWZIJTaittZmKTl3DFzHnnK0A3JKKK2D1PxUXehtRmHdjXsS4fHlEd8N90LEFSb5PqbutO3RfLQ
MIjSlw15OjgoCBGZytcKQG0p0glxidlZax4g1zMoyeflO3YoJ+h6LijIuit7DR+VxzS7BKd9BAH+
rNJcSXkuHB24PszftXRPLsgXeO1OtCL1YB1qXuIp+0A+d985rcEWdCMmTduGIJHfmzyBoo2PrS9a
LVkdPiJ9haV15RiG6Sx1aJs6Y2fT3S/d98d+zXTojWUFVea4WzDfTXbKWXhHZZw8rler8rbpsZKE
Geq2e/vLk+VPZjOqzLTZDSrTghLubXP9Kdg+yCbF8PpECxHJ8XRv2VRW70I7D/9pW7vJAI37zjMs
xFBFNXn1NxdI3nqqNbbipn3On7QzlmeIGVEoZZQwH8mHm8SD6yVAE9Jfwm7pRfJ+0AXdHkP5bG2q
N0+GW+VoL6go2fKuayi+GN+aPyL/VAiVSDsAX8z+MjWKO+Q7DXnPep10nDkhc33zpCb1uJiQD2dh
riaDbipluuKDUbAoFy/JFTl+8acxILqbTRbuLeYXrC/5paS4XZNUV4h9ygFl6LfW8xa/TO69I9D0
3pV/WIhGO//4dIsvho84xgx+tWPv9PSastfhmUNA7HgX6L4eAHA6VfqeWDoxGAlODpjg/EHHGrp2
x87BjH2hHtUTRGD8chkM0Q1d9ZNKpIXbyfDtsRAHtnVqzQQ7v/weoHjqa8mRHVwb6BwYfk2A0DG5
yGdgBqIx2G8LjMuTAvw/khSKMEbLlzF2H918CSEiIaYv0HWGyVA73TNC4Wn+3dzbmvvIyxmGtleT
x/zFxOC28ul9tCtzl+wLvel7LgG/DgmTgwcsb1mmt7UxGsVYVGEbe0IWOIZ9BfGJ/raw4DILfhFH
cCqOZ9PT40zkBb3NBcSpgGJYFd2B6+we6ArxtpvtUt2xw+PDJN6cMrVxDyXioLRoeU5BebNMmn5N
KFAz9p3vNqNCSoT0ceCaRYVCf5gaB7PHK+NfVjsiwCXD4JO3Ru1Cc5Ujyf68JVqdtgLO0LGDE4YD
SsxuJJYW7VCvx2cYp2W9K8qgL8rWmtXu22cWDd1pxi3RfE9fsiZ50E10Fvg1Q55CWgJKm/G8A85J
oFVW6itQ4JMWl+vG8SqAsCFw/n0k+ZQSr4BWITSmvuwtiV3p/MWeczDRpSdjKWWEdmYXqw4zySmx
TgKJbrY7P/h1qbcmPK8tUPp1tkTguRCTn7ro3UYfGMOfZOy8Hcj48SzwLIgdVssryrb8TEbDM2wz
hgM1TGZLFvMpppIlGo0VRIHy0whHFmI18jWauhESdNsHld+lPUjsompLnruXtb4WpQ2hgNXFokdd
1woToGzQ2EHuqLDq53L0OGNu9IBLMl4S6dJn7k4281NJZ+DOIoZ6dGix4w9GrZQhjHZkoOPOxMBs
6FPmNxGZa42etCi2h048i3c0GBZooo98rnXAWDuyBusM1W4nASyakQMEUjCf/6kN/bScg85ewccf
BMrFfNatc8/jwyI1K62LuH0v65kVHH1cUXkFv6ZK8/704MDEZ1IOFOgNPKlvzSZ2rwPSbYJu0P6P
lqK9L13OVtd9vTznAlNk3fm5ECaauwv4Nz6HEabidKTZ43YoK2nsVxDQQPd31xnYvVXQqs0qJrog
9OdUEWFsAeYR9x2rM5FsDQF+w+on9bYscn5n39jkrhlqkYCJ4a6zdDIs0i2ZNTQNbpQToJk7tHYE
uFbqz/x9deMjAN2dsiS+4dMgvlrITzcxHxD51mKk5vtTIEEHkHM5WHN4Sd0e49jmrPV/TNptaHhn
k7kd5UWeqdZ4TytIqvVayiXoqEGGNZX8oSqvFXJS+ZNM7PdZE6q+qGICJQOHJeCXpkJg7lDnCqhK
qQcJr6kNgHzDGlQB1xEeNovjF79JFnRLsLKaSQ3k6ElS0UViGg9ZYNuZNmtvVnCI5MlgaYHVFOJr
eSeoRxVpiHXY3FyqWThYrkVPp/oMC6/bVRpivJ4cadTHYsy+VWP5c+hyxRJZy0B6vJm1wgMR9Yf1
HlB0L/OYcOqT+zeOjpZJ27Pxm6tYo0XKwGAxc0xv444Ilo0cwzG84dktPzzdi8g4tsmTSF44blOc
KsOPq8D+cwQ4afzDfIpDED/IXMSmdThxZ8MREIIL/a9tAoX/fB2MIL14HziS0zUU7aLpvVcsvUmH
L0tyq9lRkCvq5TI1DL0p7kTxPHzxyAVb539iBCHF47pHYT4+69lfn8pMjVEP4IRzJ2R3uw5pCsM3
jHyLsUs55r1N02V8+1lGx0TCIbZm/+o6A/BY75QIoRWonruy41Md+HoucMU/Pr1f/PG/gCvMaXyl
pJD7v52BuClEZeR/MeNnyEhxlb7qBSl6iIQfQ6s7pNeXXkVYQz6bFUyAx8yy0xdQUCw26qF+ylTG
06cj1EsZndTx36AmqidG3oSKIO6yzdj7QHr03LsIq6I7W1Nb0+A6Wb7rcCG9gnmsgqyT57WdVXjj
ZMOI+N+5syjUT3A2frfB0ybZM4TUM/95IdhiQx6HFTZF4V8LxHFzCfmq4APnM/lzdhT+sGZ3ASxz
ty4VC91gKuji3AKoflJH++jzfvIm7Rh8q+c/KrysEFB8rXq4M2ROGfIBcqLOuOSUdJL3ulH4XEgs
JaMlT2Z9sbRnMoSXLa3+Lw+y+7by45HkjMQqD15qVc+ooIaw0o0b22QpNm5pW3Y508eEUx6WatTc
AlY5OtlMIoah/LKyIYYOM8VSfQmxin7NIsgzm5Ez/BS7HIYzYH/L4XnW04akrd8wgfP9PuF04d0Q
eNOfsnQeexap1CfZNq9Ro3WjrHHaOyIJSsSzhbHmbwexZtz6LOooE+wrSlflsumZiS6/lGzATnWl
iQCrWGzdIzClUtWtduv4HukuKIzKfucEcCDlvZYmdc9t+bfsPJ5nkvAd/MEBkb9vSc07KfZfQayy
w1/OU1RBI6HP+7fSITX56Fy+XO5VhqFeCQGjtmW7KH2h2Jb6ACxSKkXmUpUrgpiD4s5UawtfeCGD
a9kzt5c/ZzGl8O7oxf0PHJDpiAH9V9LvbfHjnZvf/BbGxZK9DyhdJAPqvu6IWHaUBhEfJOyH54yP
GDcjnxQYqPe0tOxn0ClMyzK/aHs9JJllrI6nu4V2ntv9mhaQ6iUjH+NCwpkiPiC+LHuH3o7sbDiK
FtzNDPvpxVaiig6KwCUPwt9Ckv8r1mz+Kt51OeUv+6kH1d4jMG8X0yq64tVnnQaeAkyi0wxNUCN2
pLs6IVBM1vLnSQWYuc5PMRnC5A0k/jHh0FLdtH7mjFyL5zAzpDtG86ixAnxM+t9gl+AFNO35+EHx
+ZKmR5CEDznf7h+J7XuEeW/vZJ/s0APepVDElvIUnRn7nKSPWz5uFbHFCMKYXT4hRaoJTV9aqdm9
/3QRrh41Nz5omTgPjDDKyQHe1wlpcCjrkaF2kmrJDmL4D/VdOkuJuvz9bP0unDRxxclvXvRvx1IB
zX+B9ViucaMK7mSGDthILtUn8BHK1qZprrmshDrLWN7crhmVpzhqQj+uZUXhgM+M12zVYKnrnYwD
gxQ/iGxUfdUGeKYr5O1szMD5FZw7xl1xHRhZWqbnHg7jX9LkKQj8f6bufXAOzyd1wuOakV2F52aS
LyCPoryzx5XhN+ihPXwFyeut2CohbR300cKcCKN6def3DSxiATErKUsNhOoVDeLOHrsW8Pkst5dx
kvkkUpzcqZvTCfYrEFAmNIy7qi/vBD02hG287zmFnuMf/oGA5k+nnl6+VQh0CgPTyQ0jbVjP00zC
EqwZdIF8ZLszfLotBotms8ZADHaCMsK1wJr99s7YBa5aTpoK3nFkC1467zCUzAHhwnUEbbWxCS7C
zHQX2BBDMayqjNnUH8p5vtao0RfR2kdjbWW7cKptev+QCb3kGwWaMXUsWXJeHHnloXk01Iq31N0s
4BcsS2Or+S6h0uHmG67k1aQQin8KcxkPEJxnr3m3avt/szDw9eK3kQuw6Fcz+bSk1Ea0grm0ZX/X
Dtsnjgf6ZCLKOowlWHN6BUxpMs6M2d5HlVNprVH7fz+l5CbVaojzLHV+2dMuMllAYaZsZc66JD/o
pvgifCrC5xklmq51fwfdp/BsoXycAYPBkWKOd+rbz2xl/DZj26qItZpI0v4AiVu9zSI/vBHztQX2
N8hsjTYxCF2JUH0Qf9m8iYefl/fNXDm4YKWAFUgasOYZHHDlnjPbrzvTi+QwubUXP6AeVXgCrhsf
GPUtbJcNWxSrWSArJnyHbUOyv0eutmbPsX7WepbbzeRvMa3dZ/8ndtJTDBpQqffaImOZEMTd2P1J
L73ntlcN+R6X4ohOWQ5WlKxgWHivoALcaP71qtYkQj0GHWSTfCzYeZOSgpMXC0Ow3fbLlu5OdnsY
64aZk/a9g7YJxNlXZBP63WN+Thrkq8kud5wl2dNExEUtLKmO158V8l7fK2hCv6xvW60VCt2rB5fy
yiCUvYmc0SzAZvHvnudWqFhEtCH+TrHjmaEyVsui5RGQbuFDjNwFXKHFB+aX+HM9s7gCFvoRI7W+
UWJw2jUtwb41X0e3mCyrJ6W0icn5sP//iyfBy7lxj91Qw42FbQ5Y8XpTvw65QvRGVxEwA0DFQUx9
agSxUyrql2nJKjxorU58jU6NHk4vLzF+hELZ3TebCFAw+wcV96udWGKReEVnbbJED6+zJFxOVPo1
EqMR5m4GDf1DeUAGTm/Tw+K5UbzANTJdcv1RUrvOZ+FLOaRGUhXA1jkOxi2u4y3bO5LiCn5+v0eP
gcQpDQvew+xxG5vyjjSq//Hbe9XhFHm38cEnozmCmJ4LPFpLbdLDYtsAQcw3dDa/NZPPJL2cedw4
8ppHPWP98di1ik2NFBHnyYhMqlNrmXq1JpTuXaaFI1Yf39DBhVJ1PP8LavZLCGOazoX0F0u2J694
nvWY6aKbqmF7BAwb33uRWtzKcaTtG9yh1DpX6sgNNR/wxZzzAFN9v1C2qa1MRK1fSCNJHm+e5KGN
zKncWgmeh5BzQxTcMAk7CTmryMVk24plvOx4GFPrnGWGh8Mj/vybHcjyKuqb17FXPMtKKdh6APlH
p9RPcXOlpeIgIFF1iLcxTiIFjTpsKQkuVd8VT3hhnEaDisbdNu027+F6RcxEgnnm2K4QjhZGfwwe
nFcR6ylfFQlQcLd7nvxPIkwEK4ksPY9U6jhCApF6ixpw2r6WGeeVtavF8hS5Ri7mt/smwJU/p19c
XNaEmoSvtpTOYQih4mSEXcv6OtMN9MIDJuFb0/fpHr7Q2Wyld6yzs7WY6t1vnAkeab6o6G5JnyRR
/OnF4TGfzgx2restz/iTye5HyfQwZevBi0tvnJhN/dp2LgrrkeTDvRdqkwVrnNTASMFFiN3+OaTM
Q506qLV8L66B2t0TYSikZbybudkNDp3cPZrcNXpkVA2WFAXKepimkIfwYDZPctSJP8nQtmZggAAs
9Ozeb2DF6MO9nD47yiXo40kHIBiEYBx4ACMtjADxpKbz9kd98T9GalMvRFhx7YBoE4HRFXT2it8z
MWoHBTzaTMSBDVMJVgojnrbpR4Y9+VMwTHNyLTWy6zJ3tjFwsuHqCu9kiRsiFrpP0Da0FJPj6PZe
JwR8PuxQZUC4Xk6NtQ/jWG2kQm0EbrXkNLbU0bhlIWdDdnbAVuuOjLmRfAiCpJUT6KYrFHc+QJdU
il/J9BrbX8IZAPr2a4/+sTQ/HIG6lULydYgHPHwkLiHB5S3lpPphDJo34Bqil8U7F1VM/ofsw7Of
j1jSJrYwIgts3t64nMl1e0twFzkOBX7V1wZIvAHZvilEUdFT/qS4Px3r5WcHVuLSIMAI2vLbaC73
78LeMEfYNlENj5tiYFldpn4A1iYChrU2u0pm5+Og7YLZOhNo0Hz08eiU4dbLvUaDLJYpXqqDyvNW
g1aQ2x1Zo9XT4g5CMP17ImuQ+JZYJU2grIkBFiVX+/w/y5UM4o8L/5BZoC3q7hm0Ko6lZuEks7Hp
OzMQHiJPGMgkCi8vmNKpmwao70Zmk7vTVbVyfQOWHrJuE0+m5DMQq0ZJXmsfi5tURwSJsJbLmS/g
UcFVJBaasZsKqBT7zwAJ1uzyNg+1OpCeVTix2vnrX1H5Dy1arzlk0JLFaJ1leAISmnj7I5crjs/2
wnNk7vgWDjysiXsvbRJFdU4eRnqamuwauj0ti9270jMvoVZJ6Weg8jf9A0yJ0ee0AWpgEWeRpj0K
8VmYHjk2YI9CcoAsz3XNkaQVv7U4g5U++TtI2ZYRXUARnQPKvSG1wVftI4F52UyIogJ1AEpOlApb
qRK5ARMVu967bQEK3YQIiwgH3KiIr0489w7WYXP6sbOS9nXBA7ogyjO/ADTDNsgMHnmgzjyN12Ng
GC7UpR2NzoOCNHL17/AyfrDBMYwts7zDbdZV3IZAFrUHmnBwMVDoRbj+n2jCgGBiJJekIZ8eNqlG
3VuSYGl5H7b84U+kZDsMIsTZmv3O9eW9d1mqrM6Bvi5aWA5q5yebLwKuSEUiV607T6rMnRW9dL+L
ez7AS81VIwM2bCFRZrESvseX85XUm2EjcTYs9dTJhhjSXEqttrmgVN7tvc9wbfTInRsSAUOiskb7
CZ5sC9kcDXzZKzg2Q2of3mF7WS3uUe9VP+eDr2TGWFqqgdX9sbM8fwkiPxFv2gr1IHJPOU7k4WfC
CdhQKJhax7tkUySkEicZ5S9PyBBVttAu4jr/zJA+ZPnGoZJVEON6fShiqpNjEis61ntMlgqO8ste
fLSjeNZ9U53v8mOvVgkjZ+k/v0FeUvTC+fdJ/lHf9bJmlKvq/PqfKUi38DHWnlzpfT7SN7woRbvw
O7eTqfEcAopFqNgmOdoLXf6LmtqZ7ubyTdVga5GVKt+xJEjvoOLKdyXdoI4IABWtfelk16ScFGwd
nEaSPpidUKkL4d1gonATdQpXC0dgkMq/P92gCUU2pEGjoK95yrUX0ACAMvv4Ij9KoWlZnhDNHgOF
W9QlEMRatQ7BtPj6uV5ID2IXzDDqsD8K2j10nbiCem+807VGgg2c2XamnddG015WezeNJDIDYL6Q
k0ndycyUoo1Lm3/wJJZyeOr3ij3droAR92dz5dSoH/Ys3EMAIy4UDmPHBCkzTNpAbiE9F6LsAwPL
/WCVOU2ntPHv0q2WA3Pl8YEnofWl7OHCMsD1eY5RZNWNNh4oE3lTqjWQOSlO+ednWsI8cujSa0pC
ix4wVQ6tGEZXBfR/f53mv4iScl3T3Pj5gAmTvnwsj/z0BmHe3GrGiRjkEP/d07uJXjnsE/sa3Nqu
+Tqaq5/5N21DadSIyD7pVCJRqv4/BZwYNpsSu5H98KrmN/pbFsgSzYDDp+mDHFTn8aIiuQ5f7qE4
wkW3tzz7LNaHnj1rnkSVlrrFQmy2LnWhjyTdxH1PodgLzaDOLIagq3GpW6sPxkPSjH+reONzSdyO
k+AG3MjEF83Z3XOl47TBCuKSUfkSxah/CmaEXkKCnVlddzQ6JZULIQVzxRaew+axYteR6z3lRWNQ
R0HopbCTbgC5f2DXPxEhoXn/Dlbg2cdVO6CHHgm+gttQZIxJsPNVHpF86da1Ei8XNcGUSx0XrU7J
F4pjcNO0fORdFB4+qg5kqGyXcl7ppN8of75PpIOYxKDx/iPXhGtDqMgli8GRE3gg9zCl7DxBhBeo
DzVb9YTbllUs+SE6NGDuI5hoQrNuq+VDM+LbbBRWbgTEFTZiVt400FrYwd1sZQB/+LSf8nHPG/IO
2Fzx7i1CTtWCUR7a+IRiOx/nWuwBJdTXNLWW0pKK50L0HMimEehnY7PZjUwgiJyFd/jjCFcjNYRr
gHgXdyjh/ylFcY6jQBE6GiyV1NgLJdM0Ll4AllGailFHVeQ2WrI2GAEpbbkQ8tqs0a3dDuOsGEbK
Kv0iPfq5baSFMMOrOavWfdD7e2XTeQlwR45mlSVS34JRSfV2hTYxz6akJv2ONDCaAlUMrky8+UAF
XgIK1selFYGrWrb9D0Z2qxkBSAuu7NQwhYfBd50cFo0g1PWa34K3m+2AZtAkC+mBPPIseL+R8vRE
F8oz2HRQ2yTEAlREbFm1rmkfIWaRaXKPqDP586SkW8B1h0GI8cH6+7fJtKX93wLzrfgWb0rGKmcq
CjVfL+qJyC1DBD+TwecNWmk3EH/tA0dv81W/UNihT9tlliXi2BwWQFBiINJpv5GK3aOcAjdSmlNi
P+Ew+0YIqJyk9wAtbqH1Z4ee+HojCTV8Z8wOJNRjPWuO+ioNS/MeN4yGgzZhxXxjBjksq6QC3xpo
ooLsd6F7kKQcfZx7ka5TEvBR9EiJdQH/0/od4FaRg5R8a8dG1JIElpIWU9PKG4YZtj0i1iGki4ww
dMSIuu097za/UQzAg/8OyhV+BgzqSkiimxNkTFVA2/3l5KWnkwVHXJ6jl2U/j6SfdNE68vS0kuW+
RHtrq4NVj3ykNCrez6bhHjeRnyHKOr8FN8/2Y4mj9qTolUii0BNYTNR3eiqu4GUMLc5JVePAuJy4
R1ZnF3sRxQL2K0nDNq3LnoMuhNyLhjq2Iyx271ExZ+E8YmbXlixgkxVYXZhHK0dXs8y1qdynh7Vh
D/JNWso7G724dlhO0tg1h8c0nY2amOk6wZO9GXKxvmoBA4BXsAgYhStfsne3U09gPKH2TEboEKj3
OgyMNfkKeQ9YfrQ8uXlJ6NtuL4hiWNvMefjHGx9tGByICr+ueKbYlgd1ZoJ/wwmnB259j1FP292S
TjMMNBBzCy5bsD5moJ7SP3Zbq1vzmm8h+VcMOF1VAYAaRfsdXD6lrmQO2ABnRMbcL69ZL23vJKga
05n9nZgrSAZq+AitgWf2XzL6TzLjDqVZr7mRiqc0aRsIrfUN5gFAFWwfGpL1/kYv969K8A7vmzMc
qEry+Nu7OJOQ1k6Uf0ma1shLPsvJ4dGjuvQC7WBPRQL3wu5+tTD5KTRHuDFkD/LSfKNs3CfhDU1l
zqV1ragqrQ72sEb7Lbn8C8P2yHZy3eO12VJyQngCZqb4MiFWsIl8Z2VcrT7zEm7rRo5sB4cx1RXS
3XIRsFNjqynDD4+KNEwMD98RkbocKVzrmCcMMzOuzKdIv7PwdHt6CWx90ZKh/pLL2y2uUgEEAhmS
hzE0YrZ9WWvfCKqm+HZYZ+FW5ewuJ4ZJvADbwk00op3ZjPg6XYi0kr/LBSRXw5EMOc/AUyU6yeJA
OE8wDDrXGRjAcVVUITqqOWrNKfjaWbDlJovPrzDMpjTAOyclbUfQSOQD1rjIyQy1n6+z/x6O9EGs
pF0NOf0uVo9tV9L2XAqiB+y56WimyWre+AWw2F7tdG2w9c6VuAaK35dxgxjDf3c280lawYpu3rUD
B2rD6Vl+MWW3Wu77ORWQF7N9Eyuso+7DIJid7zeoA2i/0xCrQrAGG8CO4FVJb2nHnv3ulRKCScAH
CcA6LlNJE+dKr093f+ij/R0RjgMX8MXFPLpj8MRyrUW2iHTnqYUqjtojbxAF0UI4DcLz5g3GanAV
8oGvpvpL57GmhoGLH/CQipC2cqr2NmIs175f6095H/+fF0Eys8ANacKDnhkbopfiGJTR6q7mChpL
nHc50YlVMe6I0J90Iw9v5I2uIq5p6dM85CzLIgZis9atoDoG+XAltzL/8C4gNS36OLLhiK6Ntaux
g9E1rSifrtOQwl8Y5KqZxB8gbGHEZLEQCzlHhygjIilFrfg67ftRy3+YtoLB7em7xAIBNgke04ci
SyEpqD01y+3ZhA5qnZBAbUY2KRuM3MzwBUF838BW3lelwyInk3i6jp1KETHOykA+YNTSVBw8/08b
ndkjcOm4u/usP1DHE4uJwb764OZXU6LpV5P7hDtJmVm2X2OPUf/CFpI8E2CLwU/nfJqjS2N/X+TD
nyvPKuhFm04/735Vq3p8WpLll8WxEQCTr2EgpEGu5H1fgMWd9B1Kk6DDw4aJnEjtHONStWD3/fIl
NpMalP3fyp1rrCJa81HbauDsWn27Q8S4Xlrwz0kyULbhx1XmW6eKsvlOsHIsLBGcGkOH9bCVVAyt
MDn+szMCJun5DGwxkJOtrqscCO2ajRPXnoJGWBhhrfhRm2rA3O8ng8Sq9uC3+TVLVPhz0lgFibzO
VE6LdpzE//NW/3KHmB8fFZQaYUI8jknCQj355StI19LzhrBaIbmxs479D7O5dIGmbmDq3toxG8F2
3ZXP4+2QXxHdUc2A2Et1d3dn+oz4v5QxrWpsJv0O2ReaXLKZYPTYhFeD1bVh4IExi2ScQPJcspgV
1EhlAnoz2aO1VmGQEbRSsGlrrqEDk6DUaNX0g04EotBbhp4y7o7HqgDU5aCPYxfYfIF9Yt2OyQ4E
JW7Gy8xPSeu8zaKP9qKUkGqLYxoMTUps5nsGSmhjnsNmn0gCXEoyoWXuZyqnK7OmPJfLuDzdKoll
Hb28GFHl4BtgYy9wh0v//x42GzJKsTWS77MwVpsiFNx1ixRJtcNa0D4eXRXV9Trd0sRa3G01WWrh
jNDuOaocvX2EU3vz7sJuOG70MK2IrebnQ4SKX8t1PJTCVC44pzet5z11gkrqxd0ClO4XZOi+Prmd
MGuriBABXY+B3Ug46Uyd1c18kqa1I1ROImjYToRc5CWalS3l9GQpn7FyRH9osN1mdQ/z3nmAz3To
TtHL5KfNOnm0+X1Vnr/iyFCB+OCZf4yHq07mnXX1YN+2yh7u0kErllCU2TMsxhbMLRZMjeJzcRjV
vrP8EEwlmg6U3itNzdrBwLLyQkJhhwuC1mjUivMcc9B3CQv0qHQFFPfWIqInFA6Avz22SmPzbgRE
sJmkTTCi923Eay4Z8CY+46pO8mCrMIxBJuuRcSluVv1u16OpZOUAgza2uQr5gx9Yd5FQTCYQ1mkx
xwAMgWMkfzaqT/5t8Xw66Tfq8SlCSy7LMVEP29LF3UBH9Z9ajmt679SJEBH9dlvp8Ff8o9EPWWmA
hanVqf6G4Z5LhhEp59VK+QjVvei693vdLby+SP29fJ6+++oQ7IqUV14SH92OpogK/0BT8V/Vs5ck
ZaHEGWbF84W9T02Uu92tyVr831pUeekiTTiHuaUO7GSPCx37VcC2WyR3WdeU4Zi77mQe+5UCuVkP
Y30AgLSdmPrbvjSZAtKmSxUYvp/1tW0sELW+hPNs05/fV+DgbCdbvYY4jHFsQztmvpdeS2dP/jZ6
fyhAB8eARZKgR/R1Rz9Rub63fQ1AEwpArkTRdwGPNBm2vbQGSdArRYExVzhCeBvOoH0efYt9tYL4
p3mrIk4L9tw8LRa6o88Ru1vEF/0/UBILsxmdu5X6qjvkxyYv6V3bHRuBuDWmyx6uYGwkAvtwQngF
LzmxeXzBTML03o18ZXehbsGP03SGE8wnT8xoPLOiSAN2jt/9GBQk9HYawixn4+Htt3l8J5dRgedo
/Mf4NFM9ulBexmLgNrM4NebsfP+CpZ+TkAr2sYm4wLw+MdKwIy0W1HfBbuswGrZ28ucwUlu7BUay
3g068/o4liG7i/JomxO4gfxShW4JPHUc9sblkvir5ZJKAyeK0VVetC8UHZk2mkpz9sdgimkP3qOU
zLejaygdLQ7IsTP3TSFTBYbjfzT7Y91M7AGV2WLOtOeoaXuqytD+BFtpoLxsezRUPL57svCeoZTx
FgsBVJFVP9Bx5ki34f7Nu/sjtM46qqeRG/9BGwye6zap6V1xwPCfAkwlkP99LQIwrxuJ1Qmip5KD
drDNhzx1n9nSR0o3Ne+vxoYkKbvc3BZBZg6kLxeqk8ro2qvTcPLY+GuumMcWCyOEQ78BUjYP1WEQ
+7Lg0TCZ+VTNi48fzvapCeyI2oa1YLrUoTjTUDfDkbr+qFNIwKLamCrviAd78jKOUJtgjdNSTKpN
o4vY4C+NwX2XXZGUND2ronxkcruB1EJMosxWDtbyttdl0Dw1uGeA8ZmjuXVWO2Ci2cPBQvF/p5Vc
bFqQhkS2WR9Uy2X+OjLusQ5OMEM7PXE1X0FFxbQiGZoE0siIdQz/ng6rrqyRFYrq5LIvxkbmB54F
7zHqq8fQYr6pj5drYyc/TsLKzyCCXZZbMfEsRuU7DO5KlJzJOZHxjCBw+GFN1RgufyckDY4Lq2Em
fpA/v6FG+utmjdWVUxzCRejxlA+EmGBxdLASaJ7ebg5S3fnxtTn39GIZ6LP1oh4JGFlQDq0Fdkyv
WFa8ZBYhyMBGqtXrCjqtLBwq+ILdyZTw49aUHxY+iQx6YyDEtsRqt10kbmlwGHKOvQGfkbQjeAWS
Ipfz5WC1FRs/s4D9cBq/S/769zLFYSWi2MLnPhVQoVenPnm8A5gyaiiJkJgN59sC6q0OZ2VKpsqz
lrEDtorfgj4kZlUzVkX0f9YpEaf7o7ZqkS0h81/K8WWZZYgzTcwA5Dy/+iudet3pIbygo41LYNsb
963ngKVLDkFd7MhpIurI/ZGxjjLjPqiuQvO4zQ4mSkUHVqt5go1YxzBvGFW5MkcY/Z/6CQLJA2aF
/fgVO3a9PuX6Dn8rNSJwj5JqtvMcOu+wpDIQSMqp0fn61/aD2Q1m1ZPZTjoQiKd5iaGfhWV1SAQ8
7TxWrSr7n/S8NWQs9tcSPVjxVfCC2Upyq0UCRYRdz6Fz2m8UyhWSrMPusKBerR7XwAua8/3+xiEy
e8ukfxbt1YY1xGvxM2pY/k3Lz8CZSyP18lJ0rpAqLkw41OyiljNAdi0J4i1tUS4AFwc89I9XhnPl
FdpFc9L8HfCcw+lT7JDmffdjFMkvlfMBmolF/0XtTHMn590sU2mTg7zcVHnru2Pd2l3x3Uoz5twd
D9cx0FvCuX83qS2BfJ/cOZFS9jmRvToOVm9ficijHMIb7X+xI0Apzm3Jx9xLpkP9S3jlVhOzorKY
85nsjXU6HPHXj8jP2r9XDQ7YzJCAAr+4oh/1u7My4kzd2ptWdwoWTS4ey7nhfMX9/MOyxDmmrdwQ
IqEwGfzgzaiEmt3BP++jf1irpLaYSKURrfInmd7Z6iSV25irhPc356iqVcMfrz68I1oeLeMYyj8h
saN51zBaVPoatb8ZZN6r73wspWBWUUWxYYzyrTr+Ef+r6zy2t2LFyPbpMzoPrE8XBBDCRVIOjpll
NGr1XUHrPDS13rfJYeAucHEWpBgbQydKqjXTxz+jZyH3d19X0hNjdX0jEiSREvJK2bEC7ZTl5Csz
05cCg1E5AMJrmklR81ulVQpjMJtp81eTErGNss5+f4Zb31Lg6VElks/dUSESexTZxneW775o0fbM
A0yvQSjN2ZZjT+UOaKoYNo1uSb9IkkwJRfwFlNMjhWqRckgdjxhhFr6TMx60airuLE0DWO4CGXjk
bo39otESzSo1Uqu7UVrZczvReNG6UeJbAvYiLP6ARcFI2xjJBt0nIl8Z5LbO0qeAIEtqJXCVtHF+
Z5CNvxWnLJCjfxOrfX3iNq3k+Fcdzm/zZ1fbblHVF95dIQf9LOnic3snxtE4O/QAOaSyccDLmCqF
vrPrhjh+klikZwABFsROBXo+w6dc8fui/6uyQIrOiqbc+YdqAMzjo3sFlRYdMeJtRTxQSftcSMan
VvkomMXzg0iKCfTcDlD3/dWqyoq37nHa8b3idB3Easqt7bWufQTDhS+bO7vsu1Z6LvYM48FOXUve
fw5qqG+GspJtJOg+YozU9btKC1wtZd0+1IwDnwqZoMbMABN3neWSuIux4swnf5SI5WdN4VOn+qdN
2Sg24ID2lpcyZzrTKeCZgpSMBbej4eBWo303tqSLE2wUGT5VlwrjBWuiHoYEBGLtGYDiN/wOmpyA
2utc5YCfcs7S9VEAitqCBfeTC3Qn+lpXNonS3FzExvTlw+Is6dp8Gu5V8F4jvueyf+040hXiXZsu
CD+x28AnV7NVQXEUpCe82pvZdK4AthvRN5tn9I437EmAPJcsdyQWOBg07almxzXuKStx/QmvZc1R
yMKghbtbI8ML5bvxsDxkMc0JIOAsF/sXii77yWJ50lLZ0siuvfNR1R0PoxlD0BXgTUfym6zgrSrG
PxtSY6aHTJH4goR/pf1I5p9WHHR6RjgjM7McXI+ggwf+2UhogqAPuyeHTzWo/69Q1dTx8IWvPED5
Lj4DOXjRqTOg21Ex5U8Nv5+/R0vp2qObL0T7YMHDNKSwV1PpI3DQrUCTXtyeBl2HQJAuVyZ+zVG4
++GS4qeeW15vx3ceWsgmSEO96fK4MUrx9YVLBwn1GdWulsANBuqvV7A10ZiaXGC2fS4triLseU4L
O00wwiyiRjiKnUQ64/mNP1cHh558mZJ69p8AlukFO394SgZRcBxl2P4ZBefL/aru2t5GSjxKoz2H
dj0UNBnpOPXQG0ShXTROI5s0wDtdnOpPC3QpjTEr+Hi1hsjnyDuD3qPq2QkisQp9XjSKeIVj8etw
E7NVDJHUh8IQ/T7eIstmjMcKktNvAqHT4log3yf8YBPRyXwmQqL+wtkAZgi6iPz6rMcSzyfy6Wns
ppqxIgsW9KiOpEHkSeumZ31LfvymXthza0ZzyIA43oTDoRxshDe0oT+ePnpqbWzSknSiyKUSSuwY
b+uoXK1cm/TDLAdl0hy6PP6ovK+Dw3VChy9uv2IER+BDm31OSmalTZlKsr8PckoW9Wuc1lxOK1FY
8DkHUBwmjIdSNi3uomP1oGgJORT/WEgREXxcP6yenbE4IaTGtpJuwbZB5w1r7zxN36IK35vUWCUS
Nr3o8TkzhBds+4euW6DYljKTaoyeIoi6RXZ9cdTiPoycysGp5R2Rf2gPrQpwFSBa6Y7ldIqGzvgG
2wIvoMO4BqQzqsOAkBNzQ2APpWZUd8LwuM50ygOh6+Dqs85on0SU2Xom8pmcU38daYjkWHwmTPaT
ZpcQsNYowms4Km2A3JSV35ldBO+49waBLrRKlMcBBEwEt2ePYTQ1eG13IQg3+pQl84AYAjDrw45p
7p+7EqioUsBzk7e0TYl5D8HbkLVtuiTfsA4hrvDRlVFPBQH2HmPMTwBptzqpmanDBcPpqbOlxtnw
+32rOB3MOHKnSyITz6Rs0Uzf9vbPOVfaunW3FzNJK6cXVv8US8++3g8txboUgoJIIo7dgZji2utp
EbbcWzsheDJI1vJTlCWi0nNq4q6phGfsRoe5h0atUCssvCUHQr2KPvBwClUwmH07jxynD30vYQPg
tB3ujvlAMFt4ZAtdkoPO8aHjUTF6Z9TQWbi4X3IKjSOfS45ayWRRW0glpwN/OI8/F0ypMPA/PS0Y
Sur+JY4gq4juXNENBzTdYspKqJIT+C3bNkZKj97yvLfNZxIiFnbj5x68ePH9KIaKx1XUSza57uwK
AkNzDOmuqJJtZYBYpZw5ZC27gqJqRxDpdEa+aOT/ldTJOjN/5wGPMIz1QWaG5YRFM5McqPK+541F
jvjqqRhvriKuBof45ii3dHx7cg/xb4lGoupCIxOi1pttAfBx2Mg2PfiVbb+X4Z5eOxMCmODEezsQ
IziEfW5mbvlmy51ReLD6xtbic4obi7HM1x9YiIlaXN8xlQzP/24pXe884RYBG/D5+eQ899ydM1+F
AnIBcYhTl5oxyZSjWa5x+pI+8j9UbF5jxzrmUPfWarscaO/ho4RHlE0HpHjjBHZ43eWEcn3dGiOM
GkszaQ/K9iYQfrMxrX4W7suOrh3WMmzJsGkl77phEcj/+Y0dZa33cVCDgozRuFu4pA6oIzN79rK6
hic4a2dqA/KDmYZ7jBlSBLw5+jOEfI1nG5+K59cUGca9Pejjb0MrP8OHni+SrZwqSTbkL21vIFoy
YQo5VNrt8m0acEpyoBBWSre93XjttfXZk1OkslJuFDRNaAEc220SelYSi6em2EyIkFsVOdVOIy4I
rIxkOnH5BHfpCOvkjy5Gokc3rT0ZPIPfrzzImO+ZqRXTihZmoXfJs25TTThndr7kYsdG/upM/WUu
SmDUDhGZt590Cbqlbv3/laKXfD3xVEkzr4iALgB0Zot4+lW6ScuMIsLv7Qo22bRjajyNk2VMAUvF
EMlmnxlw0dp/X08t0Ou2YKJAIlWrPJYSrliYJkWic/UktIVNlLa5UCzL6sig0B87b1/j4NVr6HiY
Ac1JNacYm3/t7kwlRwOe5PpD9+i1mvM85FL6k4Km/4do7R0HQLGYA6CpvYGFWSgglclraq+e8sbw
r6QePfITH08v03la3UXSdbqRsSxukoHjsLojkrt32OiOx0BjouYwWC2HmTgUpLz3NcaeIAzUrMXP
ONiqZBGNoaGL8XmDY4kk2/qwgYFdNL3yWhBxQcE058V/nS1ZgunoT6kukn8/Hc8jBWBv/aY/L9Ly
0LgzU7UpW5ff834zsVpdKhkwDMltdtQO56mVmh4UooINnCzf0CZfLrcptVv3W+6eekAZLEuKSpy1
OiKCNd3gRs45CnO2TRVG+rIlXpRPedU6RNILj3+nmZiHnUAy3k9Lno0fAjAV8wX8ocKrteg+5oy5
kJihFcTrZymFjRnqAvWVLehgXOuV2rW0l2WiJxcMMDNt8Pk1JRmHjOPGe4zMCC2zo4OSmtI/iTde
tdagkWNHVwWSb/7Dne/eNE4sc1iGM8YHUPkUAjchfWjmqha4bTem1FaNjjgQ14mhacR8ywSAT2ph
Uh7Ar406nvH2jYIed3ey5XGZ9fCv9f73tYMYok57EMw/yMIMhCvaFnu+1b0RkEg6I0J7oKWUPa9b
mjYjU0cMk9vzHy6Zc4yG1QEIsSk+T6xr1w2SUEyJYeXS587qcB1HfEX/djfgdMwAfhkv1j08RRfu
zg6r8Ks17yVVapduCCwpjVYe3Gf1t9MmSV8h80HzIAhEjqflBDfv3pR2yUFWUrDworVgawQdBaBG
I4XysXNpb8r1/RXDhnCmF0W6Sc9Dxxl9Vu28VzvTcmjsCD9coDGAHb88wYzW7jNbalVU8YStoqik
G1n6rrDkCMDgMb98yx5TmyXUaqrk+DCJEgVulhtZCJgFxAws+RiQ+W/wuE3QYWxdJ0kyXudqF44Q
cmLmWymhvvobruLqOiEPNdHwUchLZJaEzaJzWxpEKX16vzRSqnolK5xxY/TYBZ7nlGPAGLzEnktB
eTjQnnRDFZuWgqF9Ms2QE77GMENlQKjEMD03L8WNIvFgTYwsqe7r4WsbJtbeH9A/F1fdttGCi7Nb
/U7tHHtOvUjY5Ril3fWvQgQljju2D/n2EbeggPnTFutMOh2lsnotkgCjlFl8gejWqALkcxeuGgXl
9WYnS8kzbKQTDpdL2PCOzsSJgzMtS/nfTDS2FV25++KhDmpX1sGRVBCw4UXsBRBsJGX7OFFWeJI8
Yr7yQOJp/WpOhBphAUa0SCAw1m4Y7H+RldN1u10X0A229la+7SvrpPUpelRuFP7tn6JgiEnuhbHC
tmCDwLAPZSkq54XkbY5v8ck9NrZHJyYkdnvy8Uv9dkq9y53jsECaIn+MwqYlA6/vU7cOYOL1hP7w
LffSHissfxezWDItwq0QDEpiEs0gvjcZaAkAbo88CZI9f9AYOGxqqCqFNR5MQC5KrBsJIlfHZiMI
5HvDIkqRLyZYvfA5vt3+SLOfdBhcXsn3ZI5/X7yUuDGfHJTNmnD4reG9aqLR8gvRpugDMWrrqiBM
8LMgr1p7Pc1Ti4Zf6OeyQ4moNDIstq25TxcymctD1B8yPOzDzQufurNFAkG9xv33egL4g61/+ThI
DgwWUys/Ev4HirqTccu8Ku1Td8v3m1VGUJp5KhjdkxmPn5ZA8G3u9OkjrQynRVN2qna3JslKfMFW
bg2fs7Gi8omNR1gRi5bGE7uMmDdlGrteH4uW3ySfU2k2wHxPFSifPInU8wg4c9EKN5HFuLCBfulD
BEk5fSmdXX2V+JpFLD9IMAMAoYDxNtctsryvJk5ezY+3wNnRKniSiLMjx8rmixYe7rR4Rz47Zb4s
dGYqKHIieWI7PoJKgulWagG9NRTJGgZkhp6PG76n09pHawu0k7gU9U0lw+HPEcPuspnueYjdTZII
uOi+ZjT9YPDkhHdCQxvXohhyjThF6yGl5SmoDGyyWvEikurzNUkbsdEr2Sy1KyotUke6DrZbg26Z
idIpUreKT7qNQxEwKsQwI5XSi36gpc/XHcBQ3J27UjMwLnSaS5bRub5rei2h7I6xQpVOUyptsqeP
fFN5zsRVogm9F9NNHVXa0vI5XEiJTdzwCNYc+JJpwZVfWCN7U++BqbSL92cYNawzq8xRuFxAL7fw
rbc6zcyNNDhW26KPK+Z7IDBd9VfloDekE5PqjtHho65HS5YjIRaHsWOfUipNyuo3Jk7L8QD8Hjnh
ni9fjBKe1B6jlchEaWJL7uwaYis92adcBbkcb9s2D/ZhnLb0mvOrQTJ3gUJcAbwUGVCCx9ig0nfM
RG74FWXgPOlbr9uUralyAL/jWd/ASgideSdvQopwHpQ3XGF4gb5nrH6VXXYnGOgVlLKQzJqgvowh
i8x57ouYyavSx2HFA+ywo8ER4MNxOiYffeRxADVgyHyhodNpS5gCnnJqDGb+Cib/gmwkT4NvjIBy
VCperl0Azn1J2HshlbKHaHes6QBpMtTioq0KkwnurNe2I1ZOe+Oa/cwn/CdTiLbMisuC5SYECnEN
nH0kvu5lbEeMcO6bhrcr8A+/exl5/t07/SnfGrHCQDvl8ibvyu4QC+Z8DhvFEKOj8dCHoDcmJUCD
IeMmqjts9O2qvle+FOmTKpqRUXn+1eJjv6r1hU48xgfBQ16Rh4isLmWYDdNQxz7oEPaW3Eo8LL33
cNV87K6MR0Eak/PbalsZ1+TehAV17/eCIvMJ5w1ukhwmySX3dSsS3nUbOJYWl22I9F+w5V/a0aid
RCxErIt+nJ2AdKlEspieoYnkPQJyVYv6iJ1Xa55JDVZF6eBsXUs/EOfpbKUt4XppI2s20QTArVYz
tZ7ccav6WqpJfc2cghXUl+WlCTDF1gGVd2EGii/3My3q1pXMlJ1+jfb218JaoIGqMXKPqYUcwjvu
5hVCBrBFxEFLaa8/Yh4E9TXiS6siLyp1tYSIEW3JiKBsN1YikCnp4WNHEFTdvNUdSb5C9/19fFZu
8BPQUaG7Q4odgpAYWKOj/OjeJ7qdW4EuTnaeC8Xyv7S/2DsTHuVPbMiozOY5zU1R1R2wVYbm0YJ/
Gr+VXSaVQF0WmhM5Cm3/+DHiTBBL9CwABtVLV4OVk7l9Gv4hyrIgNEcv3PVYuQDtCuV25Eg0A/Vo
C+ZZmaNPCm5Viz5UXCi1Ktiijr2LqAIKepNXmePlMo7TBMpJzwvSQsILSgWghArGx0cTCs2tHR/G
I3QofIwOh+mQc4zK+AZ/HZPWgTLT5A/ksBdUoP/7PEMmXVgcL3+3Rbc2srCgHKgHn00QJNwcabDn
goE5mPIfbTfXY9peDNR3OK9mSb7WRfKFTmpXH5N8bgMYe7kzb76ORvQjzkbGbfHGIIIw5TPKQ2iF
8RUySfNRtlATLDOdFtM3qxR++97WXSGLNeBj7ZsU3B+XreBTGNPWI1/sRG6/Lr/VGePbJeTlL80h
66cx3aQ4z6a0riO6A9SmtiB7QOx23AF4qvUQp5rMrGNSgQvxAgqpaAYeFpgOF+BS9uMBOJcv1Ee7
THIQrh7/hJc1ofwL9oeLLQzNONADs44IiM/yne8sc8cYVSb8j+2eWHNhJPzYDbMNGRHFheYKrx9q
XarCAq3kcfdKPSC6M9SVRdfdHatqjW/ktzgHsA/LPEHAs3FaE5bwEkLuRt+eipFsn3xx2x3htGBO
lVZukB0LcDu1URJkB1H5yuoryauDT1LrzJsSVZ4TNVGscZaEZL6OlE//coUedumn4+cwbCQxR6n8
GdPyCIAuLBSkgw01pwyu6iWWj8p7R32wRyFUdJEhNZCPfJtDx9F56viAIBsCF5u7Uggtugz53kH8
h66gFJGs1F14qTz81WilAtkbhoUp/+cXWpN/PnadNclkNQ34GIcq/ti3kDD0CEJapEB2vtOIKtxM
kLU/AcOKPU1MRUZfw0nLT0GFLxICYdRaV9Ca55XRpvkypCVSCetFBG6d2LzFWbUlPN27bYdqKeE7
74V3n7KM74mldvsyP3yTrTFqrJw0/OgCRfa6avzBOPMcnBlL/fvsRICL6GaheTGlq9a3FvVy6Zxu
qYtUXHLaIUC6wB+xOJxlZ7l+qWNlWyV/2FYC3kdLYaKduH/S7wKuc8K9qfBcQ35HddUX6iNY8dEu
0SKuNOHxoAcnQpN9L3FXv/N9tVo0eTVDo+rWh1Tdf3lWmNXCsu6AvAxrRckUaHMuSzTPlI1SB2I1
JE9h4Lj8jsKXpdbIAWDhU5k+wOQFjNgtRV0hbS/yAkuTvwfLRAD/eHn2btINgFzoaJKR7FYKvRZV
zkmqw24VOgK7gZCN3LzDMIs7GBjmI+/GMy/DME0EmfixGqASsWmgYVMkAstf1kkVK1SgXuC89ReA
1S0rvRb2P7BNkmyUKRLGv5BJ53onMy+/eDVU5h859oInsQC/d8Cvfrb1VPL10a0zc7RqJw2uD99g
hYgDgJMkMwGnvDp3EvkmtqplhKnlQjjoEBzbAA4tHlbkoVqA2Q/eMsae025V0GTRpSWwcqnyFha8
NOeCia6+pEDdmmj33sjctCrZfwdcGlQN/on32QeD7bY8OOhMuxh5m0EYWiMuIxjxu1k13PM8c8b3
jOD6DvNnlAuXABtWXfeePjOxZGI2nSPOK5mP1nsWe/om0tFattDwnDM5nTdxWE2yzPU1ZD5nKA1I
r13P6UNRfRqvP6uSeIy5Vb2Ae4CCMxa6UGcEKx8LN3JAi+ESbZi/QH6RsECrrLot3LwAoktWlKsh
d1/wE8cyvb6C/w+NjhkV/lYj4I91zn4/viXEnRUgCT4rpt40XcbGkaLoQjoVncoGeuPry63fNk7j
NgK5Tlz0TOc5SQmXanh7DtFJsXZE6b16dt6c6IogpeVpq+xOMHaXWy9tJBQoo8nLeIS40CGd+qio
2QL2ZBsOXpLYe6/MzeGU9PMO6NEbHIlBrHs1iLBVwUSp4AE9jmnZVdQ+mEthJjEH6KwQcKM0w1Av
QYIMUW24Ubn+G9LkIa0trVPcwkOFMMYI+1bXrW1rsFK9w0SCkRDiu5dhgFULRAMP0j/pLgxPm6d3
s2eECjWjaiaN/Y5iICBDNyRMiJO4weLhYs2KEBlMLMecNdEnmY5FLMjWUoVkKddp2USW7fOQkLNQ
F2Avw3qybOHSW3zU4UvpXqtr7DjFavptbjZkhxmHnQfGXakwZ9L/CqbVV6u2577cTryAKtncalB5
jUClzSHD3fFLv55le2K8TKx3XomTMNQQoUNnBp1HnP4thOLiY8jodUKsOAH1eU/b960PLX6qIByV
h94HgOL6DfVWGdI+SeTrmsC9zN8hzK9UNwCjOnApGale52PrfjtkLjt7LJnv2Uk/DRDdkNb/QQJH
q6fyRxwQTIP3kAeDGRfPtlklZ93TxAC9TNYToKWYL/Cjn7dc4nDMzl18hRPMRox9obuACtnvr1NZ
CJxUMEe/jCyEoH6UurtcMbWKznqnzN90ng6Pu+gPs31PrpUEfzB5Xar2oVOv2QvobAnB8/Y/9uwD
p3Ed0ENvEaRzZoGM7H3OtE+UZ1ItS7UHKj/nzJAJKArl3HNKsgErVIcaribfGaAyPRe4MjgNZLrn
mf38+p8PwIAgmKoSJramMOQkFrh2opYud49mivP5uFGfxqi0NFInsk4sN2YLnFGTXS9uFweIJ2Vx
UUx7n2K3n+gkWdyC5dwiy/AHZGKwNAe4d11dkblnPgoWtZHS/ixrqbhgHwgqOP4yaS4h8/AeeqNm
6JzKmbsDAQz8Fdr1/GXrOTUd6WsJ9RiADUXjgXKaFfzXX+2jc/7SP+haM5aXfCzdeSMH9Gj06tcg
K83ROjL1xnc8Q2l1qc0vBqSO+YFOXnZDiQ9ZfJ1bv+/pVUhwE06r6a1mXT3nF44tDWOZSmrT8AbV
y193q+cfwQJ2Ve0z1ACQd5qo05km9FsNvMMCnZuyyRe2XCp48x+6dJ2FtAA35mzf7R6SeidRWytg
vhZivy6cMf8nnUbOO3XZgc8Nti/1P5gxitRqHYV8C6jhC3B3X7vnGdnlZHKcDNF2XY7qLuOl23vz
0WIz/EHmsgpazrsqBt8b4pbyElo90ljQeLxoRZdBYhko21K+uIJsYBxwWIWVIUzG9jp5OuUYYKCD
NHwKxkkY3JlFGTuLWNOJ17aeosuRAJoxoo80yU6GuJXMCqL2QQ4iwXaup//y+XZbfbuEslOu+yPg
8Zd/GbTmurVLfZilYzGgP0OBi0LZyg5sejqj7GbjWyYRMj5psWVYoW/VzAD1ww6dGbIoQwS5heix
CEE751HWhi38xCL9RKrk6EsqAvYBqnZpK/j0xE5m7SI8C7fzjcDOnTwLJu/LNOtKVph39v3WAdKK
R6QfvcsTBz1VkVb0Lp1k3ui4eiJUawzPfHcEuBSl2jHYl3CVCYktDFrBo7yXlyawB4SWgQz7wa1t
O6PZ6WWVujKS7FWIjnXqeSHMPu6clkMTwDjXxm4FwTDeWSykEyll0zjbdl9H94Zrc0ogHw9dwyoa
SICJUAy49MwT11MNvkTVxfOYmQ/Ryn8xPHUWKpYOYaA+Ghl9wukDkFVMU/jX4YoUagFt09BnnzhH
AF0i5fHJPsN2eRaT9dN3tcgm2DA5B9cAp+buRAhZX/rBj2yy2eG25cyA7r7J3Mjqhst/xLblv4Zp
xPg3FPf3O4UlKATHSmMLbylP9cTXzMpGwy0+SuZ9z+cW73pSiGChzUI2Lb0nMXh9xbyYYaBV6KUb
ZJUcF6d8a9jcNxhyIDWkfOKf2tSPA5PsMi9DggEvoUAj63COi25OnC6YKf6FpnCsGs0jiFHpYvP8
LJvSR6OZbb8+6i35nXl8HayFRh+CwA00HNZsO2ATUNE9KGuMIaQmzTgep54fXYd4gMSRoJrTk7wy
XyXE9wx6rWut5NYE79s2CugqHcgpDUPQt7KMD6qAFITXbLUz/x/IBXnka++j3eD4j25sApqWcr85
5CCiKSh3X+lkm9uaTzrUw4qMhT/VyMgG0Sk68urzQXsLcXUUSTq9eRrQJZ5JeJ13BVzHkXsz7fW1
kFMSvxxjhXFJX0hS/y4kjNElUR8AqMiv2qKgcXWbpKJE0rbN9hgBombYFKgn54QyxaLIqCGqS1Za
1XRO7Hp3bF8zMb1YuUjRtWERO2YNHYIO5dmnbuQeRYr/9yMHgeHvto1Khrf9NQW5cIS5mx1Ex/7E
WzBYYn+xfTZc/+MtDyEshKyqdpJt3d5I0ova7qPviS+BljyzEahc7h5JepyXtFYpajEchOCtwX+I
y/vtYIWtg1ncQpoFizNV/Q9K6ItO1/VQqCp4S6jUw6bTu5rmYxxT097ypSNcvjUg+sP66Q5wDOlJ
qyPO5y//ApQtvunmjC1ZGuzcHQThTmu8fiGG5/X2mkOA6wjcbrjNL3DcfWxEq62FuPo+2YKSF0Kk
ZwuUOcyRueEh90czu0oRt/6jX2TlaxqEDtliHRzm2GDXfi757gnBHnB3ZdTR1CE1zqdv1yFZ+JeJ
U8nnxhKVjYvBfhXmwKj+08HP42e37Nnmvx/zFfOobWkK6Quw2MO50jagixzJB3NCp9VpryN7mHvM
B/19dQBLb938bQvzpAW+S+O3eW0te4nKsJjsYLIRnpv+RkVL0Y0NIlq+W9BrAMB9uEHK1jLxR1i9
2v2HawS3rclhKELK5wDeSKH3a1Fi78hfTOMbeyx5zavrXspYFexfx76UdjTy8K71L1iB2kzrKiEN
7DgpmusY2ftij6yKNdPi9W7iEBLkN4PQ28lc0aGz6amEaERpIBJy8ZTCMFf5hO+LmZSk4vtUlfR1
0b/yRQAxYt0/10HefTPMiFwpLNALN0S1tnfDT+l3UJ7F0iAaAMj03CalCp5Qtr9lWvKDdhuP91gr
me8MaJKV/1XOqQZq8DXeTsV775lyuRlp/bTZKWoQ0gxcA+Ng6F2Pcurh8yezfQVSSyKhuenMklVx
NVoD4kpaIQRdXPtKMN7PrNKNoP4zIjWuRFeKjlrOCy9JxGWZ/D0SZWj1s86jDLT/LLhEJ0dAdqmG
utzIX7dQptjopJ7JHq4YDK2ZXs4EiwHAn9EjHcmU3zC4ubTCKyJJsUMULmHW7plFGTJYs0MG5AvK
s72nT2TxB7zD0oRg5ZEhfyG38udG/7dV0ffqli/WwMko2NkwkjLfTFQh4mLfggrytYp+wJgo0YSl
DSyh06/om2GAW5z7wR8RtBvyVTc/pzw9GF2gQBSneZ8ewZcbijNymRrVrCdtbHIP/pf+l1SoiRG2
daDmqZ5pnlvE6E3XFfMVI/F9cXSwV/nKkcfal5mjf5FelSgdmixlz05mJAJBbyd778mB58OAiZFj
QFzQ8IuUoZbcmOB6ZWMU709rMbddMcN3qrGO39OjP4BeHIF3DH9X4UWXF9WEFHull+4qXgZCF198
3w9uj1V0oe9R3PL5oNioZnr9+WaLeMmpEBWh4+mtOfmI/3jE0hCg8L0uwyHpfyu/aet7KzVIDPFk
HrRURHnMQK7eeh/wuxt5g0zqyapg+avg6FhWchBNpnQYPrfRzwfNmwIZ3Z7TSb0BW9lOy1A2p0tc
+JAwMnDjWYtIY0SgmlueLr75cPth4MOigYajQmafJAJJ5HlhCwt2ezClZ0kHLI6Nc7iocOJOzh/J
L8V/Pi3epiankEIVTnObiySKAVos5G1hL1UZ+ddrL9FbRExmiHDwnLNnFr4Yz24BdUIVvVnKn1nj
otCpiiWdA4rd8bLGC9b+3hTQkngUKhEBkyHZrazjIpwyE7mUPamb2RUR+TcfRFpvkPjEiJYQaxqJ
o6k0OVAic1ZjJUYESrb+nP6K6f0ZaQJ5ia4u0qakKz1AuS+W/MqoM4HIwGFBU5+YcgeExhi7GSwL
jB27VAzkex/EWox68cwCLYcWPr16U0I/+7NdrNCEAVGty5FLuEwT1g/Jm+FSpSEUUjeauodRMEKA
6E3Pa+AEvQjNvmC1UziWaPUpUzrsy9ByrEzBPNT3YHls1Xyg0JkqCwVB95x7ALBck+Vnak45kNaU
qyGr8eRx1417bWW0cG0SeZrlSXHlyD02QDAlq1yUtogqBfS4qLSfnm3yYTLx+5ORxmfsvq9ems71
6q3sHHzhqINnmiBPhdNizYZLcZorDv9OStKkvjD4LJveJui1x63Qyn7C2xi+/6dfsvVOuBHgIgwX
WiQJSgh+bEgoEX3WMm8MTlgKiUpFmkA4j9t2x0y3O21LHpoFhx5bYxdsgIlT1ELdeiJwiSwXrcfb
Ix+C98neo7OkY4T8AaSu3dljRiYUpTyqjyAoPuSXpUeSWMbcikS+vTcz+0dg72pBSM7A1/WQWKY/
Jh9oYK+BOddFtvIiiKl4js5NGnOTdeNfJUxRnOSv1wI9MWeAKmBBl/o42GLJeYazMexwd6t5fUTA
XIXTfFVLxd4PZ3rT8dd2J413BgY5pKEhxy7nfthAS8rU/97p5CKFd58CFIcEepEN4e/Kv51BBEZ1
4Koax2IwUdzDR8xTVLuJ0ze5iEPTiuK4G3NN22PEXhY62D8ng/XEyO3J3sqcS3beacI9k5k41JOA
kZ3JtB8IXziPmw2avzY60mP/7VjpPghdxj/3YAa2PcPy7YZRh757NG8q8j3guM9CRgbHzfGek2cG
lB2zh3kEafZ7r8CwWOGoSXWBHk82I7SLRCJCZo93wQtEXB10A4ipomm0zy6RWJN9jP24g9DbXcaX
ukI0Dl+ALvAeFFPAmdwXELUK+GeQYGb/ZGdK/rJiDINkrcXZatwv61Od4r1Wpkhu52E444jOzjEi
zFfkkLy008wT7kjz7fKKL170G5R5pLk4mjKSfRVls+kXLtcnzxvQkIYXqrYLG0uVinFBtwC6gpLF
jQR3Xd7dkh+Ye/g+MEa8zV6Z/+kx8M0PhpOy/vZeAWdWCDq20D76fR5eeh6rtPgd2BaGa4m3xjxJ
UThLVbg/YTGgFcuuc62/HhX+88Q3KB9+SNyS0jVMRlr2xCOtVYE+AobYOqCuIqfoSqS5AFrfFgdA
nPLl5t57LWE5e8E7qj0yt1acUZ6UxYCLy5VGJ0GReIamoTEFivXouAI/l3Dtv7tFcZbYn3a6vRd4
dWQuzB/wdr+INmty/tWH5C18rcjrWBarUPJRQ+II28Pqn9yg991ayvyNhNZLd94k7qA32cUD3NRb
lkJQdx+/mVsW+RZq/i6PfSfgwCKu7W9MmwEL7uVPctOOTfaUf4w1r7a0mcvyz/Z5l5EHl+chqt0P
wnuovoV/cSnmjKyf/T5NqdQHhQLqqs+MJsXFSuHAGUJYwCn2Dg6LQH9sKGdp71jG0jGCS83vnfOv
5Mey19oejslG7hc+0qM0LnwWBAVzDestk1YO0lLYI/xax1DRhFFmD63jtlCSxD1dfq7vJlhF7Bq8
pDuh6FoITN1sdyGQ6FL3vAnBiEVXQgmGNvEaCkXRC3lcH6Mxh6VglRCiBlyObPR8/wd1N6XWVsMI
E8LP2UVldt49qT0m/3HJToWQCBIKewPxMZSA7q4+gx3HD5PPJQ2oojLszRxVbfhQJQ+MmUatXPaW
NsjZhqnwRQ6ISk4oWoICADQKXsFWAz/u8b5SD8FdtNdgZLiBqCyVJiqFySulrRWdympf/+2RdYKV
3We3Z+zItIZ2v5wDoPhlepLEwXGk/OGsGFYaCbR63AlERc7ElA/W0ME9ewypjIS0Z3ABIsqMF5Lm
GmtbbVqlCtOThdwpVGDFOnh9DrXozeUe0eGLV7Uac43R+xJ3Pk5WcaSFgMeRPQ4Yl6GFfv3TdMJh
RMkhsQ6/4903oypRqVfJeM85A/VxRY/wuR7BqBEHU/b0ADZJN0FmvnBBmeSiM+76J0t0tgqU1kEX
NWrMgvU9wAKIgSUMTu73CvuTsWpkaRqQib/YmdSBEFFv7T2vseiQbYJltebsTQtSMF8+bi+yi0ie
atSrhpWvwiEcyohSb3MQnH8jSZHp3BxHm3wIgkZNhz1qjHyN69UYUuIggiNbGFtKB4vxjojgiHU6
qzI6BXV6la0TIM/YfMmC3yk9QUU+OkxVKqZqYPnU/+WtHKMwzXobhKz3SOvvRXBFDdVm2id5BtRl
nAflQX7gOzCCNwclnx0g+YhhDZoVbe0As8Pj3EO83pKDwOWOAmvdJyOk2YtYmybBL4LERgiiKtZD
cZw4nY9Kzi1lQ5F5uNIMnhQgJfEPzjucpH+XTouP6iFs9ap0Aqo1ar+uqAPGz0dUEffUEpvkJeHI
d8J3RvOMVaGkVil4RSX9XmpdbEKFTqNO/qHzVCU8MEMwvSXGKcz7EgkLCN+AyAkxV478seu7ujM9
7mgAq+8nbRiU4xR2nxscQZw0nJDpe4zbAIuLeXEThUy4sapmlGgCr0XKwd6eH/xuF2qax6HO37md
y+msG933QbcFlF5q/EMKAdybQdOsnfkQYq7v/z+kAVC9hkfyEzyxzPdX7qNgCLq/b6eRXGHdPSIS
HVSTaT8VjbZetHC+alH5BznYoRhbAMltH8lOM1ZXG7WTGd9b5lzqpnYXWR8Ys+wl1ko5LhMNYLPA
ck0O4dTEKCKPxzUgKetxROTf+zGvPV8FrkEQPd85UXSzgDDPv6cgVC+uBiFuc+aeC5EljAVR/1UH
PbtQu9I3S1w5Hrto3ClRWeKTsEq3TE796cCT5rKP8rkS0Ds6MAo9LcegiCyIO0HLq7x28IQon6pz
LLVGw2/GiYBd1sPtubscMTK3rShaxGL8xRi7yPEG6w4Wgcs9Qse5SX7iHuz0ikKyBpJgISzIiq0w
guTquvzz6bZAd5/hAEhLu0B2NWtHpNK2qqP7KUEBCU4OufEX6sZ0N6JIjDM7ZrrCaVwJEPnaMLyW
NRJVRWxbrhJEbTasoWRs85hBtcLQ15wY/uJ4BDhbE/tTASZgNR4ZTbdGpqxFTCrsetnvlXt5dVp9
+XxL9FBuS8rOiCgwdAZuopLXXcq1lYQFYJb5l2zrGAsMjfAqNZIhyI2fCVA0+QCTmM+WUFCHMC5v
MBlXF7dBr+37kTXJVnCOQ2TGRhph4TDMLrSxIcdRaEuweJENFL0sPrzTEWEl14Z4+y2J2trl1MiC
9OPB59kbjwQZOPmveg9F4xHQDUaPUGaKjkSOHucsfX3S3CWX5tSGSKS4d4jbrBdMaB9w6jPLCcjp
UM1AZpT3edFFB31LZdgqssBC2cFPjNEqsQB3c9M92tR3Mphm612i4WVvEn/Z7nJG+iWQReWT/kDf
27vP3pOo71+Xu0LrKIMyxk+6q/4h3Ru/4G1tgoLSrDb8do4YvEmXFHb+93hABTfaZn/WB7rsjQlQ
sjD9qOrTY+m9ffrgUdgRBoL2w33SYb5qIp4iwFPl8dSF6gBT8NDChfod2KvmHM0IUBvRhgp6x6nO
8lHyxFJ4FV1Vueo1ZtAVehupoNnLMV4utABAFoT880u65IVXsNP6yF3JCN9MrbFmilGmLSJtOWdq
do+pe6gqxJxx70E5gEG9PuwCNCldAscltUI0O8POnJIPTBD6AG1bFpRthATgVaLG6gK64327pYQy
YVh0vH9ADFTnzOQembWkarE1ZWhmEU4jIiXXCphf7FZJDyY30CCKFmEBhDmS5+s7YzwV8605tYwc
ALMIL2wwWPQuHAOTDOZ0G773hYbg/y3xPfQFMMhF+kDp+SdzL9bVnVw9KUVuuphtLBif6FBsTXBt
QXKjHyONfnw/LOwYyi6bFxT2U4/Lbe204kdMzqhlduocb6O/a6NBS8xsTz8vpRfcaq43vFRdZZ0X
HtVz21obDwmZdL5DJP1fYOwvRT2cuhK1clcOn5vRV/gUsfdjrxQcdfAQJupTuSAptA7dRpEYfi6z
BP8aN5JTBwembHhMBUV8aRG2BX0ux8s518pX1JBXxY/GuVHNOoQVhrevoJZW/cYzYlsAMv8gyRAV
ezELq5mDP+E782AiMpQWqrsc+kpYiOhOWxNi+DibedFVkAlWNiPHttS+1Nvi0BspNheiHAJiuC6M
/oOmW0ZL/nn/L3sVdf2uoTjMSQKheKkEKsKD8PMU3WEk040lvsLb7afFCO7UWyebLwZ5+w/Hl7PF
1X8aajDbAxW8oCEcf/Iz7vcCls3ZNNA5sNa8PXduosINqTM/MC2PPD/jmneH+ZStQv8oYetZnEKZ
XvBuLlOq3n9c+gCNQr6RXLN146MF3NzuxeUbrmGXHGqOMPQejtBDCINCXRVx2XdSqpEZuhbtem8a
xP5Bj9n5oX1ERP3HJtMZQi8NGf/vxXL/hBAczUDA6xm06Cz9pj541q7EqYV7/KNexH7kVjNUzmcr
g3ews6d9JMPNa4mNecqJKOpEuu9OvfFRsZuQVvrwULkzFLG3K6GcfGvFyGHoFtOLo60IvWJeuTka
gqESvymG+rUeF1FegKLxPf1ltJuvmk1KKtnJDsV/PFY3xiuoNFtouyoPRWKQVd8wq2RvjG6ifzt6
VyZPhTcSzQw2CACsEkC9y9BoCjV7PsHVOh20kkBj2oeH3TwXdB8kHC0ZnO2QGAfWjeJ8KjyHrutI
hDhlUF7PSOaUwA+kL5/SXSFmahi5zbYyOkkiOj1GwhOXwG29ePdBrTwdIbec4mTV8nhAYe7z+C38
VRCI07ArNEawmMlbCfVi1cp6J7rKbw10y8sgv+ZmkOdO6BbuTIl625UA34FvMi8I5A56W5dtXE0E
uo+3ZVfS8xFrv1mJg5Duziy5bVLiU0WTXYc1dY7m/esbfKTCfh8ASDjq11YYk5ZEIWp0S9sQ/C1m
aci/Pn7E/gbI4scU6cDIgvM6ghxbTOTa6oVdHAj3Oq318uhAbUdsj/S0Ebgb2w1/q1btUuggYRgf
5LD1kOiVX7QIcEDnCxUcSKrcrhaxN2dRnSaD2S8AjgvLdy9RWluCNkw0ef6kaGLKiswjRm6couC4
YXE7ItDIx2EHNFO1y+Ea+6bCQA21noNw6DoBQyC+aPni/4kmmVLmbLunt/ZOSaZ11TxbRRJRTyGq
gtEWzacbFhfoI5zS1I+wIoJg0VIbbXOPEymgjqhIgq4u6QVmNQxMamCtwvbFjA80LrCyh1BPYgZf
J14o7s9+Dkjcg2gOfCIF+e4WtwfuBjjFs39PtI8Y40HB9L4VIXBebrBWjGaN9L55Mo9m5p/G1QCy
S+eTunAXwrB0an/ogOB1IYv2Rl1VXhZUkm+/yeFQb7UvMMfBZFyh7ec4Bbh+dnbzJu/EBHZs8qgm
SEJ2jl62X1XeWgZ8Dla/LhPAevW+igSQ3byqgA6Js+KUm9xcdyuSV08LzCBD5gRhr9NvNpVqnIOL
2+Dm0dTa7bETsDleMsXzVTMyJyPqyoaX4+EIFyMYNYq2kOweOtaoG0juo8m4f8EgBYvF+SLWkuJ7
Lf5UCcuGDjT8vziSCQ62naHpE5YFEvNf/MXN1oaY3r8yOmqFZ2SVqRJ3s5X72ILLfnrC6/KDRcQa
naSxBKkIFlGd7s1XQhkG7Omlaq98ClPEPc8K3y351WZjmOu13a1wwiMWgw7m9rmghOMAo5LdIPZg
h9sWk/chGqaADoGAynfH/sSOsIQVZYg11rAQk2uTYaL1AUTJk4dKH/l6Bsd+DePkycNfzFtHLtrr
PndN94Lauqf+Rhrr0rEIpc3zpGOWhGr+3STc0cajlD4UDghPgsWyQtYLBSXZXoa3468iyJmFPzoQ
VPEVpjNV0uZ15nsCetb8O4xJmURjEU/b43fmlVbm/j6WUUXdavUrhwsZRUyPg5qoRusD2x8p8Ftq
7Gk2VpfK886z7SzwojCmjM1pj3z5xTKXc6c0ZPmFWJ/yMn09mOI+no238x5ZbblWllHeF+0VoZ5s
d+/MoTU13Mwvd2Y1IktgZPKFRN4VTAjBgujTXBL4oFRngn1Vqu3Jj0Sqyq2yabnXsEc82ehWHHNG
FX/TMIxOjRvIFtAuE+iVRs294orugl0nVEqVRJoqyAAd+pNTyf24N0Wn2N3tjKKGk9uVeCh0keA5
maKULivGhvVNCvvYclsJ6WLQDcHmgT98xFex3q0z06ss+4wm8Q/kL91NIodwvhi6j6Fjyg7xTKaM
lrCb7aFguV4D4dg0Yv4d29M2m8+8SCl+ccYQb2BgTM75hF/r+cdtlCbSweR1SHzV6YAUXbWTpl7Y
fr+tU9zRtqGemaBCA4wMWxiENEfjCdWyx777sKyoQpSYZsRVV5dqOh/axdrv7PrzKhmCrhpCCPH1
7MpB1xtrVtyCacAi85qg79mvzMvpxl6tRTId/l2SwYdUhBjPbpQ4fe4xvQQVpUAHL2kAajM3Dt2X
byi0eRYWZMDaElnyOVUjhm9IyItSVsRXA6hMqdrGUS1/cmnPUvjq5DWvwe7VzmfPFQkFBZORtgeP
eF5MWoA5sZRgGbkD+oXGs6dIeOcT9FQ2DWEZZ6pBr45hBstLShdJkvAxaHZ3HzruSOG+JeuINImD
oau8v3OlfNLs3u54ifHaf4qyvCKnmY3Lq7YqFvvU/C9GWBIjBiwrY3YCOs0I8iE2jY1ij/zp0dV1
SvqqcNxRVDV+dtvYrG+6GvyhcsI76fLnkxolwWs0/uWSW7qQKlTwM8FCLIcIgCWWEuwc2QwqvGqy
nkNkylogtAfmJBYoIiD+n8ZI7Gzn6uyN6/n9uaRCMJwmBAVEkS5Eef0B2WMfc+yINPMmz7VFwFps
6SzW7UDoRcHYHpQOPFE4Dz4Puwv58AobcmY8CdDvUQew6X41K8GbmsmNPGcEvofxiscO6qgWPoMd
C8FQ01iM5pGju0R590ldVgGkH6aORJMktC08Nga6QuuYhukmgaF0tn8ywsjxk5PFqMDZwtWy1CaB
o0Dul4/X5Aw9UJDBD26CLrCTHinxSGBjAIvJXX4N1Mzhe9ulnOxJ6tCE5Kfapc99ihlctnPG6RjI
pO0KCgslfI6l+psiBZwPoZJooRRz81yEUVnmmBBsRivrrBFNPixHreug8Obn6kgHxT7WmJ8qk1EJ
5N7nacjb5NpgvjmsPOhU2DY9cLVdqHdBqlQR6HkZOk8gFMtQIwgLXA2jDjgC3hhTGCiOFIh+pEUk
LoTtZ/PP004KBYkSKiqU8hTOcEECaA22uM1C34q+1UhWjhwqVYEEcq29IhyzRMs5BdqZ8C5hiG4S
GMJwTcjuGlw6RxK+4hfm4M7HGb0PS2xdJ358EDJdZVWLrs9s/AqQnJLPn2q1JgFbxYha/1DcfuYz
U2jAa8RI7FfnmM38/WtNkgU3ZNSN367Zf08hhG2RfjJ7YYFMJntzkha9wTYe8XqNaLf1bdV5TQ3g
8R3F06j/pSxT0mCgwKfUpFrDE9LeO6xRo+HUBfK0l63AihY1Jp+XjSMPORNBnW6ZDohMGH3req1M
NvzRgu8hfhZ7pDsPc6jeT1+LdNv9DLYiwIZRtfKkiNs9em+dDYSyGlHcMgi1F7gEshuixahsX511
weCp9OvTyK4KJ+XnGR4dJfpsrdL/MkydPbHX5tV8Z8lpVTyPbbzGvH84PGxUiSdN2VBN7g1bxUCE
L1+VwTBikHhJ1XtyXRlUau+HjM1MFLFSsIzQN2RWholeZ+m69GAiMEUfCpGr49BipdjW1U0t9Va8
6GeKB6VDUZFuebMyU1JmmPs/BOrbn76VPLN6VNeOkRSZM7fkfGbsmY03b9/YdBBgdcNkgQFuEoxN
6E//vnjmK/2qWiKMUOLIP7lO95Ijz7tdIEix8fiB80J1uR7dwCQyyp7qMVnVZBjFKyxtUOR2vde4
zcHmcV7QR8p9DC7zyNVzl/0Gc7GmXRPQu+Ra/CZ5xmpYUu2Gwk9TMXOaREvQpQWzQXNmKpVPVMvd
LQiZ8d/ttE5LIDS0UcLor7ch4HMO1J98pYE1gXDb2OoQnl+8Vbb+45RmJdrkoWYsmt2NcwT/IIfo
CYjeDws0fsRzM+RxnYZOCvx08r/FdeRcYl0/Sh1gZ/Cntybsu6uJtWGxr47XWpKNRiNWDqxnFSWN
WZTX+jD65YTMpM9Fbwl6fy89HG/bEBpbAhu+7+Xytodx3epNItK2rTfdp5j5D4fXcEuIshbDUirF
sgNNpIl7UPIyomlBgS6PPZq3k1c8aVcetkdLEUNgPwtwQ5Hp7B649T1nKqxK7VHGPIWSTIxZtrGH
kN+cAoLirnq7w0hLn65buVaE+wDUJkAoepMlMADA6xvXZUEtypS3+fd7OFJwpeNAGdqF1OBSOM4X
CBUBJsGX0nSDn2GpqgMoJaz19oZGp4oq1f5n56BzFhT6oFWnFusY1nPnZ9HdMkEa/09bY0O/G43r
AiCYBrXD84Sh73Mt9qWhaXMPCwCyWxI9iStQ3sZUrjGFKnt22uPoTNpy1U/od/qGmEpfYaewkwCB
vk0BQ85AkIruSTFke4IJRBofLboiTOg16iLlCB2Jz3nGOZhFm8m427zhs41ifArQV0eMJxiLAs7u
POhH20htMUdXuRBm66QNs/FOBHCeWCVDIUakMgzTffpDBPAsInx1LSzbh6UUz4PNjnSvaZGAthQy
1EEQOBHe/rSoaU/iMgBUJ3FXF2es2LLI8tUc6Vuzi2idhahJ5BqK+4Vc1fhUAEPcLXdmjxmTTFLT
kL7hVGvUCpKpE8Ki3A+cDTKhMlPfDzwJ6173BdNrzh3pPwN48q9VX3c6LKP/mSoggZ3ILKGecqYA
uX+1+33H8gGkNYCdKHv448tKfw1MjpctV/LE6++3f4ssjUukkjQNxKnZsyAT+sAes7tHNcscIXIf
E0bbHFpvet2WgQatAGlsSlQ9Z7ZBTkymUkJNTWwrss4hL1YMPfMvaMaHVkhqeWm1PdYUEAPjVzPv
OfPhEmGBMNE7cRQiCml2qeyrE9aPQzVFFu18AMdY8DJgPsyyGBHTjQKHN1G0UmhsSPI5JLnKLDMY
9WKnlKzedTY2+rdwGq8fWbh8vd8iAUbR/hsSQsKYEnG+Pakgow23bQldywaoHsGbMqSmXFlqn/Aj
iCeKyJ7ypnzsHl8HxmM3iaqmM+a1BN9YB8Y1qgEkTh7PzNxUpcA+Tfb83McyNxYYNry0cYYhkH1i
ZzL00ehBgrfs8GHFIEK3VrLJ41ZMGaXFduiYl0nHZlcEvYasVaGUVFb/kADjltcbn/ZoELhxpwjy
FKsWlbiuprau5st8FY/2dCGDvY3FMYlderH5uBMOQ8zbqoWWjlbOqWBMGZKkry5teuDJyA8hSDCS
oiCQGnZWaBv4oVJ9CKsrcZmWURk0gkeoEZxGaK/Aw75KuRGV1LPwkshGfUf8WKZ8t1ain3Xvb9oC
XefoiwuOHmbkdIw07YYsS0Tun4duryndscXCcjarfKmLdcbnNU1gCQyThD4O5ImEw/hHEJOQBQeq
UrSpr2WMp0yV1ZHASD5s+hLsPmCBDWe+AjHQ4lHiqxbWk7kQ2jwseyGZB6+Ecc/c4g8/fzbBmOHM
rao3qBmXLUSDtlwfJd0ws23iieXlyweyT1qUnxfrk3iVkjdINZYr8y6LniPsdACqCMG8YSFnx4kz
vq1q1zlpZYOdGQusYZ+e35XWapUgILEpo7WtbQXT+AoNHR8P8NC6dkFk6TOXLCshTlVITeRF14IL
S+9ezBEdaDv/wvt12KbwykdUNyKeEKYUBU5oKc7SwTKZ9kRFEyTta/dV/8V+3SPgaH5sDKohGCQ5
6iG9HUsUXITPW4E6Z4CjWLjAnAv7CCg5iSLfHYqNStGKRLrn/p6UMiAY7CYEnCvR2+wrFKQ9faWV
T6gmKvy0wXdc4InBAqIfohT7IeoCQWWflfcDhFH9vUBNngBls3KS0GU6B2mNPtNdgmG/cVXqhnZP
IcjDZ+mbXDjCgWt0DOfWR0FNCXAiG+3Fp9vEypEgV0D+/jD3+Za2g0uyXXGwLscVajNksdjzfqXS
VwIUaqNiH8jRK5UGHWhu/AMDiUQWIxEtezXcbuauVt+LnUkqSIJjsomx/q6B+Ya8Z71/94mXWnVN
oGoAEzXRdGPmeyrNcHVW4Le0KrlJR7ehLsqBBkjtBkOIiJoc6GgHY/bUEdVtu38iLI7Ow/6foAsq
/jysZfbIA0eQHheb8xgIMnz1Qj2BfAFYR1eACDAa3cS/1AEy9KwNpeqgzC4pL3fb5UYF41mwL7dQ
HvcYNY37aD0yBNODXmGPcywesLYtSinx5XqRUrK6sNPffli8lVnVgT+js9qOBfPsJIO5OxcH6vxr
xGSlMVbM1A1EaH7r9p3ZuVBw8QyhHp3WjBZ1qclvdWiaY7L7dmWgFT4gpb37RS6LLyzsj432rogL
2yEJjNA3OBGGGCNsgZou10/2Gcr32Z62QFgfwq07dJlfM9hH74qg7WDgudNvif/dqyNFtwELKNpI
pwcVPUYOufiGxAiU8R5BXOOWBZyOygT5nABn0PlXlKC1k1zUC1OoKBdZcubO55hlUhRDO1xAND2F
nufAhYlCss/KQoQ27rHZaGM+rhGlO1bxTBXjaYcbQGJVQ7f1vkQtnY00mF/oRtIb3MBL5BptDDye
YQLrfwmueniPU8o3NplEviurh2Cm10U5L+GtaJBvHrCyLvdIb3PeSPgbo8NizcQkJ/24aEzUkt22
zRm8XmQWhemIQSYY16atcjQWdlQU7SYtUEKVadBiSXmVc82GuPQavEfGAII0RzZlKQgMN6iDjtIp
eZSoDzx8HKx2DcvG566/R5EMwGpjWPlgRvdKKqQfxy0R1cvZCMFSvxXuV1TO8z4ziHfff+SAxUnD
VYqLEVGufmamQTUU9NKeDHjduT3mHmXanW76OlOQOwFmcpXep9qVEQj7SZhL1yOqbsjdUgu5eqh1
nlmhW16lVdVg0J9Y2n8li7n0wt1eZl5YxDb1R3kyZsJxzPi4NLIJL+rZOumkZ2DRjiiXo3DBXLzE
+cLRdFmRH+JllnxXQEEnmX+89lKfuePTFFMBavSZ2+e8Pd61P9Tp/U7sPpEW+Yw7pyy6dpId+Xe8
MyYAPBI6ajWHj4vDz0aQJ3uO3vhTyIPLcK/mYXJt+/kdFoqRRsvhVSzjk98QMN2tegg3mJFmLeZO
Opiyqi6Ht4ntEiCkYBHaqlzOOHYcD1bueAGYS6ic3s4kJnStg5OayDpxXVQZ2ojBAEOIx3FSBAiV
watxPQDJ1H9Y1O4WHYx52NFRA9gpLPkLCSIVfm9yxWMVwMEM1N4DX7M9Nb7xNU6j3gLiRhnuXF+I
LGtzOFzmbvbnR5CVc94F5UTJPcmvkKhz4nwvkvR15Nmox40LRYHG+R8Z3LIu4aNOJEuEIFOy2GSL
XKw5My14NN9WLQKUUJ/w5A8xk9ZPnmIETwa3iLtrLruEnVk2vIQq0wNLxL6v2GgVgBEuTuUWXeS7
3mdM7iYW3Y73/LIFQmY/aV1Rb1MHqhpcFn62pYr3YPhLi3ntDZcRqOalRyRsgy8ZQ/fxOvyWkvak
4l7iAbwOoL02I80GKXVc4CztR0Va7aJLu4SXMXcOU4EIg4yzd41Dl6Ikvt+IVN1hhn3JGQ2ulQRU
PcpD1UB6dYnhQadRB5I+cyL01l1Su6eaTShJEji9dk0Dc/9rWymnHL9Sjy0fGYviYMHaJr7s5Hid
qfpRSv7v0IT8egBrRrf5sXCNVmrFIi5ffVPCtjB01y3VkOXBm3699SCdyIgeIjHpICZuRhGF3TY2
noX5D10uCJkBl4e2Vww5ygIp9Vh4okIZM5lziY8xVDvYNuRTxh34m7y/4a5xYMY5HBfZOerhXZq9
oJapH6rBnh/pSV0BEyNgw+yVp58KlYzSgKtQVCrX+EHpg7fg/wzZ/PrneLsmkeyMvNEPg/wuf55h
Cp5mWrTodF1f/uo6mi80Tq+hZNf3jbzzYvuD60nBZYsJa9XSs53tcv1FcRkNALa+GguSEPHmQOba
vsCY1Y8bjQsS/uvpCjvRhLBEHSxM6MPK/gtrLX4xJkBwDMyLCqPknkpmGQZBwOdpP4SGeVqbs3Ls
DNFRLoA8M7b+NLFjni4M86eRQ6058TKXtW2ZLiAGyCol0wzXtAbdVcjeLY1KW0hP7xvwzrSTfNjl
/TBRFxZDDE9vSFpQFBaVm68Nt5sA43hvlxPV5mYxh4a2LbjiJ0fYE4QmuOAs0b1exSWXncRCOtFF
aJlZzuvp+abpwy3juWfFysB/+uBDtdXgJBO4xiustvQpRLsoWur3Ny/8FWbVqU91fjQMsuYEA8UI
EHZTORho1kNnqnLwYuRrCxyTeO34PykKMUPZ3cmRNzsv2oRAYvc+yr4CBMHQiUDayVD/TjKuPoTF
gnIVOUU+53yMTAWs1a2Km+5rf889c2oNW9H6zms/w2CDcfGmb4Dgx7E4Lb4KVSYJEibmuG34PBXh
/5yRj26Vlqp1OGFearAvCheOyRzqAObIWbkccTsqwPDCPXn9jxAzoH88QwgqGOlZYBsKTYg0tk7G
5GlcIGG6c1/qcJ7ACtCHkrf89aseMDFdvavmHoPVII3JQFPO7phy7f00v8DZVKcaR8Xk5dR/r6Xw
pRY7/ZEWZpZ1wnTpc/gUs5K1DhqQ7QXMBU0gwmHzAgLt1CpqIlB3Aparq2HiohHJe7wrUqRt6582
L3hzaCYTkzR6RXN8UErgLYvJUxP0zhaOqKWNRhPAb6xbjUea3+J5riPMB33HocXQHZsDRSxL+rFB
0/fuDL3kwIpOdzkFhGXcD2cCxojqWa5j18z9bgjJiA5aX2wiUyw1xUaefPnsDbt5L4aagmg4m5LP
+Zp6TTrQScV7P1wnMBQpUQl6am6CQMxiTep/FGp0mdm1EleurOGTJz9d2Md4rtYMVjFvKizL8dxe
fcBmD2BYjGAR8XPx6ylmaGJ+Q87x/o6v+7PlcrPzoY4YwGog0JtEmizbSw6DtjXgra6ZwyR5XKcv
vyl8mdTNp0YyXOu97Z9zczbzC2WonwbLwA9UF9A5K4dLhnOnF29k7ML1A4/zoLWwc+QlWN9HY8lk
30YW1K9H+00Npgu9ziu2qIyn4rAhuRkftCvCIzI3BQaQ4Kcn4rmf95L1MSTyJNdS+NHfSs1w5buz
sv46MDER4l9s2zkiOTsnihc2mmig822I+7JfBa2wQcSgMGzEeyobT+/dBHANRsbPeckk+tN/xnaU
XZrchJz9Y+MaNbS7W1zTFb5R+1kjHbcWZTWeDKSuxPkTy43i1B4EPniLVJ3g+p95FcYoIg1Uk+Be
ykciTY5PRy5kQaY8BrWyYhN45sXNNa5HRA/GL2xgCk7s+tkEup2kqWiZ+NzE4nE9wNa+X5cnr50J
BHEirTqShWCHqNdxNgYnL9rogdmgrFpLoC6KkRrQs39KIWeHYRfhKpwBALLDk2xF6U5JjjqHF6k2
uimXMYmrJ3bkDGmHQbvKzwldJaywQBbmNaRGVi6DmLwZm6XzAHcuuW6GXDgvDmvWWadN42QRZWFe
bw+jJHKE+m/up/KarYLaQx7LZ8+3uCGPcQrC1CCeQl891wUof1A/IeFelZA1jojPpx3Qw9qSdEV7
/rKX/asH9+2KY8Ug23HNnwEfXcAEXxdYlX5lAnfOoyDEwWHcnYlJuBOF61xEw6Ey/s2FCOHgBkDp
AIf6T+n3aQ5ZqGWTnhKZJCQ+nEndCofyDjeep4MPZaWDj6pArf0Q27aM56uYsKodKCJdJUtXM22+
6P6nVC5mYGBxmuOTde8P6I39JlLjWKT3FcN+0gYU7/WFyQwZm3+bn+aY8ALUB92d8VUhWVd+1IPX
wAotCdoBE3lQCzaFGDcv/jceo2R75vwj2tRbmLU5vbsASoIHyXRAtaV1SORydVr+m2gLar+Ik5nB
G3/skFFso2WPUtZoEeFlyA6Mxbavdl3tALeZWDv5C1X4A36YkNdV81RR+LcyZGPnLNoNezvzEl0h
EAjeQquje8AnIQJbTbQ8daDIPBwCVtN0olBit8i8lPtd9+iJfrtBxOPEYrFXLie8nz/2UOZxWSBG
EvyZygBu3bGZV+tTF2WKZFPVI3sPqPSyXF5Ovs6oJfoJ8Ne/8LyHNDkJyN5wEE488EiD065ldmcv
AMPiHurYDxyVAT/WJzwmxnCbY4QunIcwAaH90ulSgPbKONnXeUtT9KBUV0JgrOi3y+uiRMX1WiI0
z5h6XtmcWbXwGn15MYJycpdNWFjg8xbUA5Ddk7+Dq4vpN/iExom+N40q/6+N9RLCY9QUHwriEo+c
U9HrTeOJAZLZkFb7GbFh4A02KO7I5+DuY9kUqwKeM7FIjgpVzE+njHG5PItJ3uvN+udikSnhXfxN
0RxXXxltzGC9ei1ZxBB1n2flBQwEQ99gEF7VrHyg/jcx7NWK1e+HMa+Ts8xr0liT8dwYP8I9ihfv
VTUZlxUHhO82BWQoB3Lied1YliCMG3xED4vcd+mvvJJfgwQ0doosZH6mpePPmkomxZkYpYeR1KMH
yYakRtxsau2/tCOmr1g1XmU3h8xa0zR96Y929WcmnsjXyV+gne61A5QQhhPb1IRnYPYVIGSCXfxM
Jnq9IBA2W/pqX9kLjDa1Yp+QuYUrmDGleXkZjX9y3zU3QW/cuwnyoqfnHdYgFJ2x9bHpcV7s8AZm
gmoWEiaH3GvvPvhM2vI8BVIWJbaTrqnw1OJb3Rut8Ap6xn+d9Jkohq3008adF9QpnIuX3PiGNPQG
MzQbAnI2li1GHVVN7+hIDSHsFddrN7fvm1+Q+wEZo4/fS72fj3rr5jpUPwT/YNsxfF/yunmMDbEC
FExx2qRkQWkjsAuIEcjdo2J+WfRr3l/7sdhCAaM5VkWkfyM9ZDfGkZBbSrBbxMsJNyR/AQgszYRR
krGPIXo9b+jZ/JmcspKuFrZTwc1XUfBVZvnHoTvX2ou0Kj1cTOInfKan5sNNEtd2CYa/cR35/G5u
jwviQknWwgmy3/+z75taIhvkl56T5D6GLPzklm5PYXHhltH6l+G9NHV85jK8S/IXbZtX3rOOF2U1
79JoY4jaEPt4NhEDVnDcMJjeQLH+ZX/J3rFKUhCcaxZEwpPrntRHeZUUTwjndcgVOZbTAeY2S1DJ
THlznnAkPQ993GhLylBkkfGkZJ/7Kqp983mY9VvVULtiv6pNBC8JhS9UEsh5+EN9qQQuDsryRM6c
YNo7iHLUEQh5nLIS7wepdTTIgUaPX4e+vMLAUG3usTIvLdHnZMJpmu6D6bQl6utao5qwIMx0htyN
4WeA0jNSWzaMdGGbjBK43dBZUxN/IiuDMyJokBBU98Pr57HA8hzKHvYwB+O7FmC1lEuVN9MhzFkU
KosHjNneISo85FduWuMTdAL7yv43r4HaV4VIG098bGMwpnBLDndXWrdv/JrXp98TosXtEIcbgmmo
DfBtQOC29nDg6X1NQZ+p18J7CANvALi+cYLgOahSsEnqjTVoLvc33TzOxsEvSf9H8Wy/6ItrsZtS
Um54uAh3oz6624mFlgAYne7yljzIVc4x/vjDzLfjeNOuTFjAP2BindhNLW4RdbyvrMKWMONnPnEJ
PuJD8lprPHoIt/8ULpdS9dBtCTW61+NWq65HQlVyLXpaaMVC2O5hvHDwe6ul9iKDIzZIZFzrs0eS
ituTuWxzx65qtqI1HPBVyFEclFo7hO07gZN0sk7DbiUmOn9Izr56eG1HhwPZkX1CxaieDr2EwRvx
opFZ1l563wJATDzh+8W8nLxddDwcTF8Z/cI1Us+FkrPk2aPVnZEK4TV3tgHG/8ZojHSJHch0qH34
jdE4jG66MlSUb3T1C8uK8m+Iy0DZfQHVCDelmg/zKc3qhjHQCyhV8azXDOj2GethU3MahesFYirh
YvDbymChFPj5+YV4RDEohyvlbjl90RtCtEafVs3ZoS5XOpbWibgbrNnQK2NFkweMiXWmvmd6h/wQ
OgmwFgN5nlz6x3JV55/p0Csox9AeQ0EEDeZZQAXpL5wS8Gx/l6GPtUYoIEC643Akm//x8G69t8j6
VUEdqnR/Uia6pK4LBhrXD7jE5grs7j5NMSBpvVg0/kML22h8GUFE5ihKzRsvkQwEZrLYMp9fK+gl
DyNQ/vTcLvUtgSPueTb/pB7tKR9RHVvuQ+TqFtdwJbiB3+HKmUiMc6xyM2c6jO3cUeoRZnIXw17y
y0TvycqzW3bjcDN5j3ePdU9f+RJnrIgC7HWpjT0ZjjZz2fqt0jzuwNr97WHdihQcMmY/kri1vMF9
pyB60k5KWaLnpbBC+fFjyDpi6KcoAHonjVda7nA1J6xcvBBVlDISMsdwe7/9iKuw/kpehdxdlbH8
04OWe64BwNnRNN9c6Hpgqeam6kzh9Wr+uS+UQRB+RVBrjvkCYD/vO+rHkrYd6DkpGJmRRB/BcEOq
WBjzdNI1bQBQbXV63o8IGzurvyG3BDcSLFTGR4HtHEm28QlVcoWaAgrGA9dKXcb0Hkp0Kgrsq3aG
NRz+0sLNTk58P64Q2+jTjQZ6TqoOf6HToTpjBOHXLbBxO6AbT2Keq22r0HinIDTz2jrlKf7MnHTD
nrzN89GfGntK+rKBAWM8vUpFN4l1Tyx72CAyWS+fW3JWwOu4jchoMEWW1GLj0BFKwPVZJAG7EMUK
ZiDKk92P4PsB0qlNvarZWKx/UIOUcH881z+pAoXBJeJQD5/hSZbEF1t0w6wncDHYpsoxkPUoKZaV
LxncTf2ZD+hvBiDtgbXayk0n1wgaDX2/TESovfAKMNktrm11k0OYZmshBAyr0gSvvwluegulNY+U
/uSr1cGCTQ61IaeDWUogden3Q5jk0jP8PdP0mC/SYdTJrk6nicv59LbsGUhU0yhmri6q8MhAEsTI
R4JOQrALm2gcs3oyQSCzfeGoYZJuoldeh8o2Ag4OeNazkMfnk7oPI8mHO/oJXtVUGYEyz7jvo6kN
0hL5i/UH2FC9Vbe4lJb/2zAH5WmXJ+YiVKbTPJU8k3TE2+Rjjwe42f/jmrqwicfmlbY2whACqbe/
oRnGFTGYehRv53eWO5ozOX8gZOC77W4El9QF3WbvB3tdX5fKkMilf7oiVhwG8IhB3e8KKv2Yefgr
TuR1b1Cstc3j8MEBqRRyS8fGt2O7TeQA5aGEwnJEupIhlHGtD+Sy+WgiwX7mlzoVXJYuL0j6aF9W
4YPXc6lWKWk1+rWXl8pks5JYfcowHO/9AK6fFRlgKyCcUWOehKTUlW80PwD1xydK0YLeXTw4CwcN
Ec61rvFjasSV4qtqJt2sPG6E6MAgZ6mGo3HcNdwovBkYjow++0Tr2NorSlaxkjtpUG9cgjLWixhF
siBw7KzTXJLmqUQ9JDga5Vt8Pp1srlYMBsy0auu+C3b0r1WcQyShkWRPJORx2vJm+M4HVxQSaglL
fGjtbOYtODVz8z/0SZAD/zkvrCHknxu7YbbzIGJhYGBxFV0qFjz4E1IZ4zf8T2UbDmR0zt6ujfTg
kYbUDhj+5COg5UPOlsNpFTFSHzbxXjnftxgkyjARJDKzjA72Bc8F3u1K86SAJZ8lO4JQaLP9mIan
B+fZsT4qYqCytPgF0Apvr8yFtf5oNZJriOs54IfoBKOwAit0WckBo5pMwl0Oj+opLqBAMOQ0qpm7
OzjBT+HcZjxDEeFjaffNf3cXL8vaBowqBJa5QFw3bcSMOz8n/CEs0sESa+/IAExxljWlHo7/nI3d
+ikFYF2XgPistROvebXaRYyPF4ItSF6LzBStTaW9zyn5fY8XG9VfX75BJvPMtbxCsfjMlCps/b91
jdxrbHNsPavV+fJ4J4tLzFyFIO/SuBPZ5PV06ucmxqxCV73rDP8y9gAdlkYbanqrBghXXmT0h/Ie
P8mk0XJzbtpN2yXgti6Y9xyZGr8zrcuTF2kmQBYp3CvatR02pNuATggulNaO+plKBNy4E2au0VUQ
jkeWo+2a28CIhlrv0Ed8EEse2mE+9pfQ4XKXAoIsfjk26w1EK4zKyGLkxjhxyVEN/d4KtXvZGkCX
fnqWV1LaJ0PwkPLMyPI7RogCxjCWUaonORSkp08Pg11OrTX9VuQBplAGh6d02dus9DXMXEzm2fBs
IaxTmUErYIXxKvRBAJaApvjlX5YElJqpr0vsBmUbG0e7wKZZlQyomcVMs32zUvVVh3W3FU2j4ixt
UBLoHpx19k0GoVEIpdNzC7kW25g9JsxCq6CmmANHpOTdcRl5QcO99iBhk1m0EtBxt/y7ut6RIdBi
fJRgL+P4+7qDHvAu7oYOHgss2bid9hbOfKtpqbv5o6nz+arKMBmM0VJ6JkvWKC+Q0kl07Zv/FEe7
iRyOVgFC45HjqhZdkUnZKJB93YxvOKb64vVjkrKrG0jx4cyt2MwPKNZBQk/VZYOWltI33cButtQM
AtYN+RcGsv/gQO+rr0P8INn0MMedKswfHs4sSswT/51K1Q8VGPlkKD8QZ17HpiJXY3RhXvn9+yrG
zfJOo7k+H0SXcJUTlZxFxvRHrf8sajAPxLvUaMgndZo+opfUUY9X0TA+2BV/cwxOCfVMBRhJADRa
n5tNHquhDCYtrOtCUCJO2XNCMFu/djBpIEnOkUAvS7f5cURxaAQBnT8+2STTJNOzoENjdOP9iA/3
cp/0BmrsdSwyQbTXO7ZN9m9DjqV8KIzwrj8nDTav4MbT6Cn4TIy0B06JDRcPy4mN/elRMGdlpfYc
h9LxXdNj/ecjFc54uhBd124DHPRfylXSKFh5itS+9WTSiypVMTb6ajbF/IBnldtJobvqdI5a+G0w
JnWFcJMSRl4IYoHLDuNIOJ9/qciMN58JDzsjrPanILHtuNM8liX7gmYfpTajAowoTBudtRDeofVd
AiKlpy6UgERminX503o2G/StEccSv1yRmk6MX+E3BBpWDhVy2yUTMWwm4G3YupCsm/4B0SdUvnpB
jN0TtDujZWs7lCZ1crtxz80cMHJ0QTqa3CZmjAhkbvDrp1ca4AIioxWteQiUIAAZ3+wMYrzqPnZG
rY3e16iWGAhX3vWN8L3ipR+35juN6FSt1CT/iWKyA4dtEvmmQTIMA+SlAPO3KVRkx4bm3UoxyMet
lm1NvoEe1okrZnBxkuL9pnU8eZITQrEu2qUW1s2Aq5KJx1eZWip2fAYtldbB3mWNh70Rh0iVHiUd
mHEbWyIBv8Cn7GthlGTptpIzE0/XOfplXEbUhAJO30Dw0N5b3pdyIzARQ6ktX1jRujKRPuDOD4lZ
SZqSVfASB54mJ72g6O+1Nknjw5maIH9VLPpnR/JUUUhPziNn7jRv38jZr7PCs1DNTjDhVDvzWlxI
MKNHV1szQUCAojm3jD/85gMbDICnZtN+/WrIbHocxnkYWQ3R3rYflVCrU3w1MFg3JWMedHjg+mY3
sHqGj4W7hg+AZE62Fgft3RB9jclrKXJCVtKcD89MXhSU6tH3/A9SMpXKeDV4LF2NYpujE4PnbGGr
eO2vyV8K0Nk1/lges51CNT4DxaD1ycvRTak6kg/GWdUzVJa1tdOOVe722mecSDJ2L+VIGH3awxsm
vUaphP1zAde5YQKqoPE3kMHCDmnq1msezLN2Mi86zCMWWXQBG14Hgf3/FqV9cb2z6FG8/HIKfID5
+WB8BSoOhAXL8qboMHUz/rsFdW1y58ed0O7iJDCzbSdy96sswTmulJKn2w1XDqnlmywwnXcYp0he
33traTh3iYUGX5eHMq8oQlS0F47jYqeEFc7xN5W82AwUnjA6mzIphdNpZqytfaPv+N5+9E9DLY/U
C+E6yOXZNDf7mQ8nKeeL7MIhEh+tB3EXC0HtNBkBC3wRh7Y3LaCWwCh+4OdXwmWuqYl8Q8mIwkfg
UxZ0/5NaT+Z5pyKKP7Mfvbid/mcyySNbVyRLR3b+G0dtWDPiW78thKNfWe/z2ZUZGAxR6GKpaka/
/rzJcIxguthJPlX9+1EcV1r2YZumhd3WP9Ll2Qt9ljoOwcTKZQ/Q6R9/1wmekZ6xLG2QbBcX6I8i
ssIab6joDs/85MBIYPWP+hAsb3ycbY/Mk+h6FT1p/5SFYCe+d5qYH5mwqQoRsrYOodrAQBQoaxQu
rbpdOtbjIQSqNVM+jfRxahYJHf4ZhLJ9ZQQDl60RslXGZTwfi8h3uHhQh79RPiz0otMxVtl7vCYi
kjLxe2zq+y8EZ+O7mY0NKMAA7EvlHS8psWZO8makIrPyVmM+HfKS4qSJaTGvBj9bRlUhtU4bUQ/1
nYptBgDT5RaJIy/mZN1qj0WQAHIye37tmM6qgvXY3M/ZTzi0Z6qdORbs/mbt63jWPrxZfvhTJHix
AZj0DtAyVWkgBpcibkOZ2sPSegXh5FIAvZFceFWpE1s29wPKKQJso8H9K07W46VugaQMcx/YzkTS
IDt1AIIT/889iUFhdGL5JgzsEmkXFwq4SagnTnk2RiHP1qPA71EDjG+uyKqyqx2uezf802owHHvq
YaJV2XTxEPqaCezwRIIJgcIj1POEmrgXGhdDE4xW9daR+sTXf18m7+JqT+xJHymnNpiOc1qh2AdM
vecR1QBMiKLXoJzHy6rdQEW5MxDiEwOiNeQoqKq+n7xwCR8YAfbdytUKTWyiOczCzM2c5ztSf1sb
eHyujgsgFp0yLLNRBvEAp63hIKrRgZzCh5D9l5A1h12wFCZEB30kWjiXkUGwDH74fxg+DPzUmW29
uXs7EuVsYy9Axrhly5FaDEbGe1mYpOsfDQgxzBsSRNnJdGHHzvNdgNYxN4vvwHVaPn/W4TDYeD0g
jFSv1vmI+CfzO5xA3pz6lPJeb03Mm3cjf4vTrtPVV9DV/7jgNqeJTQXF5RRVb43A5/P8hDIvpW5h
P5IlVCSRvIaMxFP7t85hiFMuYbphdUT7hrFbfJfkX0Huel7FkgkzSELi8MInXkdAeQ7o3M+T27R1
PH89MQuS7ivdV8C+x10QFrKQYzgK0kmPnHMUJycWGQkJalMjtXZQMzwpZ6z/AfYBCY+c0E6XQx/S
q7vQOMtEawGgRyrWgHtylhEKTzkjQbqYuGqjSQAaaHXdCqEB3V8EpmpSV9xF11NetEEtLWOigKW4
xSIP74g4pCSC1toqLpwLWk+S09+0phAFQt7phLcLZBWmtU95iL+H+bBo4DbxEcn0dTRZQz2sL96d
qP4tpH7AefvptSadIXWN0RNE4YR7c/+jTTXb8Vx9/T5IrFLyHABR58f6pPTmlz8tdGNdbySdFmbc
IuiQKivSBSt3JV+RQSw1L/S/sGYONV1xg6aMNlYEJcJZGldCslfgbD5tInr49P9YbPbfhOrjKita
gaO6yxwhq1F7DKcQUnnztheSRIVDcYosjil+B69X4YYi9CnzLQtfGOrSZvBCWyc+uCNwrbG5A3lt
dfXgzPV0QaxR0ckTw1OHoyRfyCaXXSqD7CuLRuyf13AaNQF6GU3qeYLB7vSnvsclgjOA47GNZbD8
ME1B7fGD92x9jITV3WkR85y5IOS90IY4Z+OalZWdQn2iMNcf6wZpqAa30+wOGQ8zXOmZ1p1YcDvt
CXVcYAP4CyErQFAgOq/AW90q0ZdgaOad8tBhGW2JfzkOVrQ+69JNjIGmtea7Vwusg33SoeC9XJqT
YUIb+QePA9iF6OuOEtigczJR1XQF6xiKhbB1OcZhE0oU8ZglWAahae6IYtbY5v4esrOpEHuTinNJ
S6uuO3YaTlQxf2rVqObW6ree3+HsDSN9KYkowNGPI/aK6WxCpKuDBb6wOXaBIn/93dMg346kVK8/
f3a8wUlOREKwVBcgm8CSeaekI99w2AqLi0+WBoGkKaRGwqpYf6nRg5JAS5VxZFfWsen805Q5jUU7
rL1opu9e45DAcemdjluO8QHI+F+vq3sChMdSuFez1yCK6tIsa4agylj/dR8c+E8fxjZtxcc33vwg
JwCvvMJRrielM7Dkkg3NtzkzplYeLgZcu3G9gg2mFMJ2Oy9R9YGGOttLINanmnWS0xhuCdmueQb5
GF/XSeV9uaCQBsNO0u/NTJXMHqgbT6vAtYGpxl15QiJqN59uRPeEmvPGu11QB3sZgd0zfTnTAjXG
RMkA34Cxnw7REcQQhRA2NrJgYuIwFoiR4+98uF4PjK8dr/XsisMosC+bw80MtH9tN7jRRj40vlsD
CyYersvmW8pTuyix5W0U8W0QkVBUbPhxflvCX645F5/nPXk6ygeAWHjjba2sOdEJO3t9gCgh9T3n
24vJNX4QoFOzcMVBVh93unvD7oLR6qwVrafKAK2k8CESRshy01wDPpKlS3rO9UpCVbIIB5u8syZF
c82lFFPfG4tJlt5VYcF+SlmWB+UmqRDRsU/rpc9EuDDOOYOsTv4kYQF9JE/nb7UYPwoh4yLFsJ+q
PYpTrxwk6hj1qpmWWbg/HJKU9ig5Ic7yP31fYdgtz3OtqNge1SZCN0v+dGqQ/TX7bnzpHexUE9bL
l6HJ4Fcb5wrRVftRrtSrCJBVWQxbGH0Bq1qZMcgrfe5oLMMOFnDjLBCKX+tgEw/2z6/rds27kee2
rthCgRs40X6f1l2RdXaNj1d3CNnQEnwLyeNmp+Fw7JZwD6OijboNWHWMgAg5Ce7Ma0RAdZRpCgf5
rvlZE1m3s8XfQfGhjb/s/LyB+FIo4n8utAcZq3yrvri0VhkxUeAM2205ohJ09eHHAmh4KUT4DXyr
XE0XwvSCabnXYWp+GrwQzggY4WjeFUhtEI8zLbIGG5UmYaFebz29IqDeWewDhBDEXeoicFS41ZsD
A6a4WJR0zT0DEs+Bwik0nSVfQlRVrO2GPBJLOanpJe9TiObkbvEmqODdMHrgmUl6ghOm0Ykkkhnt
GAI0yIxze8ODO7bJkWdhOEMKjB4+VJLlvJrxcUa+uogMDjcAxTn7l1b/NnlADUHKX2/mJHLta2Bl
oAOakqYF1Y3r9dwLZ73LmaffcyGC0BZf+Zio1tAmfpVC/lg+JvKD2kSyra6tVJGVUYu+nDIfk96h
uWvuMPRR8QL3ExKknffdRbvYYgsQiq4/B1HtCoWqG/UplJqp90pk5X7zBLojBglvUnqBICA3xZ4k
FOeOaYPgJmBWEwH2hRJ7J0iLFDONjThjF47fmaaMjG8LyOLUo2648HUzUUX7wXbwT/ChWfFi3eZR
aTC6SnoKh7/bvoc9Ro0DsAE2m//C0SEMviKX29XBx2tc3hon4IdDsR/QmSsyVQUL0VsaV2ci14gb
hI7A2bt/6wuLGHKzxWHuXKC7auZWyi2OFa1HmUkOgR70QJ8jNubrJ+++oSkV/jku1VF/h5fQWM8x
p3juaFKxZ2BHGn+Irxq9klMgXhqZGHRUoj2Tq7UEGwPg66ZUVevBEmEbnnTus8Fey003zU8jpSUq
hJkXG0gErBu/5MjzC6NhiaXgcVXCjMWIh1tihfIdrWNJ8AB2rYscRsatMBTq8EkuKNUxMYV6etdg
oqI48yVpLcIDe5+IzdpDiv7/hUPWCJcgBfLUVZ/owxzNZb2RF6mb0OGRxiJSVMsaXpPSRBTNF5io
ksmJGoPciIzJbyuYeQQt6BsE4NYVW+CAL82qscknfaeQ25T9w2X53ilRFxvFNvNtnK+mJofU7Gfa
hvgdtEQOuUvtr+W8aIT0mmbjYKr6tpOBsj9KRKG9pOc5Box308hWO84dqaEgCFF32SfdYQbAFltt
FqI3ArHbk3YhxPWkNbcgVDsA46svqyPIYsP0eS1muGTWKtOHwDFHmbIZsHWeyMPFHpP0rBjiomqc
pzebimtPS3IMxBGqN0G6YeoNU1I/hZU4yGH7sshbedds+6pGwWjuJF6ljVm0IRfw+RG0wa4fFDz5
BLf27rfEDSgHw7NthzwRBHaBZVsUDbPY03cjvEJjD5o81rPg0D/roTzEQOchpSz4Q0h5b2JZ6YR0
T0AXztebmgU739R7JuBwE2WlzAJ+4vIeeOabC0NcsV1nE2c1k/kFHPNIc3sVT10/kJ0kmezusbjk
5glQnKoaWrk+UEMXPo8x141RN88kl1mSmviBJrbFPHRb7T0rGtWs/6fDnpvqnBKRUjw1Yraw2Bov
bwcbTER6gwl6hpTJVZAw+4HPKInGXnyWBnUXkxSOiYzjnxyC4wYcz9BLKyYSCPa0N4CM+DON65lE
wf18f4QPDLMz0cYdlauqwbfjcz6aVVZi2q0IQDYCxs+Ax6MhhUZL8ZItz36iHQiWjyT/ntDdGN1q
AhfVZRFwaeY3U9CNDYVQKOOlp3WrjWSi27j/+7QH0Ega5986rAGG7DuBl3AgrcxD7D1UnoU4dbZ/
lsEkFs23v3MWZoOEAjprEEtu4XoLmqL/+65ORv/aoGDBqvm88H7hNKnZ9hPT8/j1TXJz8e6RIC6L
dgZQUceUiVM9ust+J++oZ91XSGKKz3TSJDCFUoH7/vedZi824Deh4qD40K2RlDD0xEHFzMGyHb4G
keAYJYBCJ9P7gHkVCmyqIwsgG0H37lVy5dSeE07fojTW3ns0s0NkT/kr/N5AFGrexT0+4D+6+YO6
oJcMVOrEIiF0lg29oc7NQVlgGWp3tvuZrw9HA8NPNLn4LAButCTaxm1iAV0RJIRiP1kFgHzLY1uP
iJROdFjPGAFXF7GBfO26BJav2ZPVMczTSqvfbXUdy2pYrJQldj8XLoKaiyYvNR75+hxjHzpJk237
wagH4qWp7+xzjtU/jSwc/b1SkxyvmgptRQjy9UY9DYmagKCEgUFraWBX7hE2tuScv/3LRI4i0SVL
RHQBHpBTAybQFfuIDxJJ8FJGGJVk2uh/HM0bCQ4Wceu/5UCcroA2/6cnrQiEGcXsbSiOGyytCJtY
v9N5LOSMTuCAaaf2Aax7ITGOOvQO6R2K3Mwa1JqMm5X2GQFphuDSK5SNF4o8iRZOTSHFFcUhAL+B
dj/mLfX3kquWR4Fln3YF+u79zgMBU157VrAGkTYipJ3s0fNzRevaYRSuXwYGCPHEvo69ah/t6soN
tHZWli2v2oIsWlJ3hQ38w3eeoTvLzhhWWNDpdqKDr5xv6QU728sgQ14z3bNB0hh7F/GNtbpea42Q
OBrnWcGO4Ft22HBZ3Qs9WmdykOs7LFbp8e6vsrT4tdraxyPwscWUIab6WSsPJ5l6/yD/CtV4aPCX
v9EyvHWrX6MdhW8CRhRGFRJukMyaA6zBOgxCOjmQ6/4cLbNf0lHGAsAYjrp84oHuQfCVtF7Clduj
spbj58RxiPHeG+sDQb9Dkim/pjcQl40P+SfHu6C3FeThj9hGv3mpfpQdsBrA81VV+gPxkcYpbqbR
DyJSjBdJvyP+j1MiC12+Lck8Fhc95hPEdR2BLl54+daG6DTOj+c1l/SUD++xGe+wlWPzeNq1Q6Tr
a4b4G8Myexc7kc78VZbaBhr+5DjzC7dbvGHjjBEVdDFNSmRPCC7OOTjCvcFmZO4LHShPvre2Cz9J
ODgG8dJm5eP6518JZXa6rR28ShQu1dYOl+Xt0R6BJ4wt8kUlchXgUx1LVgvl8LJTNCW2VMty/0Fh
yC+QowRHKkcTGeruDWR44Rpf8rKZFBINycDvFPUbLNCmwWLVQH2sYbjv5Wm/EA1laApxfPLXjF5L
2S4xeZf/8DVIwpWbO/CVqfchlS74T//li+aBDKS7Dd27ZfrIrTpjEUYMRrK+FODkIysPt7PfrVnV
rPaAdmthV0IlgR4efeJO5Bi9McNGsgO9yZOsye4IYP1hWTntRjG45dH+PLNiAJVdP5kVdRHZE+X2
zwYygbtZzdSTHH71cCwEjLjlHYuN4v7ywALUznxoN9cfHrrnULDRtjt1VvtEp30g3Erbms9paaKS
v7nzFvXYQOhNfSIw6wQvYyeUMh0ow4PshdZN5Ien2tiJD1VZPsg02hS8+/JTcwj8tL90AofFooPH
cDQVsO8OPjexkUNnI8tDYKViS0XHs3Pu5V4p+2SFXZwCuULbZpMvwUSeQbzA7VUIS3mlQncpIFOj
O6Ve2SVerdBSdTFJ2NiVAxxDH5mPOI3q2rEBolxn7ZaTkRk9qF3lYlZeiAQTNSXIQQnUk6pyKPTP
9Yg8KUbfGLxt7fqs8T2NgPq6r3TrGoG5hdbs6y2yhNa7VOvXOyvutBXoyhrAFBDh28vpRiIEtpuk
1XbJIeKr3hDv7kR7TvgFyJ5hSogzslNIfX/4PPeXf+Ya2EO4LaNrgitunusoxkjGpNj/A23Hl0gg
c4dwq+xN5wA06uflSUJD9zV9Z/i/nhZcHBcLkG/9toyYRRjfEHOX+EmeEks66ifhXooEYM3jZtUH
CslveRFDA1j32/2/VIeEVwcpEw6vK8C2JJNDfkHpvTfceOfTJ9D7qJy7DHwh0mG1WnM/CPv6WWYJ
qvKsEszQdjlJd9Rdqe0XLVUjDJvmuX/U2j8e7E/S1T8hNp5zjORRn5p0uc9R0mmVxa3jUzYfrVaI
wfhS443gYPKCCR/A4g0Cqokzse7JZuatQO6HKD9WOE73reFAGi3gX8dL00aJpfpM+39RrgikP1rA
uR3lLkACOgNGS6NgVX5i3S38KUTZSekC8AwQGkbwSo+jDYIhlLDC2fK8SVoW77eurgqlV5KW8r4x
9FP9KpkIsXCkeGiRC5Qz7ixIL7wmNPvw1VeLyi+PH7WjlQ2zDt0J8h1v+Bpys1LFqocuNNRuFbu+
xDZV3wytJ/wVhMrbatbxMfjYKlz00Lhi9114Qpt1JO4uMQEtDI/xghue5L46oieKL1H0i8eknvpo
iT4mL2lmt6n9eD1TqOf6Ps7HaY9j6+abNXsIDj9p8b05lEiimx60QcmPJlu88uK8hHVWPg9rl7ba
gLQz2KQ22l45RtCFjQcKEGezeYpuzQZZMFONSZ+i2USQ9dkGjgLPaoS6MFbcpgjMB6/uonM5RniA
yaCv+HM7DvQbBVz+o2Y0WtYn/L0DnHxBXuy8l3r6qChQ3sWcueOqk0qOBtus+QjTcEpt1WZ4CmJS
tVZeQucmVgAebq5suQdkN4TRrMCZpg3+YB+GMetYzfuQVH8s3u3ktoVlg0yUYNwvgJxq0oVpjW+y
0t8Sw4UaR/6j9M/aAA2/J9nNiXGJeNAzQ8OosxM6VkmsZMXtC4+4il6QG98mMfeblrYd7b62ngz1
tP35ouS3uqsczEMjuo0KkiAe/LZpuQ9bf3m4Ghmdej/4HjYt4oDwy2aZaxtBM28VErhhzHTN2Lex
EqMCMC3PGmDcqLru1buFziHZtCrFGKjxyfK6o8dkrkPCWwBbUaCpTvSrHd/Jipc8hJSLcsfDxiYP
nFP/mfLbFEBcnvUIkgGHbVXbB9yLM8dD2pKsOJsmE9xyUVuHt1L1ptH5mgg0s2X3akUJRi94myBf
PXKQ+9KGfLs3y9HX6haN71jy9fBBU4y+WN+S7GfypQXfuvKlbVQ1Eslj1m45hboU20xBIOEIdQOe
/pZeUgQt5gS4jjj0jt7Jk+xHA5rWKtZgEVKEhgtWTXm7sRgLJz2NWfUPoDvhiKquXK03SSB/60f0
YYqm57R8WLKe8i/TB39EOej0R++26z6kYmkJdWNadgeKlGs52k0wqcQao500Y7PrgYuBvq4fJzTB
V4E+Wisi4GokvAZskHloLpbMS9WNgAXPYzRFIWfzGlWEO7v4NsPhzI4ExMmQlianzoTuwzA4XVoc
7MvZ1YTJBOHsA6sA0YDN1SvkREJ1NOXoBeJJ3k11vKRwj2yXByDq+O1PlHXztgD3r+G8hIZ0CwFl
BpSCSZhsRKNJPiACmR5d8PPHONJe1h6NmWRJFhXSxDwhZtARldt12gBMciRgVnoqfPazQ2YSb0nS
VPVF2lnYz8sIukmIhkmZUfQXAfldwlXtG2ofIG63KIvd+8UXkajwpzgtqsEZWz8I3vQswxpzTUQi
E0u7rag5bsZ0NxOjlZlNLOVnl1VEuBt0vNKTiHJPT4erbIqm8G3FRPhAs7xe74a/5S4fxsyZ2R+f
sUXwntYUtQQ69zvq9RlOwUkzRVYZIUe2p6kmz5Q2p1SbpeztAefBwhLXU3QoLENDyls99OiUFEIn
Yxjt01Skz4k4Fo9imub2zObSC9z+2KwaSAQH598TA432gcIthC1naNH/D28YriyD3xkYt058vsdu
850I8tlEA4JnkwsX7mPXIhYi/uU6otFfepRQ9vxIrPnUd2/iu9qPDOzUS9gRKNSQXDud6BjjIx9I
moKFdYABgbFOfyFY3ZNc2MrNhnZkmOKK1yH7etCgl0a3W95ox+MDfxsgkT53c7El8G6YYQSsD2dr
jKys57RqJ0q1oJssLwaBQi0JM/UgBwkVBeb41Uz6RCRaMWf0ay12NtYrRbt/FBNUrx3Pk6loeUPm
ECM57ClXzDGR2YiK+EEGzMStMD+u1fHH7qXusk0e1TZxsOwNZufThOldtoYPMWTIIBR8tUL/g8+7
CMqovxnSCruLT36G4CbvcvYIVzUB5BY2x3ciqV8IRyVvkpKpshmT0ada58i7Do93oyLCKxGlziyk
NMMJn/eVXn9aA9eSI34y7GfJcFfKcv97SD3+ryw3Tnu3HBIWY3/tehxC5opctQv2Hkgp/ONkhULO
0XgnxJAhzmdbcMmtFYSWNJQxm8AnlXtqGLxdOVVmSgUB1c1PpHU2sPegnHO+PY/JjwzE+eedLGX1
tzYbOdNbeG4VlQWHaGQrcvBspA7yQCwd03yzy1Rc3HJnNTPGnZlK8yYfvBykgzqibJ6JXRJ8DnE1
rnGINqF10JWqMClX/nHyO//UVCJYyPSLEpwmyi503WjyTcdf67UlW6M47OSPPsuB81/GBvURZh60
qhuTpstvMitFwt7VWHOmb5RQ5PM/Iq0BeuGwoMba/GJ2WSqySoUJPDE1mJ1+4/hkibW4ikVfeRa1
WfeIvLqZumLzKrflDkdXTh2Mwl+fPlN+uwPTPRe7v49GAQeRmLlZZfjXWsnp+0+87KE5paVtHeDB
PlI9q6orMt4/yoj4kJ4+f/fQonq5Kx4SOby05eWO31y8LNZ688mA6PRgOKCF8TMXrUpNoAbaYCvi
7VTlLKMk3ki1FgM15wN5h/7WeybiGxCa5dPkOtm4tPYuZd6Dml1BW3yDqSwrercvruS5JV4vdExH
bG4ElAlOspL2c0sU/4K987qfRFNOusd6qYSaVqYxLO35eKN60ZNoEQjLza9qZVUr5oX7g01k3cyt
rIl4LfF+K4mX5luLFwhxEUenrKQ8Qji+fa2s5rMmdoeS94ywumTIryyJud9n0HhTJHR7zpBIclUW
QaHMjoKafzk3dRobss5jPITIv+vUF9Y4dihy8nV0bqhHtfZygo8Z6G+CXS0LEgrMx0g4XOJ3gASY
YxoIFKtg/ap1bmfSHRHKqpZqfouZ/yjJOlDcFbLeh0GZ5iuZGm75T0QvoHnWcZqMLG4JOX3TTE08
PSEigYafZvKK/3Z6THZ9RaglKtZY2OCVnTnpjG3wQXP+Dy1c9I7Hx4Wq63vBfizfpRYASIi40TIw
5T/0bT1q89GvWvUCGHd0qVetBLpeShbr4ijyQXiJttJbOQ9ppI+4rsHeMBT6hn3SMQJ7aO4MOiBa
k7+vP7QLh+FfjimxCne21XwpzrKS5qL4dxJkfSHARDCJ58qCPoZDUWcWxJ9e5on+Cei9Sso/2pX2
RkIo9YAlNUEYGwpZHGlqlVXysLn8/nzgsJU83GXXGCqJPjB0gWXGsTI+x/zr27HlOAIksagIBROY
RJBWg1HZhkY5uFBnQSPG59ufJ5fej211yGnc9q5DLYazAjJziwZf/ISatrTnzJSj3B3GXPFrcdRw
9AEOr4tH2bnD2H4DOBLpRmCHPXOqvpwb5e9ovewIeU0FJPVL5WzYpIIFX+c6yhEpw5gpoycNFtQd
r854fdUMccxIImj12mQjfXiPgqQ44fel1CF1RikeF5jN+yTS6/oZ/IQIRgRq/TzkIVq2z5K9zJeA
AygYNvU7FDIGFYHK46YGneYQNbZs5dEo+3LCV6BxlIJwtnVQ/QTLrVcgRCF72cN5qrcOjxpqDxYg
LrzqRVrxX/0enbxqEN7Ptrt9VQnzb6fY5c0fRix1KB1mwHbDRiZNBMY2p2HVq/qvgXz95BaNHZJI
xBpxe/+Gu2BAWGYQGay//42ilW53RjGmZv6CWZ4hKDQN18ubZbkcTzKSEmVFBPcnqvMevFEEc/d4
Zg/nEWyWT68mYDc6daLgTJQpL4d6iEQOC7E1K8nNhpMcU2jh0MmkVpHhUU7R0KZqY4OWZcA8eyrp
kRxMCCENkKad6qrdRRBuh0QmWyfyzeFF/FpVdSNFrcgFJmxU1KedfxmrxxIvQ6W7artSr3cHs/c0
Pa4f/EpE7L4MCOWpMR0m3j5YqJxZDuRNqlw1PKq7/Jc8GSFPg7SSXDwv0jOo7staD60PMgvhTjAh
CB5FqYhYz+SBwTlDUJ7JhFoRy2u+NMCWxbY4pwoUkBjKn8ypfI6HNs4phnmEkgV96lp6QH6MSgS4
Kk60d19+HWsp/SJ1FG0X0kP9M3IKm+E+5NN3g2kbXylI76trQS2YIZuVh40m2CUErUTaUevh8x5p
Cnwu/B6kYzig0hu9Lx0UpfQTkcorzLtw5TA79V8+CtO90i7SE2CBo+h9R8z5mlyE3pRZWUXenMK9
NCHDl5QTxBGl8nUugvPLm9rC6ILhmoYmxjxReNf07PNW0L+Jm4BfiNbuJUuiu4iKQnP8XDkyVV9B
nNEqt3/Q84RT3hZX3jBDgTknGyqtB527ztuN17gSEO9JuQgODCGVrbkHTDoE1VIuW3wP1S0HxZxR
RQ0hwyVEFnihR9B/xYRS+KY5TSYsT4j6zuCnyhO3+dbW7O5BzOIIWEutgdmVf50O5qoyWhQmsKYC
1kZDWJktNOtp1jL3tkAT6fcWJXIiEQ0ukMIWeojg4FL48ToAj1CBt/XbEWNOYRGf3EGgOrx56fye
ZZfDM3PMkVzd2hS6NQHTsyJ98Gpe8QNzjEZI/xiC17eBEr3Y2z2WYfeoPdpLPA/3ExDwXd9IC1bM
rTCJjZspRY0TjiV2DTGUoHMfPNYiQN4fJrdbuPFG5sjPngC24AlbCHIV7pSHUaJjHF2ata1nEEIS
yUBxqufRc68PK+L28nKMbT2VvgVastYZa7K+1S5Aei7tI5XfIwavD5QwEunSIAgbRRxUGtoGKMhG
PAqbi2S1wI5l7IxhL5Y0NU8mxZcYUgJpME2LCfkRjQ8orHSXHGmZM/f9P7vuEvsGQtRW/bKjKhyI
zZ+GTpgM8N3ek8o8SJ/YlqK0pdASZAen7C0rBS7onYlzX+6XU1H5I4m0bn4K1YX587MnmbxNz3ga
MZffrWL9XmsGW1aUTR4O0yFJuVClkAidifB8bbPwkwuLtdl6Id21ZMAORkVRx0C+wKlVCOLFOfe2
ux5cAZkIu4fzbiAqDXoOxRVbuIr3hYt5ecKl6qGGGo2oScA00u1vWIjJ9ONEc4ALXE2uoodo37Kf
mN6eXrQ/GTETxuMo/IVJ2LbbM08ZzcPowbqknB0+7aBCM2gkuE6bJkpHf0dnJT8Z3fdUfOVdjUIY
DO8A5XRcSWXa/q+CEaAGky6jgJxZUr2oaTWZyAjOCkAYN2WK/I7HfCoZ+NZqcj5fJE3ImGo5vR3E
r/PFG12Wm+2Cq9lY4iNa2Wm/g+aYhl6PglxwOuCjMyiYRFXv2zX9xLxjVS9mWaVed7mJi1PCRLGa
asdZynBKeBnnJQtxwLxefLsxKbjaoTwo0OvOq+xSUvOPioJU8dxbt6XtEFyBw5ImfsxVvHJFMMuf
rv/O5kvzhRAAlHWaQrGtORkzA3lIG9eA0aVLzBtAtA0HNV6b1eDCl1WXZxDTWU9cIZGLtFeisNAH
pLftaFbddvBflzU9cXKPAYMwEe/Vssde/53G7cXyZawFXAfxYALRhj8+aR+6YJmmpXrFDK4yZpNO
pQg+wcec8qIpiovCX3nIzQnzSKZe3qzSNjU8Q5nNmxZx/UcUSAJVTpxsnOmRT0rfomRyRO/+AKq7
Pw4U3MqKzEq6OLehgO/tGywC9tfY9pqLfMXl7LBondri7ZxTuq1xQh4oHv6LRczjs4Un3RBwWYQe
Ko0Xm9jCWhv1VudOt2FduzlqtaAxFnhEEhrn7RaVcm2szRx58enOEDFF2ose7A6GVI9XZXgvvF9F
aJSwvgHWlTZ4QjQSrog7uzEH+n+kV9Si13iZLbBBraEZH0AjkyqFo/aEZf8ZwK9LQ4X9h+I3/rQ7
+hxEYSUl8S2mNJYoB21oT8SKqpt9psPkuVb2RPmdHoZPnwqvrIGi+hSajzwS4MiIc17R/fmoowBt
M68DOnXTj2bAien9F/zgbtzgdGFhRuPgHP9BLFD2utwxiM6TyKUqOd1xAXrXhT5sQp0IOkPAw2xl
NzXSMEwDdNR3IS9haaiak8hdg993FZ8FzZ+ufCYUy8uPPjruGPWRvxshQdKJ55DmA6svbDxoGyi5
dYn8vICvTdUfzzhmgkvKrfsxK5UXO4uJWiQ9+y8dtySj95hTeRANtKgoYK5htMO29QSXNpQuD6Sg
IFkSE9TdzWzH5EjtgJ8/97X1yR96jLPsIcal0GZGwQQkwi3zcsyNztgy2WMIk4BG4U2pSMv8j97+
8wf+BQxynxRmjr0ZAtXjfJrvy4q2kgZOrqLYtFsVkV43o1OjzG37l2VDLwuWM9Hs6P/OQm7sZ36I
GanDJDzwtxBnNuwb73WVAhiyZkuEjGgvuxZIVcDHupFj1C0ybdh052kEeXRx37P7+u4VX9tdXLks
yuJbVFqL44cH9s1/UUIIPvmskqf3gGwWYfizrCgeVcTKmNHP6/5gt/S+hq1ClxXiBXcz4bANQafk
igk+Ji/odVFlH+GwiHYgQbfEecQ9/FzQkyirK4ZSYcaiL2Mr1F4rNVEikioNtKjXKoxPR8woFyAG
Oa7ZvANiIca/xsCtoqTl561OopBKbdfqagB2JHXvwB/mozhyC25mLLycP1Qph7SG1oFKkgRVMWB4
iLbbWmb45kKSAQoZFFKS0SenHmW2Y4kMfpMPRlVB5WsgZH2h/4OLXywNUDBN5ZqSwJhjhzCKjj45
E1Enjh331F/gHlyhnJUxtdG/7OO4qKB2CSWvkcS5G/ubtsvg5AEiOgWQ7535V2NtI3DCsHPrE+FD
m3i0RbvJ2NVQmpvlH6QfTndpi7y9lm2XcO1Y6+e9xt3INd7ctJUhOfust1Y72xmfic5nCgSjP7kB
uJZirGZy0LMmv5UAXkVPXUFTJUApIkmZLnlVtBGSqsiB4VwOEJpktB33/fFcOa03DncdnKmkLxly
mmii7o/Yxqd+G2gps5JXj8/RyoTX4JJGnKHpSJVizlStGEvhSb8uaNDBpX5v/reOHrjLEQPes9s9
a4HopFDuxls+x1yKtAQvDFcvgJc6mxBuzR8deMLY5lvUmZVoWh/jgq64EpeFYrBRH1V2jaU2XKhV
kdg3F7hv0WkZ8h62BDgY4FBNng74NBD8Pr/GavFzF3Aiz2s0Q4Iy/7C+rBtjI2nSMu4gPthBHb0M
3Kb3Chhqo+Ug/34UyTOBLCxJ1L2lq1TaLRaCRU/heMwgBQQ7Jhi4C8nhUbdZzP9BWriCV6TFeaRf
HxdVPlEDYKmdsxfNLMIa45GdmZfSh9Ee9n8EN/6uCapPzmsb2MsRIOnTYaMiokYJM1K7kr6AYET3
Bbct83nhpVeaeubhRNIKeZwKAuJDHDpTKJDRqRF+AQhjZ1a3ABQYrJvHwPTy43gzsmqg9x4pv4qv
MfnlYVrUA3iQqf7fK8ZL8SOja7x7iZhN7zSTDC5ACNgO1ITI6tFh/UZPjT/NJB2ldswT1XDbdbnF
pxLlhi6+oiCqATNDAe75s3dcTGynsDO0MQSzbzePKuvzogE3QfUSJ/F3+KB30sysovvEq91vB6X/
N61IvvNtc+zncznUbwz+3sxeowVAHq/EsBk+z985489/ccO3HEJmwTCFQCTSG83GXajIkhIorb+m
d85KMUjto9wXQ2p/SSWcmHTll986I52e0OMqXpB8kD5g0oeTXEJ4BVutfmL3fnpETuAYTpf1/eoG
bQoCfII9tuZoRIbZUoMTJepmqhHuvIO+B6YE5a1o3E/JnXDur1/3Oo8xw4UzQKCtsR9RlajBytBU
G5OVIwXohpCQVkINygkb1cS5z2uQxOQlVfXdfCbcmWRWwbBwfXNvlOC11cjSINBWXH4jMSDfPIh7
Kf7biACnYNeUPJMpCBDYYEohfItJZ370JKeg4gN4thgSYqmVvtZap64V/SSYZpA5oAtvNL8tUnFk
VC1w1hXdu0IU4qyAMpJZvna+bQB3nFL8VA670IMCArLCeKB0t7XZijfRMO1L/yvy/OqXBuShLjdK
XV3LqXolvR75ZVJunUXc/gIPsQnr0T6QAvIc8oGD3DHhQ/tOSzmUvR3chCi+37jwSLlI9amIOWHk
6T4oE3Up6IgHkGvQvMA9kaf3CAOmRaBAS3dRsF+58KkDihMaEEBdGgrgCW1+C0cgCWYTekQU4DI7
OtrfZl3FZLpCfwKM66bcfxMEKiucRK7xpZ7lR+AIpqeIIaz5KsFK+pRJTiuDIqkpoNO0ZaMZDEN9
1vj9jJyHDTqZgmIKuxoIB++DhTW6k5PKkuFnESv45LAmEc2gzKITk7SxPDNs7h0aSr5zlh9asOae
UECY1GM61rXqAxpG8sPtklJNUtrkN09ECnOemfsaVhr14ZsbHxmpnG0srlyDyX0lpXpsnv+5poSc
DgDEyFDuutxPY3czr7nLYPTxYqxZzjR3zDQImO3FGIxD1eiEIeyzs7+mUAB96qV1vUoAu+Wu4d9k
Mzmx0xnHInoojGvriN27DNfLRMDcHZYEXus5xYrRaHEd0K9dhtCky0qyHKEOCyzp/WIs4pMuD7kQ
yf/0yaMvmuuTH8AtNg7EJxoF0wSsmGBmD7eb4D38S+JUwWdH9K/mmdF1iN+s9SJSF+77JH3OjILN
hmz5HoSLeA9Gk7sGFF7uIA8bDVxhHwHYVJ9vQM9hJh+zwt2U0bkyBa9uXrEBo9ArUl+QwSi17ncu
Izy51fhAItaVLdhknl4aHNYpWH69xcpXYXvsHa4fk2Bj3/8Wg6KlaoMrNEYy1ZopP58Q/oQZqioK
FmOnL8tQukqykC26bdO4QVY66yL8yXlebcsAKIiNR27ussrL0kkt3vddhYyN/5fOXAMTFlKVoMr2
JCyE1fEaAqxWVyk3Pw33emETanPIQc7i1f6NvoMTywOgu3YPSI6JjhZNAKpBHgytq5qEyEeeFNno
qE7armd++h6fKn95oFVO1QOmZ66f4IFpE/BBBhm2xzr7mvsCuetPKt6XuvAG1fzU+Y+4LEZhXfmS
OIJwHRW9FKn3NoPORVVNhRl4zXYolTvJxX89lDP3PvjIcDaMypYT2JzBDG0fjE6QO69AUH+J9Bkm
55lOdq5CeCLkAqclxaBaKm5sdJCGOcE1fYUR9xjcCO07Ge14GdhFiTGQMOy71hJX0I+tYYASHw+c
fyDPvQJDYi82TxKTevqtmn3W+f+EjksqAi5HVAXDgtiHxb9wEUjlPs+loFdt3EGh0qDmsJVygyYK
jaSRy3gtl+tag9QAWcbLGKdFtE6J1q3u6YTvsGByWbuTt2ZaqyiO3VPE1cCtBeV1gwk1l1egM3OC
bxqTpxxOUmd8fv2y92EbQzmKHof7U6jh7C+0zSfzDR2DPkiQuAD9wOBdpTcUCvYgzHud5nxFcV/G
E1aHSKDb9xVZEFMjh1wbjPtqGAMmi7bGl9+RS52M+nQ02Q/6fjHU+tyMy4Q74d3gD392g4r/i4GU
1M7hikkYLS88B2D3NtR/H89Igftaj50wp9sNzTNaGhKrd8NOBhsgil8iUZIksPophYSg4imGY6lm
n5KuHRFC0QU6haIeFBzP23Df6+NsRA/TPcbkSjoEDoYm3e6vYfg6FB1pXQO8uGXWXCTCxvsminLW
GVoqQgnbu2/BT7ao5evtv2l+G29ztz+eHxChwOXoF7U3+z5LJoB2AcfI3qMdgnOu4CuQUUcOH4Q2
W50+loPPHlmeh1mpQcetU/RkFRQLUNDX5e1O6kGH8i/wmgyB95HbHqDnjCLGUwZ/ADaupkoYoABN
8E+5tQT5THVzJup+pODYHeFhXCaFbBLA0tYlt+LBQbQ1KnFqPyDvo4DKt1EXxbRJejDlyoaatB6I
IPOISY7nfGFUf95lXR+WsP6eNlQ8eXx+7DNUEsTZzyOY0ZaeIesi0zXOXpxG+gwtquupByv/QbN7
t095EEux/QiKcoMgzOH22GnpjgyRP94B10JX95KOGWM0f0Kef4mYhXlCL6wUb3UoAHGU15w7Ga8q
zA6tmsRPMI4bEgNuGERrqzpCd5FrkhA61/PfkP03cEzdPEkjhs11tRXjp4ctph8YHU65GGnPBLxa
QU6PIfKek54qVKZaW4o2MtrNafyPtwCvcivlW804lgbDdsTzI660cfs5plJtZUSjM0SfiDevulC/
hgYAPFW4KwJOtdxJ/1WDGLXYRFEgGhCvcYgHA6tzovxsZwOLkuKtcOmNv5hyvslgmTQreZWHrQAe
orbdLS8f9isB8pcDoZVlZoYK+Q/AD/kJbU83aLqyeFXzBFBd8GRyQsLPS0CHQJFNH9wYDUFnrjK0
EIdnbkXBd78DMWzmZe25TBESULpqU+UBo6N2SjRnPzSQm5pTJlon+904fIhWFnMd7lqfll5ih42/
+0BY6/KscTwq9tUAwQO4ASiFTkYAwT+vJttGYMcsyxzpizA5c3UzmJGkUT8w7zuILWKoFAqFQw8z
Yt35TtMD/gFvtsn1D9glHjcfMfJkLxJn51h/sWBdD84lPVdVEzST+7m15ftjtH1U5YFPE8dOmpxy
c8WCKyYTbefKXI9/ExIu3cBUUpPiSVVj9EuXU2RZmLUGq69cJYHuB/IgxYT+Ii8xdxxFJt6l5yup
mYRhAFEgs9Hf+arLMGxLA1sCeyBcCZxIsUUrO5wrMGt8tlYyHWNHqQFxaP9xCfjAB+kTeM10bn/2
fbIciXxtG5wJZw0EmQT0uzpCbxPHT2h6E68IHOnivoHhb/hrYvOEclcrvk2w8Esynt5tOF0poJ4c
uh0t1JX9Lz68vbMKYMA94n6n4fd7Dbg4Gj34jKm/CW+ICBQiBa983ZMCj8xd5bZ3BSrA08CUn22/
9dLL9ARR+JptAm4ar8Dsc8CmBB/oYzVry3iCSDUbQVwmnjgiW1XZQPULsaYqym5okkb31GnTqahd
nG6oEQc9+49HHj/dsBKAnEg5o22rEGzyUtn0dZPrJf1aXjWZsINCyowT6HzvK9z2POTcd9iSToqz
z8wgaMOI810JJ4vR3LmNThPwJDPRSk3cfBXzMmgLAkT4Pj/n5uugCg4QXVXoquzpSxnMuxXVsWp/
8Wr2gapwoUHV1qcnbBBOopWW9iEven9aq01seEUFNccJSzwSrNGK3K9Ai0/uC+5XaHTfdV1fOfiC
IvqjyaBgIHAaqFUxjj2b4ZbddUvBdNQUKJOjuGOYrjWCYRQmo4FrwtShY9Uc2co7kKXN/YGZ9RqN
lICdarZnT26RoxlzynrBuP17hVLDj6kBj3ve1LztDuLG/bgk9TJEgXXQg+KKOvxcW4DGzDV5VcM4
ZEEoTnTvyKCom9//CQr466Am56yAvETCRIWfoGUrxt81Dy6BisD9YtQA9XNzOu65EsasFRBVrjHP
NKA9qLg778Ifx4tGe+cHVaY888V2JYi2Ix/tHluDL91/3AcjpbI/MMiFPiQQ09C8KqsZOPDFHL4w
umHJsC+DbvpbkineH8RmpH5h8dFe6jBppZNQ9n6lM3GfCtYnU5inbo0bvEbA+3WgOM9iN61ii+XN
pJvz7yMOLC/3yebmn7tmiJe/P3nM39E68KbW6NMt8Ovwr5ovLnWeITO0/EVR28jxc/p4xKmg7vWy
YEGIz1pK+TQOtn8A3fPmBx1G4utvBEjTbIPdk4gzH+UsZ4ZnNjxpwOjh3XgeEz1jzAhPcgLIwg2G
3NqB7PRb/imVMjrWnjvSs7P/8xbd3y1Waj1fRDrLz5pF8E8Sywx4MNgOQ6QhJTkzntLpdmQhkL3k
axGI6x0AGZn6S+uPUVWVU9F3SG+UVz6d82H6MFxAUNw3AuZnSHHiwxk1wP9a+ePjNDStXjujfbBf
9BXwZqFd1ihtxQllNkgI4wf3Y/3KcvU9eDgHvOoMKQOSDYj8fEAHpm+dBblR2hItUu2J4yXyc3Pp
KRJJR8om7nWs2JV5rH1bmF7RVyyna4dDGXAOxeuFms6DrEQslED1GyKXLoQk4uVbRZLegZvWb81U
L/HEySkjabl7jYGmq2DPYqhSws5nJJdaTQdWc/8x5R066l2fRotQOgi0n2+TCWG63isKsRQvVZfO
oGtF2nV8YWnkMrk3OJebTZXZHJsBGT1llxRgA2Gqv9Ol50mZA7cANAZ4GC7bffYyP/eb7eCiCLv8
z4aiFPvJUTe6Kzk15rqQVraOYAP/09STtiwvpdjQdv5R/salJlMrKBA89/8vkYkgbWTNv0dGIsRX
LL8HM0xugNj9YIwc24/KJRaTciyIxoeGyySaTQ+lwvtvx045zGuXU5t2ewtDYQnHUUjt7j0Jc66t
cwrjuTNjMEULzijG53Kzt37iDW4KiPohnDhgM/qGVTg9RfI/o4LkoopIM3YMlSfqraIDButrcCdj
fTyARGo1XQsxPzbBsRhrm4N07jzDyjIj97uPyxoN9fBGjoIOFZBocV/uOq+BKq2cro9TIQ7/3aOK
r5Ym+ZFbIzQs03nZt0v7rCQGX8KVrGgoYK0COrj6xhyz/mMMsKRnK+T7bXmFxLutm+daq1zi+xcD
60RRrihI71CgBTQu43bDKTWtgfUpFMk2izKYtn3K2Jhzv87iV9R9eFrdv04aEMkI/lSmlVmVAO+R
cXEyB1xoB/bjrQwnFMBPni1eyfCaCRFIXBpAznZN/wUVCL6yR5K0yMrziZWqG3tfGh0pRhEm6Rmr
KYGz52rGqfxXuxg6muoEK8krEMh6q72ssYvsPRDJlkRJf7zu1kP9iSu76hak6iNOkxpIMwYeHEPB
onA4qE/+Zl6ZjR3FbcE2oqYRU24TrXduS0nUmdhWmSoNIS9uXLt8Nu5EtnrA1J/lvzXbHKo9dcKt
PglYf3jlOgq4TAjrzuB2i4nmbbdaOIOYxPzJcSttM+eQ+S6pI1lQGzPIlX6R/IIEIElLknmD60N2
aTOPUwvVMMqQJDZUlUHU7j56gCLu7grwa4vlMhQQ5NHbjVnr1pXFa1WlScqqpvfk7TwUJ54CBxpg
nEzMu80SYhMKxIdfIJckxEDH2mouEZnCfIn87RMzBSn0C4jaEASxtMGzFPpBRAy/JK8OPAab+E7V
vZXi6LiPyw4S/HtBT9O41Z0BMsGGQFvv815KGrw/YV398dSLdKzE9IjvOmWlbNblRCxv2SrdqPZc
F35lCjax0DAT2tkXmw4nHxHeKd80zjrWlepJ5VZPNZsCgGW+OrDjgfQ/XcY8YrA7OatiOtdixISQ
c+uax7nK28WL/eOmi3vjY+aOH+eP4qs14vi2E+1FPDp0Z4UL/R2MERHUDR8E1ed9GqE9XJemkApq
RQV54R3xFcuuDRgHHgmqIioqfSjmkrpn1PCC6YnRpMkKG1VCcMxbJfbCDrZECZ4WroKjkyvitmw1
Yu4V2MBhPsR5YwWqQZ/Mr4FP6c0aVy5tfobmUAX8PqIJLMnmA8xrDfm0Sv3+I6nqkIJ4CDEkhgKr
OnZUPbK+pTSafoI8xbf7FNJSjLeqJYvMh8hq3QA0WjGU15LmNn78xeYFPtIcptPrfGiOD56bzLhh
gOY46HrRIT+sQXKXHEcoBQVNhQnxPFke9I9gRJGdSrLHb//FgzmGn2w2tQWjqJzv+h53kJE07PTh
qSQtvZiztJGqIwPVnEOISWp+ebR0mOLmJWZZw/vFCTfT9abLnAYhvcMxZHeDQcXc0OeSawqMMIyP
MRYgAhtXX0Oq4brQjhMDYddK+84UiFtF8ZWRxtF4LH4OEbi1pNiWjNEt5yqV5ETjx9jzrClewGUO
9ger6ey6cy3BDp1QvESPxliCbnpVVg1jpTWjNMHFcpp7wqiDmdSMNB2XDfErachgtkRUgq8Iwco/
EBbh98b1TmDHRpi+rrCbTwvTB/FIb/cdRK3oF4Q9xvIeJlWI8JCHQikMBp0sHt2TiThTvXy9tPzX
NrjLzz2wN+opyKwRJYDOn+giuY0LpvNXl+86i8lHf9mzMeMWySkx3TTJgrl1H6BINlgNF7L0zl+L
QmOPipH1SOomoNFPBiiZbghjiF5HzxaMuvhXMJYam1I67xLnEfARaIBicf8L2u6n7UOnamzgnQzl
IOf2fHuocJpTXWlAix5cnFpaWhoUY6dCghIOHvGJJlSeZoFwEOWq+WsnZy2LcpoEiFnkeWxWi+Tj
DyZaHlrd3ib6dPqXs280RPehuLuRQMg1YDy3hb1Qmj1SzbPjGtNg0J3sW45755OuBAny3yXuyXHY
MxLIoaS+byUEV6R6DmZD7ibBfceeyeSe0XilD+/SrHOfIJ3rcMecpL/bVPhINcckHEaqhwYmSusd
KUrERbHRQ7ecnjjpD9WUigKNCSIgLOXXy+7h8yOmCh32ORijE+Vsh/ZdHnS9eR0BU5X+rFzxrK6v
eMfxizU+BoPfIgywLJx5jOa3Mi6PLfD8mYn9hseuUje3qZ3HyArbbXypTZdoTcGIlGSkGF0f1UiX
iwcliawiyEPt3ZYlKyDS0lWM1cvh7Rz4ZsotoMIyfzyS46iGCuaexyNwVPhpg0UCC8Iujj8gV4yJ
Nbb7sh5xRibSjcBE6tcz+GPkTBvaNs3nrlPHl60OWa2VUQXiFqzLFVNEl7bBYRp72srObhP8kzbI
NEwbCwDywM4qaAT9blr9fMvhzHsJ7LZztS2g+VylyOtQQBHtjfQqzJ9iibOO6rFrh9CKf185Gtzn
qrvk4lt2l2huxDtzIzjkZlD+qwzwVDTD1LgML53ToMmgOMmjTkcbBLtnnagH7amDpdsPbeUQW8yl
HnWzMaRMfPwOC/MM7g/ehK2s6JSJGv09jqQwKLFnfz7zInc52k0lG8bPrYQ5/h/9r/aVbO8Tsuzi
Ruelj7fuRyimf6M2fUAQfxvipny3gbxXwdnyNy4zfbMP7JoZjI18AQCvJgKfhprXmvIo7UZKh5cA
DO7xvss9HId1rBO1/j6kt0uYdeV6MDXnC6tzePrCWRiwQyjXAmE5KgaxQtd9sHeuVd3JVa31v9e4
/CWR4/ku6imYI/vOoZIFchp2KWnmMPy6nmFm7M+gxr/EvyVBqX7QQPsbR8b8qWI7RICRtRCMhCcD
7QKIx2pz7qc4aESMZeHvNk16ovqwO9wFOe8UbP6k7l0EgseAvYkaEx5thS/URm8DrH3fElXKTTL0
48GAL9DjkUTRNoHllNRnfF6dw4n6ZwXu5By9lcpSReq41xOwTc051OSu4o+0jmx3NnQGljXdUq9W
G7ixdw2142bT35GqJ3HcGxkVLZZcwZeBXM03eU+XskSGZa0fdJ6S+dY2Z8WaHKZIfaLEMs1FjX4V
C1E/OKAs6RgnCyWCCA0dvlEdbOii+yuhFaZL3eVaHnCLmY582mLqaTFzgUp9wbIDrTswIOSDIBKQ
etJBsZ5+dls5uX3noSqgvriDNC9ZgVcd7CYxO0edfnNmco5ZUFzcxv3UnV2xeU/+vTt1CM47T6EO
+6dQKEvZBeIwQ/8Xt3tpkpmB2ulxrz5jLAn0qNvz/0X0RfkYkX6ZJrJ80550ReDHxM0FNyM1bhRK
jAlbpw5KgLWoquCO5G6AkvZNFDDs0oK/gd5+tyo74Nss73+Bz+veYYx0thSNbwzn2HXIoXES4kn/
O73SFoJYVcIq3QmIxouFpvdwguK+kwyFb+OHNpOOGNTEqfBnrsgl3/qX7dKxzMUQ/ofMVFGNEBFo
EAyXdZRifUW2VUJbZzcbRHqLSv6zofPCfpMCvNT1plA4CV3udiMPxIu4R9s8/5LMQFCyQtVKMqpm
USdfFSEfSgFI+yJTqGt5Hri6dDcVCv7qio5aNyljxpvxG6RMwnrDcoot3IVmbQcZ/Id7jMxeD34h
vRc2TvHkgTu/ph0vBAQ+G+vDQg2S9/shVokBi9L8gcF+G9sksZP5IM1Iw6oDjQ52y/wVH0FxV/RU
M5RFEBsEXMFg9WEJ8rAwGSf1vwdMVNoQIvDw62tSArkuTK+OIVyLcWcSyPc+85K5TbKR3ROJvGK/
frEChP+/EKlvvI75/bJ4qTrzI4alXSW308nZgGSOn82WBFcUIRTxhXBNIDVpwAqoshX9vXBf3RNt
R/w356MZmvofpwpxB7w7H6NxQGgJq5iuGknK6xU5vZw/QWzdohiOsPhdKtQtNI57pCb8/60PITUH
I6sV9vs4VYKfIQhvrajoC+/rTiZhWdtev3b9Ieksjh6IVXi7NeRV69qeVcqu/P3XvHEnXcBv657e
qqf+1PFIM0d0+U4BkIR3PtExGn9z1OyR5IU2eQ3mPhsZk0D+NKuCLmSWj7kPcz13zf2IhUygnE2u
92sKVNdmMWFQkoyx3sV3ldUFL6AtFCjq/BW8uT73lDdWkEIEcDgK+ZnCLK4Z1lndJaanKDycK/Mk
2cjduoWhjO7Wi5YITtXIBdZXxOd+uCSC31Z/EawBQLrQ7VOBnzX4+z0uLd0p9Wc/eTywRzfmU2aN
ZP3vuqi3HTqHTuG1hoVBWbYQGSfoloDh9ejblJJAQfvxUFWTVUgdXX469zWmxerKifZlSRQxKkmQ
gpoGUGSjt0FDL/lWhkIHYTlygWPiERyTuchXIh6lj/9lmqxK29e2FtoV6KNbsixHWCuXwXzoQBfb
/3PPgqVtBzGudGoKBilSaI8PUbU/W+7SnFbzh0GJ/jcGCJ77WuTLX9YwoMCRVzeOylRuP0GcGfu/
MbGwG0CKKEeRS3Y4nvtLAYkPQPtiyxUjW/up4mb9DMh3ZSCbLLbmMjk5USJXLXKryO/w1yUjgnmT
TWSH8jsCO/DokUUykyXEE+VN5zxkWNRU5vt3rA6pPR0nOMwGmaS+PnagHlhcdEL/aiCpwljXLvMB
Ei5SLo6WRtTSL8SV/LaH3HwY1AqOWKYZeHSjJYmJdz92MefKuPA9EzWMgjWCijQm2BvpmULNdrUI
tnvR0UhJyd60Zx2mgY+euJ8kxlcIbJDoD/GGnwin7SQe6dPEnN9CfcrJ/vhx9jsoDN/0jKSz66Dg
xsbAVKnRuujst1wmY2ZcP/yeidqyJgkdaAMWomEMkQgHyu6DZljJjTkWglPkDgZdYnABs7B3aJtj
OmRmJU+2tLIw5lDR/rQM2D3JEGwKAp67NpoTI0uudXgWlIP+vA4rqYQ6dOCzzEftLa4/oyaHJGuN
aBfYxwq06iBs6en5HcesPnVAgWPhjZCi226wfhQaBiIkw86OkVfvon23Sd3q0N/+mjjJQmeBY/OU
aonnorzYuKMGOEkGZghwflp6d4zKt84g91hlqeHqmVd5w6aCRsFMmQSpGrNLf3GdadOVJDyuVqPN
E0QiiqZ2fTcAivPbrRpp5w5CVN7Jm/VV3WUrjlFumX+VrgvCVqZrG1T7SZIL8nJo4enYRM7VEBD1
Dt4KeFfV6qpk6NP5Q6HzRh+lS7k7s51Li+zMFqRTGEoz8JzkT5y4jS3YIw1EIpxEMgvIlzeA97oc
L+AMV5nGbb+egNnZL6ssv66hpaz3w8eHvQuqG10VQ8Mx0Gezk8M3GYtfYS3OlCjs3tKKn1FwRK3w
ymrWRzIBLuKZJRusc7vfI0ErwT9DQdmI2Kqwo58vsGTIMp0wxpGO5ardQUQCqrvORmraLEefWIj5
PqT4rQquB9fajqX1ozlcwdgSkcc+SVFjsPDeYCYFahxYpnOgh6JH2s0AqX70ILXZ61m6bBX5TndC
pf3NOMX4YJu8UMX7ZAWJTpPe+L3nc2ujnTlB7uplMNo+342prO+kBTumGj3eAVg2kolaEYHZNp5T
QchU5zT2Xm3nRMdpw/CNxTWqPs4uA6WHilkJlkOSUZ4jayYvdM9Zu03VbDrYDHwOlDDXNm5ZWzvC
zIeQUVFIlpz5tXZRtXJw1PBgtYtSbBR+i5pp+csRjeQrOjE4bj+TIS2tW4wLB1guqSMOBKOz6h5w
dw/BLfLioarXZnipU1fx9YDpTahmtc/ogcw+qxmu5grhUR+CqxoMkck8u2nBanVFv/s6yKkXD8ZG
gYV/gi/lDeHOiM2scyORCx7kg9AfZhEX1qEO20DkQg64HbeZrDMbE6aKDxG64U8DROc5mDksCZEO
rcxrCfmqyC1pXASZ/Z4aWeUwIDE4Nx4E00ANvmEYP4YE2n5TDrD3GiWDYV8Zkts2SpTgPGoczBxW
RJOMXY2bCSSzrotAa9UpD5ISEPKjqGUqJYlioMQ40BdCuZyvuVpjjJWupztcl1/7cb2Vo1oOQFIZ
5Wsb4H4xBs3ahtG4IB+povMAWnTW3IOwqZylVuLqZx3f+tO3sTTtpVXCdFNDaoT0F7uJihpg/hAc
2nUdwm/YWkLwIhurWvFrMNp5dibD0SQDE1gDYzWWWcpo/GqlCOo7Nrtlp+pmWq9OJzkh5NgNb55I
ARQxzyLmYr1J1cRSqRxzSTjTTiZhxX/oeIsMYaWnROboZpHnpc/aNoXRnrvH0mqW2j5dPW/EJ0VS
GmoRXC89U8Ho0uOqcRXb21+41CI2ijeVewqSebEXqZIB6bacu+dHwVNPpfmAZVSPjbd+wASEP8kW
OtWpO9iAZt7s4pQhQTWj2xG8lAwhesonmJtvBoZFXt7M3B5XYW9oflACBpr6u10G8BDU6bUe9VM1
3ctCmi+O6xI61TtgA1Djl0Ol/5UROjFLHyghrGprBglWij261fZ/IvTjTNt2oLZNNr9SldAZ0ZGk
HWQcNWflBkQW2j8CUH5nBm04t2ae+wbWPETxLbsiz1aGVO3DxqgKKQaHKkK0K5PaxEcs9vOhcl6c
vwMdMdsUW6RIO7atc8GOVyf/jsveD/S+PCUhtKixA4MfBkyVRUxlf/7JoGAW2C+7Wae/84JiAOyr
lKiCQkNjyfqtesIBvSydiRVX/fF90f/qBG4KNxtPbliJi0AaBFwiYE1DOnGSqza2zR1s7ipLXnix
hRhm8KfloDHrWzsM3JDIbA7RGKKy4i0uJo0yMmkglVpXnfIUw+4EZF7xip+JNfeExDug4uZtZvBQ
WR3k5wubkru7Pzihd3XKXw4RO52Yy89En1i32CK41j/lMDXsnmckScNUcZe/TKrjT5f8s7vxA6aJ
uaqp/MNIWTUm9pOI9+ZNotRwyUYHKyE5F/K3YN5E3qdfJftX7EvmwJ8mwPNbEVlknOaCZ9KggcvS
rtmURwr9nM70XuxYukiK/Sob0+k8L6H3HBIeiRfxpgFln34xq6KJWvoWHpeQcK/BX1L5ZYptKDC6
3qvBM56ig61gemn1tgaFS+UmIUvfmi/UGvZHPpqnZUuxJKrjlA6w9pVOSqEP43r/0/736ME4r4QQ
ktMyYwpfBFjEMUwHDCKH9enoymy6e3WIlcfN97gizhGU1bXFQ+fBKKFV4PLXDkIOLuTPicvhH4cQ
xOuUvcssKbk2Ny9HPZFasc4vSdDSdnx3lbC8qvMLkT+EmXjORqEuSRiM1MvUNq2e5IwQOeJwukUm
fPC9YbJNL/j+CYY3LOLJmcPQtMfvVG2ShYvUgs2mPdUPxgWIaotyF6k45qKnjo8qtE++Jf8P4hIw
sLA+YxrcCYr5NgZkfVE4LT2dG2bXXtEEao8XbScf4gN/0TKVEkFnIEDnDd21FOaXlO97Bv897ysd
SiDTyn+MXiF62EX0ZagqX3Qn4ni1pZ4IejQ+BHDDbjWilIVVNv5e6kQiJX33Zu7W0iAgjTvp3K+4
FDdhV+AGUeeUZACInc6nQMR65/SQVGFEepzv/rIBL9wdC5fRDtHBaZofTrxZ+tK4yJpz+jKLd0W1
cvQhzceXJZ/YCBkZjO1q1pL0kQtO/DRvsOy8gdXIk8NlTDQTpQf26JMp8kbbzCO0D8KcwETHEbsP
7dGziLBONVoTf5DsgY0nJ9lj35TRRYEZuBRgJtwlnI9zTMFgpAVICbhZS1CwQyF051/2KqjJQzaU
TwT0X7utcfnP9ZOq6X9M9w0aFG2SEZahGiFgJkTC6S7d3Qh7NDhJb/NLgpCDCetT4UooMOQwAt8U
JBzd/53Lfmpn1Qtm1aI3CrdS88YRq0jIkEgZvYJC3XEPo+Dw2/lSl2rXgcKDxpqwNrxIHWdJwGsh
4//Ms+20e68UJ2hTguW8XIDNWpDvYf6loomoAXq50uvsBkcX1KLeLO/dzG+IjErW/b3NQmnueknu
GaN34Nly1sw5ZFD690tD0CGsUcZLRmDD1Md8VIrW/qTv+8CkmJFg3c7cG7n4RWM9M9jdzK18WWjd
ACaSsTMqwHi/zj1Areaq7joOBRQOZiTtkkzPk6/iIXuY/KSuZhb8XRSdYlfoQVwSsEIuWrH7b0Tm
uAcdOdLV91DAT/pkgQNkF6Inb1+N+kgIv45lmUpA0/HzgZqq8eC6EzKy5rhJ3ZMhoacr22yBjfvU
cXaViFWu1zfXEuxNJwoX9hlhkcKW/60IytT5f7yqoINrFiUWPbymnY2EtuHDZGL89i4ONBYDtwfH
Ugs9IA+BSTJLyEgTA3GiKVRvU4i/Yv27+Alc+7DDzB8hcETAJ1RxxH3P19m3/Wj4UZe8y/EIsWiV
rkuUQW9+atDTCzzhvYCzkp85+htBliJQqBCcopA2FZX5hV/cp8TsAWf7ubfRMUgI9HhB/8rbxMUI
A3744veJEV6veb++LQPnS0tLnsrFMfWi2sSE2W4DkQpG3WYVNeef4VVttYNtyLYckinrgoTeQm3g
SOAmdXK6wQSRam5U95T8AAndgpsmy2WfTXMaaYEZZggAGFR6N6ga5EcDb1EjuQz3znk9enRQM+i2
NkngkurTRph+XlNJIi4I7w46eQiZk2qXnqggrlL/80Lks+A9Sl4/yrknqbrwD+2UomfXK/fq5ijd
T7MxCRnVve5yxsMxlHHcUf1avBCCD/azWpfREp+Iv0IgM4e9m9YWfeelh/GKP81Ih0NMADb5ZnDr
DLMy1Csq7ee6HEp1D5frDWPKToem1NSVX02R1WwkLwDjK0w18+WRmG7B+7Dfn1634gMO/nSJY7jB
LU84ggvBWBJM5fcLFYLmeGb32kzeFmzfirxT51XNpq4ZV+V3oeDbaU61LI3KFh7MFItnmQMFw5Mc
bqWDnMqHhV0pQU6q9pxY1+QOwfpwualxjm1/4mbFZtAUaQoyjtu5i73BlMoExHGZmUWYfW4Vs6gZ
UQnXq4LgR7DAbU17VAC5CRJhp1pC3bAgjn4b1D2m7NJDVVneLneZoflhXRAJA01lfa0D/03UPsbZ
mXEwm0yaQyoOOBBLWzWRe63HLMR1U6ApK0tBMRs0h4wAUWrJbkej786nFPSUrfN2NhjGxpkyuZF3
cF3XyNCNnvTMdnl/2Ir/tE8o4WGWwQ3mBRigG+z0l9NQ+OlRlCjSrNoCKeY/MsTNQK4VY9O3/sDv
PNTCXRDdEtXIwZZVAdIYjV4r0qQDsALpWuTsEcyBwN9INhD/znArzyNOra0ep/xBi8XHjNJ+jlEV
656jUu8Q1rKi8499BIG7vm/A+V2qQ1L49oO0gebwSVSq2aIgIj6YSFJ78oEzMowHrZILYc1xAnqQ
IGYcDic6vAkYMcBzHBCRC5p9+FPPet5whEIyiIoII/n3aRSACV9s124X35llf08JQYLyJ7IbQoCs
OHQ5NRL00LdGSGNawGOdmQv/YlGSXfH6OUSjnMtqR6Z5/yRAUynUJIpY5+LfQtyR5MnhUQQB8M6K
ziojZTBqfy4KyWVyrSE5P2qmIoYltqFzZVWC4qL8iCPTzbDCGtedw5hk0Ea6KEUM6qfRCoL9oGru
tYjSzP3nu75kdMoMBHP5LIuYMb00nlDJPYYF5Tcl+R4mstiGcCcq8bK0QTudSDf32hCy4k6JBCv2
Ak6s7K9LYymmhOyjsOlppqBpBRdEOOyoHIGizxUnFbQQ6BCcIuPZsWJ90CCOPyJGYAXDN+Fmgifc
QQsLj+wrvbdzAmpEULU9vPHd9nNLjVVlw6LpRuVVJZDsiDUI24bdI+T9UjvoJDhtuH2/WzR4KQdk
47Aj704A/wMr/XcOlFJD+HK9KlLhqcLV/FzPSzm86NNOyXg306zkSiu/QiJFkP4m6Gfmb6pja7tG
7YtBPMKtVXHcvQHlkzoW9BEQWoaY3vn1ZBsoHFDH5lmwdTqTnuooqjp6iogzG2VN/IvRgmzFLWAE
IFHciwjCe5ti0klNI5lnzn6m31lrZrgDR0Wvk7d/lkYB8P/zmD3pKIqbNjDFB7SofcnR0U7UTv2B
E8Phw8nXz5lNa77ADtVnRXnfgQZaV23GLxe4J4jKBn+JRAmMP++CCSPlyyqGDf5L2wymtJshGbo5
HOMIleQ/gNX0I1fQsBLxlEC/ZSaZiLgpAM0k4XbL7kQjMuFhoC96kNGZaP5B1PVEWgQy6RP/7nA6
Fkscr+MTItfrczw7jkKre7IclAN97whxP6LLwQCTJDNmG1DV8JPYsWuEmjOYZqrBHaNFC3dt6W/t
h2ey6QzIkIUMD47Klh0SUMmFV8Zx4prg9+cEWA7CHtsFBv1u2JhLu5i7TyYug+lPuWoFOkocCbiz
2+2Y0zqWF5J8RN769qjFmt5/6Tq7jEFRmqXcDBe3mi86ppMfXFZb+9SEFdKqDZXobzVBQ73xDsRQ
XejBL4LoECHHJ93lPX9nevzLxRh2fgeVWwh8oOaDoPSZPYuIlL1jLP888RhIFWvc4pdS0D/WbCcj
532sxA1L7uvPddCIdNqPwxX5w5aEsOiWrDpuSLjLg9BEY+r1Zc+Bs7t1XA8mWAV+TrSkn7Tq5GCx
sJEV/gqdaQLWAD6OuuyzXxE8ipY0vrQQGq1pnaL4/imUVz9C2m6UeslasWXlGD2/k+0plU0lA3dH
ITUBC3dofAI1mxMqcvhwtx/0+XL9wAv4EJX7Z+wQ6otwGCCAyAXCC4+37sdAG3Lmhfhwqlm3hSRp
hWu7SDm1Pau+CJRLOKJhZ/x4QnhN3t44YJHf8JZoImtuRE+O9LBiIkJcEsLSb3BhPjiAiunzZEVC
HqmqqEoHZFnmMnY1qALZXl81ljqIlmzTLb3d2RZIGcG1A/pwyv+Ba9TmXilxz2MxCzCaTUslDsKg
bDdWX0zaQG/YU+thPTlOgShEWV82EC7HsGX9Y+hf8jJFqzegp/O7RT4EekNa586o3KE73JgQ9ADa
po7zeHfJ6ngNVbYh+micTDyqiphwlQtfoTrJiRKX9k40OMgctxU75L80NXS8F3JZ1Ti8DqQthffZ
mQ0633BmXs+aQlSeX6vv468D8le+DyGniqpwQ7OCiJfuJgcEy+a47YAWUsVNwfWMtvQv/Wlat76L
6G2s0nB5KDBqO1r0/H02a0Usev/glJma0phEOKZInE7JTJYMrD5mLcqJZPKxWz5xesSQ8CORKnyv
xwFpIF4QpgmBT61aBvuxTLqGvBu2PGD0xGqtKN5L0BF1n3Ba2KWTLmPyccKcYbY1BicHdrUB2/fK
Ixbm72ukSL02J03Eejq3728NQQOeCLzaPq65AfSEvJf+im+wq1KZ7yQYVq3s+HyWqn2IdxRuD6Sk
iVfYPoMJebQQK2vHXPLCFEwBX4NvdhmL3HG1dJJlAJCUrxilSEJovugLw7GIg0MVIK97nRIsEtRM
iBzHdq+FD+h2BbcyTHJgUQvnGk2U3NJVKiIgdjxO/b7+ZcRsVOAb7cBFxIjJ79gW6wphpoows/RT
y/smeQF0gh7wwQ0mJllNMIkJqSccTmHLGoitymV7c/oet7/K+ifxf2fNvfPvHFSS2L0pN3/aQkDt
d7EDoAMJdPjySvRi1NXB+pjXSCkE/VF4pBz+vIUqGHer+YCBUaSUhjR3G+rImtBoQX+Ss4NXAg9i
p5AO9w+hXrXyMIodZinxl/Z5yTozvCclhEMwp612RM4IQQmzPW834EgrCAYKoohYv4GD3WPlw4kc
0LnxKAzQ1HRZkAr/ByzbrbF0fBdXE6ocWD7fngEb+AFYmv6DS9unbmhihxkfsONXaUWciM1g9vNP
PpXiXpALvMOpjyr+iWetIfk0wsW0rxVxIuDhZBj4cHx+V5MS/IZY1JgKk7MTR62Fi8WUSH7VonqO
SVsBZCZX4oUjyZM8/ufYNJAyH407CeiEoF37QAqeEstJrHu4VTgvfKZsl0wE3z9rMhdET2dAhTer
2DUNgNkpCzzBBfhElaesPqqxdhCZIQJGFUgDTqFc1Fmh8Eucu4BS6PnAn2XNkHoHDiVgzIMzjXP0
6Cyc31Z7RH6Gio8+1TXJKqUaWNrR0JdwyKoqp9ysVh53cZ0CjVS4lr5KxwyzPBIeKoNaURJnM4h8
d6ZsT28STuzBHTG+69zwn4vyRMTETS/DUyfpXPW75CAeTClTP9t/F3tHE6htHzrrQ6VqEExAJqMZ
/5ZXzJnNPtmWFeFpaI29J/1uQmtttYfTD+KRqgWaNhdzNWYBKB5uZL+matxqCnR0VenCWABwAYoG
0YqtSfLoiOTs2hBjAIgDdZYAihhgymeFdy3aGTdxAppdQjz+CN2vDnn0q7qR6hY/7qAPqFhlL98O
rEXntBIruDfkMwGKMkGm5Ts7WHVsNMSM3cVWRHTvVhrHxMJ+cn/LwFSioMn2+p35ypwI7+qP7aDY
sIid8hjxWxU0HtWyAxHkc2RcrnYsG8n2ZSLzdhaeV8b01TIRgnXUisez+ziHfVpoqWWA2wTwTKp4
zrAw817yUi8jTAuAYpMPXZz9BeeiXx5qPsvNS25DAwM+XvwpQcY4ThqKmFF4rzjm9hXj5q1Hio9A
zNR52iBpBl/zXS4NSa7xyHaI5fIIAnEX7JYhK46tPup91Y2OnDWLOt7bTTzBzViggXtatKMVeI6D
6m0Ium5ljtW5ZOUHvRASpH/BsC/w7GVxw7deSess14pXhJTSobJuGmUs5nqjW1HLk+TszzsI81xO
4NFalbLTrlOHBbax3XynLNWKO1VpC0askjZkaOFREUx9EiY+jWeKuTUphspEa5SRx3TWTQqJjqG6
jW9msXdX+WSyHqSxztahZNw+h7Xn8boxd4Err6w3l8FR4sPOiEvTE+UJw2kk+Cq7EyMazolOEK8s
n22UBtI+Px3B8Yp1PB/tDISODqrLMapf/rPMIjzUsuFUifHeux2lRtiF3cSi+ok8/CTRDHL5a/R2
E7L7VjNnlhYM2p85t4cDSELUMnNK1z7+CKc+v+/KNQcBZj442lqTdn2Ik9+iOMP9UTxZt+SiRfQK
w8aUZ7/IBmADvJyvIcbsUe5Ls47b0NzYzuCJWZiQL4eBjbHTYjGLWJ87omHOHIplZtvRWJTO341y
Dt+uV/LpILHbES+1fUGvLkxh2RpECR0pWXXWXghUhB+XK3VSEBwT2EbI/R6nPIdsPZz/spSajDgU
gqd4/RhCOzkNh3z1nFVQJfIaqzmlnhfSrxmSzkl6AOFpFAe1fm0LmPqy06HdSwJzuyZBhGNDDHsP
jXfW2+N7ZHOEHhOZxglD8F9OKSwKLUHWHBBMzJZvVbN9OSaU6ZBkHTTjt1FP/XeZmIRNZOoV7CgE
VxofR0QEez407duZ/k0CXURDZ66xzZTbFpz2xe0CzzBUxuw7mD/YMT9kcJ/L4Gslo+Dx7PbIFE9G
iIjjSqbiZlBdjbqCzKenXCVAEqcayp2MnmRQkI52xYwWjWwqj4oRnFKbGkJsTvtyHXTQPZpiWdZs
n8rbhDy9I/SRtZtjt9DB7rxodDVXVLVTuG3g5OyKVoE8wRSF3s58dROcyubTGEjZFZx8h8P3upYL
z+/codmNqxiCfN7ydptgXNhDG4vETU85TGKwZ17Qub/C1CoS9T7iUSaruHY/kSbq3d6est/h7fg7
q6qnb9SpOTg3PoT+MTg1ftYjovptvXcd0PM8H/Z8sEjzYMzMaZ67ctG+vhKrRPjzyWGFwHRCWqQx
WpQm9dOAPj+hDFmoVd4r+i01NY7rEVMKFgmb0vmIy82OpUUgZsH+Er08MJXU3LesdkvlAL4/7Y6h
VsnzHo+NFGbS0VYjCrCbyo6k7/+umcQaqaH9u3hvZjHfGW0E/6S/peinWA80PZJh3qzjmSD5Z79X
IOueERTmanQT1VF5xS1v8ioiE9QqYcByqKF3goYRCN8rAqng9+BOlFWO7eog7J6GBz4adWkEQ9fL
hHfGUyyloDkU86vBVP0nIlpfE/Hs4a/EnFltTZskXKHO4Wd/gSt35PcORPzUmob9V8IH3oiatibc
cbru9YPeEEckKrC1sV57R7TIDhdn3sMUyTm2tcReCWefA5/YnrnclPSOqk8huMegATrJSGy6uiYl
aE9qJddHiFebC7Nmi+gP4XhB3yepM9EtttERWVUzKf1OjewiuoXhWuo8+tnvcNRwFdQ60CzF4zZa
/SSv0jN9Jts4FCVbmueZy8X2+L55T5kq7DombJGSef2rsPqsE5sAJaRGleDi+cU1NvZHHKu7m4YH
SM2CMyaYTl2tkKt+lhVfmnAY1JSCpGZLSdl2/+Rm+dvNBYxl6gVVVfJyiu08JouLcY7WNBRmD6pL
ylkzXeY6vb4+h7DDzKaRiaJ0wKCIada81kD5vevEYwKhIGbn+fSGCQfCHC/0ZveV/PioHTwP7csp
Uvzrst1itZre+vTmGymlEQq7Gn28slpvTLNZI8/lCRhjKzdlin5pRd44LFkTyoCC1uyZT7gB/Com
jyIjePuoV5x1AMGdAf4U4dWYopCdMBqGlxAnj+3/wsqrC7X5+YLXfncFxwQSTb9tPyds1uyYfSUu
dmDLOVzbwPxyKvKZ2GF9poIgiQYzf9+4c3Lm79vRD88609exuXMA9oea+TAuU8dX2k77kDGSB9fx
MfhvJkMlaVt2z4O7McgjWI4ymCFJOcyW5YurrZuBuCMyZ3+4k0ONA+42LqIqNMwPjWfm4bpHeghY
AnT6MeNGeffQdjJt7dh6P+ogj3w+L2TpLKRpgDbDoVl5BFbUgNjR1IcP4AEeacWHjqfYgwKM1ZvI
9phZaLOJCFY0RcgDEQlF2EbKptg5WaOIikT3VDUaHQ5OEYmRYUtiCcYqrj1SNDa3leTi8ttIfxEU
xV9HONKYxphDaC/8JTkrhxlB1X2lhUFgWfqxf5hVm8Gzlzr5VQ56pvIPNtUsvzyyE0p37g+bifTi
suLCdGq9aQo6uzx3r7aQJcm5AsS+Rm2wWCOYUdia7CPU4yMDmsx4NuehWx7DAXC+1cLw2IW5BJyy
XQBSDCiDT7uWuY2jgkeJ3l3eD3yUKJfPKEyd5CkUU1kOGcHNGygPqufErVHcEfUP9MREVkDf2nGW
s/EX4a1i4+Z98sV54q4wcb3wa9ZMISLGD3eBzwhtpQ1ihI3nDDbq2uoL9xJqMHdSG6tVvedHezxx
Gyx95gX0eZwvb3se2EYhHYxKIzZ4yJMHpPjZAtWZlkolWAtG/vV6JYh5/VB1GI10UiBIu2HxCweD
2nKCr6XmjZHH4YXe0OGFa23Mz+ux+lY8cxH18ElLcCQlIh0s1Xgv5VdFlz0fn7ONvQSg1wB1DEEw
LymLmjE2TTImrz6MQ7vZWc9u/4tsM+TN5CA6sD6friDBeW4BjjcfMmNvcV76nCXSCQ8amUepnikg
OQS9+C7iTDHxYThI2FyJFAwBLk5QBZg/kNgmWhv1Ug06Bgp6tYVwAZ3nf6jC6eb9XHlovlrL4gH7
qCMFE79b87O8B4THsxZeOlOTaB/2oTpD4IxtH4w56TfKaRjt1HJVXnJzJkdpYKbIPqZMMWGhuxMV
h0u8is35GM084zhRbChlEXoT1wGRLft3Ab8iEIU9GziJu2KBsGDyaNjxGVqL+vtAeCsoizJHQ6nM
WF4TFxVY1JKoZBjby2ISLyb7G8/OPi1EBRF8pCQpDZ6RlkR7OlA6DI2re2kBCen0DDA9D+ZgJx0L
waVUqeh9GywKJ5CFtW8kcz5+V4vroN9tBnbzXejuYAcRxnsgiZl23EqN6R5xV6awTUX3YE8xzc87
RviAoyUehMKdktkvRYrtwnfZmhRQNzTSksxjUlgBl/moy2r7zj9IoUzpBov+GYYs8BMI7FHJGfK8
f8seos2dlfON0AEkPK+XhcRTG2AjCEFRxKs4MMzDEa/QeDtJ/21h+117NzX3xuzAQeCwbQd3dOx8
rShFlJj5mrBTff4y55fy8uhTCEyNKdBLoHFm2yD9X1EEI/muyfxHbTTQXORBPr3RexP8CR0pyvL1
UowdO/3zQd813N2MS8QpQ1kdnvB7VoUU7u+UiK2Fo6+1LSw2xq9y8B6mwS7jH48yIYLrcGWYo/Us
DBEHR4eLK+D8gYbskxGgx7zHm6Wyl9e9V4rb38d9h6iw2FYjElRsalzGNgkaEAigTg2trGMq3rw3
oXhPTYGA+RUDnOdNx3rut3P9CpiFLFUAku2rfa4lvwD2TAhsz1BGNUlMkAxajQHfo9R8EsDVi0Gh
KvB2cSHSKWKL49fnY+0/2tqEEUT1E50nFLsdXwCq8xfjh7ydJc8hyv5pC2KiVR5HsdzM1/9eWrg6
0tU1o5z/8GJpwNnO5645jafG2q1nToZkogpdazaW/c4pfyeLUwNXHaTyvaLAbIrBl5bYUHF3Af3/
cELZVxZWezQxOiEPpyFtRWT1bjSj1wOXr66jPXQvx6PlPxECTTnXgHrxnW+5keruSOL4qBSKII+9
kJ6Wgo9zjRaH8bhY+hgP9JLVLn9CB6Sgk1FPn/JJb7wtLl0yNyDl7ZrlBSpj+fiiS36Q6Z7ViRZ7
4/JJDguqY4VT5xwZv3kxu5DPxBhGKnvH5hNhvsqSj5XZWVhGYMSfYXlYH41WADksZayecUfsmnzj
UA5vMK5eivRxdm3mGBW5YoT6fj/1clJVJ3+JGGfG517OSQ08ixG3ELEIYsyDmgoNs1XTkD4DbWX/
Qc04EDU9G92kY//aSskLoxXfDB7nQSmXa/ROtUrK+stdZbQgdeRrqJllW59epgaDhpmqf4G7hjXb
y3CtDdkScnYuRFn6oR2rHY8MlwMHpic/0v4BJ0WxCUKEJbeht7mK3InKpGdV6FLWEZG74ub8LdZG
Jlf4EsPCbIVMbOd89l3AVB1kIgie2bVzzhEI2VKvsyEKvQspdSDOuycoAtmXHoJ2vmQ0ioYnUyWo
F9S2vO81Tl2do+0GRVNOxkI3AOGxKCWyUyZqtX2ZfvdB90bZZ+7HBFtEgs9PXZF5lwhn1mXrzlwg
5s/8XSB5E/maVg1Irk/9yXUMZyMz5+IYoBAAyNILFQ6mdpo4Qmz5YAXRwP2GGsWEuHcWa2dTh1C6
4NMK/o/0FSKpGE/At9ZIub/iyGryRaJU6vUt7NDoLgFHyR44hIgWD/FINxgLE+fwoXHKuJqqTJ4h
0MN/TC4RYl0Lr1/zy/GkQapaHuW4dFHfLxVS8LQ8fbTraz7XHFrTeBleqsslzwYfW/xWRH+M+iZu
s1Qpm2hNRS7NA5Yd+sefo0yhDltfP1Mm/amUA6vef5FBIKV77r+KG/6zkckbckip/Pg9qPYdGIHB
gYvOK20ERnZ1kfOdcQGygrMTJ/6BpgFaMkOX6gccaXZVVqse2nTO2W8Y+9x7ac1h12LibMOn9Y+w
GS4sCWuBGBuK7v/klPOm4MDhKNJ6+5AKqfEkJtLyWaW0mF9rKCgHS/oVP6jlxB4/c1t29A3qd5jj
L4ZNWEHi6Xfk4Jj4Z7Ce1WZch07SOF3hChHWISUxZDi4KwMel34asuC2++PymbFuyz0M/PcfS6bZ
ILUXNGbQKO43m//B6Ge9YK+GE64/a6n77MYDyjD6flp6zMuu2EA3qWmruJ+SybgOCGy+hg5L+0HI
NEN31FqsrfAhndip09gmADLqTZycrIkbE4iHE3oHEsCuK6sx7ZIOT3imoi99RMEi2sl6ZpsFnUVC
tdgpXv+onxPRD1KVVJxP4GcxyPrvmuHU7ApYCPze6IIZ4ekYjnsVl9dKMTC73XGhvDyowdwNkjiD
EAbdwXiKUkXrsI1g+hTZ7beLfMB21eT4VUuin0nZ99LhES+5WKSDWRX4foKPRyqMKOIKLdh2oRhC
Tn7bWSIjtf+42EktVus8mytcIxjRE+ii6YR8Ax8Y7iPevsXhAkyFjehvsd8NoSSilyICvt8rqxat
CQpCNqmsCCNxdRmlc3xuNguLehW7zB0z1mEuVklYvAfo0Qf/ne8ZmTl+0oIp3Wo5XAX5VfdZmphW
seLKNU5IMSq4lYQH4VeHLjGJXcxTcvd0B7bs7OmMWLmNnY0yJNYKEaPfS0M4tPh7H9KeDaZfosJY
Xmku+FCLrjh1dp/Zpf6g3RF0egiwNIsUC0ipgrtq9399+e8m54DYeUbYppwml+IiK0h5rqNm9SBb
5VCde3JoJJfv3/yLLh3CYbVQeY9NOz5vjhKR1t36f99LjGLJFK3L9GCgNEX8tnBeZYNSOarOeAfP
KWXqHzcJ1z5UD3G5QeetCriOqvWAEiwwlEpQk9oEe8yj7l4vYrsmRV2Tr/fC2MocxlSmtjMZqjqw
nInuBv9d0o9Cs3pdJW4QZCRjzd8xoQagejB95otJoAMhwF0cqa9HxaGa4uCAtL3+zrqH9mKru3vY
2r1sVbn6XbJcyRuMTxXc6q5W2W/KwdjK6yjnw6kYO+vQdytkphuz3TDBzedwx0oUxg/DpGFLH92f
SQQkB0nWd6dPujXEZgeQl6EpnnrN5wOLZD4jbjTbXXGMnlx0vSIEXErOS2nTs8cbelrnqYyYrnZl
WUQtdjwgW99mw0/NrD6GhiTV+IHRZHRZZcZrhgYbPLhmqseL/4n1tki1cW9DHJ1Z2VHHD6rGEd5p
9nqVVFUDozMCiOy9OseaVmlId30EJ5yU52gVL2ejlsT5P/6f4Wn57CUkq/Vo3NNE5cRwUYDmg06d
gVW2yqFtsGpscY9RjadC411Z9d6Z1IItiudaR8UyTrfiaTBU601ezIyrdsiorDfc3U/skD2FUDN3
xQAyvTUYCNmCSTet5O3zeHUHSc+T5atlJwJaK19n9xxq+e9YyiDp9BS4lVSClX0EAUyMQMorJ/gF
3WF94NApcI81M8xlE6q79GHzn4BxmYZuG8yc+PyEOGo7TKiM320DQs3gFVlHVLhqYR1y0b/zQ6rL
Z6yGpWV5avftEcBp4VFDs/jQQ3hLdq/dLwlFNYMPaPemvVHGhO8jNXSlQ3+Z9HZmbzYnsk3Pm19C
BG/PquY+WP5tVIv2p+1EOteLiiHxgZg3PZgsznVhBQuEd/9KD+pNhMG9ppQgJ5mBfp2yz6KeOiEi
2tLwdw022x9siva5lNtohECTscoAbwU1sJe4LLY4USMXUikFLPxEhtlSa0VQSuDQfOhytIKl5k00
iAlhCJZnoZ75Ufib3KIDd8NS7qysfNfQth5SkSaOzNfm4uU5pR1BWK12br4iASG80cjqnaAEBgwu
oPT900MMEHSxCGdBOQyJoXXIARsqy3x7uYrFZ/F7CiwLoOJ1rBN8QzmA6aaDmtVBE9/EL7SJymqO
HIRHFdZo33G2wCcw7mV0dx3uFkKsYJhXeMmh1HuLwEiUpl9dMmzfTMVU1dFvNw5bPLYzweTmeEDl
ExORWuGzjPtlf+Wa85Vpq2eAiUyo07/YbK8YUHzVkNB+G52yoH2WNV9kkCIEhsenGafk7Ezie1Rn
KjYtHuEmJW0waAyXDcEctdi8kbprbYkDz+k6m0JBZKyFDX5SdTirip8/3hQ4v504naxZ+AGL4tiF
H+JA1jPhHhKuxuxjO6Lmz70wQqLvh3PbmcvulTYKdjyTQbp+otzvd6ShhsFAHcKiRInyqJtl7xRg
xqOB0xpKsZrd7XUdf120KZroo+2Ty/5gznrMsTVkiJhTzno2bb+u1G4wkofO2MEc3wKEJ+arNVvJ
BaPcEutIR1wLG4lFydVLdbQ/vPT6sMR1nAargkoitIH7d5ovELiPYq4nQ7pVIFz8G+1pfH/84mbG
Q7hK66P0SgBmX9SL/q9ZTs6n7VGe5UmN+wVAe4ejpD6CZFMI9pWBS8gAzBinAgnOY0xfGa+R3vSW
R8uktGZxw3K0zRX0Xxk7qDj8vYDKJEAqFg4gclQn/4+6jScVYh/WQqxTiI4p5UWTZoqH8Hh6PRcc
AzpHWVSqodAA6Z2j3ZwQ/ivZbJm7zKKM6rh+CmaqXLgdH8EAyn685nO1rLA9fto5HFfevbAiWHbq
ciXacUPq7vC2e2A4GxdBwktMeFFMXqHVQpak8L/Zbev5Xqqyn63cI00qpuvS8bg9kx6qqCUW/8a0
/oTJMRARNq+MEY1QJ/77g9PMJWnxX9lBcZzAOozP0G+opTfYgGLBgT2TJ6JP7kVUb/9GtuQdIMPu
HGEcwBB6OLye+sJcoo9Nm0dLjIBUDOkrN+BDuTJGtishRQ0xfQbKJXyLDY4H7UG7zV/2/hC2B/JX
NOpDsEB1iX6LIuCdQgIiB9GAQSpWn1+hX51f9SuG+6U21Y61IDDYqpZCT5gU8RmRX8RVS9xkd0Lv
O74J/dWhcQOdRdYcNmjY/9DUODlALBG31QG3IEf67ypxagKkFeUG0MjOV5lMwSFFe8mH2n6+KDlB
S931i2vzFcwiKZ9TkkoreERFS1BUux2z9YzklJ6tJzNxGNUpgYwGOiZjwG046RnJBhAZ6JeosteH
hwdBa3rPYcTKdqKJP7I6v8oc0bOFpAzpR2VpsiIeZ5EYiua6l5lmgxAZQTbnLE6glTKAEWfSsrCy
X0M6G75hIjnTwjcfMp9G0GOWkSXYQ+98m5QXispaWcVEHEDslV4uuJAu2cTqFsl+Ahb+SW+lKTNw
JuTgeNFCk1FBQ6temHEwM/Dsmln/23e0bpTpYAMeBykxoGDRILzQy4t+wJELVhPKw0nzFDq0yHK8
x+uVNxAYxPrRfoeUR66ZmJ1fIdr+y6zYktpI2FB4Psv0bpi1a6p/SKVrwaKRpCmOfJTHWNS2gXok
FqpS59ztOGLxI5PihclOthFqXH9x3Rui5UCVMgOE8EbtW+KfEGOmGR4NYxVCe0CWMcz4nSUhchk0
NW684DuE0ivobYTp0D36nOJtDLey5NM26zaq3Pmrm2bd3yazotWB5yFzFmVwWwTII+IolS8kn4NE
pLfPyQnaSrEbWLej8SPDSDjmuuAncyzHLjFblejjjpU0fDRDx/vTbiRNlWKy8zmoeCXDd4AgIczF
ngTSfnGHeLBAa53iUiqyDlC90/RyluiuOWxLWe0eDh3WmKWNLxhdHU04UiKLGnlU9W2mGJUhmljP
nY0zoyortIwv/77DuhE0j75K0ADQeG2yUX7nhj5ujqpIH8YGvfSezb1mWiEYLGVph2GoThTs2hs8
bRAmLwSN63x+wtnd+OcEmF5WBJlfJYp3Lmjc0EpqzWl5sKWth7o3T4z0t76dt6jAqqSh3hGK2p/V
ooYMhjbYxLsJ89XGWOmhQFvSXpAlWegBVenfeXn8r4r0XrgRiXakY0ZRrg0VqQImRdGRhUWeB1tU
qHprQW6ZF9lFPO/N89bDT1MwI86obJya5H7lfNmcLLu9GrormgXqLCj87o69nyBFw4r21kF7OmzY
rmmRm6YXV9hJWxjO21zElAKQ+SnL5OcllwCnDyVCxepZB+kogz2tsnraTzospY5MMynFk+eg+qAS
Zm4lmH2ax4HKZX0Ut9K/aWL6cXdkz+Y/ofq5o8EUq00Jc/37I6G8G27FeU4cBQVvE0GldQSVlKXO
4E/2W3VIVurw//5mI9ZL3Ts/HS2TSElR49n39p4Jc9IeewB9/rAtCQywnirY9dYsasNl8t11A1Oe
qV0+25ru657uT0DS62Y+oKD4aXurb2k9cLKX8OVZ/ToCxf3ShRyJ5AZCSX/N1XPDWjrETFc9gQ1f
9MYocKo8GrFbey51p8fUGiywg4A8ogUEblnQRQP18G786UDWR+lmCmM73bkXa99e0ASyd+rAkL23
NfuPjL4WYG9pX/yFrox0+I7U8we2OYJTG3QZtrJ4XRZFNg/oeP5JXNNK7jgqLJbmyOrkTjuXBrgB
za9zelG9MjRk30PbjROGWc+fPBMx2WcBswvbkag4OdK0XRv5YG5l+pgdmycs/+G+01LmuOhSu06L
JgAgWy0+h08BCLC5qYfjxnFI2ejzg8HZkIg+wLiyQ/CijxJsDJIqjhs/LfvafOXBmmKuxlrPuAK0
Y52VsUPCWqHxQUY3R89QpDHsqMjccoTcq+RFVbOhEX7vQg5TUZe8sXEJlVQBtHsZM+OwKiRDfzWf
PGyYwbMB1BK+BowoS1kLdBgyt0r3aXXk8wgm+B4+VSO98ElIpHCRWyO4OmxGX/DvIsqyeqv7Hsza
YLM3QXwTF2IDhkBMnctp6mG/pnPQepgfmP2k6x8GPtoXD1tTOB2B9TZW/BA4HP9Sy1NoND2W7pdo
GR4qZpgR55U14iEsIL8Ib/Mn4P7Fc28pW375EQFHniXFfHlWZc2wJO4OR8ZVVGs2u7OQQBEDVVXp
jjYQaX1XMQJBTT+UnAawDJPJoZiwlD1L6zrVcWevbYgF7d90I57Jucr1sR+lielYeeBElngIfHpf
avYiWoU94ZJZqUe75Py9NIwclEuKt4sNiHUT5NKP+kq0396GOVjeFM2Yb1mCX/NC6z6ZZryCJESd
oaSaG6X9L9QB4rRVC07mii8fl5y9mMjHDTnf2WHH466bj7HteWiZjbQG8jglNrtBudUSw91fpvrn
HBgJUvZ3hdtyOyQQ5TkzySvbiL8TTdsKbepQ7BY8KkHvweyuIFcoiQq9r+Ti8Z2Sc5Ll+qKUPUao
G+sNu0uTcv9QGcGpDglrhdRZXw1hkTlhEZ6M7SWkyorLM3bh6X022l/Wy/4RURyKgZMUnnoWIHEZ
FgFWKP0MinnMSD4J9RIgcKoJaJJAHp3kcWMy38x5IXrGmKpM88dwUtLytIhMzjenhijQXYcoQJqs
tv9a2Ggy+DmXzPR1i5Ls78tHm38qvONvd8OXv4CcC9NI1CNkk22/kaeyAUHKHAjpPjZZMpQM2H2m
tIZPyz68f3pV6CZQwn68mMW4iHetyQAxKBtMvT1HlEw63SAkUQANOax6fOaZk/hyzuFWH9abdFD/
NWyX5ZN9Ns+uNuw7xcAkjR/v2vbytll2bbfHzEPvseIOdn2u09H7AcjfNCbzefRsY33PUYMyUk4M
g8Pcpzt+1AmkWh2NR8p85K5ndfGllrxYslxDsZt4sYJXrPJQ9KTGsf8YtYhJ2fUA4PnzPPVH+KDI
/BB+4rd8vy3cuodf8nPKXbpQLK2zTeX+fH4U3b2ByKLMK3qRi9BD2vTMwhB9BJJpScfLoSTgNrxt
2d1uanv0N0bPv9Kh7UmjblVHQ1kF3SyQUbFmJxtm2/mUxmQpASXJC4N3ZGcJtrHnXCm7P2i4x5wK
OiXZTP7jUUkIWpzbq7zlfkf4B3RHKsqLiaj0wnm3ug2fGq8FRfS42Ci9gXWAu6fYXPfTMMEhvSMR
76kGOY4UWj1xcHK28aThrr66wBa3FOWHV2171FckECGChH0MgIiJHV9zSWtHA4GfSctvDtNLnda7
fGyAWIK3bXshSp2cJ53LRzAUg9jIeZhUxst/pFOFsTHLth8PagzZlM0iUY13eru1Dvm7ZCsFBC/V
qcAUjZW1/xZE1iMhYzZgBYNlA5zufQSJ3phm8XNvfBidU5+YT9Va4r2G4fR6ftD6eMcBKRGM4vde
gZIR39xaKdBe1KdSFhpDjAR5juwShVVQghvRj/jbVuTrMMj2iemrWAhXjkcbt05NqqgEXmRI91Nb
xPxRIBHqSoVe+Z0B054b4k5Mx3FH/iuQTTNR5dH2Eti8sbGfCIwF5BCp7Ypt3LCJ9ad1kU2oxBzS
BB3TYbkET9if2zR2F7D/v2/jSO37DfaLnz0CBJJ2RxybFtYZyaQRETnTArUgn3YbPdI8VlFCvtvt
0S8Ro2786AQyYCOQTF3TE+I5wfADyVQwouKV4s2Q42DrgbaTfKuPF4rg3Ng/pRZYNPj9q58at75W
WZZwIruHVjwIr8VfonX/bAJ2xAVABsGQCMwTLfpg4BHAldnD9+skFFyXK937qtJjD6ma1sYRkg88
hzpJ8zrR+yDlo3LsYAj0b3Jq764vea5pWQlqoHXivrGWKL/+WIc1ohKjXNRkwpMkrAQEhM0/m1Tj
rpQilz9l//cOYKYUIv1hugU7mGm1zkt2Tdk2wzLQfe/XUY4GBTCRJzz881mfEmBkiT7sq6WRKVwH
vkV8cS/faIcYO5rMxrw0DUJ/15vJiYq+CGAETkOnNlhJhT9fP5r8Akc6wD5ZPuwKGmaOt4nMMEgU
SIC3OkubO7tU0ZED6Zz9VQ6CYNfpawh9hdVMrSZzJwfll/kgu5FPRAKTFuBf5dQjLZYL7YiRz16e
+a86+n1loegV67NTgyGgPhn3sIuT+FlXfbZ3G57LznAB+IhgXbUltlW+2q7BgCb+5P57BbCqLi8P
isVfDSivYI5obsQFOn+bIzpSKfLOUd0GikP+lPbeBFQRDhJpHSQdxcL3UVC7ue4utnakpaMNF8C4
TEr4i+Rqdf4UP0psgtoXG33iqM/7O0eEuaFV3GF63Jpnd2FpaPxmuPg+DZC5t0wEceajHNtgBWRE
PEWhM8X27BGfo+3DQGwi6tUoLN17l6/VNZgTg5DP64wEj/T2waoFVS/Ja2Azrp0PMih7kX1j3fFw
CctAJpR0/fve6Crjblhr9Y/igbd/6BQEXTy+7pPSjOFCy3nMzt15fhoIDn3PDPUAtxohBcs54m8B
9+jmZl62Mt4970yhKO4tVc7cd+8Vg6WGLFuVwqWdhnGMZ3MOnA7AmNnzo1uGZWnwBMhS5Hra0T7s
sq0WrQ0vYvevrtvBt/OTM0TcT2k9hWjOIBXvkfFg/Ve8gkSYD56yzqY4V5qFU+R+Vzv80amZcrAr
jQJBUV/8Lj6+zzhIVbAGObvyIqYdzMHwd9xRFJ6u9TgcvTqtOaTSjBG215v8kEc3gq9KwLx7ka2Q
GBA5rSD+pkv2i6swMXtBOpmVX8ORxeQlMU27igTGv1G2ixdgOABZDE9MoThnJQjcD0tEomcERVzU
Z7JmRahDhLG04fciDBDGehQlI/G25Yv3/fEVLYxx9szejGkaGmeFEkLCh/RO6KdQ8ZWdztlpWDZw
B6UKu0S+uLsP1ZiTpbqs3tvh6VELBt36oyP9a5yrlyAnXfA6SlIG7v3CxZPcZkt4/H6lPOSTKCoU
NyfTrDpisyHQIDx+q0tpXvBAK3HO3Dh+QqMHXN2AbES678Cqii5cfF8SCm0VDl0RRxlTXPzof6zV
i6msM8Q6Po8C81o3JtXOENeqXMQi2wUBDkensXNS6BNKGQBwUpah5qpNBd+P2n6QXPryo6TcCYEx
Qg3VzbJ4SfI2al4LEnQT5HrrEnJlJbtxqc6Xwg03c27c/ITMNClj5T4Yn+99oPB6z/cttoFn+BZX
h0LVZ1FxfxXLH0+qIVUKY91EveN0DSYqEf6wOGO/Ev4T4+hoQ6PmuF6YGWD61yKpRvI2cxNqqBDz
zZWlmO0DKGHaueeC5/R0scpRLAtSLHQKhLMVI8TebY8sMvksCwejlJkP5J4YNnjS5aC467zPDYHt
1W+DilsYCDUW5M2A6sLfhlhmoEFgtyYW3SDmbNQPz3vhVfN33aDL6SzfqjxCsMAnsUzL7ZEbZ06O
1ytaShLvAVlpN10l1sbD1ci6HiqLyIMnCE99U5eahc/Ofcmh9SyyVo+gELWKG2a3Y7MYLmQ0wCqo
KyymOOW3Rb4boKr5T6Ih5GWolFNbubF/mzsYGFrRRG72JQ3DUpAmqxOzvwrIIhUfwoUN9QtE6yBB
Vk68joJjplFGejShrz4HGee12uarSAhINi1tT99pxBxYFHzH1HZVTqsnulFJahZKFohPJ28qumNk
2wl02mG47yaR8PwuNwHC/aH32ZBJ7jj6fqaaEUTxEqZ8YFqtG4BlLHKBzuGCmpUhFRBpGJPfR6hK
mvV3mxL2r37ItVGOlGjgYxqJiX+AizEXl0XpPjUMjkwRRGMBxLmwj7Riy1vDugMdskkFYSPBm+UT
+fvpZmF7hgBUI/vRS1a1khZv+eVT8hMi6mZVjvf4k/RnSVCqHF6KgLgKVKbvgxmmrXqjH3URAISt
BUE4ey1EdIvxhz8Fj5urmPUqfwamAxtxTWdQMuIAr+5K3upgX3jxze/Wd6J8tTUbA0nbpUbBdGns
qCWGn+fimUjc/mefyEAS6+k0iVm45JGUIxEx2axK2Ns2Y4zOtjZEfJVxYdl69t0iEqfFt2s40sMm
EgHY+Jpw8+Vd4MSL20uHikJ6um/hpZ2fGPotgItwOeP5UtQt1kqI4FMSGE2ZjXwXZW0iWBgnqPoH
lsL6S1zHQ9ANIjO0EPOsNYiFTJmHQelXucyZgM88dAPebWxiUivV87hCUz72wf83HzrdjWgE5i8G
YiGOGHE5Z/uqdzAQisEzQ8QaWeLBpf/3ShPuPlSPysFhUtn2HgJESawNXyTt8AV4t9mkosrqcmc9
k4KyZhIh57dGytZ03AMZF5FO3EuLEkkr6yELlBm1yeDyHJ+VRV+w5qXchjLMKy5V92oBrOPVLZBD
XSuUgTARAAFcUrMik+Gs/qDyYwaiyx9GkBj3iSSmPK5XSedpBPoFMMOHCTq4ti5IASEY2Qka1gGJ
EtmZNdYKXSGe8aKVUqdmCSbiPcZEfjwH/YnAtcMFtZoGflZb9m3iaBAmxPwYJcpoKpRDV6nu8xn8
EbDdvLfeIP84XPtv7HG1upDOBcqKib+kx2m3y+g6Jos+vEJpk88i0T0lDrMdDlHrFCPrEXI4yjqu
E8AKhO/iKZiXMvGGkxm2pJiqVncgamnSt5TYyvD/izjEe0Jv09OOIZW962NBrc0AnIzR5T8F5P7I
Z4sp1tD1TWs+Fyz4IfEKCFyhD+/DbDUWQh1LkyOT7nrz/SGLBGk+Uo72FBhIFR/d+Ic8WaHkL+E4
fwLeGF2U+Qk+JThohV3F9/Hlmz/oUONgsXOzKnboVGAqVnpR8hvAIZ8FcjqR66PObgWIN8vy/DjY
5vMfvh11aWAw/IoSld6OQnpUnLuXhXj1DzDgcGLfvZaabPbvybLWpz6/dbFZWHhItH9HXgZpWzU3
MC7j2Jxfz3aLILV6rdIR6ErzgwH89h0++BwODSQ3ttpaDmHtwmEZsjDenbnnOghB/R/jsxYpct5n
LHZZomeedCfU0PvxVDKJouPXAuOSFNusNKFzOTxNcAoap+Tp54OwXjh2lWf4+WT6+YVLs+nmFDeC
WjpayhoAV1a149Cv8vrIu2D1haC4ZjUKU2eLVWAg7jxc/pBtnaw9zXp5gpyNoorHM2rwQ7sejwQK
Cbmdz8CZReo/FiuE9Z6XjTuVN+eulC8hWvxHv7ZogbxBJMPS8V9RjZ33tfjGYowYg7Wc1mA/etON
c4GoMZHZciyi5XLrDO3AiLerMSFGGx4LOr0TLvJ8pgANJNvyePR398xOxCq9FOIbpcB7v+ygUL3T
tHhxHoI2ZHO7PenHwOzf5ydIpywLA8wiai4aJY9mBqiwDTD7FETtisOB3TSpv+I/3aJkF65dFMRK
QyG9m+wzdpbU4D/fS8rutOx/03Xzgu7wv3PaZbOorLqZJ1geoQXzYW5Yq5Oara090335s62SRIBe
2zYc8j2nSe4GzOfEYUyytJ6pWM2zi7K1LaQFQ7Pk7lzElDLH+DB5iyX4ANWOU7xJj6HLh19rnxDF
cdqMots+o5+Hj9CIeYAf1UVnzp6sL3JhQ61kSCxYStJJwGPh9Vj2M93FS60CDjLTgW5i1dxAR6ej
aJPLdVGUXrw/bqtOvJ3YY/PE5wIR6dij7Q7IqcgTS2BbG3w1TXrLCwcJfYPe6eMQnlKmS18C3O9g
AtubC5zp0rpP4FhdLFWMrAGKNg3iMaenAZIMudZpyBkFJPJhkVQSrGabvVCnqevxFVDJtRWgrqe8
iXBA+mX7qDSzj49/c51jvDLMgEnJgky3D9MwXaGgPmodSvV7Q0Zw70vyKp4DzqMT4RzghtTLH63t
IyFT9Y3boZg/3FrfjG6aS2oa9Ja4v558zesqlOhzsak+ejo+D8cfEg+g3i0YCwfMk2CF85HU/hYH
2137VdtQ8IaI8fAKehT5ruozO/VU0Zh65mhzPim+CWLRwwULgompFf0O9w8qkc71nAArXU6J39oa
EYZSP+m2LITA/lFHSVw3NNw3r4ZJNBZtdp+IaOdafgOD7MPR0Y1XJ2Q1RW0sDtmRr0TmnWv3rZWq
Nbeb8iOR4wAYmGl9GcX8hF+IiR8G6Ue28i8AXSxgmjSIDYHazsHcnsSe6k+Hco1A5h1uPBClxfHh
FOBWK4OtHitgM6iWg6OnmL3Lr2uVcDqpmP8Ps3TxDMCov93sLxccBKRuK3V1okdbuuaaxW8/+iSd
oU0uwCWojT+aKIyBM0chbSS+axzZD2L1nPLQSK0xhhpRIEPjVlq2yD+u2XIZsoKpSff/U1Z/KRR1
adWq+aPrfz+UW9zm5UlxKiWBDZzKELFrXVJItiH5KlKD0I4qZE5kqCZk4kY/pTggC09pH6oHeAoU
fvQRhoQuKxAH2dkwN03k6o8+jk853xFi2cN5mYYc3AsiiXCol7l/ZyCK9IiK1jgN0GqcuQqxJoBz
vN3Ms1KNmqxabFxxO2Qu+JOKIhVvrMH/3UcLVhlaIUw4fWyI3tU6bOmW78TE8ZVjhRzjI6KUy49v
jwtXWU4NAIAtAeQ4CvS0De1QJ2vxPVS4ht8/2uivg+aXkPNfiRE9YgZxAsyuXmRkzuF1sx/yTTj2
F71GxWmdNj4JBh8oA7xwmfUcFQAO916Mvpmx1R11nPoZx1TenE2icpXiQSOoQsZktn6/Sn5Js7DL
B3QuS0Qv7SKfzkRP0A+/mp60wWDJB6/g9WsiZfmdysaAQHBkYDmmvU0mudcenx4Fh/yJQK8DYk/y
gOQfJJqmMTzDgNMP+zmTvVHwCkR+QW9kSfuD8pjkfD01VkLcMqTrVmDmmi4tZ8dYImy93yKdjHAA
s8i3nwue8P4WvtVRLJIzS64Tk12pA/hJN0VizkJ5S7td2K7orOiWmZTsb4SzfdNT9Y9BdeK5FVoi
DmE2WZMZ+Va4nh5W6V86KrBG7vEMG1Paba6KSfOnmTH2IyG6Wy0uG+jm6Lu9IU01robCpyrtZn0I
qs32VZJY9pGrXTLduXXdlxxLWFCsxvVhfs3Y85LkZimLyEBfs5nNthOG/VrJVGxD1VDAlP6pkpeQ
Q+mdblYo4IwNVKxh/A64S+NXtZ2inz58uDUEqWnhO021mEifvkqwHmfX3bjRnb1XauUUql6v3D5s
me8rkytESE/tp+0ZGgbzhzzTP/6eFP3SiSXxPhJe/lw1/VclzYg5FhzH9Vf2nIs2KwEOAo9BH4Pr
7mOOl1gMyzq+/flIChMYe5Yd7TLnSv0TERf2p/dDXYNomHh6u3sUY2Pl8063p3ZRFaX8RiNCbIlM
+78xDa9H8xz7wdyuwwO+2TbAKc0obRG20cJT/k523a/QGJpfLZnhTcHfeYNR5k5aAdgc/03bQfQu
cfcFkS3uI/CuOhT+AI6ZthK81ry/VA638hHT/Y0tWJu+riaAasGuq29Vsylxwquqg9rUOhGmLzYC
sjolnlAfHYLC6gdWCDSyLaUu+uf+rdz/4WfE/xK0viGhm3n6A5IKFlTlJFDAbJLUip7OI6GR+cGE
4TLjE/Ipb3RstUIO1zOF+HJoOEkCWG/itSfERKsEjnVJZBnzFJBTHekvU85VI6W+EoJBc+VuVRj0
oUn1qKE4JHHZDQGn5R9k6I2hjJwPC+LNELJ6pUUvPiw0cLoh8W63v/qx4VkxvPnvEUoUmgnhPMAm
PgW6aZQaZdwzTHGAvpBE7bwas05e1JdycvQI3vTD2tV6GmiUWrQys6B4dxKSP+MKXZ58Bijse9l/
HH7Ol2RDuxA4Ugalco8PVNfO65oSWxnzWW3pLh0nQyJU+phoVp+lqUf3OLzwFBaOorpsvhQann/p
cvVuDfi7puG9eM2Sm8SFhJ1m9YieGhOTH3J24cJs4MsIVOp8C0ZH2iIe9zvPqzQYW26sDrPUtCmw
pF+eRkjTCWIk1Z+KQzddLdwaWaSA2OlsMOerlrO38m6YzHFaUzncMblGZGJKn7z5duWPtNHBZr85
OOAnH+02S481Adkr41IUvJ7ODR3EVB1k7JSgPdZuPM+rFHa3IYx6q7pkyZT9Gdgeiy2d0fyTDomA
cW9Wi7dR8ZUysKSxj9KF7FLFSbmvDJ5ahMztDu8sMB3KQztROYhNkLD/Xf5LRpCTJTRQiNH8lIgy
jy6wLT8qg1lBTdl2wIF+VgCMbGrkWEyXDi50wtIeiibM2qVfEodw9eTXLsHvvfQIyerk1yx9Ippa
9jkIkTr/4LrwZADrR1nYreRkiX/fNuxhJ8RaOBDQtK1YTKCfOOfXyV6ugc7poObk5fw2x0OvDjWe
7UcGnMkhgK9yRg1COYrxf5gDG1jdQqOb42LrxS2zCoKTtE/5QHLYHS7z7cHPacBUOdgC7ixAG9Sb
jYbYyGHMSILU5cMM4TegwAf9y24dsJaLwhgFuyfmXJMVPTRjmrzw4bsFWPggAjBs0wG+TdFZy9Ko
Os2cM3uotqx+HZiQERI8eAY5YH9hYZASQFF9H9oCH1mX+KbLuVVI6CX4Ys4D5VmotdsxXRKo99GS
OQ5IR4LVouNKOrINvFKdiAzVEuL9MTm/slN//F7WXlEHOOyDRyMH4LzKac+1RSgyhRWkZpjACAnm
Q5WbcT7j9/fStygZBad9jeJIBoFq0vm/RKAbq5CMvb8JFc8vmi0Q0qdi1wKXavvYebPgf/NQTSOh
CRWBmvOXP/R18ntztWhrHFmq4xSPFIeZiIvFA24lPrmSh1FBUeUoJ/BaQ8Nc/+fviAbGk7M0HJUv
RbxlSTDbTBAa3/5y5EvFv1FTFVMWx1LpN8EQwhdupnvRkwohL9sw7l9VEtKfdE6V3V3vYW8oEY3E
4BAJG+8K98rM1kTcEOa/hrIcuho8VphuMc/c9z1D/ROzIN96ehYIAHY9+j69pmQ4o8jbrFbXmEqx
cb5S3uSCEKhC7AZf+YFjgdqwbD9BfPTSzJjPYpLV6g2DTVZ1j/EeL7Oz3DKeQrHBGKBBAzQVQaps
YP+zCOp0x/oIqMXdqj91jyBwNHwmBeIoWhOvkzpOpyvbcuKLs/3mQ5jyufgolFo4drsBhXPtcbfP
ub25IUip0DHi1PpbLZ0qO8nxoZt3zdlMHYuE/4BKaqrtgZb6tcjWIvSfahbX9OoU9l4WIDGMhCoI
Bl/xSjSM2PfGr1d6TQEEWkVtTtSug6pANjeNFKewkJ0JxOhnoOOlP9t+2QI9rd4lbP90wrBw10ci
b43a6LqKsjYxePCBrFmhGHujFbsn5Q/dYEXsa7SACrDfxTltfF3vMqq62uY+61pLpkM0zm+IFWIy
sHKuMKGzfvZFSqeKObM0MtakaZpVBNp7yvVbePbTcFztKb1DPfPd7H/9w2qsOhKI9V06lUqHxkyP
F4xhZX4soAXXuO9qR5nJqdurUzY0MaRlI6N0r9hyCudjDUXx6p9FTiTUufco8gHWYcih1NZ4PxtM
b1rTW7ucxN46/X30YS4gpn4uVvUfdUYcdZhr64CGGIPBhDFguJN8y2rXqW2WVJyaZKMvXmKw47pB
I5aDyjxBHpOj3LLK4TmKRtvRBtvmQ9lXO+AsGxMuPw4oU3VZQ6CGew6S0G9y6poQRTnzWe8YaHZO
HZ8PACffIZW83hFbshO5EAicofvyKuexPNo+Np2OrjHSVs05Prn3yU5qtIPhVvPofs7Jin6Q5jJO
AJxjc5xQLff3UW3ExoayLIIX63hfyyP1Glo4ofOhArIYsnlLqStS4dsw2BGpc7DNcu3ndyCdhegQ
HDyanPl9gaoDRzx+8Eko9mdXkIaDmxECS0VZ4WWJAQa4abLcbPOQqh7PS40kvkxw/WHdsglckvZv
Gz5+CCREh9UU18CQzQimktJzeEl9vYgsK8/FA26ZL97scB0oNh3mWaqrXNBXd+5fbTlBKy9RQka7
xyT1Pr/Iuhs21y3hqTwXfAcu2aK6pamYJk4Jm9pJVq3RNjYUbD8ZjT5DAMQN1tTl9oB3P1JyQFtZ
EYH5Dx+DvN7XVTwgKL2Yzu9aIoi1p/zuB2WhsoR1kTnvCxR/EqrPjmAva42b32CNt/yuO2fw+GHz
41oQghl0HCdPNBTy3NUWhCi23DlKyYKwZmC171wIYevnnCaLq0WZRHnxTUS+5uUEzNpoceO0wVUb
yWl7Fnf8659YlUieJH18cQ4RaZLu9HRACdzM+Ec8yOhJn3FfLpzd4PSBsNoKhpsSKSmddQOVqsKz
IWtSawgKJ6diOnGxQrjd624zFE/CaD7351NUE5mdCg4u2HBWZFzRjKtTjGjq8Rc01PyN3xgIh/C0
tzLe0XXopzNqpWMr2r4b9qY7OvCX6YYKDtZsH4TM4roo17pk08CeSpwPlvwivws2Iiey2E9f9UK8
8NF51meUYQVMazc+sB7rhfeqd22dmgLB+8qsLOAEpE0NmIVKKQS31WiG+LP9KFgh3/JcePmjgC0o
TpJDXKuTjvqMHLVZ5cJLBYGAUHfDLkchO/2Y51R4ok3QV/bs9OsXR+9Ta9ayBV2qXTL2R9rPQe82
TYl69YGtW6ie/itl74w7ZVLw5g1RMeWErMBpby02sgorFvXeBeixW1jpWnIf/xyojsaDy11g/y9c
9HB1G2TxjcThpd2RoadSusQgkbhKgLmwPe2WDCwG2ymEZwMZ0bvViN0IYctbY13D8FyfEID8Styy
gCoFZgqA0ejfdx1AvldBg7po+0HXK0WF5BsfMeETku8pgHK337vYfhFtPQvm9B/HnSWZ5PIuTdED
K8xiHExAxFX9VSj6Kae5X8MIdaXqz7nMiNUxglaLAsP+VbcRttJ528mW6K0bvEQx60bu087/kwJB
S6GVOLayXnPYbwvxd8FOVWMV+FUabFevkKUUIGnE0WaZD7bUWwbYwsTP3ZeM13q9uvglr+eoaOX/
Z5XjXJ1w+xehICTkfMBSB7oIhDkS6QTnIZ1d5zdNkc4IPXXoG8bDe0wfMtBT5nOANtrhhVKskxq0
IhOb5FeazYfPxpTu5StMkXrYlZbtJPLGfmRrbeY42wLMYlcIdmJgWJZEDBSWIfPriUU30ifivIJO
D7yR9oAXHeWCF3c0c816R86pIomxEPTA575iN8M5xT0Q7yM5Lvz4kiRqEWNrrTEfTihLno/BdW3P
O8+ZdVITsES3SKj1H9/6gvbMe/tVd4604Z2C1kNGTXvbbnweYuDChoXJOOW6J6Robb42Ldqrzehn
taWUaVVZ0ZV19bYp9wlS3jtXqZx/fP0L+qRoXOMzXxy2B7D+MUHtw6KFphVHhJcVAxh5uSy4mm6C
bm8zXr7XLazJ7QKPCBIASozBMWGzNjDTaqD5maZg2MhHYJ7mWH/a3BLeW94Vb6B6qR8qdeXO31D5
9+Wlhkp+QCnF1uuwbXH6NtVCt8Gp+f/nq8k+nu8epvNrDKjqMHpWfzbmgFPkswFrfsQIcfS57LDg
QPCtFJrkoM3joXBLwNCtTyK8yCleI9y33/T7VVHwQ8zRnEP4mFMq5bNVUeToX5xtugtbsk/Z8GGr
dx21ckMytIdtFO0g959xYch8eyj0yueBWPDnhvSwx9Qy+Y9st//9JS0xpbWANP6Fgn64tSUQ0PFO
P4pEEYB0liy6MZhRusz2inPcdmGe/IrYBa62n7IHN+2ZJ3Q62g1OEX39OhQpwCCF6pMIn4g98Txl
KNuNptp8TRdsn/plcfyvmKQClxGZNdREJFOF7Vv/KrPw9zMtI0k2n/laOky4jG5x1+9r8045nC/z
cGSYtIczawpfuSQQ5GSV1I9EFDkt+MjRrfhPcaTzUHb3DQn41JrgUxITvuSJcUe+7XUX8qXrboEc
DygtrKbnrk1Q+/EEokdvXyiXQea9rKQJhQdPptJvEod8c2QQGgnxKw+XSKjbOc5fRy+y5ne/CxY5
Nihoxj56d7OvHx9bEw5pMl2+Ne+4BSLDEW5EblAcODlKQymoUz/NK6uaLEhIB/RKo231Lo1AYXjV
XEOIjWgVZeugQSZ7l32BYWmfod9YZbty6oAvjPKTXbxCcWtpOERYqMMmw8U5n8PpfuWGhb5SaIhX
Tuf/I6vawTemNnlB5iCIMK6zHamUFXqegdr/SQ6bT0zhSyKkmrtHeXBphc8yqmoyQFptL8jUICcR
UH0+6RDWUA+IK4qKW6vPDmcVwzgL2XNPsevju6kS5fkoFC63brXk+cZnV7IvDrSAJ0PiZxiPHhu0
7pSbRsAM6OL5lO9Om+UErHMNqpuc7rUymcZ+fzk7VWpvsji8k1wNi5m7hxUbqAxDtWb1Sfp3TQ9e
pe48+TPiaWRUo03mH34sK7fYLoFX/IFF/Fk3qiucShkhQ9zgGseQFDcXLYiW5zkhcJ2O6QI9KcIe
9JNwYyeVTdZo4r1IT+EUG4bUpw7ePCXED6IA+0AE6SxfnwiMv6GcvMmX9zaWPgEbSdJ4mOAjGKvF
4m4VKge6E6P5Ta+pj7ZpMHg5lBQHIgvtLFr6c7W3qxc3LtJum3XVsQOK1UwXghQpxgfJgwW+HUBq
VtlMt+fnELRmSeKrTZcKfcAwIQZ0N+zOVAWqMVjyEEt0IkihIaJNJHHU5t7cDbjtzZrxwRrMIKIe
WrkkUiyYnsReqv6I3iXC8h+ZfSFgkCshsZkbZubUSCtYKI6vsSSw9MLCCd+cDjVl67qqe2v8ifnV
X2FAZMpykd/FhA/lEdY1RF2RUIh1oBgSEmJKqF8DRbMdOi3duRpG2B9AwN8wBI0uE+8Xf8UJs+c/
e/D0xWguQ5OJLa9W3s/sckfIRc6SzNjxFtmEnr+L36rUJRwfKkDl3wnWoQuBn0xWNfPg6qsmoZU9
B5LCICdle3vS5gX2p5+rLY0Go1YMVvqRqK8vx9t1Xf0fQaCzsVOvI9+BFLRxNGJd9Bjtlk/ekGun
v0uX88AvTdLPEPjR4MzhEnhPU4Uy+XSdqs6jUvTWGCSIkAu//OrU2qyJZ6OsLQ4aT2mrSSkMlyON
MC5F5hX8LxTRU/FRiMRUdvApp1GPxN7qJp2MpNC0TKBl1wQJZxnaa6ocZROR5poqYkIVL1Z47Amu
BmFrOqxWpqqUc2Jc1D9Pvu3F9YBOpkLZbzLuGrVE71G/nu2NVKE2OElrPdXJQWS/vU6ksEmYjGCU
kAm40u/oZyY5xSTh+096PXSi1VZv5RuU173UwL+mef9rtZFb5Lj0onvZ5GXH8a9NWytYy81Stdja
QRjT2W5HZqrFSeTuoFO8WvHxWdktwlFe33A0tYMmyprngd8dcErIlSQdZ4US0xGw/+ueqoX6ORtd
iiaMCZij7VgKthOkORijYfjgRfxaLh9YN7jYsI4oyoVZLg3PtRZeLRAi7TOYZ3c89h+vUhQNRArf
tnCsPu0gpvr3mRsgXm24iWn897Z7EXM245n9BEEeDrhRjDQkzsZqtypyTbjhzX3Jna3nPOadWp9X
nGwy8lY7aqAELZInMxTUJNvzaBPpix5aULT3c4Xw4kl1QQiwr4EcA4SheTJoUQdxodrNgORj12ax
+YhHVH4ThSXC79UI8Ze+wv8AdwFODZFvlGvZ6TRWpT+c4gAp40DwlQIqMMikjvC0LgJG1T7aeAbJ
60bsVgoBFE/4qIQxYC+msk12r+augL3z8zFk4k0n1/TqQvbt1gGSDQu5FxviWBORLS+zl2GTm59b
k1GDoEsFz10+CaPJcgFMoXzAESwfE30tTd1Etoeo1q1A3rAZWb4mWNQowtb1VZHdagXowG24ZMqZ
q9o8A+dq/B+aub5yaJjEn6B1G0/V6UbaTUv1zCFXvPo4/F6qr3MZ7Czc02B+x4seaMu564TsvnYC
eQHLTbUHXGBzJYZHdJmVfxT+v2NJppTAarqLPawVsCwtUHVg7CYfZqxRDHbIQkny+EyOT9adHnzA
6vcfzPv+Qioku8BCUb/t6N9+G8VAvpD5RcfU1ULqDw8TutxH7QSCZ6Kd6BzumpvfURi3ALyOLMZp
xwL99PIFkHGGyHqdZGNwciyF7DUystyuYu9tTgdt2+Dfean9Tg8JG1Kny6lfRrarDPCY4DHqf7F5
5AarQphbDFcxvlMZeQUcWfzRjJpHbkcWHzJJz5RnU6cH/O6shM6fiF+mE06ru8em+gtZRMR9HNn2
09wry0KDOSbHQjx05I9yICh3+QAw+yilBi/Cl4cK75DwmG2wqLKHs2NhU5O3+RzFQW9gQuwUq45s
/GUl8b1UoPvI1GykFqc3uw+HysZXGcuI1DcZk0bcznk73zT+R42kkLgLuxMhRrooehVqD+7Vj9Dx
/iFkwq0r6ytpIYVkZp0mGwiOwU3KGlc46thYyPDO70YX4J4aTMKxtG5Lk/3vYYJNFAZDqmmyHld7
riTfASjMuaDWPo/AcLTDbWhYZJGuflKy1qdLc2pP8jj7jMXQ+bZU9IO0utTfPgNslJWtS61js/Zu
+PJhgjoB73Gprgbc6eTzCVRtTVDhUP5/oUrjmjcHxrMDBxpbZP1YPoeGOWZG0/1Pl7d6eJLdJNPZ
lRSw6tXS8O6jAY4NwJK9Jc3k/uyMJjopoAFFbuQGtQfMPqER79Sox/WMQoBxuZKFgY3JFQB/DnnQ
+C/DHIegkgUDp0hAwO+CvLZZHDJGykzyjT1rPPQKTxolCMUiHpKx73MH9YbyQt97wRyqyzERct31
9Yv1wOpjJyed0uNlXrV0Y46kGwiUQVn+xtF0ISCz9XYpzveNNuw2/7aSnCkz1ZtWKh0O/CepmtiH
OJ1rJiLe5tVvIPgw2RwqGuEE6lBQDYQTimZHqND4YuZD+SNRFiPleRfYdMqkdE8WZh2l5PNLdcd2
G7GCeX1quJcn7g3nJcx8sY3xLyLH2Joe76mu382FgCqUf9R5AEV87zKNtDD+hBqqbH89xLOkFz/2
KvxDFb25TITNe+lZRm+x0NUfwGZolgcwkUyIrJimCDZ/xvI41s5TFhEmFKR+UtDRPzjw4sM25xzk
G5FAj/6SExL2SXZ5BY+PS0XuavD+inYFlS/EF/oHFyEuc13IhvHnytDwIT5pEURFXENwVpKc1Ni/
46eRIkYSiHwlZmF81BRwhA3X0M3ThKKPQTP9EKbydIseGsyV8Xfg4S7bdavaaYWhWsaZ3MkMxZHH
RgMTEs/a+22G8lZ/ciGogJZ7OHKU6KO5pG/95Rxr0XPxnyJXk1d9oNOufO5nTwOYXqyxPXWvTc2S
v0TuK0iaIue7J3ApXy3f2DUnvxC43q/3QpMzJFOooSenlDG8fyfwHW/a6y4n7uCb3X3bPyIXocr1
9vv1dP+eEAy8BYYRGTsfGuNMbsW5JTz8VTmPTo56tbZJnQo/Dl1csM0ogT1HRG0s6/Es6kx9og5K
UYjo8Mzj721T24QAaHMcgcU/ROBAv7rCZykFxWlYW+9krREUw2/cYrkonCXPlBj9cgDKqyRocwPm
KKdZaEhloy0m3wO8mbuOhUg7cr4yemfAlmUuKM+YPAO+lNjrYuogSFECVpTSgE6YEN745K2iMg23
gqLXYcubmULm1kRgvet2vK9zohltXySBitcemUf3dFyBHkA7asPdqPNwYTCmhSqdrrKVd5x9F5Hx
r/+n3TEuyjFHx/A5q112pRqMHVYJe6Ru+m2sBc8A+Ax5k2g5Dj6DP4WrwhJS71UUnWAU09J7FbUq
HzGJxqWAraNBNsuAKA6OIPJ3e9SyeFrKQyk0q31PAjcbsDgE0SsGh9vGq5N+0SX9GBbhZuZNpP2C
lEaIxUPCwYHimpsZRzNOj3ozfawU1shh4cYh7VfIhoMm2GzInClqXDNu0d6FVTXiDDWwMFLNIPIg
eHPWs0n/FOYkaN+zmiqoz93N50vXilPJo1hpeWswndXujv5RKqKWLA8cqEwYlJHwnIOppBiLlM71
eHeSMBKxriZCHK2OMLXaPusIvN7AsGw1Vn8Qh2lFK412+zH4tU6Muu/WGROjeTv0IAUwVjzlnfgG
0Pn7+7PwZckBDU+1sm4JxeO2aUJjkLj/YZHl9v4DMF8haejTgZVeJ3bON44re3WlBq4nOge+DJLF
jRMYh7aRE17x1JxaaQK8OyR8DzfHEam5QqgAsN/t8BIeaRIFuQ4DoKfIZ7EYLbayCJ+lCyi49tRu
jIYHwWR+6ZicMWT4HfWuMKa5tE591wFuwtymk/S3hwzeiUAkRL47zMS1yIh1r6hMdjZO+7Xb540M
xOgnDsfM5GSi3CQOZCzU4g99RA5/6KM44nZ00ty1D9xMmeGVRzKKjG0gbu8tGQY/vv6jNMs6q3aC
3MzTKt/s/bd22GHnYQ/FxXU3qCCdVMrFdEXbz9wGJQLI4eQxm8XDB4Opx5BFzA/+G0bnju28Ku07
T8+p/74z9G23WjSZz5U/8WFtyPqG4+wyO57Qw4dIf2Bj+tebUJLGy6ZE3UgwIIhnHi8V1xXGg2X+
sShknpKmw90pqVnHsdPh2wk0aI3BW0+p8Gcu2KPxspmlSQeFYNtf4oWMJKwE6W9h4+RrlEf7BtdV
RHGeUYXZNfS6KqjsEE5yUU3Nfn6pNmgIYGyUY+DVnnR1okvbgqoNAtdVy1vL9MZizOw1QgjZXOQ6
L/nQPkyS0HrfluAjwwhGAHBeEL1wjijW8ufSNQ6y5vc+xnrdP1t9V/NffPF49uhWjgOSP32SvIj+
9VJUxn8BXBKMoLXLIfzShTQZJZeQuQN+0v3XFrUlxMA3RbBHPmCbRhr+n5idN3rVvJRZkoOEwZ+B
QjeaDRniyuT13xRB3C3ylpMyJve1Z6nmVBgzMrL3bfUc/r60M0VPSehKB2ThUq4IHU1xgxezKX6W
+KzgOPKepTOajo2PblK7fAd2aCzTcv/p9Vwt7hZ/z4Fmqg9Pz/UoKnyacBxebHVdYblf0I4YKycE
5jvaeaJWk12xHFrbNRWhrgcAq8utoFOAoYI3QLwuZ0O9PDCbAvmkzTlobcvaIlcEvX6Yse/6pS4r
45ikSTTD3yJyTyHE8DlctIkdxBJlGp2QdzaEnX0y11emIohY9z+YZYZ8gCwzJgPfvIZYuy0MqvBl
w7c3uo8r9iT5E245wuR9r94BUwdwDgRRKmVi2GLzIGY/dEiL0RqVcGzEtNoyg0APmjt00kjLNYDB
6kHrTInlPmGVYey+yY1q9BZEsV83pqpGeTAtNqADpJl9dm8Hz/2D9JscDxcRKcoZzhgThk8/icFk
9BcIidMpMzfkKQaqUEOj6sEnWhkn20TbDcrjj5DlPwf8i4yKXy/y1NFOnspT0T1xVaSaUV7YQ+FL
9rh+BDdQdSkqXfOsOasN85xPP4DeOYzyTV/BV9qqi2GAzGiHfe0Ax2I3EI8f0Mtdms6pET+2A34r
QkTw4VA6iE3fveajP7lFMwyTqjbrIYRa60QgpMra9KO495WtNSsvo+JEXYg5MtATLo6ELe52kLn2
J13b+E2oMAeezzg7BDfLBprQ0FF9hrWpA3UweLukufWXc/sngnCJxtIX9OiVIFr8A9e0amPwgoid
CZHCZ2oEugt53UgTT/c+gnl744UA9fM6Lo93TfyUGlVrvB2DXqpVqsXRdkVEqrCh2HV2vlX+pQuc
NJW+jZSeIjPkjK+vzi5b3cGOYywKRnxPdWrJIdNOFog80+SZwdnRCFS3u7t/qdDKVYejzoCP6lDc
JxBuIg4GmTnrSn3ByM//Us2Bh/Gm2331CkzAjHchEKwSS1HGaPdZLG9lzXKHkvSzgXWC+diC+n/q
9PH8AM9e3JuYcV5RQSS2x27fJRd8Glz6gHU0wXXBeALEqhnESO3TIf6sOpfxC/P5vSvvsKk7OfBk
uPYq8Lt7OHqyL7V1k0pZRfy3jAUQFV/j2UAs9k9uLOS0+jhjFZJibe3BNGclFqSJp6U0Sh9CqdWk
x4Mr2ZU9H7NwzFUxuEC3Vac5XDVWPihwWRiW6EEizpEQDcQZzNz1+vSV/bC/6uVOudSJnK/hVvGt
A+N1Vt720RJQ9LiRHI0sc7/5Ijw6zNVhoGBAiaiSvD+fo0LYKGOkjzapjT+5OEqJBtRrPcxuxNYi
HGzftssdzwq2RGTWs+Ddc8QQtFrA67owHm7PICUz8DRjffnC/8lVQV7a3m2TJyb+p1o3hMMlU53b
Pk/5sP0JL4VTUFozu3zcnsiZUy7wpned/19aOkM6VGSQb6KrGp77L0kflkDe5vLbaBA+P9Vruqm9
H/SIa5gAnehBRpRbFThSJ4czmFhYCtN0PvxfaGukHg6Iik/SkMgUdcYibUsjFlxXKZlvg+UuPApu
H46qT7xHnP9Z43an39tYL/Ts55PKAhtAlXx/k33xGkxsMMr0gHo2M85gHtbaP023tgfKwa/1N2QV
B98jk0ybQ2hyFaBdMFZQF4If1s85GRh8mx2yuXftTgCXCiP2uulkh18MH711geUGZMoG0ey+c4KC
W+BUZ/mcMVcpHoNdPE+KiZbY1s3Xt2NW/YTBtT7oj0KM71WAko7k1jnokQi3OW31dbC+TkX3+QN1
2wY/wjyWSSN4vL6PnPoyyVoqSmoE936tO5OvdpaADnGjgyknC4hqt2s1LfM+tbk9Zgk+Gqc4yUpx
P5r3nd2W76jOgV4UkhRUV+TdImnlMHyrU0dP7Xe9qTJ3nPsoXmHW31JadvffVtmLviX57cxpruc5
0sWKAZjgFxFjHIs9XIwwjVfXXsOKGizARi1GZS1HcLuskDioHx9u0X38Lr2U2XQ0S8uwUx/gAlqw
QkrQBGmAra9bOfKYHMxlUXwiAUeBixXT0Qfn+7xvlp+1bwaRgzuQr38R92KuiD8vdAiB3pJqz4v8
z9CaHcQIx8JwNnhGVXPLfpoOxiM1T05rAyU9AAmUi92MV58NCKNYW3iuOg0WOfrNxn032aKg15W0
bj8Y1Aaclr7gZTEwaYsCxfRbexMe0QUalU/YuD021tAvfGj8YrzHUGOY2f3yuOScBUckcBvPP5Dl
3oBislduPMRay0RcAxRcWDMuFL0CVK25m7VuIGLmcM8EamTO/aKBL3RoguCSONjrzJhGto6mdO2h
nd38D3f9qy1x7866ggM7DcG2sKYsN1TirVbWXdDOUn61pbiIHMg/J7ieg2EqryxHn1DkFvicmGfb
ZRyJoWv9OntNPIldFXjsKCDWM7cPqUntGVQAaZ7RUR8svW5GuW8KISiu1rrXMFjj9V66O/nP6IHI
E2MKWKRsJb/ROTauy09/Dtv6yDRuzVQYJyUhasGzAvWN56TVBIgZTFVZCbqqIORCdfd1sb5IJQN1
02x5j8JT8LQhJ81GUM1nDVZt2nYNGBUBVEhddpgNYztirxyAAiSqu0xhMRHM+HXhwDwsoOMGouI4
ko3CNgV+0efsVqTcJTlI6F5fzR87SuDb7qq7+XY5mS8QD3hn7qMVLsJXmJmZ08nNfpi2hyGznPvT
vI2qWGqwybgCzCxQg+peU5TQ9V41z26XzJ4Q33CKfHeO/9NXjawHxmcDf4ls2sWJOH601rTah59X
CjordbIYFgOVKR1vEmRUAoIc5Gp0u0x3VMTdyzeaxk73gc7I4ktj3/3Z20eoRcHdG1c0qO/lqSHJ
sxDESr9s5e9ESJKDm7D3Zt1ttx4/6zHMW6OPzFe5nxQis+z0V6NVB+g0ZP0DnWXve2sjimQQpfVo
m0c5OJqB6pd9zdnGwSux+jmMbvCXd1qoBlKcKLZAQNWU/Pj2mnTR924l8gefdsOP20+lM+ZDpGjQ
WXyQ1OI6dur1hhpo1H3obAazyhKCr6p3kFtnSD1GvEMsGdHTgtKFEBDJw24gOqsL9ECBHvzgx1Hh
FtP+jAgToSD9Gofsqo40sgB/V0SK3GlqHwMPSLmHUDwN1y7K8fwmjQ1gcY89r6QeZ/XfR+amboH+
ILyKkfguZU6oUEqORTLuq+Puxq1V4SpWmvGmFnvoXzI7yraksd45xELqDTZoYtYGZuF0MS90sSKU
vtGiLsNxScxCkrAmK2Xph76YUyEYrOwsHHNmCSqvx/TxUMWnpGSp61k7pEVBSoGsDUjJOdSvszFA
xHjAKjF1mb22JNzBYyVd3b/kvX7MLDQ21OqYKCIs7ukoAwQrEW1JElC3gkee6j31Yg9uq5G9zAjj
zfaNvgDwrHZXa91Y7EQvaCJqdqnmLukvOYRuSTgjb6eOhyDkpv1Ers5wWBsEiesTW6vCs/4d/ElT
ujMlJbMCwuAHVfQshWXSNR1uwdw0OWXwIP/ybl1ZXQ6dInSDlHNywCM1VjuPWJcZret+LGxOLyDS
zMA7A/jhEKVkfq5PzVNJ/k6NrgUUzuohP0z7R4wNg5jIbH9kLyIto0fN7ThXJVRgqOmYcNEV7bA3
sfbEfa71ihO0498Y1vWGWf1Sa63ZZMd30ABUTufuP8vpxkfa6YM/zwiJZ+3PFU9hEGu3B1jamZcO
U9fCenJmLSIPDHcjm/q5p5zqEdgQnuA7EoqD6z02mZ8EqZg90h1y+ch4cdqhObrzDfC31OsQ3r01
r1Prmbk4aVYmX+BP+LES5P1EykD4lVr88p0UlkBmIwuUlxCkANBFVtoWA0LUv9vZwqwz50NeW7Hw
P9gxLx6UzA7/rxoqSIV1Ngsyxqm+5T/YPOomUtCzuJI9G0QMUAj51+1JaUZ3BjIkCN6XcoS5nsCs
Jdw5xfUfzfRgbUKvOafO4oz0eaosppmS81DDy3ovhX0FBxpJgK8eOnrdUbFl4MjA+73DaDPNQBbS
mzJ4zEl7lonZJgA/HIL3eUfSK+ZORuYKkgPkhZ8H606XF7Bcy7Igit+yavzrgqqRkX08x6zAh0BF
LLk7u7aNk8DIOC8zccLVqEpEmZ3QGdLlgMixMuNlKLgi09x1WI9QfIU8tBoxLZUst/OzHAK6wxqF
0Lz2vSGJIlvR2cm9cEAZBU72jFJr5ddcLAeO/H203zZUL86yg/RdE4yBkXloGxe+O9XhUo2WBZFy
LvDX+wMu+GJAs0SvTUfTvdnCZr9uvM1EYMQp7MGhTXkKlsF3gibCXIFNdNEvHclpnooQ1QpSYmp0
YoHdAq+n8Eoeeg0T44w5DWwPPDuSwLRf4aOxpGh1wVCia+Z2ycx1HOkDUxjD/Qy9AENh2Pj7PlV4
L7kppuIb8aQaBDTgbSwyADNHYKz7TQv/5rUpCuWPArrVm4YQ+M74IEyH7/cOKa+6Bbjn7PSty0H7
IxJ5BdsXXH8tzC8aZRr/c/pe4IU4ZcZCpEBBUGRrPYzpyqZ887E79aqThtgVMU5+ZvLlOMfkpHmp
Ad4ucIjsV04q7Euy3QC9myHl5weJeG7peiDBepO1VHAsxXNZOf5JfOHiewdae6FlBeISf6EUr1hn
h6q/y1OoEaeEisWnA+RotCBSMBAf5jOgOtGCEs6xnWM7Tc2/p7Eq4r+FhbDwfO5gYvBKDCstL3il
Vf0sVNG5aqfxiD73qyT2fuApyMLpLqfhlOruFraPXL79Weia/MMBZjUDT740hJDckgzWK/NAixM+
MFai3TW1TXjKkVKB7nxXmk/VSgOBm9KqLANXAxk4HSGO5MzEhYQqdKanbPUCLQ/LGyRFd4p71w/s
bkXCLdGD8o+Z6eykSeZoSimSB7B/Dc9T3LoRUWkxurEbzo1IqUi/Wpho0gqfdPyQ7MN/T8nL9oBI
vlkYYbX48z/CGXBwqPD0tuUf7vjhGrFugr9vdOSeSXj7yRrjLliWHza7VS8mmPm/c7eUOryAZgjK
YN8ahQ9C4qfgyzxHDL9MWFOpXiAeCj3YUelHA8A3tWWv/6pubnwrXoLuuNerj5cNuXvr3t/ZBW9U
DAvwdVG+OXGzXwcy4RCjtALdbL4zO4ZKED2BARrBvqWCho70vicMFpXJ9EZcvdLYV4vUEPBL3Udq
QOxcTQwGer0uwUnGG6U9c3G2KkgwyqFT7UmlcgLsgvGBh9ITOYz4tWCljw7ZTolj5bkPOFuFxagO
rSuVlxTNg5Dk4HnW41KBQWwmbgT//+ISEJQmF4vCTe7Is2R7HKGPzF2E2n0wPoJ6f9dYEajBNMNp
NFYWYKH0GwNChbE3gVzrEL7acoAznQxAilv+Zo7dTLT9lWwcUxhacGutt1vPCV2Junf4Du2yD8Yp
ooFiOAXHm1LNCkmflXIui+D985AkfH8nr6KOPWTTKObun5jFJBWpxH5sFb10zVlHalBukkk1AvPm
Xp8396DI4VNQh32v+89XJ4Dqygh1xI23wgsJ3ndJ/OOfSXuH6SlRoODuRqRN0PhJVYzb4nUq0JjH
YxB0rjjh3HPsdgYwmFWSHyR/hk6yGIASR5zIcAHM8wMC0f7g578NbYgMuhDPd0q4iGJ9USGLWlf1
3spEamowpv4ZLjjo5tqtsABEPHrP4jXBsOFEkgfrt8sueLw7gD87FgQ3wX5pQJocGPI+lxRdzPfs
xG2aE4RzoOqilTK9xVPv1INxz/INDduszu7OnBQJ3lmWYoLSKI/fbJi50GvqwrsgVcdXg6C+DCB7
2/zZN2Wfls0GZQTKgzZ/698oDegvrLD6olxLQhizBFXw3HYrvijs+2kL4yn4XFB+7F/USnF/aBUw
RvvfQtmh1mfqWJNjz16qKf9hBxOOplX+1oCLsb6ogwEEvmEvFaUTwNhmiTzOn2Lmw4G3Q7InroPg
mUt/9eYQlSi5uZNdIy9qLAxD321tifdscZEDbICSKu27SnurfvfxpG7OYR0Y4Tubl4iwsd2CEFCN
cJlPop0hlTnP9pdk6ppkxRgjAw2cplpPAElbGgJTTPpIAHwFOyMos1mVyYO/zICcIO2cmv4lC+25
+s/yadypxEwlyMOVwmLW7FzSbZ4kgEqfyJwGk0KhGV0rHUa6YA2YBM0OIsf173nGU5Eb4tjDlpPJ
PBwdvNRfU8/FF7fppgsjiGPsCSmVGwg7WVtaMHsPFpImzS8KLLaamZtpqzcNlDWBooW04plYjHu4
qjFnOeEmqS6rJUr4achxD6dayW0WEjrGv9WliyD6HSpIoKw3OC4SZ2aNUbwstW5BS3Oi0nH3GnoX
NIzogRWC49PQ4vwRF1eHG9YbXKaRdfN1OGuBZubZl33uozueaIBY2s7z6DIFLTllaClmj7XgTh1H
1oM5LLybrUYckajXc+bVm7i7kcQ9uP8y2WzOWO3SzgcGlptxfrgnv+Da17vg252cTEtEjg+XYfZh
DPJAVfGjoQjjES1bbvklSnhiu/2NUe5i9W+Mfs1B2X1MUCbjoXPYajPQI8lBH+QhyAF7+wta3kSa
dOrlAsZkhDnFMF79g/vyrzxZlTgBglubCQWYly7s38MYRODDnehOD+4MbKG6uAPM7+KZ3nUJERl8
N8khiKdTOY6E33/Eol5PRFXqyB9Q9btgsof/msTlTsRIgtHwqZ1xDkQHVwE22rfzzkUraklhLf3a
vTRg5x/jt7x0oE3NLODT9vIElcuSlMhV13FFoZUirHCwyCTwtuutThEWz5ydsgtbshQXSJ2Z6RFZ
xc5KelO0CQOGmgcGyfqnp/RFBf50Za2PqcNMbXvMddiGS12Q2qtS0opIRXFfvHSZXuxRAAI4aYRs
72QxXIC+vSQrKOpfTpkeirV5iqgnKLaOO2xgyvuB3Q6OtFQltD9ELVF9XgaURuSdrSqkefGK/6LX
GVzd22G6Eo5zBMKVH9zemUTLKXeFHkFmh7hF5lWG4YRq//I/Ecz3scTEKUrRa7/SU3ohkXXS5Cz5
3zXek38YAJKiHT3HRs6ilGTAPYx5qDGfBbY16WdBzAsPrms10SIjVa6De+l1LPVA5zjgxCTosey7
AUhCXfrlQozQZudK9HOqZsTcRSPo67CXrwBVT/rZVKlTJwDoqADxLmlkuzS7Yib0ojaYF5nBJbf3
4Pfa93+6phlntjDdrLOq9hWaBooUTkJVBkRRpgiBXvTgoec3fdkYf1BLsWOpGEUg03Rc21by0GDD
w+NC8PJ+jh+8jersIqIJxriQqD1rEuV1l5y8gPfvAllXz15X+JE8llqrV3oLRD39pddbr2+3oTDh
Vzzn6CNJvzAE0XaW7dMeuWLQnUra9qrVRWz1IqtWAQU/CPzlGkWoNpDrrIuuTii0z8oH7Rq5sXE+
/IHuTi5Qmzskws5ZHI91aPGEiV3MkoIs2Xj2/v/4GBaV1/V58qbpl65xkWf7XMtrdUW2arc9Od4d
RWiY/PwNYOU/CeG352fQj6XsS3oEBk6bymFvEk5heyLE1zi2pJKY4h7lyJ1dS1O7XRJ6mAG8jO9v
g/cOlXdAr5Oe8Vkf5Oe/y9fZ6yo+4GroYSTzt6OXvqMXjwOfEyR3tYu1ccuAtGLVN+Ltxhj0Aziy
I2PH/ikBT4CQsPjXlR2wkspGZN63X1oAf/D7ATehkETp0XTJjZ58RYhI9dnFJ1SfBq1kH6Px/1Dl
k7skCSgDHpbDOSX8A2svUVeNW5AqDzbE6Y6NUOo8mUQcgNuVtnOHRie4JSPv4birXLDAE8hoxxrP
mQiHkDNP0iiuFjTzO1Y7hTHhJiZYIJaY8+r4oJXrwzSWb/rxU0AKZ99HHFgx9E8zGeNajBXuICoM
A4H51v8liIGetjl16E8g41R5YEYaqwudvZCQq04d9QIphJ84vkRQsVeCBFTyBdH3VS9M7h/MCGex
UuM5oMAYqh0T+qSBjjELX06H9Wp5pJJL8yY48KkhUkrzjqaEg3jbHCiXunhfKbO43NkdAuiJZOpN
KY9yQ+iGV1SYUtTKdFKRbabeaRtkHZA05TUghRfkHR2lUGr5QjduNnBLq8tUq4DL48e+WBzk+OS+
FU9rHUI05vjiCGsn6/kn0r78a4e52HwIXdHucZNup5X0SZe3USofPlvLvrr8NS0kF8QpJRHWSpY6
s8DSdQGUk1pZPo0C9tktSnw+Ni9RjBgBsYQl/ReT/RF8RbMiPa9/RwVljvTo1lRGOO2P2diYp6uS
CWRT1FDi/nSinxRhxxQH2NYGnh/4MkEdZPIb9lqJozA+gdy9YF453S0f7D6y+yyvk0/M5F1PgIud
3SPF1REmGX8TO3OIQ9XMuTriXyBB5POMJ9gvqnEt0wFmb1HkJ2EqbP5dSm/aPk51AEq/W5W5r95w
H8WbZCFm2dudgPO/qDkVp/sqwl3R7bG6PulrddAXOSEAdEOUvTUJ3H6VKDEKZG6drxLnszdbnJu4
HlBKnhm63B1Mk63HW+v6AmsTwNvRxwdMLReQOLGI2jxHqTAQ2fFvM6OHcsaDjXDgINQAMKyN3qUK
eizDqOvkclls37ESbWhelNUHg+d7T9CpqxXAFMufqLi5IwpE2vz4KmkMUaqaomi6ZfUwOzn+JdLl
Wb4ZTwDMFMZFldlLe9SSdnLukdcKo60ry7q17F3czqeTauJbSToE81J3ODFdpA4SfV/uKN2hDBF2
PUVP0Pg9EjA6LgneUAaWqwQnyP0PBh0+QfEoj8fhMC3qFJ9IFqo8KMpyIR9/SQG7AwJ59VpTHjKz
vx/tyQUNUHakkVW+JBmnbXAJ/rmh/GfKPCpL8d4jvC7pvncWPZ/YQlSEhC4uWE9UcAqv4aMfoACa
6enP4xpmuXPgCTda94KNDoUoh6wX6qw5NBCwvJ2WUQMaWtgtArojv0tsQTScItNbcR1ORmweX76Z
AI6btCx2pZJ33NeW/UAmouWje5ugxKzrFsdH8XnmKOwzzzQh7kOGJ9GpV5yGD/c2sGiOHjeQpeeZ
G+cxL08QWlvhvwdV9IBXVL4pL4cr7BgD8ha+8LK/Is93sN8YuqWf3rnMq7v8VOgIVgD2DExqG1TD
KrsDqpluVEIO1OwGCPXnxvLJ5n91IL3Xa9cI6SVgJSyeGY9DmmIgatsAKvGIvEhkJ6o6jlTc3lqq
fHIwIXT83CBVxNiPMRODLnWI1eQ24iGabOy8jYyVTwZu858yJ83i1ETosxtFxUW35h9VoJmCJDUm
a35qnHinf3D/wjw9iDeIFaPoePnCGWMYbYSI0SuchWDuUlG9J/8vaoWJ67gtvTmFmcyu5Y51mEHi
da8lm3gd8ZFI2q/aAUCsh3y2wKeUiH/p8aru9AfK0XzBbOnQxObCsO5pY5pR/05oc+95H1H/h5Go
4Jvqo2Egjhc8MGxN6HqMPPR6BMTP7v3G+lgyh8Rky9tfZdss+AlHI8pfIu3Po5Z9HmZ/Gt5v7P+I
/aYgxAeoNUfdZe0QorjG/ROMSNWADri5Qe41mBSJzdKQWbL+OyaKyCtsU4A4aNH3vquA7+ekcxE+
iEW2DEUWJIuHf8rkEtXJQ/cA00io/TgvhkJ+fhTO+Q+SY4Ad4xwpUCcWg4dRp19jKAfMdjtRiC5r
MqzSxgnCxfwO+TQurzIyaIT+7nOkXyZd0FV+o9tMMav5jaah8R4LWIyOWAL0qWgd94TK20Nl4yYu
3Qb6UST3Vo0/jkavoVFtgyXroDxdZFw8UR9wJebCPj/YTZ5iGPgKNvi6rtf+kweYpFH3ELg4x4sN
9wcjwMaH7WgSxN1dbCqWnja2Hin7N8/CvCOITNkT4e9BY4QA0To14dj0g0W1Y2cRQBZxPhGMBHHC
S25eZNBn6vVBKeoLIprRmVCMnHb4oE6+oNprLSmSWBqtX+ab2WuCsusQt68DmIQ4dSQsjDLZ8Vgo
x5wbfvMKzTulmD3T4ncjK+NboPpgSehi95o23kC30oRh9noo5M4IcVLL8ciq5OOYh+NWWbmGNOHI
7KJOk6ihyym6Ki3LJgDJ0n2zXrr77WRh9ZiueQxcHo0M1z4xIXEtMg/BrWiGyrvQeq+yWB+AyfpG
JOUo5UlveBNBSVfQr+WpRbgdzFkJP0twAVhKGpWuCF5Z32E3j4Hc4XiAOquqXpjW2YQwKC927q5Z
ZBnDFC4iMYZv5iwjHuH+i5xNOxZyNnHC5Lx+8KxHPdfh/OSWhu4AB1ghlR/e9okqLRHQEU7mGm7D
Bjq5RlS4KQNB0FpEyynWJVNfI+WLLjwfxG0233RdTZKS3zaw0IAVCeUQ9yPet5NJeDluMkk2wO7d
beUHZMsRqmvQkf35wKeFLNo5IONssvgTUVeGj7zFpaQIQwDYRI0MIKpbSz9WdL5Mm91fuVwH2Q2J
edxiudA7UOm57k37QWm4nIIy0ZHq8BWj4/RR0jRio+jset8yi1Rn3/AjBiiEdzfi8rsXWpgkrdza
r62zISkCnw4KbfoHY/EbE6A0uHInOcc17mhGhgrM1ymYGaO0qDsiUJh/u6jggM1XCgmwnx+rsuSj
6zzJzV2PGqsKHiFoeCv4+LYevOGZN4PZV/w4CGL/AcMuzpdCakSreGS6XwxUo9fIpYOBXe2nu8Iy
fsMAcyuTjjTMS+OcvfJAQ7zRX2KnltNdIeT/60IE0jt2C1xLQLOIDXe/Cx6u9u6bTaIbgzx+wU6y
B1PdeaIn+UALsbz9bQ/5saeV6ktPckDLQy3PeMcRNayMTT4JEocLRVkTAcMGqSNuIs9LAvIdrUsY
fCh9CEKN3Qr0YyCkoKoQ6Q9y7TxfmWdbpQeaSNPycWc8ih96JsIj1nb679y0xEOcUnx3Tj/RNpHW
Dq+6xDaI4RBEVRmnsoMWSgPrariMlyP0C5KRcVN+DRiY5H7d7rSlFqMR5vSfbwKmAlhdKIOfLIA7
cY14iwPqquxrpqvLI2yPNjme+wF3ECM7LpnWJ91bNPkK8eVY0NsNr0WYQdQtunT8jWSGlnCStTfl
wkGVG9o2FBuGzfwNAvvZQ0hNmZzp2rgENwvCvDvFNFc+Qggh4sFZdC9quc0itESqoEJ+zcCdxt4k
93WY+p0D9EYChFqHkcCVehVa0ZifVDIXTSM888Cw64UmXtkmci1EyA89B8V1b53Qy3+A1GLz2LzI
kQGmlU2eU3QPwo6J+b18/BmGW0hCZNGL94p7LzCTv849cIeWSQDnVOOtmLPDrlieRyCyKCFgG2dt
kGJXIuR9q0EHXpDGJz6HyUoYjVBrOXizFV6Q98n/4a0YOKN4V+vqEpAycP/pvyEsphrK0LByZtGf
fXO/hVeDnIGQPFFf2eeELQH1COnWZG/JiGzOU8ttoFcqGI9YMw0rSe9h4l4baZeVd7kbchyD/kZE
6BF1MbKCuKrKSZY6Tx4eNxwBKmm3enqtNKxsliRyX2RK4z/hZ5NEJTvRAai4/L8yr0WOd0Ca/6Qq
mxri8xbSDYRLwhoOyKwe3f2DodHu13ylYZIY3o5unoYjWHkOAqIdgCY01y7kGYjHx7DLZxARbPNe
cHId7ww2jmnhzmwxNllG8TTcDVPVzbREc0/5Gq1yYyBg9MlRrC1xKvmz6KNBAOEIqPK8ct+zMpVF
ADxtZZ1mZY4Yuc8zzAr+rgGR6R1Ei1lln9o61YTrCWI6g9w0nwmOfsP+sd/QZJrCnHqkuKNEGBSj
Ny1hB4LTKUmdiGnY6AQqAm5zC15+qqhNjXczH3Eqk6Av/gJhVqv8SqyhiBifNa+vrKvz1VsD4JeL
4tDIHDAWGm1DGnFQrBRiOPLpc0XFU3MR3wUMKZcyGa7DfGa7I/RrLgVSFyYy2zCbJXPN9Lda/l1L
c+AHr9eMisBBcNVrNM15eUhyEFRVUwXZXdgTYCg71ynuZqIVk3P/LwSnHClOW0DLriuySEg0FYZJ
9k5aaBBbb4yHDOs4x59Ij+fhb/csshaYQy8cUW6/sYS7WNAXK7CMLWm7e31odWkrxvdAANPfP9Cj
78nhydK8OeYfCki/PgnKt4FPbK24VdxcXtkNywmun5YnVwLWmF1pKsYPwmOycHInWRAP0MkkX6w+
0pNJxjzQ7duz8m31Hbzo+yuCNOF2lYDLK5eN0E7Ey1lNj/qzChtKWPbLHIWm+jaz0a9zqQMWr2xD
4bhbK8g6ALCk9YcWBwdrJS6kJDOERimD+RACWG6GtMdMZpTYqEwHqnYcWiGeuwf4PYz17/JA5a8G
94/GwhA/03uufAW1mqzml6lWXc6OXH5nsd/7EX84mvM8MrwW78CcasBK7bM9nc0ELeQqu4cgMW32
uyAKJlc4HvFDN9jw6oRPty7ThWHlihPAiEKpXImUy1V3QK18+GfMx9boHoowzsPPRiryfnPyuVu7
gA8q4G/R0pN9XvQbeo9MIEMQ77CKgAfPvHUYPdjxSxUuSCKFcuvJV/5Wuqmi6ktFC9MYB1QWbiuK
YbJkb/ca1Ia6fV8EBrQCkkXDrgH3oOD2R8mW5niI8DqUb4qMY+VFhWR/opz9ohzRtAxLfR+zPUgX
dTo1+Y1RU8a0YT1Amm+n0P23vWE73YHHyRXxY7dToDq3lad5ZrZa4zsBCsZxi5KW0xOP0fRYz8Ph
h/ZiwWjDWiPILBG7Eijb5aoDkf8WZKvM7QGQ0VDWLDOdQ92uwQLzhxcfucRXjiHZvHUOLsigKcDq
R1FxJft/VJfLRRnlvKQnqoCL1MCiFdD2kUEb/xT/KmFiaUC/v2QYnZ10hcwaajbNdfpFXxjyAUew
LWJ2XjwpJz29uNIOvfVZXYeIHJXwBcIEqiRcvydvz9m++ha9pRSUg/xG1G0eJL8xlAd6qGARs6il
5v43loAGG0pdn759q0bwq6M88JOqvS77NQDrzZx8wXtSw3IJnPSoarqBrD95DrhLbA1fgPIQPoFv
UvQGLRugtqvIOhseyLqWlRd/xJsPdEvEznLN2U6twQY+9s1YOb3qoQPAk3fXSSMQmhDR1CaJ/Q6N
2GjMbGGpBo2k0NWtEZYWQ9UD/7wKcwMrEx4inoSRfW+qgquiEmDA8coHVI3RQSf/1N0fCganRnJI
pCMbDpSmwWR6f/a5eNI6xsAGHjWB4KpFpvHcU5HlvvgCWpXWKZ4BPNU7blSM05dZ82ZWwrBSokPQ
HjIdy6UvtrV7Q1W2xWrWHI2U/uE3tBIFAg5BLYLYJZvv2HXN61TUvERR/yvLH7TT+C9r4YeZlKJ/
YOGbfbqyTPqbSlSiVhQVEV/apjWZ+lQuOmcAt9irxJLxcs/Zk1QrYDtdPd+AlNJJ4AU9pc1VxL/W
YM97Yfr2usj2rx6q1q5ErY/kzIjqlp3VPSyAEyiDajZFzEXHYIyCiYD/5+X8i0wWATHivhgcuVzc
wuh/homvQzc3jAsWn8Su2SZvE8o5MzbidWVmkqskH3fngq9dUfisHuKmOueWrAXjMeP2nrYYdFhg
C0dtm6NelytKmaQi6PiTygIvCo7MGj49/Q5upvbw0NVqv3g6CPq11TcyzBtFyIlqA+u+Nix7le23
EPqkkOAFrc+lheiHHFGJGpQvHdKgGb+WRnnLsemoYvJk4WOqnxEHpp02jRUUmngBVLtA1pUAoM2c
Tkm5BwAGdkLaRc+3t+cYmFyJAM9PSQ2+1I9pgXTqREnySTnFraZnYlRx7Us4zXZLzuukb7C8w1gl
MC280lMNWyP7W6X2K2YfSDSQ3IeVZ+/AOzLF5K0Uq67pEdZUbZznmmjiTQ67nK019tnjPgZ+UcEP
5/rKT59agTjgGbxRNWwoXiYSd3TTdnwUG3Duzkz0TUD+hMaCrWJYTeGGTMeLQXmx3qS2LlN5vsMN
6ai7qQeitONisqZp3XnWjTmsvKladLW8eobuVmQQ4xRIQ2RqStTzxSfKNkAp6bfk/aCOclpI7BRZ
t5DNd7c0FsxAcK00en9m8HqxrN79WX1ZD8nJjoEB6MC948KFNS6L9Fpu7wTbDjaB8kDXF/DtflvZ
Ne25+A2NSrZUHSgUbh9wPLQNctMO6ki2llNYzSyVYE10LpQbqD2YAXKdiPl00JaZbvkyMKOYvdnq
8LmmnF94SB5I5k7okUZdaFfy6FWeyucL+sZubChZ65IoZg3NwCkhiBu3xQ202I6roJm4ifavW+h7
OqP4P/pMCc3hMlmQVhOnsPTj0Y+sofZG11m5+AuitiBjORwhr0gqg0NOJGpq48P4nO7rthbqDYAA
c/6jvWIhQB4r20Ll+cqqY/efNRNbPq5nGoDZnpKg8wy+ZIPFSQQG1XHs/NmIaauVUsRJA4EZ8V1T
wV7bi8/MeFh4Gm3eyr39kjhmdRYTZi1C6m2QXlpclSeKVNW4fd4oJjhteWqtxHHPiROQzAVspkTl
LZ08KwIt32wncQhgNrXgc5d+gcZ7Oyi8ApLo7MQqnV3BFvZ70SA5+AdgWY1mP+k7U40PJNESr4Mr
gqTIBao/lD7VCiI1cDh+SmK8Tlm38cmePefr4+80yZH51U1jdO0Hsu/z0SQmG0m9qSIUA9os7+7g
r+R8VC7uzpXHZo/Nva9w8FWWnRuc2LccYC/gQQk+zLSgHZEur5b49oYlAMZelHJtgdl6sWlUZgvO
tOQGecSdH/dSTAEqTn76Nyy6NHvStXEvrU9rYYqC4kBLBJ3NVvOSuQkMz9lVCgW/uAXUamSYh3ba
SuTl9XrKHIOg+dRxiyqbo1yo4QuSkgqnDQ6GdFclNuhqsr280ENZRqIPJKi6+sv8stW+roqKjudK
0IF3dvILvJtryuBDpB0LxP2GbkAuMvQ+TNNH059KNW7RlDjG7gubKrZnmUgls/Uwe9L2Fp8tAUR1
CgjTmNH8dxSvq8MF1qTiLMLnbZQ/geWl16YYJfD8REcqAowCRQD4AayyAxja9Gk/ocofsh8Fobx4
mokSlM1lszkJLmjR3o0t1BRdQtZNEWwsCnQ2nxf+1Fo2UkH/fNaT8SI3sfKGS2fuNnUh4p/3emQn
3gjo0Ms4PbSYDGlKK2VEO4hdu6VYPxn57/+CvghTzBnJv3HjAa20bHlZOQ0TJQlVPav36/IVFjLy
n5yG2TEbKVKLAvz3tvHYsg0/o1xMj8rla0S8uDhlXE+vj70Hiv21zZYPqlXz1h76oP6zslumoNzo
LFfSF3Z/3njKIkQesGdqFh9JHwMZsty9vnQrVQYugUlAaJUjS97hyYYOrkbC8bwgZpKKfYkId2la
Wr4nlgOrDMeEeEvMLn4JXkY5JidWi5Q/+YMiFEl0LyVQAUFvcTcKsmZAwb9L2myxgPv1JQsMzCZi
vBZL6yz3LAox+S5WedNSYU2udElg6vGCXrocLgRQbhhKGWp4i/kRw4y7jhj5iLjFecpIJhy20iBb
j90HIYDio/uv1k0Agre4TxYtHQRF5OLA7+vUH4JajKpl8/UYgTujimTV1H0S8G55idUj2GZwKNO7
7tONe1TGArnVKZbPgMUwDQbxaCTE5md7NLscxoCldsF6pO6Hw+/QxHD7EJt7vg7Yo4lLPK/nq5vC
kO5tzous6xoMvHGGmVmqIxyNIETUMLtAtJgylB7Da2tUC0s/6qYzZ99GKwHp84vmUfLgehs3+1uw
KRbM+pr4A82isD4p9zNJJDWE0I/6SrWj1PfpBSFyhg4w1Hq6OLne9ULHrXRRpFBrN497lOQTKkz+
tgBu8fyOWd6WVdlDGhGUVvQp03PAVutRJ8klGaktbVlay9uSWiM2LFNWHK9nN5YWMr+GpJueoHmU
u0pX1fX5z0Pt2yi0kS2Nx/RnnPaI3ytNA1ULHuzBtn+n58Fo46/FT7/sSr/fUTdnzukU+/x+6LCv
IxkpsO7NGopv8eu6sjmgWodhRgyOcAxfmYbMQLeyLNqhwdC+huGH7jgpNdUYvdRd6124gR6Y2TXF
KekGGs7RkLYi5TYl4LQpF02M8GhZQGgdw9QaSmFEeZKlkm/D2zyxp33PWN6PABIMHSi7Qba8oiC6
2qovNC2kR/9RBc+9xqTm8L7hOSAfXckodBDoVom1Zqqo9dO825t/+cE9+nZ//hHjVrDYfd4aht9t
ju2hgEErGClMT+lZvVvOoarzhY0Zi+VJvBFpRdVT4YxTpaJeYJ/ed5Ie/QFkFRAPD91ofiSP7BfS
inrdNPJD9EvMqg9JQBgkCLO+PIy3O9mWczxhyHFMf2E4iU65odQ4qe8v+eDFX3DgVabpH2HqeRC3
hFBceHTdzxEn+6zcQxBfn10xhU6YB7zjlEPlkys5cFWQUZtAv8eMQO5lmQ3hTk6gsS6dueM3SKlU
cJ3f7nAPdZDZ/Gn3sJN4+H8ncS3ZqpO8S+N8lb3RL4H2r2P+hgKdFbwYlz/7QW2MofDqdz3Mj9EU
eb/b3CE2lh772hoDcX12oJJhGrqYVSvhYKAjzSqamaLqo+mARPRkzbytb/C2eI8u4954qiD2EwI4
10nJ8q27oieecFe8/vDL2KhHtCJDzRxTiuYsrgCb7x8pxwL7btc84YiAcH/uzId2211KWNcLKthZ
pAMScEFiERXOtyejWEXmjh23Sw/djXxo0I8Z+Mig1d++Fs7z2VUeNqoUYznfrnmyKhnVjW8r2tnY
bew+eJjHcQv9yKc3z928xS7GOHQN97c2pLBjedXZOFu4l3+xf6t7rpAX9L6tV2N3fxYcyX0lD8HZ
H5yDX4ymEZb2304CXr4LlvoeE1D1NfHqRhJYX79f4h1n5LDtjLs9ynzXe3Vij3KatQZDkvTKOtrH
qYYnUwCMGBoqVOrePEfssK6UMhwkjD2BVUDccVe1edeYxs1TjLySsoiJIXkI+4fqNQoPwLl0sGYk
b2CIe9R/Mu2g05Mb+I5H9naghP8rXdguqV+gkWvEA83jU3E0wkjlzazglnjDE7oERwgNGRPrm5cS
2o6ks6GYx1PFgtMsQM73mcyal4qgz0DYpTyIZtQMpJP1X9JTq+GBRCTM0RVpaCR6Wvt7BNpOjWWq
kgzciOOBFdB94ZhUAfLbEA8CaotYWIvyfMO24SdcGVTX0mn0k7ZX9ZI0BxKfM8XACw2xFLta7Fsu
aK95scAUdTrwShpwxSYKYip2W2th/IFRpoqQ5TvM7cOcnsq2DCvzCwGA/8ClHVnAsDtNu/lPwtTe
qKwuxXp0M8peWW+CAitPVlT23Mlmn/bymxPoXsQSNmv1cHfoScVnlNViQeqLdujJkyQVLKkjIM2R
AVf9PFzvpO20OusV3/NH71LGcrhI0AJM6w7A8eJYBWdNgCZZvmMW9piwK8FYbTu0VBjvVdOJtvRl
MZdIKd/CMYaO3qmjnmRdlvJv/wCNoxw4T1nwzgJDeVvziQa1fEVjEAkT+mL3dEyB00PMhNwLUMzm
mftyc7ssRdFjgBvxUh+azg2wHTa2Tqg4xGyJkbxudgrS7pKHG+SNeUefSQaMZI0xtZMm+Wk7pp6Z
JQVr1QD89szMUrjooAuPOnm8HGnTeXkLBI7K6iMY0sWwY0HHleN074j0BvhO99KwkNhYoSZC14qr
V+IxVkZWf+qDchsGYTpoNeMfnDvGzdI65m//qeCK6ZZRlXbRmnTFDfOsoD3LI+Z1yfGs08rTndkx
iAj2TPsz5i6GQxhukVH9/jTBWLtpUYqMMOjlI0/1nWDiSRkTFRou5o6VPXAKWtmMlfLLNrFBusPb
FxnLl3vYmnwhvHKf839hB8HLKWZgC46OJaWGBRmWbifpFaj3z31HXfrgP7fWr0J4Gp6gzv5lfBEu
0CSbGf/Gzd49O5iySQ/LQZtbTKxZWjezWmorLZIUhPXJ8/FW2PddR/B3FCcp2Gdboyym9cOvYQQD
oWXKcOvhzpGZY3yK7QTHdhG24dkzcGiFbU5hhrPiwIDy4x8zOOk9u/BG0lEh09VjoO9jy2WB7Fpj
MQ6IPnIEhtAhOu797LXbCUCTwsLyx89Xedh2BhVlHoja2nNwWEojIr5EXjSJXyrqTxvkFZyt5lTD
7Y2pwz8d+7IcQIdWfWQnA9K4bshJzt5dw71hfPU4JF1ZAc7oxpyv1fd79lJdPTvIRGPADxp4YkEK
BNCf3zMt1kVxjbUxs4IQ2pP57ioZq2TBJJhcz3+ByZtvHaMtFyVGyk9W3XqtzzBHoSBsHJSxYzcS
s2eNyFpAiUGVa9yx22Sw/PDiPgxZPVCAC2IUvYPhu7qt6UVcMFD1CFMtfDNPRwWi+9upon3PLfHF
249hdxdiQkyCqjdcmzE0QcVll7YKr6e0xnPG/qrg1U2BAFGKci5ifrUTSufKGWc2/azj3EhdurRF
F/0pwXqRFPGC5MFap8tweA8x8aBoZ6iaBuFzfzQuU6tXxpXRjFdHfYUiDvBDgSV2Dishx4oOQWxt
SR4tTlsDsKUUlsz9MF2vxTmCWTgp5d3mBDqhUHSF43xTD0ucT1ZRR2qduQG3JUVkgtCzWnwEn9dj
nnP8amaVsBOUWk2CFxjhSzBH8B5J0JJ3zDNag/dsAq5xPjwtm0rp17RNBoOi/GWxaVlvwUIYZRjA
Euyntk8vRbGBkMrECIJr/RF7duIu57C5Y0RWFdeKd1YEVyhULCKSxlp/MAJusGnkJbozSzmhvkMu
tY5yxTzrCTEn/L371u2Laja3bjZ6auku+a2PZ584le3wFVP/gRdsyzmU01vIV6lpEQ5HOgWD8sC6
p7NTkJWGUPejMCBQRI/MnnbPHrYeNTH+7PlLkXFVqtqxAaMTyHDGnM3Dzr7iNI0wZkkbixcEuu7m
mQP8rwTUIK0JIMBO0hC0pKWY8p18G7Mqit7zET0gW7UeNq2J28dosNxXRhWPmT/ovX6RKKReSWZQ
IV8Q7b4nkvDpG+Qwqncc+xqOhihSPn0LjIjUTuTxpwQs/iAoFn7EF9Vkac2caMpOevWfeaNT0C56
2VTnAkzs7MgMN7EHwHzYZlZMPQ9v1b3sETNTodkRoaCvHBCr7D1+zoT0KH+JfVKsNhjbiExLsqVb
AOqqWYHmmaNh+ljzo2ptQG8tvjH8pHPi9WfdTxmPEO6JH/Fr5kv4sCwUmgr+jPrrOlbq3Jk6M+F5
fv8OhLlyHPyvVZfKxVf5vHUfsEqRuVVT8KPgmYQBy5ZIYfTTTRlT70X82kw076v6281eW+6Hlsyx
HfLHe3R/cjmjhSWxiZDbqtmTPtjfUDpFjlfgCQTNqdnnsr7zJSy6AwoK5X5TAJgQIEBn+Aycma5X
cHJjMON6L7lrkPuntiJCcO9mmmT19c7nsCvznV84mfNh/eKxM6Nrla9irk22ZfJUi7nEphVPvz4+
dH3Anq3Lc/feAQ1ShUGIQ7ci9RUTysykwwsAgdaRY3eNhLSn4sm5+M4ytG0Eq8hZydeL7eZhWtEr
jeD4vCl6KsHoCdh1xoU6gCoKv5NoTDkFWpheuppqwAgcLo9Fg6EjcG4LHWznI2v7U6SLF/R9c/ha
0uFm1RhD+egKgKQeyC1ZIjJjegrJdYx02fuY9Ys/e+GaEG3z1rP1uDnrdM25g9MrAb6p7esrB6Pf
RkaR5appA/A2CM4J1+dzOw53WrjecHSacDGWcySdWoNl7OyLtZYoczH5CQxMJITP8NGufw5dwzFD
X2AMOQZjo/nypSIBCJJEwtZtIQZXL0ucJteoUx92F4hNtrjoaDMcK1kmqANO8ZBh2wKTZEyUlt8O
GaA6XSApOBA8oPG2XWAYuNNqHCu/KRrDuU7MwwwIuhjXpPdssYPwuPkYuk5kDJj7wTsA2HfJdR/b
pbYRQ9HTS8a6Oa+hSI/A4IecIa4ia6+hdrQcG7XMTzDCoeYLOWz2vv7GPgpEudCJp8KAM8AEvnFY
HwFpm8ty3Rs/Q/pi/76jo1irlheblIzzY7+pRea9Sjrhp51tCr7bPOIicywJf7FtjuK+KSFLi0qi
oYqrE+bS6cgaDFBmpGKC96eWTdU2f0Yd36vLkFbQxYe1lxMZv41jXWsmsW7z/yGSk25X24r3JAsC
ZyMuixbdovMD5mnKai8SWbbW6kXAVfw9aHaTu2bqJbzVvsgR+WuR7zdyDrsZclK1LAoeXCfpTeyu
VhZzuOFAJQEirmvWFug+9Yo81n31nIonupxQZEjUUpvl+wUXFJH21oA9kSz8tdpPoWqJvv+ibvTw
cI9vKKtEd1wjpJEw5azeYiOvoIBu+Ey6an4NXlGdyO9CRs32kU1t+hX4iYPN9USRyooxAjRy3k2c
87l/VqlKFUJd1fwhQYa7AxFJXtkroSoH+7oY/v7wWZo5ul457iH8bNHXBHSMGc+z6pw/Hfnh4E94
xRz+PPZDIJZkZnJuvSe4xpuaSszQ0nnQxdcm9kbsbATBnvS4P/BnwiDGDbzoKW/01/jbo11Y2EEC
R2hLDZP2f8PLXbZvNJ30vMKbnvxkEh5qFmdQxDzcgKHD6sluMwCPNfs8WzEd75wdA35MnnVHzkP+
ev5hzbV4ECoPZuae6L/jBXe6etyBV6hg54fkbGuCnA3i9Dhtj++SdheOsjYgMbRxTWWBgIECvjBp
fpvc40zIGIDMb51+8YN2DhgR7tZPanBm9jZjc5o+du4QvaypkAlutq3sPhK45tPRXSE639WmenXE
+cJ51regqsVq+vs7MPX4akCRyZ8xXw2EnNX3gaCdOY6HztbaSMYFp6aET+0a
`protect end_protected
