-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
EzyU6CLkfHo672NkRhSvat1/iACL18CrQ6w/hc2+vr8Kf5ouV8HJaN+svaKx8Tpq
mBvx3tQZouMHKtUtdc6pBG14Xln108zX/QZovOB5skdnTvf/ifNeKUnAke7fO1tb
VsHrALqtGOi4fa1dhToY2sOsHwXFsfVk+3KHg/le/T55MTI2bMEhUQ==
--pragma protect end_key_block
--pragma protect digest_block
GuBuQWaxOJxBsP0esO4S73fyJpw=
--pragma protect end_digest_block
--pragma protect data_block
Vf2IFuYQDRhlueHiZ/iBLlzChMI3JMIeRkVcrENiHm9bDIXzXR8uYojjRAbLUF5a
32l1GTmmUeY6FeaYXwsXiF4lbaVKdqKIrS0MvyULhuJq0NEy2dQDgUJgHXBQDxFt
VJhVhmaUAJRO88WYBRcklwj9CR+goj387+w4Reyg8PcX5HvJcXQfyeDshHC/dIpz
QxAuMo0sKF3xrN6kH9vSfn1ypk60O6Qt7R7dCd12yMjid1RpDIi6d1GPtpmW+R4e
HmnJy1g2vhGHZQI2SJtOsfOPTAWrUf8leHA6K0i3p/LnIxo7J/54uSWaJZD32C90
MBmaG6OHQqxHcTqJnRN9Azv49VJS5oUPbCY5+FLefDnQz5iHREcav31NwG2ppmTB
NC5zxVQH6qUK/EoYqWNuaSl2tdByy9gZWapcLrNy40qW38bwMVDMrYM3Uj/S9344
B1xCEoja4lqDDhzTs+HEDamR73ooShkw3ApNqmD4zcTKJlrTejvLspDEHvaHFXb0
Enf7iQSB4IXVsv9HMAUnm46fuQEnA1h+GRwqNhQDyVGz3+cXf17/d/2r3nMx59Em
yeVlFnMheLcrg4uBH9jjLbPW1RCfRORtNMSKAv1pLe6pjq2ExtW593HHwD1Cj923
ZIIAAOjRr8D8zlXSfGrC+2NteQF3kvWRv9pZnfX8bJC9tU4c0coWDI+t3lqpAsNf
UOUapbptaE6JFk7Jzs/6QyRWHkJF6AUBuhaECO8PKKDRHafY3OI3imlyA0fi2ldC
hRITBGREfbV0bbuAy/Y67jx5wL6ncs/iKATeYnXgUVAcdlsoQliVc+vNdCUm2KLs
FJQh59z8MXTQDzYjwkAivLOzK/juubZ3WsRm45lJ17nZGTm5NQNVYanRPibP8Y8w
tBcu0C50IiBg3eyBMdeodBnv049yFrDUScLjilZ3VVRssp2ze3HPelZUclheL08n
owjjqjxM8VNCmUzrSLWAfRzZV87higpuvcMuZwqf6oN0gcENfmQwqI9C2/4CfLaP
krygrAgy1WuEOCiAAcPItFotxyn/kIV9TzNKuvfe7wuoJJAqCC0rKhnIC7jgi8AI
YZ2tjfn3x2lUPvPfF2zonCd5Xqt5JhpKPT7Ikk1AQlm1n8HdXk+CeHpL9fQyY/Vn
fJAm8sFFUj8NKU/B8ZH78ijzNfu4kUqN2dJXo3PzeKwbouzXt7rdMzHoAGXwIpMG
FQQ8EyeAFCUa156ohiy4XyDrnhC+wRjp+48TJGOHX26aEVweEwNI0WFfxSVFFB8+
PGGYNdRRW+gLRzi6Xzd9zJ9eCkCbGE7QelhyT75A3V5RGtiQPf49wa+3cM6ywcFj
p3m4RVunip/zab1sQoyfn/vLPNFpVQ4U+QpC3X/GCglFhKqSnwwGX3b7OWb5utyj
sajNZwAbgdqXDhHTVVzUI/J2/IxtPsRkEglfBiOJ2L2xCBwZSf0x/99EaRTJYsVl
1jW8WgAjCbjTvcHwtmDgXHPbWETVqybYtUxd916C9ner7yfhI+rWQDbPyECuF2tj
lpb4QSQIdZxmhkVYHneTjBkFFpB9/yADOxMpjfFmxmyLGrDgO533Q6vpvskhZId+
WKS7ieNbNPMIh4Xh6mpknsakFpsWPQ2X97fkG+JFO1YdRjq0nfCfdR3Ucins8jUg
/7VhWkEmyQ5u+Kb9UTU7zPg1PUkBuXcXJDesLYEAGeHYJDu4owQ5F7dD9lxi/oxM
/zQSVE7YzODp+95j/eHmiZXipBU7psl24TPpCPQJjL8pTZan95vm9UcD+FpwQQMC
EFBP4hQftRWaJvx+88lNapIcAj2nbK7hJbbr9Xjre9RFSpH6XSZSVudc0XKAlbYt
IVKmU8HuDm2ec8wT4PvmiT3GJHMEkOXeVlencwGeL2EV/VlQ9cmRHqWtIR98rd39
60pvR7E1Te0rjEcqZ7b2AdtgNIJSgqRxZm3qP3LfJ1MFbUeuDoGnbjrY4zXExR4B
eI5PDnJEdtMd9d78I5XEd1NHzM35+WiQlHnQYZ6iu5MA4MmeuLeimGbkWWAeLTnt
IpbN3mPDrqlWTazS3jUprj+RTl5Z4B2OqZZ9m00MboNYmlS1n73FtO9tqvWI+66T
eQADqsLr4b2CZ1DBIg7bArXPLdFjm4Etl0pYCEu7n8t6I4PRxlZ/ByhnMaUkfsQb
tkFZA0Vub5TQedHcXiCUJZNTMMmjXU0wqffS7xIM1OLNSkuTMzgCJOGtuudVqiqW
CMsDFu+ga1bm6LDitkQ5G39PHVkY1DB0K2+yncEnE5gO0rFkY/RI1EhU8if3avA1
FJUMYRNSGLY6iNHPAPoaxjfWDPE8oFjPW/jHkC6dhwsJnRHWolkUXCqJ6/DblI6W
/BSTqj0NG6642GQM4xu9d5eN/korl9bJOjWgP/1jc/cX7+pbdsX+/mDfXcUT2VDM
xg8EcGDRHpDH8sXx3v3MIDcXEK0awEx6V+uMuBc6Wv+C30NaEQwIYjAMzw4lkQLi
I1f3hylhXcy1xtprR6NSD+fIDA98RuMpjuGKyi83Obpxef5R6qO0XPgIW1mh0z/V
laYXe6r4n5lPisBOFPj23b6KWx6Ln2PbIxOWozgjh2GZK4TDaX8U8XOcP5xhXTqm
VLOpXiqbxy/OrZPKkIUatPP3zy4fTnvAMnqyH56Ad2ZdKpe6XO4O2NAJgiy1r53Q
FSgpIkQLVJOTQLqzq8FHev1NYDlZZS6qlx3/cS2B24aD60s1Xm24OPuctLTI+1IZ
ZTn5ish6J817RX0kTGutw4b/Bj/MZjup2umtxtTHOqCdsw21OkPUopEVA/uiwUAX
8cUSoXGTpvcECs/vE9EmCGcLS+CwiJUREskuQLNqElJUqWHpJguputU03Z2/rMGO
MtxouiYVXMIhhSYm/yBnlG6IwK0FUyS9ibtBTX7Or7G90qAeJy9Xsukpk002XTDF
gOtkGEexVLAz1dy1EjTLSuKW0Vo/n/7cuyIVKN5fb3AP6qsJ/3gi86IlY8ZnERZ0
c88grwd0bYtlzjs8qEVUU2/NT1KR2slgvA6i7OpbDv9LdhfQEGAQc/UMk8d5IE1B
c7snbIATXygwSjyR6AOzx/o/CThsM5xhYcfqYDaYxp9tYY/5CjoqMD5RfLU+6DZM
lNe6OVfxkOGb+MSjEXYVEdbU6/HOWEPJgOgQAFBtarz9dHd/wfFDME+f/31b1Zo1
JkkWTmiwf1Y+xBFT8PzB4odx216jHdetES2+hmo5VqJrDYsZ0ovVqkazuaF4TuIE
qYukViPPAgr4awABI43lD2oEO3Sc0IBsQo73r5USHCsGwYzQDp7xPKqA5RtOWFHP
zScO7JeraJ/Px3R/cAmQW6hUbTckq1P+KDMz2Yob3y7xRh+OuqKgthUlfkx0Dd/R
UvPiA8cqeDWgEu77zlnPlJUVSoLIk8r5TTZmGqm1DQQeR54aekBn+xsEgAiCmvIS
dSWg9eu9nZEcpe/1UwvpmA7vjlDcHRUPmhmkwbfDy/0YCh1YRcFIm7mfwDo5/Bxv
QOmIiR4asdhg8+SGFFDnDAeCHCTMvLZKio6N7LOPVCiLF5G+3Ceg+USsoANomHzC
16crh/+16Cc+sCEIJEhZBJrfgn4e9qC5xekn6bNxy2Qkk8M1To1goAHykzPry552
3zcE//A6te/h6PUjR7MYY2pJ+wjvvgfoVlvsChcX6ZYe6H/B7lqmel4jt8c9fwj0
9kQzfZ3Fe18yLXv7hwfJoan4IEzSU63/PyzZwbKjcBUZsQB9xqLg883DcUUrhDId
QeZ58s6baZfg+4FxvZ3f9sWyplrZv0LNsPJFQiKuOsj/40a8MVLXH29zbVg5PyLG
0op/j49/rvNtatCwH7MAOzveVtXAbRgKq9/lobTRhEMB7NDPAqlRrbY67k4oFBcC
R3zQILdNMzTEbPT2p6K2D56Vf/a8gQaTshG2EeGxyPPRoLtndfrI4g63Q1pKzcHX
ctGdeW8rSfKyte/k+nsfian3gnZFk4ZZGE/PesZH3PXCU2NgqRJhDHmzUoSzDBwe
sjTUDuU4SSZ1084YTJD6ySw6scsTYQbWX3s1gHNmv5I9vDmWa/lMqEef9+1XLyKx
drOby8zqrt3JiBDsgvjf53x822dSKd5bI48EDzq9si5fBXUSBXXgGtld680Ttkr/
PMbOMPJab+DvJTynnwV9TtmHfFyvzTW4WvI9mXdNkPNBUMlDTITcH+37/VUX+QnQ
m0jL8nb3KVQ48dvG1Zfx4eMBMPAIkB8ODGob206/etAeDeM3efiaO9nn60femqcN
o8dVvk93S+s94FyhNgmfMelxpoM97ufzZmor1qUxPzZSpF/JVkkAszhQ2GkyDsGh
UcV2ChE53RuUhWq/azcLgxSry4qNW7LQwjeD7cAV6Tz4lTCG/EvWZz8nHj0HCSOr
acXylAwOs5cHMdhd34qi0pYL+qyKufVr0htRpcEFaptS3ypCx/3cs2f5LGUPzbQR
lZd/5JZn4hDYQXU4V49cvYluxVQpeXquv6aMmUCDvuNke3t2W44H/ORjjdoZJCuP
RWHIC1mcZJ7SGZlwOuhBBZO/NBNyBt+jwNMgOFXKKDfdLN/LoXQFae4v7maCfhKx
oGy1Ex4FO/endTvPvC+YObVeBJox6qKt0vdYG+eesXrGXyOdrpizpJnGLpFUi/H7
qdawSpu+G0QKlT+oQJ+BrjUGB2MJ5Y1XcAXkHISVrZTM1UqfBRM7VYcLFFFaS2YL
pMPJ1VBH9PpkkJ+i1N6TTdt0VvOZx3nZg8rcoyqKc9qwXiOFbKPzYKOl7TC2Lpqa
60+VhhfyeIToF1h3LKFSGtCe0H1TFCmMaVsxOltln4tgRgMuVxn1dNYi20QgbCqA
2wZdGhs1/8NrdVHw0a1vYsarx8K58QvDkmcvWSMeAkb1g9q12zU3zkin61usYHnW
/8mjcTs68+jDR0qgPEY3Kq4XH9Dz34GcslI/CC+216bfbA80dGOYyGqWuX96mWhf
aTzeaZNVem8VZaIqJzCStP5LxtdEglqE+i+scM4vaMSoRDPRBbfF6tUx7rY0N/VA
Lj2G/dmts2TnTxeK6jwawjQO/Cz0bY91em7tdPRBYO5FMAAU87bBP/dYti0hfU+t
v0zGXllHP5qid5jzjczkAJOX0ZX39Gai3giNfkFQoEWNRelrC+poiuwdHYCnSsKL
OxlglufB9s+sAuFOvd2bxsst0XuCfO6zFCys9tyxw2tsVPI4V236MhZ78oSDa+Uu
fJTClBYt8xxVlURs0qiqUaESsGJz5k7qA1rnkPv6NlKPIachWKGzXEX3IXF2d+6q
Y4ffJImnapL/xhW9vsW7gM71j7/0LrZd4n+eWP8vDSSPwGRmGp2qeOfDTBd+p3TY
DdlbXAx9lkxZGzTp5G55doFDjot8We59gFc6uhIEFEW3kRSP5AbqLbfa8qT4bpI+
bREgWAehi6t5/Mtf1IhqFS25kpvdtn64ztgzLT5OP761QJWOxe0DF2GDSpL0hGZx
w0rf8LLwq3C4peXo3axMLeLJ7cZJ7JLdIrRQ6qDWWqSK7OQ/+BbfOlV9CoaB0i2Y
aiCp8PDYu7sIMhk3VFtPGkdCa2iXsnsaSZPOV7AYbM6L+KqOQhMSJQ0yYxQFmd6f
hfObBpNxt2VGvIn+PfObtcdixCERKv0k7EzZ8DbK1cL5p2mpJ8aQBwCGHACg8CVw
6Gszh+K0z1cFoMv1b8Sm9CDvbh1lPVX223zeDk9svG4r32cv/Em343QCWQm+hD/m
fqJu9OUUYNDHfr9whC2u7k7sIOYMaA0x58gmxghC7GrZ+NQacarn/kflOekhnzMA
puYMfBdTMNZkz8tExNWz9wIi52fmJyRromU697CgK+B15dYzNMJI4NkiUKfx8jda
3fvG+la6+4quCfFXwPoVKaxTECZcnTsBrI+YFJQJQNJ8V+XOLSieUl+Z65WiKY4A
auOLEFVo52D1mWIjLqSwqEQ97geXyieFux1KKx9znUYazyj49WFQDCl8zzBDpXfg
V3e2qSKbm4e1htrjJ74Z10lztku5/3tppmqqEFfBMbSZogFkLfCf0tEREr/b4//j
LgOQ/IOHf8fMlw7qXGxI0YGWWgwMegGU5oi0eGZ/8VayWpet68qGFGXTPfrWns5v
JV0X+GbjFIkQDjRcoFn+8IuHc+IuuyRb/mLFqGuzxsqmljW5EQpo9vqch60mDa/x
s8wUqPnNpBafqIJetgqFMLI5wkEOcpvUXyyqSzwE1za852MDt2AYBHY65P3OSq+e
+GZ8KC5wQSEpxxCct35GATeQpKON6a1NGXzF17Kc57DeM/yrDicuXYTls/dCk3IG
48RtDA93yOCE9r8Zpp31li3GE7OuH/nYpP5yCLsOWDxRWBz5s8tf6YHTBEu2sn7r
mDqYEK/Pg6KZBZUrlRmgp4UA675fLiMH/wPfEIUiIUU4Z3mOcG/5EEgU2pioanB2
tAxddqkgmGB3DLIgXZW1KZ6KZsVT2E2zq44bz1eb8IXFbW85GVxdP9duxrL7xGro
QGAl0lgMr1DvF5TDTos8sBC+SEnQEse98J/gRLfvDXwPooOhaKmNngAgtPQ7b1Qg
QEgfRKMj9Raacnm+YAqIsprvPEG2Iszk65hOaWNNA6fqAyDbi41V5RxUgJMbc8mA
LPaSzsRTSyB+ncEb2B+JBVRUAcuIQoC9RgQ7tWZ2U1CkaTDq8rFG3Cr9VrImdXxt
akgIPf1MeerQLH+BDvguYFfNTVZFlE6VhRPrPxsevoz93B5DpBdnrun9nMGe4SML
VqEnP65T8gw42BHgsq/fd2wvkoNKL3bNeGwf/5ybf/STbbKtgZcSyT/0VD0PXIBa
AGTNzCI3vYNv3BbPD8Rs7bSdrhopwDFCTu0TKkVZyO4tKVB5HooMProL4PK1WqvQ
mRGarEsBH2LxCgQmcbaWAUVbfLkJIc/qkiPRRpjlPV/VRXCRKiQjVNXOjel0AGQs
ZVsE71v6w7fv8BWRBX+0Ul0R7YNSkU7CVoiyqZmNUkTo68otTRowN77g3oe81Etn
dXrB5qetWdHm4BYnEyHe4FLdO2Z3YJw56ZFNSA+Lvy9PEWQe04GE349T7ujgU8l/
KZbteeEf5NhDE0W8vixhfrNtpk1W3DIdCRFDgtfO2hQVHibOC2K9Y4vGi0D1cmgt
kLW1qCtBIseJ3a7f3ULdUsI/1WmRg2id02RBxHyl/BlPOccOd7easqonfr/w9c0w
4ikJzpIADsAuxsIx988nhCLLwfsa/Z0zMyxFDkOoQK+XTJCiZET5WLSjmQHrqqxf
Buh7fqwIEDjysTa89Hvdt6I/golLbUuAU9Qs7c72uU7EJZIingENM70kKFMCEvvu
M1HEcbSxIymsUcjGmCM8GyijyoeB+McLZnSE1uKhgcuBW4ISSAh/EGKuGIB2txR3
9dDBOmAL5MXciGq0JtK9REAkiuqxo1+KNjJrzrFUxyTq/Ln6poUQgZFwf4FzAGAI
PwsCmitx7cgs1/UuEddg5U/NC1r3smazXNdeAFQudIcqF0pm3iWIrTSbUONTzQOf
btJQKevqrW+EAkOdiPEqpmsD3ruBoLjIhCnIJRdDyhlJoCCHFM4tW61WYHTvWWPr
L2geC60AeHwDyB+fc/WIhHh3j44bUiylKAwz8r9pr2wAEqiExai9VnAtqnJivWPI
iHBDXJWtS1Ag58CrcDZkKTLU7pWTRNw/uaBwOSYoTM97DdOuWdVIbIBFAxQmQ/Mg
HHpdaOnjVGsOQGdrYtlq4AMbIkHb6p2CYnQavMk+fkNeX3HFzZYnO5oD3lMCmN4I
pzHa2YsBp8En1ASE/Zeymxlw8JQm/JbyqnKih70Bu0csJTc5qsxPwjQDPfck1zwZ
9WTJSPtsyblKGRht+nQd3wOJwDePJozkABXlSOOfbl5nqF0AQolh+kv9+G0yoIbq
0eWC4ghXqStb26qbkL6JRWH3CSICvxEZRZeCuYbi/5XMDOD93jyM3nXDX9SqHJV5
a9XFP94BndbpaufPQHlFv2uW0byYwPP24MGKbO9VnWA7w20h/kJTbdcBSOZp7gZM
g/LrTFJvJpQoNxqyiUaTlkWz/eLzvmTDM/pUuXCH2mlnxq0VLzmvQf0Sm2a5N7jO
E+VvqevG2/BhmfbdXhAE3DXJfgWYgboFDSCgl0dtlDd7hXp6K9Mv8Ci6AeTiLaJY
uP5EYAHRVupYAHtIU/t5a/fWfYLO0+MirE/yqRuGr1h8Ye/d4YWWpoPDiX7yH9L1
5jcKHEksL0Ix84lOn312S7qaTJKJQQxItbOY+a/NV3ntNxctSM1AzOIqwSsUbDMr
BQGZAeuBqBfR4P65vzVoA4rmPfXeCkRYRBJz/3WA4shLiyqQ5Ls+EqKwxagHm5+6
li7IEfWTCIsVo3YfyTOJKvolh99uwVFrymdTNshnBNhyHi2o7y0qKavgsd/NoNBI

--pragma protect end_data_block
--pragma protect digest_block
qOkXDyfL8SFYDGp/MLR6eRPuDSM=
--pragma protect end_digest_block
--pragma protect end_protected
