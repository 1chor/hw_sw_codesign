-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Nv5aOIK7zRTVMHLLrqqHgW46HhdkbXmfoEq7AlrQRCDECmW3IM9erSZJI6xsApe0HBAv3Fz6sZci
QcKEydXMcjhbI2DcSMGTvC7n4//qOPXEmx8gWjdFL5xGYqr8KzNsraQHrmNIFULby6epQ30BXpiW
BOVgOd+Uw20jlAhK4r10FBCGmemqOZiJAzzyVIyay17YL4a5QL2Z46TiK3bl4HSLFHHAxWz/QyoI
8xMYG9jYegfJXqY8zZYc244TtkCRj8g1vyUYc7aGB3axwRrKN84Z76aZguBn/QMgFOptra/Pqxvy
zzZL4x7YG6O6USMTnDQlls1JTU/vRmbJs1mETw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 99888)
`protect data_block
8EFnFkVHFI+E77xPlVY5Oq2OqaXg+Q7fcTdnOXTCpMATcQoeQbJkXV+jJnjEDBCVUEFhbReliUTX
YUfxnOaJOyun8Z2Dhg3CVPj7pg4T8wjv/Xzl0jAzzNURaTRvB1rUbEMk20nV7chKiFGPsFjdjiQ7
5abN38qeOFuADSNCZeZahX30BbWnQ6/3b45bW8IWamyHcOR3WvAkFpmCB7AsGLuvh7gQAHUDLxSG
eZ1Xt0jK1xS6hg1GQW/LOOBN6sFupgzr/JCNXuj+Wpg5PwiD7Qr8B1FBG/nI9RQ+VkS3Jg4ETKED
dcF9vUFiCve9vMyJFioZ+t44rpblk3vUr2Nyy9ITzypzHDN7UiCWakSgS8onKyeQRW4tt+kXF+f+
8G2TyKyX0IfBtzjexdDVutuawEmSEsZqhbPTHS979ijW+vON57kvTzM3LInPObGRULROeJS+wQYR
Yxi/ylfSOhZHxPewzJ9egYCbx5eTNHD7L3sg0xkoiXo2gMGcaLYVwYJB5/X7Dgxgc/2Kf43l97Vf
TRffJ9yXXCjQ73BN3eBATTAfZF8vXeO6w9ZJ+LM6pvuUqdy4fCzM3ZngDmWRnNVnqd2zikP4RfxK
WESk4o6r0UsylVCmcS24+l5/qIcPDHBWC9z8I2L7X+1V2mfvF2Rt9wS1hhaOTD1sBJvC2G0wBBq8
uiSZK9ZakIBxcNkNhLlkiSXTzGxaSsW5KTfEp/XZTUsfZB/bN43M/Gf36KlnimBhZO7G06Zys31A
jNtJb64KAUiDDNW5GwGPc5kGY7xupef4cI+bteN3h5lR5ztZujbtBYD1u+/nVfvnOLxH4AYQ9NJK
fe6UCApGUo7U/DDXwgG9XCWpmPERNHnCrIF17ra1DmssGpKIYN2Lj654V9Mpygfo8pqDi8M8REFO
FPXD82gKrKbz1B+HwYUaRNZ17QLNhrApFPbLfkcENAZhmWULhrsohAXIOIoZLS3Hxm5VHJ5+2AJZ
RWuFCyYuLQCJLPih7Op+4Nf1MJlMHfHi8qPEr7CJrr/d+VEjJoDNnNEtwvVCSIUWbqvlYcgLvuLE
EGLLDBNY7ry48b926Mys6EiWvQfIdd+hlgbJQBn7nFlYKNvkv3LFpG+Yf7p46N8AdCefLVBt8UAN
ptrh+0jvoQ9BxouQmZDYjDgicxm3wiw8DtP4eCW+T+bR6m8uJYt4LQ1xwIYXz5K4o3nr8A6d3ETF
0qK2Hrhqjoz0UuAB5sPf5CNxsdHtO0RsZAG886bwPgIDkqJaDjxUWUpXyURrjoEiBWGszU+IFtRo
oJHrrxFY/cxyguiEDCAMWqjaEyO9aBULtJOMchXOUf7k8XHLmOM3/t5FT04eNNFCb/EbjCrOpCDH
GTYnpCWL3sbjYPunyP9jWCXG3A9jwkBGJuc1u0PS7kmBuFAb+ct5i4zVaR9ujEvK9FPWkDrZZo3S
Z00ZxiHecX0lJTDPDyNzDx2ibh9ZBf5N44MrVvTcZnhdYEl8/CXpzzr6G5F5y8sBtXxwkM+YlRKf
5Wh0vXHgAtXfFKlWhP/O9uEochOBuk6ARo+OndKyqTQYfy5YmSLe5h6oKwDY75DiYCVkxOF4A98y
1JGyXA+cCTj533wd1SNHC2ce3PR/k0ui0AZ1YWua0rjW1d9NfcE7FyG47eWpI7+1a6XGerWT+oct
Y8MmMPxjlyFTJZrCwID7i3ji1BypOP/gNA65LxoOlWzGRSDAH+tc8/zR6M9YoQmk+/Eti+2KMnex
zrgckmK/WcNqzSObciUwYJr5AAbDy8+iQgf7GkcMAcH37/ohpxcgdPA3onbIBr71YWRZyAN6XOPC
racGjHAAXTYFeie4YZUig65guPG7y4cSma2aerrs9MRpzw8R/Y360BSGVOyZuOEgvD6C8qhGk34L
0y3PUMI7m7OjW2MIUW4lL+7rYsx8wbsLXz1aA8zmEABrZvvaH71+bWk8ZaSYw92tJGPse6M+Gt69
kDX0oOR2OHR2vNWNeP6fmrdXeYusBzZobn8vY5nK+9QgXi4N2WZo8wxxGTGILmSyyHksMQ5hMvMD
oOGUHqL33xDq+BI3LgiTtygGvtwoAXtcMen94gol/WP2yF8+5acZpPTrgnDDJbxfQDRBKxsAPV0S
hh1PCN3X2UI5S15G8l5Q3OhtwcHviTqRlb/JwnUI3ujfz8q0xbkVaUaytHbAGQ4T/C75I8QqNjs/
qmDXvBCvlKzB/M9X8XZKZJRiQIMfmhQQpqLOOQLhk6Ai6VmOKM57h+bcaaSY+vPMJkIAKiH895+A
cHru1/gT7irKnrGe3+lQecWGGmUs0uEPGo0zK81dkkFFev6rRHPMSCMr2/PB/u7ncVcM+cVKK0dD
gY1KL+OuheAkTTpsDiXckbl0IlT9XGm2dagQpFpXvJlNE37XROpgNn7OzPVtY6WucvhREYakdupc
kcLa3gb0PPDnRo3cPAgNQoR75t8aYI/D2GaMLr55sJ0+wyVKvlLkS+UDUrqhDuDRKiOmrqprhTfw
exZEq3n6uxH9PmdQkGiHCJYvKbG7ZuICeBjuG8DRbokbfmhjvquXWqkli2PoN9z/uJQ/+09mWzDh
lKrWSffzYhgOrULb3REX3/lqJofVMDTejJoQj19Rue3C1V4PI/ldD+WnIi6I3fq3ym2UaIkEdlGA
WvrubMMGLaVWPJ2sXXkJ4GN4Q+CeO/wdAth6JB1ZYxTcXT9W/i+9S4Ty3C5vXoOzLkNykBQJhE9I
jj1ZhmgFuRjEHjzus8QhJLOjV8zmATorEr/2KqVvt/1qIv/ZSrA5sVpw0hhO19L4NDNBIRc6eCVa
+3c842vaHwY5k+yVi3KfxVsv9ThaztWt8afftVVo+Hvl5DDJY6X37zmQf8e+YaoDbuo79muyvfzJ
wMOOKJ1cwUWrmCoDjJ5/3rE6skemLl93YWknLIYcc0+A/jTOdW1ul8OQPjOIkOoHH1g53IfQtdWh
G3STgB0V3nN8iWhu8BGzRExa3mI8Mbk9Xaf+S+f4AEptOOXZ9Ve9Rm5NKQa0rT6Q/MViEYog+V1Z
zNfr5zT8og8yhcWQDqQVRYFVCXNMwARPOPYLr7O3ePe2z+95tNttCgdUsF9ZL/qOmo9QPX0m9Y0z
iMkaxZEvjB150rRwDNNhXiInnSHjQRXAUKAgUwOmjTdO0Mx7x0zV7TJ+bNAHyfnh8WWszoYRL0qY
14VUMsj4aR+G/MhhH8f+kkqdMq62ggxXZmyBIVOM+1uNv4PJ5zFEZ4mvyqFGMz8E44x/KjOceFQ9
SLgaxQsinlRFlAx5dNadBghvJT8Q+EzNVnMkrUXJBc62UCuD1i8jXUtCxrAMsmgqPm8KTNaoUbkV
2xRTHfJeF0TO6J22z/B2E9HQ3KzLxT9WWxNlTGdcWnHq+tFSQF7h+Zd15u9FV8E6IPssm6XZf9If
F2E49xzV7nEt8+eX8u7QnaobaG3bphbMVGPtu3s0Nntn1sgzC6qTBeSBwxdrlhVYUL447ApPwRgm
VWzeExKRDbYLrLHvQDyhtZSCrmiwMGfQpOxMFIOZrj2PYjuxld7oxc6vXgG4VeS+9hLR77nI2Khd
w24zHOjTVlMjxmWJRT/qNvqHpUx5IjG1BvJVmXXJwRNk4vliH0zcfVAbw9R19PWFCvbF8rulG8RQ
zsUrado8IOG+7zsV/Wq/NhKbI93iJRolft3fKsZNP9IBDo+4UE4+N3Fyl/X1vOomqX6kZVajnbcE
oPBr65WIrBcUc0+Kb1biqnmFcXj3i/X7EUNb6GjLzlAOeELBqrLsdjLeZW2XJ5cEatitadxGLJQz
pRAoj5EKQsjXIxiL7ndurIfJZKYGFcMG/muMkbdKoVUmvdPPq7q+p/Ak7YEX79/cLm3E1tI1dq17
k1g6ag0ZZs5BjAdR1KhesY7Y27UPMZ9adb+rCsjGdrUYqbdGo5iOjkdyt3+B5vIzpLOnW5d7t1Zh
c8v36RDFpTtmNVjYFMaiMi+KasueWT98/YJx3a/5YM564j9LtcpwTfAFOoHs3ZOk1QYTl0ou60MY
VVLHMwY3nkK4Dqm4Q9OaieId1P0kbUd1cBNggHQ+q6Rsv/N3sZHhsdvzqVu/K1zrCvM5tN0N/gxC
3rQ54nMK2ryOSJskklZaMa1k77Cc6PM9F2DylFdRfQfiaHW0/SqaTogsgLDIu1DZCq71qVo6dKrS
lCPhni3WUnAw2AFc8JMRCVW0Sq2d6z/DGvbcgN0lz7Hjv4tijADmJypqnpZi7fcAUD78RYi0uzGR
X7QAw6nbtNMYNR4qTF+Va0N9Uy4CPvb7FQEoD0DG47Y7bZOeByL6sqaWv1giW0IiF+/Kvh68B6s8
baxOo7Uxjd7a7WhzimiuOfKy/bLViX76yCsjPq1kiZH2idwAhI/FMNWofJCUqyBaY0XK+zE/95HC
UE889meSPqo6CpVula0QQBNMtrUmfvCoWuyIWa7I3O+31SPBOSeLmDndbGU8CZrE2VXNsf+js8B+
dwC1hHMeLV5yd7ANUc9Fd28lZwmKRU3dC9KHphrkynEIuNb1BnTZx7+GQACQPVZRRHL2nAG60PjF
Tiqw3j710zrKxyGRDfIffmQ1GQchXZbrD1NGP/dalwwiIexRmEnCqyKhwFufzVV16+4Z1NYE4jHd
R21tdjPivRvriI7YxozZZGsZP8dUItvzqzLO0lHkmcUHo+HTY0IKwwv1+EAofHmmMMGrUM1I66ZQ
TbAfFyBAwWzhcDR1etDSYyGX1XvQjKBayLjLwHCVEg7xAXr1MjmhCfpD1DNFukgJ6TmPxiw5TVX+
TqM1XygZ7gas2fgTKUPfJqzcdHKJXMIXMMUyDr6rCn2aqEcLKbbXk7fFwpYYu8Dg9AantOiUwdtg
IBWI1YXyO/fPHJSuM2sYz4UC3mJmQyzUTcEz1Tvcq3pyDUoFl9N4IIKDgo1v9ZfvwjWzipCVOLgq
kDwmNTFBGfovrglK2Eq2CiKaEE/qQ1Os3WeR7Q37HbaVmNlUiNHj7zWqaMWcdruz8SwdL0MC6tf/
PYbH3SVFHZn33qEfyALq1IJIobMBi5LcwZD0EMoZHgoJ0csItXnTihuWBPEmwKaizZnzfy1y+1Rm
Yx8m5ZLxWG2/DUwqoDx+stvpjBBEw1oBhEBVYEL26V/hHs3x07uA2opcQ3sT0OMPbMwotLCc/1WA
RJBzAfiffv0baUNsufMfOyAx/RNPkWD+g5/z2yrLKFEa6dXjCNeC29mU4SQtuplIAGMCgYRBRavM
qO3aIxgHcmvnZOrr71g4Ny/2yS6fwjf375QLquTNoQfbtxbO4+Bscn4TamZaWNPUc1ZH5k8G7piY
PuOIWzmgoRXEsS3376LdacbMc5cPA5EJzNsa0mgT6rKxHWI4b2w/PblE9blhF+ZehwD3AhNjOVEw
WJ6xP/vvjJWq6Jl+L3ZA6FW5By0KqNose6HftEEFCa7nIVINkELqgE3s7rUdsVgcpPkRJ7WkteJG
F/ljBca11SPzKepEpXE9iPBEAaPrIDJ5sU4+MkBny1zNUVgVAi8+2fvOEWXVL3Vjvc53+yXpiXbk
gPlUbvLO3AlZrSXcLIEPxccMF7vu31CAUGl+Q20R+1l9nzDfd659a9i+YKNKDiVr53NGUypj1lcc
wA7Woh/y40v38jnZs5vT4W/o4+p7V7JAJDmIFtPs37EEvK4hDukl2BYQvDzmLey4eqJ65+j3+SOK
sKq5tygE1il+ZlTtHhCh/vVIIR2diLAjlYcsmJ+otLz5U7QFiG/Np3QgjaTtEMTG+pmy6/FB7Zi2
4KtGvNl/i1/XYqAsHrWlBaNGZmtoBUP7mIU2AfyWobms5zm5FF2lZaG2mc3ePdGJ/pA4Bjfoh/84
kFK4Re2a8765/LXCkE4bNqgXwLBqkfeLNQP6o9IN1jlSdwU+D76MYNYG0ZJSV1d51yt8ncoVa69R
nGXRUfqMmKRWDldmus6N1ADGrn2tawmwT5qQ0pRMt1RVnBK9OZbf2Dn7pfYAuZWti04DiUN+auDp
x0mEmOtaHh2fAE4DpK+A66/kZubDMmKHaNvZR3HMv6t/MJ6MSFgElYOpnays2mgEtlFG4x4bCqnn
2LfhtefvqHp2VsAHRLjF8/aM/chybgrWmw6b24bpJJjYmiAFK71GfcDdFndkeGuLECRKTRGr6K08
7IQ0HLggxZXN4TdFE08ztqx9qebndg7NyDqmhQsGCw2gN/rztYoBG3t/sn8GK1SpCzjqs4vxW5Ub
nyqebLzTVAHFibjJRv1k6TvZ924U5k5FzDNM4Oypieo7NjHlnrIgpodrtSQgvZzC9y9Szg632KtH
ZOH2FJ2TXu0T+M8Ix+LIMC9g3HxLV5sVipTrgJUX31c8q+XvrYktbKsPbZZkRVcF1zESgGCtir/9
3+KumYl54kvUqjE4WlLyjCKG2C18fzhYgAa4+Tq66+6gn+OFh6+oEtulq9VB6p8AZW0enp1A9dFB
+KhwX6W34gD/6KBHrJijxRw8dktbpRUlgUHPIbHWqcIWV60HZicU9W7Mo67eTVRt/nHA/VoCweX5
WVdVbZ5XEE9UcLGszdOTk76u6noxRQqlf9Xn7jVzSxqu8tNRh8zg5Tyc2ApVe3IZLwsUnMpd6dPW
Wf3QmJlsbKc2cviLMk7mxihRFvZTqlzJiVas93bQnEUIZbJpsqI8UVaxBnj1Y1EhHGII9GA3E+8s
XUb7qLOdD8EnfL7pxok+ijRskzE+DtrOLhpD+0jwKE4OcLEeuwVcjVIcVqAg9ygMyyQx4XNV5UmJ
MDeeck3F1GTDA7ewyfyBbJJKYb9yv+jRW26GldcfUnK+CLHSoeUp4yw6Ybk+tDwnbDh8iAKTLpYC
0iC2TNfWN9an3O4X7fw1B1d5ql+M9VBQnSuQomoqS1qD4Bq2YndS1O2d8lk5IZln7lDNIN8B/r/n
jbC2BKrpmUcGaF1UQcKA1VKd5/zIe0bmL0NQEnq9C2f0MxhCiGRfkGUbMJgoKCqoNdLrkHOBYID6
iA0yh7QdxkMPo+daXuI07mB4C21lO/Im7GP+/5upYGrmOPlEQ9a9Wlt7rOxKPsnM9/112yMrX0Yy
2rVkJT5apbYqBZlNTmkOAc/kbSavPkycTQVdwaDeVfso5ukUhm0PmJkmesrTSuDyF3ULgvL1pQMw
apcXpzrNbr+htQEyNOoR9+evEZIlSBuJGGUyWboRBABO1MlIJOt/4Euhvxr/JnqhP+t2kEe8hsQ+
9GWBkgisMzFm9KYJn5fqtzIuFW3W5OACTnbdgkA7XPLa0mRVVtZCd+B+HIUVHlGZVjqYVSrR9Js/
XQP10bj2/Afdvi9P5AtRuuLeDJwYGiuJ/ssY+Z4gsmzO4rNV0WeZAeE2Z0SbVxj2Ybk0XGiJr3YC
m2bDqa/sYRwdwrHE9b2eum/JY2TOhna2rwc0EMZ5ojnfXrKNdInZUpBr+WzdpF5iVG153Ojgmo1L
dpyjdAjtsV6uVLq1PBtNGj3eo8O68QYhXSuW45p3Dp77e996VRc+enTdXwKem3A5Pz1b8pJgUn/7
n2AZj6wcG8v/9Z44imuQqzDzin/L4/4jKDAqk5ZuB/py1MCTARBJZUs2xWDD9JBLewvcsTsU/xfg
9rMmcMMHrxv4ZAgNt/23tAyAq8Qw5X65EAJvW2WZq8OnhV6QfmrJBGOfD7WKSrCXIwuBU+AuCasI
D1ESUuwgY+FwiR49CK/KU96X3+U0SKFXVaB3XRMnV5ebqHZ69Y6/JtxtO46vZVAFGLeNWKIw8NP5
s72shzda+CsmVY8Ch5jGFbWoqaFSUshEKhN7sulHbjfzRw1WUjCpNR3WVmH+N4ws7+w0N+UJg2mx
uVm/EvWUpGjopzc4CVuuQnf1445yZDdXqdjrrVBR8eR5+k5/rP293G4puFpC7YU2N9bNh062SFtJ
P/W3KsmEXnxi5NcRROa8d9ct2vIfJsDTwQNdvka1TQjGFbIl78qOt+lMniOX12Mo8+DAqXhDf8tA
HXy9uCmypifTZKfbB//RQzOOrrr+Ck1UQ009l+k4X4kJkrfBhweGCgW3z0nuZ9VFuKRxf1J6CzwY
EzQrbVaclBqSBdS4iaav7Awoeee1UKbESVQDd8T5k4GzxLlAM++6AV632A3MKZZofH0AghJBxl6K
lTUVJZAMB9IQNLt4OqnUgnkbqBFKeA3YsIE/lZkG2NZNvbTJ1CKrDnKwt1qi2cULA8fjIGFMKeQF
fujtIbhNqw/XftqHWgvHEqi5gTcCayCokSl36j4A+7eVw/oSXuAurYpjvFw6dwViDnTxF7ze+XeX
LUFmcsgWSxS7mLTSC1z6SnsPjReAWJqNmJxOEXp0VqjcN/0siL5THfjnLSq1kcM7+vKoUZB0E4Lm
zUD5ZmcXEEAC6hcIrqsD/Yu51qXTr60r6UgW/va1uDbE5CLGzUYrfOVXHPT/qewVEWAiai0EvhIU
7noFrF0eGcNYTbGcFX+VWySoP7pJao3BtcGq4I9+eUYG6NcI4Q4JWA8rgxdp/HDnS3PRc4b6h/w2
Agou4aqXhYle9pSteknzcpYOMgDTrmPb1F3SYB0EQ6Opuwwt7npBPeJ0xY02q9NEs1Y7LyFa4BtP
qEYHsaAjxbpBxcTAM8OUYUY3ydw+09VtzKuOt7oXMzDmJtlEcdrbc+sOt22tqmIk4+PW9MTlQub8
zT8wfkYvdNm2mKutLx6Y3ceFEpGNgkSEDvTreRxp7rzontrw/lAzw7GPGLGb9FjMTJ1Gz8Xz73RA
ETEpuKRQxcSZvjlw0BFYGlO8af/0ziDaBU6f6oXfK6CYDMoBDB36xeKbcq7WsrpFKVbFmFs8zR+4
DZHmLvDOzBFPrxAiqM9bx1Zv/Z/LitOUFQ2JzVSShKlhbhKyB0oG8PW9N3IqKVhjnSP+SmWGO/H5
yhus/+BLLxBW0D3R/xR7nGNAlLit6umwT0VpN/uB4JfC2CCxzRDbzp7kxvTGm2cOiRujqJ2lMIwa
D+qfFSw6vIZwIxndjDycRsokBJG7LwRZvP8/xdF5XBwrkrY+A1w972wK5f76Xy6EoH13iUIsj5Vz
vlH2aSNICTnI895tCrgJxVs9TcMk1OOWz7vOvENWbsJWcyzd5WnDg9hc09zSdwKfeqX3prNR8i8a
n+oybenck0CDFkQ/70Kx+M8dddXG06T3X6HtOBQfzoLiBsZOc+xlZ09+CoqcMsMFDwXvyisOrryY
3RaoVsB6GZhKs6pWUYKbigQlW/2ezqG2nYxr+Aov2YWfTIfE7NOuApQjkUaxoPkKydKGr1/AIAlC
OyZTSGiTesJArae84xs/+Xq3iUnIOQcHQdIrBn9c+ZBvsz0ghEXrT9YsFJVKJnQiDcWBkXieoesm
5TafBtMsCBRggCMcQipNKaret8lm9vu6yCUI6SH8X9sO4/snRwBUFOW1rQwTEdyQOj3WWPOrHATB
yXQxsy9kAB0u4wOEbttEYMHbLNNvAVfdGmh2IA5e+uOuFJUvRAtWUA3MXgeDUdaFQ+JMoOWZ3PLK
cSklsGQ8y2ug46lZq9J1CEnz4cepXIsdH88c3dqEacrLr9NvKAAztDTm9tfylEPQcIshR3xq9Vhq
DPBx4crzOwuMwd1g7Soa8FUn8eHRFXqsSET9FZu5ILpCAiL1T8HGTwq4k8uh0kMSrN+NccrQie68
25ixBvmWWydaCULlGfAPCXwi2FSyLQdizYAm3htz0/oPhlGzB2FtKIlfFGQm3YapzslsHTImvlA3
gRmZcrOyv9pl4JzHH4n2UtQuxKdesMY5x8tgcPCDAkwf1RHSE9UABVQags0Tn87IKwIfvJxXLFLx
0uZGNZ3nn1gcN6PqkI2wVnr/BeijW75e/vhQ9WlYWpIJjgaY7lTT9/IeY6uV0i/oP++biIKXQtQk
CpzbiDSb+28iswX1X5lia1fO6amUoqAx9ba7tumc9FD5e4dR+/3kXZ6pG8x71XZ+bftWYnSeBCfA
UbU1pB8gnYH/2OlhecM3WJKbprYelo/gdn9A4JdX5K+SAGC6kSoB+fdgIVABK1iHhA4PUf0B4NMR
eTJbaPIp71HyMb0Lk9ljqTc+yNyMvLYiqMyVwtSxRJ2x1M9eVtMpir3gLXeHgnnOnabNTTKNzF/K
/tQxBrwPdfXT46nBT861UbhHE/jmKNBUpIjv3486vXWv58RmSXgIt44j5lzeG9BOhzvGiVK1DubM
uIJhH3rYN2DqhYG7oyuheiHz3O5EM/3IrvPniSG2RP1XKjvuBLQHgr9VPh6CTPRWxzAfj7uV9ZKm
pkoImQRLrwPhh3s3MZsWpn8Pl37+ZiXXenNs/JDwlL2YO++GkD0U0SPmRY5Wzj19bakC7cEbdqme
hYOsRZ4fSUBICzR5gmx5tJGK/yweNBLefN5BGvAKl98AVCr5txsjp0xINznBAvkOVohjRNIGINM7
KbGKEGoVuJXWfmL3xhXHyP8CfkVR4g+BW+ot/o0IPuh0GxUsiMCcK27IPZKadgxyhch2tu3awEGF
bt946PLkFfP+hmfysXR2SJo41t2Z69eKZWXniv5fQ6fC7LMGe8rruIlsVi7lbmjsEwqqc/RWwC3v
i5N8/Riwob09IWFkX8HQTML5JRycBqlEWHDewUjmTbuia2SRQnHIUVbwr5BclndJauTsj7Utlhco
e+vREgylhVtptfobs3gNq+kHeVnHIvp29/dealEQKWjbAmCZAvlpDa3lh9ENc64dHFleK+dxq78H
nKrVSfqzB5s0flqouk6IkW5L0o/DcgONUJgBRH5ppjv+4z5ieg0EyvtMirYApsgBVDYujSu4FBv/
WIRrc4RHN1biIPkpsaU2ofGr8r2/TxD82YccoRy1dzt4pwYt0q7BwomHr7TMNNszpc8b2qNEc24o
kbof8JwRxwENPJFqn6ZebRBjc5lD9xkAMqgg//g5+W0jrtmKYng458VOMbnD8NT0hCqoOdWzG4TZ
kRJ4pAA1T8AoNNsGtO7zrFugLhOHNcJO4n0jkwvcjHMmO+SdptBlcJZGcP3nG0aF6AF1PHiuX3JI
6MHNvHjbOscHQVSJfuta1b0UVgEr5kgFPzMr2y2wyKTg0vANho3yiUrzXfZZgWxehyMoSsbV7lnM
0upF3ESThw8qMFGMiYGkDkXlguGKqLFvRvb2ekOQWu5hUa5cCpC7nKKPL6tPyAW2r0mY18vNvCKr
Nk5CMSk5/pxJH//A2Bw6w788ERckBPtOCUL8uvP4SPvJATc37SPf7+qdDVYdo1qZTXbz7XqWHKxI
CrX+i2gNrjDtx+SLDcIL8la+O/lw0fFAJiL9mA6um2fGzB/bTMXpmJdsEpLuz+4uRdTVMRDQ5r0L
e+YNBCzc8sR++0pkDQd52qZBOEbJGh0zZC30ufA9FJ0veG15vppRwi2jor5FmTbmr+jJ3/7Iyoek
C3lXEb7C5+LCvHRxfGcltDnkbWLu8pQfMIBmpQSm4hg8VEohI2nboswSD1VQfGCsG+EtFVabDqSi
TnYN70kPitB1U5z1dsIR6Q3W4jYKUxwYc/oTrM3hEwIruGRJNXau6lnPfYr71N/41HULCBQpb6Mi
a7ebtUsQxKDcu0m2dELycngAM+4cud/KYoaIUGEUmtg7gFDMg6l+zJgPWag6bOaeO+7EqWnP6vKK
RdDYhUqvHGw2gBcH4zmxBfuNUZNMnn9s0TO+8Y5I8d5hh2WUkau1cP0FsGB5ieeVe8nUAX8795e1
Y930gHFoVj4PrPGIpWxKjOnK2W3HZherIxmAOLI48GKyj59751RF34gmfd4R8CTswq8zCISsp4CO
yoRmUTRLU6193ndUrN30/G+jvdt5F7PbY4Q7oJ4zNTj2tdUGWCiyTgtjPwI3sbKMhU6zj6FkNSyC
nSXXuXknP1xwl0ZV4OYVvV7vHUSShjYHFRgcBPcwb7cm6NwKi6Lco0p2F3xYzE6aH2ZJfRpyCpnq
CrGRVrUXR6EVzUzVwJbO2SdBpEZfbyFoZgjEL37DOX+xUw2gmR7A5I2va9H+KGz+bdRdTRPSI/tg
PR29NYQmKVfI632Jfcq+/kCgPDJzlxYFKKts1rdFCLp78GlAcntra2KyUexApMSq37iDnAzByie4
UPxWY27An5o9+ujFiZ6uuymHelKOOn/cihEHeU4+0x2G6QxMrtNIOdC+O3AgQseT7VzRNaX5sVr0
7DomXQkyB3ObXmsx7mPW2XXOlDjPwIdGzn4AhaH7RlhAOSWDrWn3tknjgzGjS1OJosX9/fnZYcSU
tV9cAu6zDnrUwEutkSfRK7ASjL03ip1g9KzMEhZhI0Zhxj3S1ZArB+nxNVgRvJsEr4PhoDFjyZnc
YK3n/ODdHZ/nOsSWgSOv/Hz+aRDyOfN8xGld65oP/CYOQPHWsRLLZ0Rpw113jCu3aMDTuyT3/251
dBAWuTsdR+EDR4EnwIy97hTwkE7W1wOn0Qr5eW1/Q9ulcR5CsLZVQWBdwggQ0oRMtDW36IjyltF0
VSKmwzQfvN8JP5wO4jKGi1jrgNPhR40k5wJ3NRoJ2iU1KYvI7+e0RC3LDJ+G0afJehDE3E3ttxGp
WJyDVQoZQVxNLNztCIvuzw/r6IRGNXMVG50L2TvdjSmbhS4FQrqoOq9ooR0/ZZLGL/5V5LHhNd9z
tjdOFjQKalK5vkicb1jC6cnfjFrZ7+vXC5pEfWKYseq0dLhqsPzA3ISkWSkXrJEFo0PiMmI3+HCt
vEulcYIZwjD1dSUuvTU/UaJ02YmYfQtNqlEbPxenZTMt8oWNbfT6hs8ovnoSFHGyeQMlV1d0RyxH
qRacoGJTYVIOxI/ZbFFwDQyL5QUxbzRwYWC/XbjsTvY1ZSzi2mbh/9WYcdVoRvIKDbW6mYxAIKpM
1JQFZsyQlNN5EiZ+dIQ6wbTQ26LA1yc3BIUiUdsXqAdOzP9f7gfrQ8BKlziPIgsDKqrPI/5gW0+c
CUCgqiwXn8dRtP2aSIkHbv62wh1XFlVBJvucxVX75P7YKYWmaaxhSdWrh7PUkpVhRnc1wik8W2cr
ARZBN736PEWW8T+27q7f5VIOqfIrOI4y7O31MzANiJODagyJvtHGRzKnoCIwdDJ+i6puPlyAcUcH
uMZNq0Ba9mgTdaPH7NipkBn1wEXTGj0J/pF+6Qx9OlrQIt6+V6O/6qNfsFKH97G4TNXbwiFsrKBZ
j0M5WuagjAix5PvdWkBrYzs+kZHwI2AAfWiMudePwnBYHqdL8CtCTYoohUodI4tctUTjRGvK6x9Z
Xz8Nnt38vcGIM/ckXiDK+9BdSDGjWtiK5yr30YUI0cpqoIvfaCnk68o6ILeYwpfWWWLGYiX8ZA/3
mQ2L6L9PbQqqUiHVeOeXkrzTGC/zp/tblS3QnP+S5RQno8/iYgbjIn++3AF2utFRBq9kCJIRvNL+
dPZnOkpQ0pxS+3VmGo17fxEeWGV/sb/ocqZUAEazs6GNxHgcXcHPSHcCYOj296yEw/cO8b28RZgU
nVXYDtSov6K9N9zhm5Hu6CADwN5K70vrr4t0EvAkZJSKzQrC+eslq04/5IYN6C/vBir9mXY949Jv
+u7pWqDgzzEdnwjLcvUOxFoOCaQfg33y9ifXWVRaTypbE4uJ7M9WUnSdAZgunmx7Y6AHqApuYKfJ
q62xtyPx2EFfAO0KRFeUSeFDHtx6+kTIf3eNByyHVGCUVJhydDV2eCNQ3oTkitEsUyK5te19XW4R
/9ugoqbsXtCWSA3FKsprZ+cHA3UjI1zhUC1HkgQVXVgXrK6zF3tGmR8CMh6ua+Xpew+egSEBU72z
rp8h+x2jMPyqbfEY2pC90Ck1BWHnioXlrDNbIyrXqMNOrg1g0ek6sj/w5OZJ9RZqB5kx2Cm5oPUI
Klz+ZN0aACNuWHCKm7gbR4yfgnQDSIBYF8a/WK9Nuu4mwu1vE1CjQ74QcAl0Klw6zzaqEjxU2bFl
DAe4/voeWnOMR2sC03lh0YmjUDLMTwNSZgk7BjPeY3V8iWIXcZ3KNwnxuG4iRm8u9Wj1C8Op1RsR
pIrQ5xs8vdtd2ziCx8NJxe7i5wMq3jO+UOFbQYFugDMw9NH3/EuqGxuGLliRAHhFk6w+qql3rJ0i
66aA9e+/xNf21jOsz80TJ2DGPSV2EkOGGhnVezmuO63UgamDQCpXyQXq5XUyGIbdkkfWEcDBc2Ez
DH1tEA5rNSHyjy+gjZJKsiwAPzkGC5s1y64P2pt6+RmEtFMaKwCZ/3IuxP7FWohrK9LDNMVx0e3J
av53/jJKsny3T78xNqBKvIk0QhzY1ccD0p93Zs1YkLssWfm1bja0LwShb2nK1YqC405VM0cM+OmT
qf720ZSH22OWERi4pZgcc0V60+JCYIl4vWFcX/14/WV022VbV/j+VnGQKo9bzVbL8uIEKUmcI6oW
CQGE/sDr9iKNZxRqxBujvfUh/eRbhGZhubkQMrV0U3m0W5+y1M6SSVHD/Ck71LC7nhL7vH6H1Z7i
JwYL9U0UQ7L7YN3o8bbvMUtL2kxn+K2j28Rb10HpCsmgu3rqTQSScmIvkAZUFZ3tQWVx+WJ3WKtN
7mGjTattf/lRztbVK/9LtaI+CNvoyr1w+jBkPxENJYFIIGt9Siux37I+sl4NuFzJk0I/3qN5ffw+
O4R3fg34+Pg/UBsaPeTP314wJmVuBlsjpYStnaoGd9IVzEhSXqB2vVr6/ZScmZD9zFEMJTpj+vFd
Yz6125JEv9+xIzFrBr8saKw0FYBS5UpE971zOAHBnCxmaLauhI82D1Cq27eJDGS3Hvf/qGrLFn+l
nxhfg6zlc73brjnl4pziA9+fruW2a7huCy70+sBdr8pM8BxNi9bX1EPvTFpULbxVroIVib16gjQP
wVjbNVyh7bJIuOdLHbmJ1COkA/Eq9szGPYJ0qsTrIxA/9QpTcaxEEwRkeMFUZve5RMYtZtRgT1Uj
Kun1LMgyJKB88wCDo0uRRKaMB3UXnP9xRtLCLZ5mJZeZtm1hZlyM7mbPZe/SvVghrtLG23FUiNVw
p/uAzfrvYRahWEumeFQJGATRd5lOFdpnXWClP1UyWpwrpGmhEiXALA8amTx4ejhgyNs3cI2EnTfV
Lnp5PRm+qSC0bNpheGWLOsjd+rKydLBlIahc/CweoH8u7dp+2bYfqq8sgW9Lkert++kFM86SGKdr
GfEKSeA5LrSTFQouMm9C3YDb1uK9S5uPbNg6HZ2MLl11yWwJG590v8oLzM9PbBBoujOuCs7YJg69
m/Eycf1h1Zg2IBgOO2QADa7tv55NepIGQRq67EXLJ4xi6Ftqz2jf6nn6F6NI/fNZvBQRO6s2d55D
seOpeiMzhMs5b0+gbvQC9khxwWEuLTBw0bd1JreJMWbGjYz+6tULIU9nH2dV/8CEjLYtQ56g3ZmS
RmxiE/DBLFFhifPAq50uRzaNZ4KT7XJXCYzVApXyBpuOpWaCeV5y/vHUztM4/k8EP5jih/PDlmsE
nbX53ggL7BzSK5njV3Fqs6uTq1aRWQYDZXtrIhxHBp7m36r5KDT65ncl3v9yYwgRmwyff7UravO6
blGRJeGh47KGP3gXOALb6SzaHNGFrtkg5/3CWJtT8yejMmt5i8kmFiU4/2aEQuxH+HGqE0WnutRj
mQnQRh7Lx2l91I1N1V3qfXajmX3+nLqC3p1wv761BvFDVoymhJEkpM7KF4zQd3uR6l1RlbQGhPNp
zWtbOqhdQuj9xx5N8CNCl+Iz5CKbGbVaEDQjcdSD//6WvVmKI9MbGmGnjStvRW2r8daqUmkBhXCS
Kj+ZrrtmiaphwgyiAzttSkqs9KsywrP6dl4v9SXNCyPwH1B7WxFBgojwl9+XOGV27frmvN4OFM/a
Mfw5vMW6hsrbBHUxsO2Yc3w29vw0EFl31gL8GAWEf27+Bxg1o3tdllajJmUBMoTfEc5y9/dtfcag
ugcuUBsJLv10InGwr28/j9FYipG7sLJEQzknEW47uJTqpiQQAveRC/20EsrraNdNNQyNoxAb4lkD
XnoulUUpnTnK3hbI7qf1gTaAbLwpgiGEdIaxcUHhfPduB+zGxKj9AwpoinGqP0nbkB9cmILABDsI
2IzkNgo9UZaatzZIQWCHEfXqaiVVQn5BccgDdp1PnXNJDpGc6zJhonTJygDeD8mdKe5lugoxLJic
cZ8Zs5c+brqSiJvgwBqS74OiUH7C1uACa+KPQh7c5kLmOa3CvuYnj6wBIYXlDBQoTzfdvdPyPLkh
BFIz5XW1LRH7UYwGp9IaesNhikCzmUi3kYBDusqSAbkF0ynKjuAkWRHbr/+X8x9hSGytV/0Srkpr
KwfJHhkkcM4JO35EoCcyXeyDnYwLcvdk8rXV4kaF0BDX42sBdK+GPmIZ8BMO0YMw5nqUSa/aspJi
pfZdgnxI/2sexBu1umcLHIoaObTvYAZru96zxHesjXZtgc66srD6GpllmpR3U2B5YaImyxJ4g7uS
Qz9UNweoV13Wpv8xdshNU4LZwW4UjYhmXp0SVP/RApMS1rxXw4A8SYUDowAZBoIycHMVyMyYasml
LWbdLIXcYoI3Hx6VVpErsVnkZQoSzmfOphozBfAE3r/67N+lTgS+NQBPQQJSsyFVGimnFLloJ8HS
AVNEiltGtbZPs1vZI3qtYcOxPesF15yp3ZKym75+NnbuQUgIWdERkbq2IRpsWbf9lrFRj5H8J6D9
Rczm1i1BPeLEM5A9jetxibCyLXJrVFmswj3Qv42bVzPAQZmKx/F9isWK1xRfUL9TImi+ISh/sAnn
a4xPsGOTQlhKxBxmX1wM8sLGcSfmNp90j4m3WRhaeCdySDChY7gczUj6YTumwyp8X5O2IWmYoeks
piceI6zY5KaaspTbh7GsTW0BQt1h5hQIYT6ow7nhQhmcv29GkRRpqhstt9wOWwJATIsKwGOSdXK9
qK++Zu4eKaBz1MtzgNF90GmwA7RdUXUQAHLw3AzIObMtEG8bCZmaozTjlXV2baK3DYbdtmDEKXts
7kSxM2htIZ5aMCP8s1bxGj4bzZmN8LQkDLUGAX/r8kpjmX3jBdARk0JU/O2pBClYX7OtGCbSMAgO
QCj7kruAcqVZLvvzRYTAyrQM9k3E3jT7sKiUBHr3Ptj2VjlR6Aqx2S3tJcx/8lgg2M3zDOib9rDe
A4vskH/RpY8i+mKnc65987lT072nFK9vI+A43sgJTAnEpk092NdfKOMZ74n0Zs2eT+GubJuoxEsh
aRKMxsReKviXt0eVRp8hTftX/nQvqQj+8R5snJ3Nv4z6A5SQu81jGZPIA4OG1UPPqL61+rdjtRac
qDfbBlt5EP0Ow0dlj/mRofyQ47wdY3iagF3uLP3u35uwCmHu9W5mWoFmuqQDFBELUNHa2JQ3lOfm
7bsrxDzmzU342M6D+uFxkEvKtidoOOtixHgcNuTbv34gpM5dD/21bvhVbCHODz8wZQReipQDqqrJ
BYZIx7tGnYL2kxipn1DW1zV3s+Rvy9d1mMsIBbPtXacEFHZJPVW0oupYA+qqILGUrHDxrfdGHJEi
xhQ2ysepnCHPhJHDKP5JUvJyno+AO2ObdCCYT2Et7whG5Oca5QvCqtTfgRs7DZvTJ1uHAaVC35Zc
ooO+UCFoaUGCurY8dpvd5d4m3wYM2eGLyQ8LXVXsyQyJR3F8xta/tINNL5HmJvvMypsxK235mmtC
iJodkApA1LxFRgPk/QPEkf4SdSGmS1h3cNWt3xdwNyiVG4nXVDAh/O5R1Fgzil+isqVOh1lG52lB
Rb40VETuzlWMX62KEUkMvr0E2DYyitWJElrnH6flDA/RPHOopoj4ym8Zh58bWW/MvMBhPzqLsjTH
tgOKc++PS1OGTU+bxTRpBUJxWlsFX/5xa1HYLykVxa04jgwjDzdneUY7AhOjk+padV8sW963HBi0
YYa15tpIvLOIgyNUBTWjXM/4XA1Wircyxas6Aw/+Z4CDMsR8urP8sybgiPiVEwXlHx3oTaKeQuXk
vNWNSLAmBR9YYHX3pS5cfjljGzBTz2tY9do0lWD1dt1/1B8Gy9+re9R5CQx3CrV5/Qh2gk+fFvj2
Wr1oSfUEbbovJze92kVNfUPVMYAIw5gm3D5jW6Sl/mqR8Wvlihv+s2w3uvJxVF5juuyK94TTDZ5u
sMwVgYfGAL9HWya5X/NFMCjbSZv64Ir6F7Im8srBH7NFZF5nFKEm3WrSExEJSjSo4ITcvTX5kR9L
rprCOrYb95DkU87cxJgPObtJEBQhW/RoDNDmiYX0617k4273iYLLItdEZ9NWvPZKha0vSN21n5aa
CZGGeldKweYFddBOoN5Lf6Rq3zxzhG2FWg5mx/nvd9efNX29RDTRB80Y528txvkLUra1SkOI6cxm
j04G4exL81Caa2xKaD/0NcHrXhAQ8knJJGSxg6xpE0x6/fUHg7tbO4DdtOx2KneIh24gh7OykueF
dH0HKJcWEmCgkg/v0E9JdOhAE63/Z74jxqB0f4/BeIywO1OXuJmXUIhrPsf/TUHTSV4DskYGelMY
rFQ8BMDWphbd871Ai5qKJPKTWO6Ih9BQ5pUTCzRlPT3YGcLi72Ga9deTFPACExj0YHJAw8EP/rsO
Mzoig1PNwLHl1dY72VWYxJfqH3yeQLwqogNwzU9Y22FWLCsh7hZ0OzAMOvOF0JZ8FubXvadillxV
fZO2EyveaG4NC1+VbatJSPEBRNkGeKpSPcpCnm39UFd3h2FzxCcS4CH9dx1WV3qfsXj2xbffPllp
ADJuwo6f/NyaIsmF8Y2yXLrOxN1TXq8Hgq5po+SXZu6UCgC07cFDLGmb6nV5yPkhiiXyds72PDsc
szUbWhfxWLf7VCaoUcMhotdVzWce9CW+QiSKk8fX1vXj0PXY6XYzJlqCwToskGDe3Rj4f8t2CZK/
7OxnFI3eyxkns0yaz4o5OUnA9MbI+/TlyNOjf+A+tyCuiHkguQtf3ejJYE2ga3ecuW6ucn7SqdED
elsduQpEBbGNRPLT+bf5Swx044gC6KYd2BY20XpckSyqn/o8FOLgmhu8+6ni+hYgvcRnw7chMBzt
aHqj5dkLRWlRqRNtGapHnla1esknP9DSU8pNTEGItXdtCcRJ9hWLozKqbUdO/+A3Tn4NTf70nAEo
tjuQm+2xwNizU5RfQjdLo0YDs8oYrYO4TMf0YVp6IaHIm2CVrKSCSGTXBtpDircqWpG38VmkEnOa
DhEPxZ/dem3ALM0ETGni6DBRtmX3OYngtDXc0A2B1Hn46H6iokRh74MbAMjqooWCl0M8fAIVFcww
taPvpIbbm62fJhx3vAQ8uE6UPox3gvPRLK6k2QKKluVC7+Z2l4Tj3MyybHvgOD/KsRdHbRR/oeou
wKqkKkC9hyJ11JsAesurraegBiLx9X2CJJmgJX3CSGQr9A+TxoLVOArDxxojmVAGlOXDq2MUwCYu
5tEqYa2IQ7f3WrvheIisY57fa7Mu5+XPwkiyY+XS8whSlkKjRTVS5WxKAAY98KUs19IzdJVw6RKK
oyVgTmyCrO1ztfJpU3UJblQ2jStbbOMmTirUNGm+a/ehM6qv2mtBRMm0uw4eFQSneUXTqX76FHGh
kxmKqdok5UhSuw4Q7/PNEApi+ZNFbtTWcybxboZRzJM2T5WqsLLtJapiLNa1cb+nGIlpEc/JHYkp
v9WeEv/pw0Lkt8ctOuAlXjKLgsHLl/+tROpR0mQnqwyHMKInSE2HmkJ9jkCAUMZpw5cKVtOf3io3
yMnLAAK4PqKcxp49YrJNvhreQWGu0ncS4IGuZ9CLwpLxHu1Ti2Bc/4t/U3TLLYoaorIMQ4e8U0to
3pqRmMU174DaF9++wVAUovlRh/mKJRes+KJBZbtzbq3pQYJjhXc2LpVdyc4iZeHHLk3b7DTprgrw
Op1Dt/tL6q8c8nJ2tEWjhKWZrN96yo+s9/PHxkPZx9lQrpdegVnSUE8wF0l8oAJxlV3SNQ7WuKAy
drPYeZkJ9GhySa2CQtWJZpEXsIA1bDjTsenPQRHW9OimyW4JWbb1hsFSpzuv4FnMOsiISyeHjZJq
8w5X/euLLC/eTnC8tmNWQQEszKV/qY7ZwOZrmbfLrCdpoyDrpHYRUA94P+3iq1OIiil7ymwC15iL
ddx+PfbAS32LTpBUQTe1VnLq9B8x1x05ISqKOj1Bm6omcr6gGnkGRnW3erNIFv9j49YWYwPsEXN5
HpJ3vL8VPu0PDfJ/RlgAGIvd6rgc8nXMOJWQurvOk46Jhzqug3vQDEsH0r4tdAFfNOUMoABjr5oO
GshSC4lUF+1Z8GxJNOGwIW+hoo7QutfB+XmJbYKOv/ydRKpnenop1g7avDI+gpXlNWEd4sUV3Ytv
PIckCyOwb1F4613swsMKlwLBD0mH6rie9SwoqhbJLPZ4uqCHdu36Uy91tm8V/vMRGYtTpzl+tkwg
DE6Uqm82a4xe83/b+aXm2qxqUKgEWaAfizHbOvIBcxsFAH+HU03MXT+9B9MmJvg+z1LKHzGL5yJX
hb0T2N28LJaT0CTeLOxDNEo0hrFlA0C65ItYB3lSCC9oweniV1wEvwjiNmCY1IIeRdGnM0s4PSv8
tLXWecFEJxGYAyKMzzANS6rIx8M72/TBD3dRjPuHIRlgH+s0F1EqMqcmaOdrkVKU5+/E3i3hjHTr
UsIMdjTGgKdC3mLZJsotke+zHVOd23fFAUiLbhGO0GiqnsD98oLpTjAZJNOvfwbcD0uiXLhBd5CY
yrZ5Xm81QTZuFFaUx8hxvSoprF7LS3x2NIbk2KQpi3q50rkcWlCFFC1jaWkPwLCmariDGsxW9VHF
Upbuzbk2gdZRIYrZNF2VdkVnSAelKE+Nu7EPbh3I5qxnAoWDCv2Y8URHocmLltPX6dr6KLiq/T4m
DGvILwcz8Sr647wAtm3GNfcy/EbgE9FvaKVQVoHEqVmmhB7t/7l1NyVr6m58ah0DuX7XZlWiqItM
1sjjkhwGGwmi6kBJBpHmSbb+ALzkbIfFEi9fLpp1bV6IooNpqFvlTmngrsbgVjjv6ChU3b0VmUPx
Q93JK3ys6/sbNTOnv4WoT7VVDjAZNAXFr6vVBevs7zg56jSSmYVEDeDga/gr8sjoMrPxPaoE0Qbe
7jUhqUkg/GTHigWkhh5+2Mi8qxRC57UrhXnYfJ/AUH8RDpprAZu4W9DFFQVs7Ig/KeW4SN1VJJHr
pOoenUO//oMaoKxvmo2Q+bcx5rtpwZb3mBh35QqX+J9cF3Gk0vfCv+yeVSAKA9PAnCCqfKHLYhjt
IVszfQtc+b1/LTIOEOUUZOirHVu1jPYzwwQj3Q4qHAqfiA+IMCViXKiCfY4y0ZFjlRQc0HVdy/GM
0Pxa8/PaCY8/lJyxRpnHfwmr5ATJ/9904llExTH04MSOZPH7S5UcTPvvFtqd01/OrbVi0k6fXCzr
IVOax967aPy51yyFrnQb3OFgCgJr715yJAfEeeptqt7AVPefGvTNKWs6PWZwPKs4Yo5SoGCxHb/o
a0s5bWnL/MnJ5H+OxJzDooHFzdvrLQWzTFRq13y8hkOam9oS22HG4uV8cEP1LaDl9mN+zPbZOhA5
J5CE7aXfQs64WG6tKcgld3RpJDUOMhmvraZgyYVN168XLdFhLL81Vt4EWN29QeHOoyo5FAwyTz1c
IjMuetqX09WDLknAxIOheg+Li2G6YdbJoxDF0b1dGPfFikirQQiUIpxqm+/nnCT71Qbf657GfFeD
5y/kBRJ1CBW+yu++H0kYtQ9NDm1f+WUcYP6NPaM0z1F17Ag+7dKV6L5GjoAZP3WPtJp3djei2JKG
H/PZbaGkHzI4c0qcot/DbnseZi2LDzxG31nbJ7h/VU/1xnRWgV21sxsQVR9NAsgrc3KssaHDa/Uc
0XoxAPHc8cjjkxwg3giV7BaSc2Lbv953pJet7ULxBe0LwNf92igLA4nE4v5zaSxEuWg9JKyGnGqv
XL4ATW2lT3Q6WlyPlIAJl6pokRQ0DYlCu3ngLazo5FMVqBQS2W9Amj932UR6BHGwnhD6iV0yky7t
8rwMJ//ViKY4UsU1ClAdqZYwK75XZCZnQy8ASgMjoRlg2UJz2LFDkcPUFQiSGCh37C2TaB8ELI9S
+TU8TJHc8J0Qp0jK8eHF69KSWzn1FTcXYqfoPlnP0rQVyQtXYDjilAgF2HYkETs52L7crj/qKUCG
IP+c2Bt26km+oEEm1HrB+o8i3rtc2E49rLr422ZlPdoMZaLMNhX5TFHHtN1tGLtspfRzN7/WW070
tbVAVGF1DMje4HlG87/p8iKiQLMfdeBrvzZNdKYmP6p39Fkcv8jCo6FaDooazKYewxlr07H7Ps0o
tqwp9uqppXa2L69ibK90EY51yD6iVInE6WNqLe9sC26ITMePg3q3FIjOT3+tbIiq13bvtaWPIKmm
Rhsc0eYWWolgDnouI2fKywR0LVl4LKSvxje34tRtSIB5e74oJV0tjSgKDf+D3xV6edalzTUJfwxU
rLp4i6YbqEwQab7lQAz4YlBhxOFTc3CDMlYMrcHTxfAbL++A3tXshl1r+jcIp1ZduLYz1n15pwsw
VgRHQX0ad2T6dZErF/e9wmbp2pDX86DyqxJr1aSHhV39X+FqzpjUtCj5WEiZRJ76tSvHJg5h+1n9
EaOvyrCdh2yrCUvBKfn+BhOUUXiMsGxs8ytrDorudrPXOLeNkpujuflKSnNSY9VBOHVrZQZBXGmy
ui/5DLIci5smIrnPljHE2uM8ebWboXVd764HJvEPVZ5Bo7DecrmW89fB5dlNtB7f4HP0tBl3/pPy
uoh0/K403s9Kg6WpzhZRxXZ8I8pka0EDD60/hLLa91htFcnkiZMnsIH+k6bUZeBow3BgDie5QfMK
oGVAdVDdQOOnbpz1NzpiZNCvQ9pPOMBUayXpykopTX8O/wKdjof4p0dhDJwJrtjb862hETusT8LB
WNFaTEc+AOyta3Epw7+46f8aKLkvp2TJHOPJ1SjAUtsHJy7n9kPmuF8tTSJ38HM+zkXG2DwnHVQY
/pJdnzR7SC265lqObENTTAACrOQSkuhyNyTxZ+gKYaz98ygE8vO8MBceAwFn3FPxksZQBy0UCn+1
Li+sp/SAGOBw3sulSxYJebPq/0RPPyOJU68NGEIAp1tUtwlKpZz0u1K3I82RC1CNPgID83HMa5S0
gdMpDD+csFffpSZFrdpaXytbITyHYYvU8nkbnRXwATzIxarGk3ugtg4fTBewUEYNjxpjEnP9awHK
KEVKAAG7OKwgrxWy186zZWbafPdn3k7KSQTR29M/Z138ks0N39EeoNgPaNtkMRrXWwj49AItVNBd
dnOfOZkjCRR8x0IbcbltadM0Fop+nZz59YG6+nAo2F6G9ZrZdEtjsMihg3/nNwU9CsvmEhF1MXX4
pjNEyALupZN8EF9/fSjTGQePiPpg+O8vdlAD8YErfCPHJTiaoekOj243EL7qWQqvPzFZG+cnNbPj
Re4yQv43x51UzylO17D1LPW8cbTlDFAtfoUXj952wao934qdxwXC6osugF7pnHPEzYEB4WFFuwkT
/GvHyaryKHekiC8P4Dmx77hyM0BBWY/WUwat8pyVNBAwYcZwIbXNo4op9VEsSffcLz4M+tjeTLAs
LMzoL/2wBTLN2UXf4LIGWnKKg7vvXR6M8acLqJqLC65S85CNqp3BHQy9GCJFGuCVyyk2/0whG8Qk
h7stY5QSNjdP8Gl/VzR48kdrnjDirzkpmHy1O4HawKown9/jcifK/9DzKYsIBWQYuzquYPIcprmN
o3UFTnTS7GvfJRTjLaZ8WOdH9orwBMsxC2JyA2kzEmUV9WcSTSb3eq8V6vl08sXVLGwj1EfynQd5
OPxuM1G8aFhKDLA1MXeIs3LraVakvsytUxEL2ZLN+o4ffD99A3uyavYW2BIBKnUeNzwaxd8qmG53
56MRVtFwg/qru6qrimravKejgk8DKBRXKNvXaQ5MoGC9c3FqjitDmI/9k9OUkwvVeWlZJ1hJvOKK
eGdcE8Fgwml2TO2rutlUjMR1OHS6Fa71K/wog7MdehmcDCQZR3AI16beIVmOpEuWuX3TKUUlQ6EZ
1vv4oo12+/nTwXH59Se5IbkF7N2N+NJPbFyoOGLRfOL7chPJ/6LNxN32St0zhOmeXBjKh0maQT/E
nkvLEZejIDGxlUvc3Go0u7/WTPWvDu1Jr2JMo58KCuSZ533KRE1eXzgSm+1FRPqz6VCIEKnIl2re
rnRlDl/7l3lQSbTXJDyC7KgObCbPHLlPlyjS7y2f9oSBHsuCUJ0DCt6RMj6c6ZCy8vrxbjDoeS0H
j4Y75C5goeYaFOME4/jjsRdNkCvDvdojaaEvkNgIKe6pO9KIHvxwKztfsV3drVVNRqs8kYGSvWOX
2VyraAumzTnvVLN2khHSpTdDvqzvb4AfFXlSKFSfTtOFVGxxyPFERgG7YJ7Dbol72lTz8QvDqxyL
bvNBWhG56ZomOqgXFdB7fiJ0dsfqkLMO10ge/b13tmGlPRt2G2yiCL2jBALxAm7jydm8hv+VCWZv
DSmTzl0GDWalqGKhb/7rOpsJ4d1engERrxoxgTOnvnPF/U6iNiKr2NToQKPAcxOltlYy2ZTcmQRT
Xt9dSrtxuiafDI1MOQTrRwdOPT0gilVaSMSJInwNq/BpFUCEKrc/dpbdNhpU8PIVP7YEWar/O5Hz
banRuvpJdrsWiAGD1G6wj0sKwsX1c67s30+wymRSdBKuYobExpqlsSYH6nibyyZTKwQvAE7Y+uV6
DUE5ARwWzZxSaVb+6kl3AUkeqFP5ImVOdPZKGKX9HNJbtn9W1kE1Opq3WE1ZhR38bfM0jheUtSS+
wIKnJH+fmhyeOjYOM1sj2R9aD0evAyJYgDjaRncM5r5mLnhnBu65O3zFQsqX2XJj+7ACiNIcCWHr
p9wBdu4EOZcUQ3dGjPtFqbPqnb9zNRFKhurFg/LLry4XmQkf0eXQLepBGtvnNJJJ0sjRKn0R90X2
0RSfKJmial+cYc8BUWNpnHw1w1aOzn/UUWH1cFeBJTCznGYyYKpyj2KX7IwZNvaHJx44N916uvn3
b8xKw8ZD76C9cMaUGelXemPqyJ2w7dwaGZTEkgVr9HL+6vqzLdxHcDZfPbNFghewS7e8sja2Ntoo
5F3RW+ogKKSWOT7RXSS6AkOiOIgfecAqIFWBN8BMaBGUiZGgx3t61ghzReNXpXlmV61VPH7gOROr
k9c0j8clRDf6Pbd2XzS87aQdsb7p+27e5r+vOySxAL1yyOpX5iqCqWwzfg1booYHZYhOdhCZOjKa
vC18pvqK9U5EIWgY7vUGq4/vzOgFlfQAjrVc9c8JMKPhLPX1wpcpmNrsz07I710+H415xt3RsSPu
btqqNuzWuTNaDZREv4Dty7wmzszmEUK/krj8D0Gnt01K+h7ExEsAVHpl0nYUjO7FNkjsH9rtr1k6
QrZQRemvUFU+RxUhGsNoE08UFlrQru3YV5fU+6RtTUl9Egz0oHGR8ay5nrQMbSzvPuZg/kFqcaxq
WSIfzUIE0rEIMNagzl6MN955QkFAZmq786TreBpuqHoGA0qZm09zQIfO3q4busbxYUr4YLaUbCAX
+BTIWKlCHw6UPb8s/4Z5IOYDQNp6ZBrUkZSZ39pVhjvWMknTdlLw32NAahRb99b45YSfSTcqNdeR
g+knUTITNztwH0TPp9Sc50rChRW4iz0GOUZZdA4vhbYmsnKkKjt+RJGFkSYK7Hf7MGh5RGScVA1T
1wCoSyNmOaVAo8CTHBnGGSjBqPNGMQN6Qw+PW9zsIrBXAmeuM/SnIka5QHmp/nodlGbvfp+2G5aP
djOapztEeg/qALy++YuaStEgQ8KBrj539jnZdFB6v0we3zq26vWH3wW0/3dpLSpZWO14SmR3pBSL
gV5agGyXn9vV8VEpdgNby9qSQ0eBcD0Kemh5eb4Qx9u7SuhOH1NFl9oy4yBL6+IsvZn4h7ziiCmA
KG2gc+2OLaR7XaOvAi6jKS6GZD27dPlr8VTu4gZ6mlQ7AlzmvFxe4y4lmRMNMfMVXNURj1oclGuj
fBIN7p6cizb3uNxcAMGGYIwc43n+wbdnYOV69jRVyhBIGXlgVoZy8sY4o+4toSGOTJV0+HqtPAUX
LB44KZH3KdMaCIQ32Myf95WVU/uWkTlDFCGxToGlicFx1FRFBAmn8iIF2qJhyvvLHSGZ6VdCUEIV
aczcj6iCjfWoXAPGmMhLusr94LG7KzrejEzQr9NUMbWwHE45a4Q2s1kUaDl9l3Pu5Jujzl2igy8A
d9YrzgLDR5wifPZyjNOHNMdynBeLqgUq6sqlYZF4gIp4EobhjQnmt9of4Z3WTMWPob1gWaAKAb38
Wxss1r7snTEG6HfX4avopZxtwM/NwTscKw49n5rQ283rKzW9JrHrX4w7XwKjMDCmA5/R+dkCI4On
JK+F34tT0snyNEAvR3KVCbKu07Ri4qBp2pnCIukPMiMBtVPQ+jyQsC2+GxyIGoErYYmvz2WunXz3
ZMUW6RlTcJOeDiE6F6BEqv6w+abKJVTTE0FY9Jpvfo8hfHK7Mcx6ERSx2MBfQpOuiSF7xn0n0/ft
Q8VwB2MiUE9kJeVGmw9nabz7UPu7D9pSdqNT/pKitmkZRzTW2qr4z5hRQsEZ0hK5H6rNv4nBtA2S
IgIUQP68n0Lfa6Z2QabUSjdqWinVK7vnJ6gUl4Gq+Z8hWKBkMGBpjnTYMG1lIJEQrrHacUt8gnHZ
9U9ZzmWLcuMkfA0hgLDVTHfie5T2nlHT6bnSYkYEF61Sbz+VSbCSvvIOSyTnXHmFstCiLjdVUiVG
mHaV5i4bPwe2af4i6bdRa1Nqtm5J7ykrHHfzr579IRb9jl4f5ydH1Vav8nDalyNw8KBrxTv/7pH4
is86mOVtMj0+RjFaajP+maYL0qFSchJQ341OnjJJRcaR/vJQHsm42Y6JW+mlNKfi9JErxu/VVPKY
xE7NmZtma9HTgXteEqjvF8nq3lYyouZ6tRjq0jIXsYIYFSSyBSXza9lfAPhnNRHtWfJA7ogRsKuL
pYxxN2+9MZRvUDk42RhAEHpZVrwZiVl6KnPudGA4O1L9NblkISSuq6idtnCSdZZdD4ln/ozVfBlk
+0n1t131CVMKuD4XDowd/xCF1DM280XvQ5e9mJwid7UjvQ/oRWcRI9n0pjKB5YHdNAFkkouF42KB
l+vrypQcnK6lnYR61sZd1+6BTuAdbr0paYmS9uoWAmOWMYn6J+hx4ArrjPsZ/d0Om3+xc1wxxyLd
PUyvc1toXKpLKg9T4u/vHab+1HgN7fzFPJw8MD230CbkghaSH3d9+HstB1Xw6rpMhpamdBJEnDzN
nyUpZalB4ZSUmnxmWE4sGXUmQoK7ugFyB/ruagQJyNFiHDtyRnJrOPPsAXYRXX3L4d72bWWx1w2s
bxPPqjzq5PzDD7ouW1qhNnFqQ0M6GACSCDlDrcgX2LobUCVAY5scsm7xwU3ixfkIGseGi23TMaJa
h98fdD2tR5R0vIesZyeIlchXl29t6A+6D7ue7LYobV+wUurnYxyR7TsffVF11cyG0d7F2EnWUuvL
Uwcme4ylitEq66Ic+HlywQHLhfshzjISRndmexxIZPbNcu94mgUGLNixBG0+FpoWA4s5OYrr2b+t
lAUDtCtEXz3T0X+OAWCj0X3i6PIAvdsBsJXQGEbqDt/fFUz7MHijDc+d56rt/L20/eOXddE1jRyt
uCzwF3P5E+/rnDZVk5LGXoSpkcAet4KkzXiGxVyEezoQvlO0+gdP65idVjJ0F7kksEdRE6N79wwu
8nyW3PpFvtI51n+vhPQuqp+3J2txLutDBuC7nBqSWG+ve+MeyIhLRDgSmg/jTuAZmnUwk1aVxe3H
gAgeaAI0s/gxtu6DUQeMylAAe2Wp/F1gcjoc65+DDjlc9653oTDo/3+alPTsSMbVBfrTHJLa16lS
WqCMmHbUWCpBsDWXl0iyPYwdxtR6pFONuo6ccsMlH4+IwteDqWUMWnIxzz6VTTcD+H8jXtmMozXc
SjlydaHiivqrOqlAbzPkDMCxiobd8S90ZwqzcQaPqO1hfGPXkRlmd0yK0UVRfVhPAXOyaA6A5qPV
sGM3atnUlzfTxuVbf/RuPhHflf+G7Aoi1rn0LAqa93ElfeJM3dpUNN4mAdljBgqIklS/+PUdRQ+v
qmXdC5HiBCOVoOSYaDqlAaZMe80EucT5/pGhkfd2xB9wlUwDcu7ce0UCAiPFV9AiW4GksBdMiIxT
RH7F3wKX665+K3PAJdoyWdeVICV2/fj+CNMkm/UDQDrLh+s3d2U1voZEkCtqimM4qeUPCnDDN9sO
Wcr0x5FjBKd9DiO1Xv9RA0PmgRPW7S0W2+1TWI6H6Bf2hkPKVraMm6xfbkWVIZ6AYWGwFAIdA+Jm
D3dh7KLu4CzjKSmgQZM2hERpf52ukErnQR3WqjQc72sNV9+pro7W2MQPViJuS4Bk859+BPJCTV+A
hrIAJhEAi5jxc2/gcGLl0KBS6k2KCF8WwAYhxaFx5jjWlA2uIO+BXa8GVShjZMVZu5V2MxvCZHpi
c3oJgXxil15TupEvyxA/+QQtKF90ZsWNpRXJtOnuLrZOk61U4lziKkO//gGV4Palw+gTvFZB90DY
2Q8/cVN4/XEQvqp3w7oYnWFowBq8LVBm2+f7/4CmngVn9vOyreD/Mo3ffHH/8wUbra+180Ce629+
TMs4sCTe3PRW9XYN6Aj8tI8/nB3trUaQwKVHBW9hTPs9xqi0ktwa/e4UkJdnEf1G3Pos0xC8pd4s
njNDU0fw/uQuC5ALbU6uvHK4XgDsaYa8ioaZgUCJFyohpbsSNWY396IU6JmJJFVL7xujIPt/4snV
Nw5zSUTJ1TjJdeIyDI2cnqtVUrsKnhmaRS4G52IX5QSGwTbsUM5hYKFyr3S48wONlWQXPpXgrMsm
8rgCNl7fEyNMt1J0cyKny2Bt3rr85PxDeC0FHl5HypsFL+iHv4H5eQjXwo1cxNGIN+43b0raN6N5
/MOLyeWKjjESEFz2ArkuMBSDJoFuTgbX2zc8T8v3j2QBP+vlAneeek9PCbTqiFVFYqaBvw16B17r
RCdgp1oCOUgZ7eHE2uaf48RXqhsUDMLmnwEgcEmNJc3hHTkfxPgqm51j/16CzN4DHnrZ5X1BPDii
kUYKBdJnlyqAsOG929UBTgVANIV4vCX9ar9KLBk4Hnd7MsDz7J4+CdcgtrAFjGnzfVOyd/BTZXwo
yey4Zu/jF4DTMh+RH04unH/qvjVIOWAA5tWUeVY3x5t1/bIzH+VHMYpbC3RUQawhn4vQA/8kx6ZV
GqOxs6r7JTbZGv6pTVMhPzmldJjcZyTFIIcNaR+N1/3BLQyqsVzYpOdcULcKYG8rEPVRW7WfTwuk
mo2VajZDUQRYIAj2W7sTwDTQsRbJ+bWLMgjBYv6EPH6RGtW67Bs1+qhtvbB6j2xyDfK6umw264bb
RIEaA76d+HMd1Ee0wWZrq9yt2x3SqDR0sLZjTaP0+1vaZdiXchkRsrhO+sy9unrVJMmL4/6OZ8FL
iMqc2mzIShLJLsHdFLx8kgEPH4HWggDKW8TsBZtMk0IMOKyBkA40jeg5cW1pkrhaVHvFIOkOGidW
V+r9nIXpW9S7wA1NtH5FcWpiAKGhVTXO6H8xUxZbft4EFlhlSPAilVq80vnqO5QDZnImoMaFMbXC
l9IEw16TV/FMYEKLi18WhAqjlQ40eGXU7ac63XZFDcyqfsvVTHnUZNkGBsd3Bk+BRKdbHc1D22Hr
0QR6p1xFh29RdHk7ao6OPfcwyqpbM/VZn3xOMY9kMoJvab/R4HVMhaE8YzS5LH11pynkqPEMklPI
2LVm3qdTaS/mmAFuwaWXAvxSBl5KkwCciaX6xTwNnIaLE2t8BF1NDlTsFfHYt9pEAgO1DVlG3b4R
Kg1Ldf9KhQIiWLDKeYsyZFbvJ7w8WK3fG6GLHGwUl12WALQdb3SFTTt4i6cuazXs9NacRdlw5Jpo
HF9NbOwUD039b5t9suFd3MT5pVaVyxTebZY9uxVN5Ub4+/KVEfl05UeDg8hqL9zJRtPw49OF1JVN
3dR1cN4NrmMfVjWzjs0pVnfT+yqXfb8VIM5KliYNuUiEug45V8rBcWg7wsKXX8Z1BhQhW7wYCRGf
wjJUIQACNp0tOT5PS6YKM3aq0ZJI0/TEz7eYla1xAL1SPSqv7JFeJH+LbXtXjP0vSgXZ640e/Wl6
+kEAWd+RBKOT+E6TzddocnOdNs9HKWY0xZ61rWwABA8ObCFBSA7zVvtDW2ENIS4V2i888bFCxFj3
5K1QAC38ihrBOg2qnv6UPLmywUmTF2e6e4iNFyCXpVZ5EaAFevTLA8puWekDai0c8fxV8R6OJJYt
RRfSo7Ne2zzhBKhzZ45saeVEgY8L4Do/vJJi6NWbi9V0IVywSdwK87QluW9yG12mWlatGo0lAZ7x
3yuRtBAhCAiyxESeXdXm37mw46rdRDBnbs6fTfF4c4tHhs6sMLt8TyVmBYrk8naeoWF58yLj/7Z2
+8/5quGSkcdIUiFHYRH3ZTltlj49pf3O3tDKuTW/9G1SooIB/gWRwUgoC8jrOQO7J4egbnophaXd
siE++ccAt1Pjw9UAVgPTsYKx5K7bLA9fgMSjtNCIfTSpUY6xc7mo68lR7YIn5jcBnEiAqg4hVcKQ
gvAIolIUN8zJ8/QZmfNOvetx0cO/R7wv1qOfDDpdGdgcqTPzZ9OaMmdZwm8WrOTyoUxeTtY73wZ7
iCKy7G7OdNwWLIG9LTdLss7K9ofAj4nYQoryshAgsRjMxNyvzDqyd4J9D9+sSxTM8CMPrju2dH/4
2rlc+PrnttZVGuNqAGifI9XDACWUixtycpuJh4XoP+b2U0kH3ZRaVUhawLudb8XvjnPbQhpzhRSX
gwy4nLSeDL2/RZD2/X1tLxCfeKteGU+NvE+6hruS73JzRZ4urH6zlcsJ8wYqbxKZVDVfbGG/vNW4
e4moRm0pz8YP/LB1X4BnJ1qptBAHIcuObH/vP3za88sHMAyF3O/Kcl6/diH3+PCckQ3qIZ6iKepB
zOJwUvsfQ0vWDKiS0nQ+Cuw238W6dBXBbBEU9gkmTyqkKVwtyJMU71ZsvYLx3MAIDieZY8avhLcL
zxKAPZN1a9e8nJLaj2eeaKH0EaZs2Y9l9JBlnW584YfL5vJHZP5HAl9KuiyGRGmCaXpvTOQplMMD
zrvP6AgMMl9O0hUU8Ut/JkOsVQZsONRAP4MvZBYV8xVLfc+Deiw8gRY/V7/BXec5oEcx5lgpiePi
qVk3gLw5AP2NuYo1WlQkKgar/9fhTspjHjiKtUND/Ds7W9EoZqRYu1D6IoqPkCzgF1i/hgbpif3t
XrWqb7gh9pvrXbcIuTCmnwsWpyeUomoIvu8HcotAl1MA4MMKTTHwVl9pJvNeMTy97r/jsB+9Z/JY
cvRNmJMoCEsYblgDfiht/X5wxIDQEy+RTZWnkfCseK9jMCueR7z7qJI44nt1xHDhbS0SUwyUh5dq
HnMJudR36pwArmcVDYlE85+LdBkHeSXS5YshJM2R4W70IHMhmlWi58hq0P5Kx/75ce5GJY3R6fy3
d41x5eNRrAWRv14A7OorC4tR/1RRpXzn5UIoGjBkF/Ju2Q0jHv5ltaiQJQH2rFtW3WgeJTtd8jcq
wSF7hqz5xljahKOqSykXgCBV9LX3hLkRdHv47HAMs/+qU4qpl3hn0OMkaSq1fhEOOXo3H8sn8LG3
lz6DTb0UYjiPYJOUsJBN2aafkqjszUvYZLgW7BETcjfHXgiDgGKx+iFqaWzRlV5ibjMmmhDa1jFd
WFZQ5vBaaQEnbqgcdf31aPjSk/JKCYfhV2kQA+Gu2i+GxbZwPrslEmvaWgscU3ANx4T6SVdvLPmD
MkqpxrIgARbRiWlRcb2sEeshXFt7dNhBTMWt+/rqvcg8k4Mwnr9ZbAk9Uz0AkJJ2OemV3E5/DZtW
liiOQ0a+EZe/GoSd3489FkFPaWs5F58YyY7Dfsazd/El9MTdIaxqOwhBAjCvajehHT668V5Bsj5+
1MfFNjISGJvZBx7LhmxODaUW8FOm9FuqSWN3Bl3n6v3+LQHa+nsbnhcnckT3L9kfmt6yLK0LU6HF
M+NYdsOeMVuzaZfB6FPdWM3R9egYt3VyfpxEMUqI3trh7zejHlbi3s8bna0bzE2SQ6JUvgTt7dcT
aqjo6+w0YaPexYcqFYzz4vdD5uxxW7aqtYws8vpLqim53pNScDLvdf2uS8/ebJx8On9tMMqZOfq0
TgDposBqa8kT+hNeF0MqlMabsV1nu3v3jIbJblL3ByyJaJ3jYj6H787v097gWrZTUWKxIovSavp4
/pOa1xcrtQIP0nGNY7T1qzw76Vy2jqPWQRnUSWCIbpgjpwbK4J6sBs8U2qkN/0eT3BOMAKC1n8n8
FIz78FjMyCeH77Dk2d+HWQl7B/IdFC0FCiqLyd+gwTtPggmkmeRV1q6VHaqdH3RuK6Rg8CyNAcp2
0CTohCwNO5Z5+In9vY3UhXo8VLk+xQ8Kus7iNXLYxCFl2PNxHOw5yAKmoBo7NEq21SqucnkMTATM
ZA04XFRIf3KEN/UfddDtwIxWJqwTUY4aizf/AKUkGSQYXk4w5LFzy+VtPgof3+9dM0Xo29nXYH5w
mfAWAgqp0EtSQ4mYHzssSjTkFJXKF5Cmn6J3mOr9JpvMjn4pB3TQimWi+sAQgGENDEsQlKFf6+zS
mD9cQoHhS49rm8PrrG0AneP/1TIsEF+rjtfajKntD9eQ/3RppNKahaKbdr46hsbQt+p6sOqr7090
5d6yNWjGUsVYZ6c5OlLLXo0LclMkYK7uL9d3QVI2Px5+fz2s1HZ4fkZDToxhkazjFlSgmYBjZ3fM
GsYouFnpnEEZYOw3xQAwQsupiq3Ula/VuqjmImVEdsT6iLjRg8dTx89d5MUB6sn/0Y46CaakaL+F
S7jRtGpFFQmo8LZxFaNA7sWkhOX7NWR2FAM4X7i/m/N9/YhDR3kePQal1tt/7x5+bhQtU0f5XAyw
1qOy3Vn/RY6L9YOOVaBgMtQFLgpA1fkxGWaBMw8+2F/CqXthPwh9HrbphxPcJE2v0K0rbxPb0CKL
W9/khFISH+AizTXfeQhibxjrewP+xg2S+A8aB10NJw6ncSb/IZEyeiTP4oEKKxFJap4L6sVvwfRZ
1vhuOpFNhlj7uzi6V69U2jRhiWuFHc63KTRjFyE9n4yU8BEWeM0MjZTVbmU2y/DtWN4DWn6z2VIa
ce8aTVsPcJNAaN2qRZLiTqltH3V8FCT+vk9py+f2jkQJI/ARVQmsACDiZcvGf4VrsC2LRnBzZXOF
xnZn7wS2v4/FcZ1TY/I93G9sb3JOT+rImwbZ4qDCv2JK8XqAQVhlTBootrtUIOvf5P6CM8iF9B4g
9qhkE8Z5pLSjTRRcbOdXGDIYUQnXhCL+RHxArOlttlPgPSy2Jm6Fb0F09CuiRPvCjpXM4kThJ5xm
Mn1+8lXzZtM5SMgQMHbaMT/S4ez2OmCJtIjWnKD1A9i15otvdsS4VemseHwl3LeCFMfCSPzyi779
OC7ZXPOKmKpNu5dF0uklbu7lAUyS4bZZi7Bv1xakcD3ON0IJNb6VMkQnCAOsBMhAe70NLU4dH4Qv
MKN9KwK6IcDrqZtk7c/VODiFfQ0mmvGysGHZ23ues2aCUYo0cckqP5r+tlMy3bglyUL08XgPxkbx
j9c8Tk5mv/kNgaoMeFpr4k3VA/amdXo+AnaLkcyyr1uWJexEFD0yzxipB7XI6fjSP5WQmaOqIWCm
+PkQbriSkgpwB229fKZFBXmQiSHr29yfXo50KxqcqnGWp/fKWqSAXkoZNBxza1bp4mBWX+JBv8v+
ghqPSZ9pY2/gyS+d3G9iDZvcdJZ9rCncBRJplAEX8e/y82xOsbzqLfj7rU9/En03vii4D2iYjghk
NDLFCqCLsuFr7910Zq5OFgtiUpu9lGhmKIxZEPQ/O3bACfw+dj73q27NUOX7B0RMbquJOOB9vD7I
Q5iievHkI4/SBrKGTVf0sOe8JR/24e+m9CuKC+DDt1a1a9Tdtvg/8OY94zxWFlryNKgqCORDVY7a
hz9ppkIrC6sbZV8zf+DHYOfI7jldvWwy+8jIGpclzQpBZPCdEvfON4IsYXwi+OBPOINta+woRZFn
Zj1r5vAlBzbJJhgtawk97/nLOxkxReJfdIqm0FDf4Z9ZaVQHyxSSyPrvSHq/IzHMDzYVa4CgpLaf
RcnBlshqAUADN3SVusKURCeH/JhvNhJoN7jknvGjK2qe+5LnksIS2QSgvN4tCvjlUQyIE40sqZUE
31Xl9As4eIbQRNnn+ggKosVhxDKQ7MNGOCBap4VpVgMG9nLaA5asjGAPtM6YD857sVG9HI3GUdl8
wfvgnuo2UjHAKwLk0prS5cpTiLiOjpqTGvD21P7skDsf49cb8lMWq1Pk2ltM6DLbDXs7Zh+b/5fQ
fU9LnIXamNj+g7hZzmWD5tSuIOsPPJlECG1K4sAFpaCvpOS3XeGkwOnNbJpbfvaeFPl33j8H+Qre
ZBMGVtdMK4tZusVkNZepl8zmTjH3Lo8C9KDkRLCAvYq7OfSdOaTbgt24VHHP2j5yte8CcydVN/Gi
T38y+deVTMirYJ8Ms2R2JYiYXUDi/sMH9HSpTYoV0oOKe8t6lojQLoVdjJC5Xfh+1cI3B5wrLZ30
tc+u0OeBhozxN5WE3QOsd5hgMpWE6yIt1yorhqJX1Kwfv6vKY76k0sDxBKpE2pq3Ti6pu/vrkMTt
mjwNuvDI7en5IzydA2Ue+IXg8Z9DA0BQLskQWKZNsZxrKhU7gt+UQLikrnmHAkXQiEx/AvmxEpAA
slByDEwmoTff1lYzgKIISQ+Hj7Ba2llrMUpJlhzZKBxquLZArnkheVYZZ63Jx+bb1g68IwT/NCWh
lE2cXBQJ05c7GUL9jF/298jdp+nWpUT2h0mbcHnBnEPr84i2pbvB5qklUbLBi0jkMa1cBqh10Kbw
nCTW7FFhme5Sy7Oe8SH9j6XC+nVhAPDSMP1L9CjT4bfc2VdodqKBzBiz95RZirKXnkdPLe0TCcVw
ic7Gm0KmbNtutXye/HNCoeRs7suBn5rV/6wdMZCxsJ6oYodG19kVqM+ChwHtywC4sU0R4Re31GNL
ut3683x5HESWhBiSM1YsOkGtfMFuXGucXlouZc4WiEdKej3V4WKmdBRXcHm27MKR5hwFFzGHHISO
cUM7xOcPEXroftvCw7UFs8kjnVn2K5FgD1T+3pBNOOojNP1DA6SBLYe/CsP1JlfmWtW3A95Gz9ue
kYJXM5adbM+Zin2S9vb6YukPEnk8uXJUSRkkK176+oDxMH40QGqdDKqNYlFmurGko4D3CHcdzenH
YDdbj3lVshaLFoyEZf+NEjHaEuANduLKTX4DgGLvnA6DDHc8xSc4TkFmnE3N+uf50Pqxr787U2GO
snp+SaBKLYjTdt5lmbivMuEEXJczGTiAWBXSTTBGP9/sqggSZK1xyBMLRP3w++iZG1PNBdUgCZ70
s1wQJzYTxomcvBNLFAAGJ6T7RFVq3v8wKb1cArp0N9GS5wvsS33n12qfsMGS1oqv9Hxk+aJEHz/f
J7TSz5qSFv9N7UwrQrvVVYnFYZIhKV5eV//qgMiXqSEETjlZV96bC/nfyt/qfDE8qb/sIl6bJ+k4
gQFmO64BMZ1efp0omZ0/7+JfugpfVoFdP5XCC3hdSsqdaexHhtDlPvaZMHJJoSW/NIwdTABIgu+k
eiR9IUbSCLG88va/FNNKJeU5jVQjkXu4v24p9OehiEzosbF2jylNQqQOLP5W/HwnlhcW2Cj4s95A
v7F/0D6u7ZOdsKGlpiyB+68NUr+6N+sRjQSHCgSI42c2XgIEx2KVz/Vo9vrhuouqMFCbFgdkBhtd
EeTnaxBbiVmWCjR2a2qD5Qy5tRjvF+lOlTa5yM8c2eqYeVPa02VxalgqUJTVvNKIGYjoUWwq54Bu
brJvjlfBcI9gaLcH5zvUfTCLT418jJtps44j7IITU1YVAdi3vLzNmgGayuNaISyOx2HEZxDspdeU
QwQpb+F5qvl4FhW7vyEcNhHMKpqph97XQPUzKQveE98CpanqhRJdOfu7u90e4fC4yNHd5lcWjdVW
XKsItiVWUB4H38rcHBTIO15ur8gRMn9nxZDXdRUa/ShnfZbH+TfChlPO0JHBuW279LZrmRjscuwC
BLLiwiNtGEKMtbKtrnpR8+lJxfPqJTjws7mRgPdohTPJS3LLVTFh84FNclf6Hy7IJpOz4p6wcFHx
D5lTdbANujFTix7RL2Mj6otLUfEmGy2Lyi5/aUIYP6tLTKxDVfxhbn7av3ryxNisUOBHB3r1eQsD
g4TyIvwvoJf3fIYi0o8SKkQsjjt6VOsy1WxrL2II69cY9+dshKqnWOdEuRHJmZAV/uEv93WZ8RXP
lFqStYUzPROF0KWS8YCIQPSyd6OjhoDt6hV4MzqxzIv24AOXzX6n+cmhRX10Sggf1GT075Rcoayu
/qCYknSDqS1dR6awUyw1b4DKT3jTvZgycVGwsVl4ZCa6LyAYGzjQD7bNYMJHLFbDE0yU3QnX6Ylx
+V7llBTZagkmcaNt+oo60ilYkD6my+cMv0TOZ1Yn9ln3hnTXhW6STBhZvzARD5YR22cJuAGjeqLH
HS492H4qDYdkcMb8h0MvJUuh4arg7lgWTpKbxXgCCzdcewmfE6Q+aChNDTQRuJRLXGYgxWvCD2u5
aB8MqKOCFyBMRFbqpgOm5v6kSKtAbk6DGWk8y97uAqm6QxLjrY6DjA74IocxK1OWL1wbhh7Mf7IO
rRHMirmg2BLjAyF1rQFnfaFVKAkbRBWKXYGIBeNB7AlieDQvmlrf8bbYjBFKEBg+3JEBIm4d3shi
5/IWNaJ0GtsEsfR0iYU6r6vvAYxDk4qwRbscBBKZWApuwBybjYyEXKcA98ZsBuDs1rpvUQOgq9vz
wbXcvPhHJJDUWISEBimRepJFy5wDkxyj7zroeI3eh2dgBZPcRI4RGwhNbNwjG90EJqthU5YtuGPD
xU6mkEz12r3YoWCMt4Fkfxex/+GGlGsXUPiY+c5ATfUH4LFJrPyrJWwhv8TkvsualVXwY69ML7mx
bwZKcUO5UL3un9wccjQ/cJQxuvDj92N4TxFKxcsaYJvgLp1V3PBkdHZc2ltGluRHpJDTPzZQ/tU1
g2TqtuMDC5kPuLmJQcxesc4LcWsPYgTWtRxksFIeEOShrw7NQ5W1Zo2UnTeqT+eHZXm2n7tB8tO8
J/sIZC3+U8UInt4Z0MwxL2bw/1GXCnjyTwz82Z/QXiENXNNSPEA9iGvjqAmTUgyk5gVvd63DpIx2
MbPG1385GYqcbcUD7wo3UmtPSghe7iwP6HLnmySvYpbgwo8/XujKCX0T9MvKG/ngbzHiIipnl80g
MFy2cAJYisOX63cs+EVkbRi8Wbvsik4nWvPwgUwv7AwWmc3bNOyarkkis84EFQA/tmfCrQz8XaCe
mMAW8KSlupPcXYMglEqfP7EUH755Hd8AP7O67E5Ocm/z+0epekVeLVZ/2Mksp2X9X4jauLa4bcfS
E1VIa6TAAVCJ4NtmstmRGbuscSQJycLCC/aBXRh2OMqpTs5wpAeKqxCosL3dQUiC7ZOBsaN+l56N
1RYHmoTdBnFHRHZUPlKUyE8DPszvmYURzOtSp9ms/TLoEoHKaiszCh0wZGMRT6F0DsMCmPKrsILK
ACFKlPaHh5xo4XaI6jYnrA9w8lLciTmFwRlcLlAHlOaAnYFbovCsD8nXy8X3L9wPGcJg9iXKaIdl
SZT3a/rC0fkrSCQF/Vst/eOTyIJ+HBPbo3SSLmC63xwXKkKQzhOEOR+R2TcsGbXUu5FZ/aLu/mPm
xV+3LuZ5TSr28eeJ1IGHFAN3POUYs5hMpHbMbkWmDpq16XEqnNxXAI2tjxAPCp0SBw0BE6MiDAeb
2AvU8HStUE3OvWtANhqLJ5lzXHmSYZGbjfDtp5iN1m30qBdH0UF4hkKnkiMSHN89StSStYmhfeTY
ZxJjg5Ubj6S9qFiFJKB0qrzWuuU44sbIYzwAGqjai4e6c7y2L9lC41UTTOv0mB8Isyp6iNVm3Bbc
u0K780qGylct0I8WCdoEseBXLUuOsv1rexcvXYXD6RtH0eJ6MXyfM0uYDojkOKK2lUWTDcVDuam3
nXZ4uIi26Ww7CrbyEWadQHOLORWOvA0hJwJxV+tJ0Owg91+7KXlqb3/AUKIfenEx8wYr8YRqzHhX
nxBldXLSBN/Zvaej+sl/ATtmGJru23IX2T9Hlt6zwemzNnxHp88sueiEtA5QtbbmVzw296yl2bGJ
xgKnmCt/5zzBfUkihjCGQb4tJ8jmdMl61JF8E79TabukKJ0Ah0Rf2LMzS7xt3bzEP7PL/jBHV0EO
MXn2FiYK7HEUlB0D9kfBjnsQi6T9yzeRt2CrFm+wrK5VoqskVp1CD4/28mJ2EpMRabtGSbdpPgZ4
a7y0s8gaKiEzZoAo5O0Qa6hVJ293w87AbInkUGVYX0qqkrCVVo/pSXPQVGU1hf2WGTlwQFB5NPXB
gM/bs1mbGcFdI2yptrnUNTCKfVDrk0B+9GepUl46SL0yiLcrFhSoqGh83b+j5g7Kq7eVRaNTZibi
oQb5g91RdtYf8uwK3u1kBBr+HcyzLwroYy6efLEyYkJG6kzJuiLLvbXfdy8NW3zh+3GShbx89bci
E5sa2oyj0rJrkle1Yn28/dpfxl8Kud2mUdVEYP0/EWtWRSDuBcF4YQ2Vf9ICKjkoLYjVZ7XyLL2W
dvVwvNvNWbn0ZR2IxkUjkjEBbXyUabGPXSXr74mzO0ARaZ2ulDUyZsj+7u5+XpF9jQjziICUlyyb
khmQaCjVFsqiuzh0R77+khJ0S5sjLByqau03eBzIcf3alIZZ/B7reILDJDRayPvQam+rMLtKH0Cd
JTWZ1vSsj6KUIgFFS0ZI/Ua2IAx4mWB3L9yxx9ONuA4P49k+6ZCMqVixi1BlU5ztCygTuiYeLbAU
dxclyI0E+q2kqyaF1/pDMXq7ssfii/pAf0LFrFnWFIHEXbTiJyE1uHyoeoDoz7yg5ug7IgQCr5e/
Ox2Ij5DRfVpVFlgScwqylaX4ffAMLNnXTP0D7fufjk6ynPclt7BplqEOOfgvUK11OY+PnOLcCfb2
yS0nn9AWh693FhfQ4SlNOB0Q+IDdTFtpgS79vQkWn7xcyRqsjEYSMJyC/2oJaGcQYYsDtWROjnch
hNn/bIXV7/MyAHo42QTg2z0yWnjne7CfDlJtyRyYeN2eaq8C7p2T+F9mfTDA2uFy+bVZFXLHY7M1
T5x+lv/hLHogePQ2bFMHtDrelj400XYYqnI4qVl1qSKCK4VSgmNN+60UH+dGvWP6g+FoFp9yq2rC
RoNm5NicZy9kYYM2k+nCyp94Lf7A1ie51mov5ntUJ8dYN1+YexJE4hoBcveEX1Ox/Y6CRkr0vWQG
kOVptDSs1n13OmX99a3fZL7c9guXHnG3A5Bvl2Vj8xmjK/Z+zKvR4KwnnoOby38GuGGyIGWgAcB9
jbf1Js0yJEWOMeiw+Y6KJN/4RdrY8hF/X5117JGUR3KvzH+8SdjjBn404MffujbaCIm97SYKXpLs
gAgpuEaJCH78wq2mxQKdWIjiXglS0A1bHvIdqm6InfGYTsABL0fw41Z2mxVmBTtgP/mYf4AqOA3F
YCKyoLG06ZUmBrvEcYB0ii0aERUgZbIPiJO8Fj0z076yIH2ptmZ5n+FedVX++WJBfipJw/2JCq62
bnJcHxrqf5sqBWftce89RMMZMC0uHtNNOQjOqHn7BjT01uUEFB3AiV6i+dnXkwa5QGCaDUIE44Rh
E2iRhCmOw8XmSEDZe/58PAW4CDTUlswNcwwlqIH3Z8xkFNp2ZuOkATovxUnfD9pliLXAa2bAmIUl
U0sO0R/55ciOtGKM6qA4Kw4SqEj/9XlJBqDVHqzWYhjBzxKwyqE2KmAEBpqcQS7od8+eUuzquYn2
B8w6GOLfeMOQhDjn1vyJHfbKW9CfyJYdkHhNutB9QeIq2khULwZJUkLLKSWcSlnOmqmZhkvty62R
qAuRNQnQwB78HfOrjNL4N6ooj+ttzKInAaSUrhH/4EmNGwUxC6wInLp/Cz46Br7R9cPUThjrnCVX
evwMgtiE3Yf0QETU/+fIsLtrAciu8YKl065ho6BMVl36xGyXNtQzMM1Fsd8dnsFG0deZlcFiWQfW
w4YPUCCOYNs+23U7QE7SyQmnYMWNK6X5Wn/RMUzvs4ZEM2RKmwA37FIpGkp3nrz4iSGc38t2vw75
U49nPC8GaZvcnnIawnlN7z9RTjPiXN9ydVMMAO7/UTTEq/2bYwBwIcxIEwjG4TcvNVa7c9Ok0Cpo
vDvg0n2piQHVJeqEXwpVFyBCEL32JaQd1d+HQHhC/T+KB87JNf2WQi27XMq8qE4PnQ5F6kMRiLhB
/Dv/WRu9R8ZZMIGgrSAYwmNvximAd3yu/491gGJOs6NjeWzRix+lmfYgI+QqV2BgXYvwokGmrvMK
5myjJyF8ve7wL8CAPBU6kJqaGto9M4oJ4t/2ALdOMbjQy/KZw+BJH7k+ACeumTnAnGrosyI0fV1V
41I/WGS5CD5eIiPfL729rrS6v774RDpCcshsPTVs3PGoa0VHzzO4kLjQvHlBt8wOZxCTY7XjD3Uf
AiYdTMr5ywr9UdABJaSeF3DBSkmyqBkqtX1UMpR6GqBA7ajLfY5uo0XA26d/kNLE7Cm5Ssa/BRbi
3pjBu39VC07ddMdUlcXn5MW4mwXpx3Kf0tzg7kqWH6DhIsbfrnfgSCoVuEb78pjlaf9OsBk60WUq
7Iim4VRYtYyQXq3TMvME+G5jOwWImvLFoOyQAZd6BTmQK5/618v6B3us/pHQDmec3ak+6U6tw4hT
SeFYa5WG85fUIXFSucUIavNv0FLd+Zc9I+KSvRqSLXZcU5zHYAcTTV/iO8/YxM+A13AQuLX3SxJQ
COwuO8i2n2+PffpF8HP5M5gAWjbwDNV5Y5ElhkD+0KudGI9hpJkit6YE4AVdlZTI/pnDDOkGtCN4
0vRViT4sha4G7K5QlFe6okT40miEZV91HbqH6wGyZ1HZL/1zdzv9fJ/qcg0jmULqy9dtNlxpWjCW
DKhJQyKbjOj8EkhPoJq5gh0rigVbjUd2I5isdWWHcs+QCi6/LhqC9IrOYKTlasNGD72HX8ZYYvrw
519PhM8jPQnoZv5yDjV036LvkDwdrIxcI+VdBFfQBilDgKNtk6J0T0FCjl2VoOvXzlLFEeRs7lPc
FG/mSnxDuBl4raw4G8GoVLVvgwvFfjt5UGQzi+i7hApjS+SPb1R3FLyUFee5px0ZgnC7vKePi6uy
g2gM+S87qlkji5KTo8Ez5k/Ywmt6dvU6sbhbGdkhWkUjKE6CtPH0zd34Wu/iEmFFqBBXfFPlw6uz
NqN3aWcjyvL/+ezPmAlfGKmmxCL82Q491zHAGg4mqnQNoIrB1307JMxQfJ0bhzvtPtTdmHv7siSw
mzSkp8uRXf/f/n/SnhkFplQcSuIimHrC3/f9Jhv1R0Pwpj7HLHKbkB3j3JYIyZOXksmhZ0w+DQb2
l2vV5uWU3FdqxxlQYoGvdpRCYTX9H257e3XE7QfKdcEJTDZqsLxscqlDm6Np1Gw9eaUx/vxxGw/1
G0khEa/neQuLO+IUv2PIypHqPqGNMnaHuYb1MTbdOPrXxCuo5Sn2lZS1y/o2KvIhqi6akbnxmqgu
M8T5hnYqtu162BCjLBjxRlupHkhFBg8fyioqbOrBz2PgRXPBf8GLQ5hnxG+CrC+rUlrodhcRznCT
SbLrlB8ErLvk3yr2oj4EYaUbQTcMdngkWLSUPcTfH1T0BH6bhyHYZ4lnW2O9WI760Xb6UVXsAGYM
tfw++Ujz9YV5Vkepv2LQxRRUNrX6cEYiAvI5cUVyszb0buHm6mY3BGIFilh/ElscU+NgrWv18dg6
0FZtwgCNVcuMhch8JCtfk77v1mrOPRetl3AKDZUkdZEjVzN07yrmyaUnK6wCRFW4jWSpDLwxgNfZ
/9jaGDIk2JJC6HWq6iF8IVu3ODdIm/K4+nYlHwMEYxMSRUJR5aymH4EjMduCqj779kjif0PlyZm7
xljeumhbwxYsBVn9xjfNhApzAuLIlBxo9L1CM0trz6w8wPsVcHr19FdLotpPX2NcNvjG1yMVT1Yf
05XJd0G8McToaiud7m/WFMC1IEbrfNcJawRTo6KNq1yk+C9DNrLFvWCqRQk1r0ZjuIi+p8lQNV8H
C19m4OOfM4ScLl24ZLhg/iCK+FTWiLquHY7jgYiGhqPdF0RsALZlTcDqPznRzkK0IUw+5yjc0RWo
iS+cRyewiTPo+zC5DWMJiL+hkcwRLN4s4X+FDuZhkbinwZNRhXtsG0oVy3nRK5OOsVlhW8Z3lNfS
ntu8mEM/SQM2YrW8nUNd1LqmyhR4Qb1y+7UkOCCcZ8KYbXh7VKZrtX7SGBM2XvUD9CiKKv72jWJL
sE8B9/YDF6Hr5Fb05FZwCI5+kaUtawv4yfcAcYGuQcPG84I0Dz1WOVVd3W7z7OIjxVSUCmp2upCR
tJdFMMrvgvz1g5N0zq9t/VyliIZjURDeMi9NYjSjfL8nG8l9qA/cGlz02SnAltAgfilDb6zlad0h
62O7cytPTGfabWZIO4k8Ou8HXxdl84QBq61bvN/hZn6SvY49DYLT1NyKaMMg8F/N9qO22FHrPZWY
T1t32VWLoIYy3LtJpaQy6vswb96ySIX//lU2Vu3adFQA6owT8sucsVc+4xRsSDOnQNMGdGjkfFSB
VTfOKfpEqrJbTqnIQs98cQn936dmUAUjoo+nW10WUmBAYOvxHvfIy9xzgK8nss1QYmUcDj/bkqn/
/LCOnhQKd6B6NkLubASj5CdyMw2PSUjLpyxnUwHTXh6tZhEtdgEdm/mFvIsMe/6QCJK+GxcfITRU
XQCnRFybWbnQJiwMMZvmj6Xyhlz35/c4Q/gZSj8zRNYdx0pyXWIgdmkVMzgJrZrnsb/HvcN4vkV6
YvpWbMBkKGcWznQunM6wIQoj5QSqe+L8cGg5rRdJtfueJTJBcVvBiblX/8IxnkRK2NqM4g/b5TeS
bBzBuAUesR3bn8oQ3C6Eh2fIwdeeqlI2W1PUR7y2JsxCxYfX2wpXIIr9NpRLxuubHJh4UyfXhtgn
34pJ6LJzlE7vjwdN54dae1eEewZVWbJ/2nLUd8gOznzDtkuf0bc3ZDUdT2XB3/k4K6/dKGzliIdh
lpfSjbio1V42CG9YNDlC6hN9dzwkEqETsVX7Qy/nKGhkKVdJbiKbcbdoEycrLTQsrhbKfrfnNCcS
sYiR6wo//eWse6po0u0ukC0kmkHyRftH4ahl+pb20uNLpoq72/dBrrTBVGyMek4c9z5UwAFyBHq5
vruqJKnMagrFvznEptdoFRmkdeqFnH4b5xhLxQR2sLGRl+TrZgYGojnMArZuhmZYbvKGPk5ExVHB
KoZtCKi+bYdVBacp3oCOLGjCdfJijJdbesWQMqPzSCDh6uciaHLjzZKhKr0wDV5lmf5j+u095VN2
B1zQlmdLkTS3MaA/0PUbVH/0Vnp0znOAF01ahlOywVfhkTB0zgfUhrbT3cp+IBR3XIz+IQEtbXty
xwc29/sc93+m+1PZ7HAj5EQAy8BhTFIT7GVCMzF9Fdd5/+3j96V03oR/J7oerxkcPB1i9wcUZbvF
zHxqMLOplxpCpH+A7Yz6+sUAn+hTkDwqFANoZe5jLHsLjHVS3Tj1WuwI4HO6RyN8RjLAo7pveAP3
KgbxZZ8PuRvZDBJDPJrbBCGSqWrEX22zxyc7uqThHjC4ceKlcb2Kl6ePZfA/Yi2rB3lkHN/Ct94x
yZx+3e78I+SahwBnvfjtEnp1up3S68m5PvhT8X7pJ7kxKL/Yh1QOIMGh0Sna6m5D9F8RMAapEkX0
PtTgxPG5+0AhDQXFYc4qk4bFfwJ/e2xhleK0m/d1YkfjLu7qME+aMzAmY6o8LfZMiWWUlSM0C6hY
BOuEbudNPKdRIaq6aYnGEYYcDnMHV/ZPO4lt8T5yvlarGZfe1bVaxKME7MXI1oqCHDFg6umAs9Va
9V4PZT+3kdpSJ9KnEzUz6FFMg5FaSCvIv2KgbnusvJZ8T7If7UNK6egs0mTWLWhki3qbcFQV9XvL
286mEXvAORsvrBZLsVHJJLQviaxr3TXsSX1SqFCePPDRDpllg/qD/zklN/ttH5f3rPdT8h97dOiJ
pkw5RqKQtQNv+LcZ4R2KJ9RYJnRqilpJ4rC3BybiJu9eRLKWwkU+q3IXdmWaDiW5Du6xjFJBUi+a
r25UUUYLrrqLlg+X29oddjmx16W8gqKSk/nGeJdGEag15yJva8zbS/sSLt4GqZlrogKcuHVONrTb
Asiz7RmOrGqjr4fgwwo4DG2gb3EZoSpXAcecAlO+41fS9q9i6t7sQzHxdy7kf1BxmjHkaB4hrGHD
LoYk0j3rMysYVVqOyVchZklOwnc+UvZp90qF6ncvwngusPMBTbL2UUhP6yP/vIihucOcYqMiGG9p
GDya+Q5ta2R+nZLFBwhOlTarMVCJrzUREeCsdXT90qmVRt7jM5QJmrrIPM9u/xnXvIBy78zCVRyW
swlw9T2nIjSHPEH1lPW1QeukK1dT8yDou1lz+okchCPqsajY3TEQJ7ned0umWNKL8uDTlNgT/SGR
YCZQcsGf1mCCaITlgCVKHLTO/tMtMsBNxOjYzLvQQbtmEozgcXG4lGimR5QjiZut1zjSj2wO/jjh
RjGMUWpT3V1KxXdf44VgI9+Jqat1AwdRy937jV+2osDKli0LELU9N6taify13+yGBiZ6WmyYnrsN
meuzohXd6IWCXHo5Y90YbVLLDcvXyFpY+BW8MHb9FAG8um5kEfl4fqL69+hZQgjcx+/DnAb2y/L7
cNOipqIDgmHRru06CWKxR8iH2c9hDoswXWRjxLQElZCZSwRxGCMV53tTYFNOAIJ6E5GbK83quFKK
aAul+wDIWtJeLmsHY0YQuw8bjH+aQ6vgkZCZGc8YplDrNg+v5XLywmUBbuVI1opRX/2YtHdkfZLe
nRsQa/TwcU9vfPE10ce/E45KrqEKxj0uYc8mxhr+ETDWMpMxoyMxRzSfT6/FLZ4Cr2E2pY0LteIj
03cZWCh1OgEQSnArPGJNynLv/3PZS42Usl18bmOwAyhKpqgRl6E9UhuhQiH+WA7Hy2fKXmJ/30xF
LOCVLM/gXfFiQtJaS4TyALf8amZPSxj5Fk+gqKX+gQA4PFP1juliaDQBKVhcHS6y7CAAaJ3JkU4i
Fzv2LBu2PH9YSZnusfx5JOP3VKg686fNrgCAoqXu1Vx0CgrY10HZ1U81je3V1unNhbpUgx2gMQvu
E4mc0khXR3RXBQt/ElALcEDqlXlHQ3IEpCyUb2ZZTHf+4+UMpJJvO8q/NmeT0GtPpwWmCEiOJ4Ov
EisPp8O8Jjqlvhq5i/+6aSsIJ0jjkHaSyLs1Sts1FA2kjXTosN1pqNmjnTsLoCvUhbGVjlpAB66Y
geYySwq4yRFuPXAkLKYG97RbWXe8Q9nXNuHQx5gLwF76SSk6FerVx+XvUdRXyJTE9N9yOviXdeTb
NhdAWVfUCEHovyM8Fk9TVGfomJXH6i3plAApBwEqUYK2XWABMjza28K1HghsO4FThGqDdkpl4LbI
1qCRdgYoQlv6qUtpAPKX+VJ7eyANDmqylJvv+KVY/t4SD1qMWcdWEG+SO1f7klXMaRRhpej+Bamw
0IlWynJSa5SlElA0fHEdo9L6we3UB7I/tMzcrGEoXlgvPuyL0swIZcFHcnK1L39Ix2GMz5PiTGSe
No5+sZOJCuJE/PLoL568yUhk2vYHlfMYzknKHzxolbdLHlCMiGjdqN2pUS+U1nkjRKP2k0r1oEFl
abKlcdQwDK+Du5M5GbX1q5a0D42gOtY9Q+Ueov6dZejefRz3YOfSZs0qhaq+ORz5QupVou33kDbH
eu06V+9XTVfwE78gkXdNYbcv4fsKjqUgNSp3hKZF5SrJvADmpxxsb6x1a4CExeHYzqrfLmMwA+pv
+qR5rS9JYjDxKawgFY7rCb1jmfCYr+jzIWDc2e1lW8mtN4JLiaHD7j3cvcwEXkpIp/mZmWXDJHkx
jfv4pbO8CTJqYWJVEVdUAj2ea7jJA+nk8P6hewf910ER6gapGn+Ve7TYd7WvmGSTlp++cTlAUwQf
31gBzahy4PjLIacYd6te12XRbYLK7XrFyUbA/N/sWKdKBi00weDsYo5teQMrQ7XooeiOTeCKvb1W
VvygivDUrycqeHtZt/rg9+McDyV0vtcrdwWOnzWJM+mhfyqETr6UapqSD9Zo/g+wqkyim3hfcPzM
XWVKRxTdl3MubBIflovtGxuh2/5V2Zod/Um+qohefiRD6x+rZ7Pd6O0F4CdDaab31fNAFJKpQNLI
obRWuMpnI5UMPycrutmjjN5ApN1UCwbm+kOT4q2CTkbFRqbGmi6U6p88/pE7XjjyDox9uPBxIrqo
mUhjd6i+LuAxExzFlUDxQMJWnqwEjGtXa0QrKSpuFPLgKM62KiazUOaIIyOrkF2JQKaVDG9uzgwD
Hh2gEy+RpzyiaSjpNcu6m27z7+ecyt+zSn1wK0FniTP/Kvm2gCQ19P1BcCrqmciTDev0Nmb5ovGE
9/zZyDETIZf8WZU0Lm8+S5s/nOBY++QjPqxzY9FJjOzwuKJqxJG75XR7Duh3HlBVla+bXu9VKufM
Oq8vcBh2NOJJZWxQZV77hVmAd3gAVS23X2rI3zq4tdg9RlbBzXF5oR9eir8xuuOwEWCWGN1+4VYf
FVafXSbMdAkGqX//xOQnoU33D61z0ziBXshPBrsnnYFZuOx69hqBxIZvoFiDA+9UHYoHw123eN1j
5kBnhLfZ0p23K43tVD8hq3QPN1WKuxO6BvO5KRlksRK7Sinzv3br9xqTk0rvoPiz5HFIp78oQXP2
wahWyE2Ibr8pqiZxLpbVdm2vN2gKaWhIw4NSrWRW7f9Px6YTUpwLkm7T03X1mc2V1M/mbltNSp2V
GChQviyhwCm6oMFjcmfPznJVTMBueP2SH45fiv87fyLhA3w0kyG1H9jvODo32yx8G7qijNys4pra
K2lMIVhupws5jCqBmMihV3k9esn1jerH9hcgQqWfWBdP7Yz3mwqW2jolCfSz9okaJjPEUN4n+CFv
C5CMFLAR/TIzFyAh8SsibpmTeBaFx0H9wyKkEFK5IZvWaVzBByDkqbO50lscg4YmSgQU+fisysog
Q02qhyP/fFBoTTaHeLkTbogBYgEra2pnGG27rZjlQr7mshLaai5JznHj5dFKhl+jVYA3/XlQnVQG
CHnmD983ucWSFNutWctf0TvuOcGRwL970ZEt+rKexOAyjxR7Oh8RJEixoujrhm63j26A87HTrsQN
lgDlucmZVhjQYId02bBFqvd7Y/wcULuHc5YoOfj1kinw17YuR2TMxU8k/PeHZfnBPLFD33GRtrr0
ODW9XgOp+OLz2/P4qWCJhrg5m/pB/97Ne2VJxebm6CAxTEba6ltyA/sVuYzdMuycUV0gohjqlQBq
3jC/xY+hk72k5ZKR4QP5T5sA158KeaJ35d4qA8/1oh6pcwwlPHFPV9sOV47j0ZZKjzWG5d4TPLYh
Wn2ClKrwBGIsn3MpkF/3rvyARgFqhHNBLvtyDWSEte/inmOEwePBRaGcDXeD3BQ4klD7dclhHeaD
cPIypGKJWt+ALs0BJSX6fUKGm3j8Dd/b1qfcYTgfaY7DYRUVJAGdQJTUAdshgE6cETQsYMnG3rfz
s8/IyCdSK9RY41WVKBPmTMusw4nyRv29KWRBW4NTqBNwLHlcPKUM3HB5WQm+HvirW5a6UDt5Nt7L
NOIz64UVgq2VV1qvDGKuIItuO3th0xj9U4rngb9xZMwMgZ0ZilLezRKzmd6DxtZlXIHJghddNh6s
eKTIWykVnJs+h0ErnVkIZ6VZ7rtp+06f7Wh5byoUVNqicfTOMwOK5cWba2yCQR/OIRBWop8g1O8f
Y8t58BrcXAxRk2u2sUBHbgRWq/G7X7TlOF/sHileSCy6beno0K+n+BZWHtMogC+4upkMikr7Ed1r
OrDRwjCesgEoIw0MSWKhD6VFP/milHmebrCRghpsGfNgqQ7v4IN/4uMpdbojyeUsWttbn/Z3eoTc
EJ4MDYR0zUe/ubcu4zOPWgnPawHcNYXFmb8CSnHAFrd8r1ptm/rjShUPgEXylVsW7bJnlYSz8v7T
qYhSPNN8Ba67R3oDFODjQ4OViXAuF4kW3OmWvw7gZ5CXpRRkiuDQd22b0w6TED9XHZU4P1lkLiMY
JI2ifbDVt9MEtK06nbzR0r46rDTJwBQEomNse7FrsAPRapfVYO/a2C1rehU6+KR5+xFLtylrMzMa
YUV+cKuNffF3Aq2P/ksF3htXDbK23Pra2IqidEl0mZZ0gORfrddCeDD3CQ9RdQqtKoj2m44oIZCq
9/grOlwjReR6Pk+vjMK2Ccnn1ne+fX/ihbHSMBwm1COwjXsYUUQ4vLoEwMhD9YFZ48y/hHNJ4202
9hM5QgzL2WH1+8NnqjV2AewFtpGwSsnvkjFKuz7ZKBYSEUaA7+Swcx7aAUuDqi3Y+ibtk34+nd/e
v+WZg6loMWomwqpssbGLE89tgdXxm+cCtBMkax8dDf8x/8g1+NcByRLtArKEVCJO7kFL4mTdDFBe
Wqpg2hGiqcdknbRoniRkz58zjxtBAE0hXDvcYDPtI4PcO4JF4f7JhR3ADhCCMS2bLGHbj+FWGOaM
Z9ZC/Qd9+6seBf5gWNGo2QO52x4LIeJsuzTCXSSgW8zFcmgrP1PWmz8N9NsFcWS6ecoV0oIfDc0n
CitUcGbcg1/HRwz+qudtFEOZWdL+36UYWgXpqXUANIFrqc6jdPyRB8KmiUwwNJrUjDQoRmNWacUi
EAxRudj3gbd19U50vyrzoLNuEDZQtBT8NDQ0VWsIDuCNC240UQ7Fo/FnupPEBjLjCJpwWVwX31Nt
6zkKXUe8+p3wS/Y5NJBtrHnqnrdJHQwLS5Jpo/9WUkwmcHUNQhxrbkQNZekEWK7qjkMb8V3jo3hj
Ob6cMiu3N7YRM0zkiTCQxmXVuYi4qSH/QlHC5rPgNxeT55nBZILW+y+HomEgbBCVciE58Ms0Wcch
OZoRnl5yTEjMtUPakScE/HwrdykA3kzz54hT2ugU9oYa8hQ8OMkNDA6o2FnEiNs6SX1dVuorat5C
SLbdArNa9q2d0DQBkTAd8ZDXbWmlEQKSiY5ovLqif5aelp8nt0BA1ta8YGQyRy+UkkdYghO5jrWA
yMqBNaXE5LRfmgo1Hc06LppoMKHrOSPzrmMOROkkkq6SXhha5L70sgilDT/Yjq4+bkVokTVXR3+l
2UZ1O1bHOUH8GkXjYNn4RSpBaSv2fpnwggPdO5OkqaK3WNKKl4wj7FS2Th89ZBudb8ljNwaN3gZo
YF9gBXPqA2o0+r2H8j/JmS/6jSxmWHAgY1ixxY5uDn7GeKUP9DAzBhlLk3/ESC9TUv+cwQW6h1qO
aRHDH7GNBbRmP6vunjELRN/wwi6GvOzwJL0+paLuOYZ+a+KTcWHb38QiDY+jK6xj4rnxdzTKr9kE
7Jg/kIpC+LzbCTSrqaBhitrsqvxMmxGXOgqCoQwGYEjiBESeMmm5iG7SIzAAbnrrKBZC5xihaMuk
6B4wBs3K7OXJ/gKcm4hCGCpQxDiv+iCOQnLnmJR6ArwgTALrtn/myzOmviHc92m59jUP/vvA3vui
nHcw9FQzL2644lzlmDNnarKqV6wA0E2vAnflYr2DvZobRHJ6N5HV9i/FmStG2XMiyYeCjfe4wKkV
4CnJ7YMniq5rYzFXJ184H+kkA0LmwynznQJi4eZuLkWZKvIfYXsgGXjubvwAoi+TWng0ZjViFbHS
oEds8nrXuL1ErZA9c8pMLZxiKbBZJP9QW5mOKiy7WzyjbzjgEymUGJ3lyCkjaBj3i3f/a5hpVuKX
fFB0aoTNWXprk+6msZWBKKEai5SctxpTVXDVpU8OW6ZvpY2KxoXSVdCOya4mvAR/EIBehhwb6Cvd
aG6qzs31X+lPP/eZMWeW9CR6rwG2J260D/Dbjsfb0MA/ABxw5xPl4th/feXUV1jGYXRrMoIrdPte
z6YgBTIgK/ympoeRDY9IvVBwEnqxaf/Q8YnoIS3OzM4qQiZGPMQdey7Mj59Rr7dO6eg5z/BHKV4/
/m5WCIkSo9LMYmzYTIZOfv2TxCgvWswgMxE/Z6wHpgFQEjy/SoTod63asQcmGte3m1LBgXC7948i
as5h4yzfrMF/UEQsoTEQOkyIPf5pdtRrvg5NI7yzur2qbaeb5rXDf0mziuXiIlYfNuSFmCDSMX35
3jNpDW0maqf1FNtyPudmoBKzlt4AxvfhRYm4e6Xdy8+LQ247WtBPkMpt66tmBaBwQMLkMOSUoV0C
5RQJVUKjN0Go72jqOgeOAcy/fsbhzRygykjd9MH7q1BBWXwj2PrCOdEhKQgDkdJmfMS8OpIaBEQs
7BBT6dG/VWNp1W3HDCoCAn5lwGP53L5ZEld0BaO6Fm57Ow2wGGdr9SaAqqU5fC50Qnpq4rMnaeyF
KfuGZTC/9rGQCBmg28qhf8QfRyaVa92q0hpULhGdcFm3dhvGXDZLy4gPaTk9nYH2aEAGiHMOt+Gp
EOCHXWmahnafUjDssl4INjCOu5RrtlwD7ISK9oPr2TdCC74xjhY+SxNbyVpczbwMiX2k3tg+Us4i
34A6VvXKrPLbMipqfryAzyJ80/m9bG0wbiPNAPZvrKdGhyVa/ZmX2uaBlCJ6aznklfysps5TKcBE
W/oh2SwEM5bU10cOOtqGqMHwDHxVb7GXsQc5VpBMLDLeyvwBlOeteyZKtxtsz6NJ64OnJOzVDx+w
LckwCSaV4wg98lcfKc5KBjOQCpToIniBG2Qd4lf9hT5jvhEF3YYAs5CRq3CF26Mao3Vwt1D7TlUT
VVb0W1jDUJZbPOiZANjAMgJVIPL2SFd5mejhN8//UcBhOpbnuo7HNUA9UthVySFu6IYYO94xglJL
Bna+PZf/R8XUgpV3YxB5kndlhPwoMO2r+iPu7WWWZm/xsorHDj+WHTTuWfASpk1oQkR0v8f57uBL
bkcBn6DuqtULr+FKIPQBOC8kKOKBCHtpWEjH0JXMjBxxFSRkQuq8aoUu2aktAUw0TIlDbm8ZJR7P
l78V8ewZbiiU2k0L40tDn2XIMSWSpRTXAMz+oDka6Skq7psdbW305it6GClfnOVW7KpYovD+FH3I
kRU5DGb36vfWwNmqNxbHWNGMjBSwCXpkpvxZdVmuhbRmPCZW0OgiT8ksFu6OIvU5WBxWmJvs4ETd
vwsboMC8uK+7AKvl3C9Eh3RC45AAR7DM/EAcOa2+QR1NNlvc4JzVDYJ1sao+yt8yAprY35tkakXA
Q/fYN3ImNtavfFoio4PHNUyADhzg1BNmRZgf4CaFw4C6dKqLr8FCe537ShAeUejtmWExxc/IgNyA
mzQLa2H1OxNfEjR4Tt0cAxic8YgiiTAUBRVK6aW63Hmk6+3mofqVxFH79b1YShczv1teOQAeclIQ
G9j45DMF9pc88gfcTCKQLa1Ohloj9GRbSXij4vAFh2QC1maCc2Rbfr51ZNCEOX5C3m3/rHiGaYPf
tz4yUoefTar52/k+Boght8YWCzVIbGzLGY42gFeRxnIc7Qbz6/ILbGueah98Scgo1oxZtq5gOgB3
2x5ALEvc3Nmp+Y5x+N915jrXbr9IT86VjwXEfumoucoV+iJcYUNNh89rz9VBkZWaie8DzBRx8JMS
SewvECzIUE0Bc9hQOQga+vFQ+MrjE6QxIBBNUoAb3tuVTcC3wmliwntIXOOJ/yzmgHHH6hpkZT6w
dd8N15zAMfFWGTP5fBitSkH8x0XeIprIhfo4PqfUBCGChn/mrf8jsbavMJ/2LphIvMbDsOGS/htq
Tia1TZENI9vXeWONbSakraVz4iNAho58QrsHUjB6PsLlQppIlWKI5xlrJpU8jGgyy4MglktMRso6
ypwlVMXVlQZBbmeYW2zyyTguaN4MFPgNhzqjw13ISFU0A7ym7lmwB4P6z3M+r7ZLlxotjoimIld1
pcOGv+PL77ABcN1KXYAvrqa9V6dcqqkE8N6CuCKjfWMvKqa99doMV1jGfWTSjo5K4dypfZ9m69no
wbULsRzEAp9lQbr8P8FUunLDUFfjJaxyZjoRU9wkLNdOFi8ZwKytrxZRWoULfoPuet/AAiqO7WDp
CVrjC0OTXQFw6jeut8xJ/6fXH427LcObfh1oZGAbvv+BLdBq64WEv2HWIV39yZVD1hk7nTMLk7X+
x/8JTY6td5g9efwyjutzu/MxXK3n+iND4xajz7yAVDQBCw+RpMzb5MhcLib8PCVaXamvuTVJ6f4Y
zlEexuDCJvUeM9YWPOFuz6Fo679G44R36SH7/ggEkKsx9NGgsoeBUQ8+tJ3ljjlmEiex35Kq2YLz
5pHPs7YPpM0zzS4HGVl7BMpwuxFBWS4K/WUS/lMTmG8fRncVQ0Zbb1tTIyMdACE3sr/snvW9em0F
UzaiueOFKCnWnwjyHz0lIgIOJsCdIwM+JJg3Mo1CAdDTDeCuXbA5syrsrM6YjgvNSbxNilQZXj24
c95nav05n4HnRLAQWTfNJ1wFBDDD8rrD2OROuzLJOxWKphB55YCSmLjW30fkL5uBJxermoavQDNK
k/Cjj0PgbuIwXRG25gpq2LMnj0QVq3wLuc6NkDGnvUFAjGPcJPdGddUClTtOdvfMsYUGIk73o+XI
Hiyc4PrNXZ3UADlqancWC3OLAfTC+d07qmP44TlCXSFp2VglIhk7p2A0LK2M7BX4F8I9LC8XB4Y/
7gHRUnUDLgMtZMxAMGxWf8UdlqFNAnWWRj7Amo9piHeBjWto05RQxUQBfzE7N5HY54TkjajXxpls
JxjKqc0klsy5LKzL83//65LHn7ChBtEkCz8dQ3e1h/+VvbG+lrIPSMgzoemkXgXAT5bznIvqwoGo
ADagW+pWBgt6xx87QTu0kdDkszXLp/+KTRGwtFt65eL7MTnGNRAdeaXsrFRQs7ZrQ5sr1kBvVKR2
SmrGmmjLQfIDhayWgR2xfhjkzU+Q/89de9TjZDtgN9txfhoXYSwMIBkKYUsF+N6tgdztTCPCCpEd
pxBPJ7EUJfPSFNl0IKmif2ivc+IRWtML54tHTpSt7woYX9PtSXojxV/I2DzlYOqmyz6knZUbMTPw
bPP7FqhtSlrJ6p0rys1pS4KBDfHzVHELrlZTA3owxprTlV0Bkl/Pj5Jqxan2t354nkj7pm5IMsYM
P8AKe3uP5nua3J7KsMJHP4O4tMw0qzBz2os7JEO/r7xvKyngFTxzv+jsYsuLkr87ySA88OSSL3l6
6HLE1WB1qoopvvPkMMIZ8JPCiCX7lUN6xq7g2Fxl9LHOTjr6fViFQE1cfaigvhJRCn0VOrVWRhjq
jr0sWIVi7C/uYy/boJXszltCUUs0rRJj+5ckDVRl7pKehm3fLqESd1fTiypsX00Fs3kX+4W5R1UP
aBxNNufyCWkXwHdlC75lLJ4CzhhaIqrmEyrLUwsfoR8mBEf6EkpWdedYUgupk95jswGur3bbVeXB
C93b4uSIWwwFySFT8asNt33ynepUK94URgv5RQ11nilt4CkKqkz7qkX0PQjRBEBdYdPYeAYOneJQ
eMS375fB7EQ/VurpZIxJuFxI1wxnyeSN+tbczHknFERfsH0OLZ+b6SBOfrgaPxCBV5dipAJnrca8
bw0g0quVWOTJCHpOxPHPejv3QL1dYcpw7gkC9HVq6r/dG9PiOVjWWiMNRX2nydmPsFlMbEvus7X0
Zs4AuwNcs9FOg1jY7gaW5kZzl+UwLdOgvE8ljRacHxWg1KLNg6PXitAgpSM2xLMR5iGP+zoNvCVh
mSNqBT4DiY+26/5XMv/yOHGmOMv9xD6XwxZAvwjNyglnej6/OEieXBy2603A+/8as+8PR6lJEM1s
GMQl3AM2vG9jF2P7c8fu+xvTV3c2eTACnxqlujJU8IoNHzV0O/AbxcNJtJCbe4QjDIFqYFjGPJpp
KwJF/BIizU1Hbo1yYzNY2FXt1UgVxu/u7QccTBn6KtY51f/KvUNF0iZ8yQsvVwd8mXKZZCkhlTKj
i67Nr9SG3X+u6sR3Qk1kvIVytwhMo6JIECyKWBraG0bpOujAmoMscrk0/AOOpzIsNPxRkh2bd02G
MbAD92Pmqt2CmnH74ji/xTXH8Y5o22v6BnxuYg0kK9vWwNEbu1cbfB04vKFRxiKG462WtrYpCC8N
Yd4RwlexuhL4GV9hBTU+JtXJgskIrGlDLTjZpruoS+UIkN+vhrqZgVhvM3OyTmonH62Bk302/yQw
cUcn2reIfks8JpZkfDWx43AhoEn2s9gJKX3T4QWYm+DfaBAlBOu199gYDktymVK/YEpaIR8oBJJ5
SsVaE+lVFcC0IKTv33Pjj3mZ5H2Qnrdi5GpbPOHSgsYlsf0+s3jLrs+Ul5h6zFK30zjXyzLnhrxx
rmpf7rL9LgD9bmLs3214/TILBvCIqMfT/YCaPYZNwky54MetnmUEGOgFq6PaGsz/iV+riHUDcdMc
1brknCBL6dcMzUsxO+as0KrzqipUhm7MC0aMBa9EhYLGRJWrpVVemNYXm2aGM0/7g8YFqanlot8Y
z4f8H/QjCJ/FXdN9PBfWvMyFYsQ03KUsV8sa2tQojNY1ztgFSCi8A6CgNLj4nzq6mxM40zz52HBg
Wgma2neI/XBVdDLBBymm1VG6O+0d57Sl+Aah/xw2rUgbNgZ4tjrPFR/gWD3rgkAAUVM2Cxh82PN2
y8rkJuhBCi9vUZkIL+CziGBtG0oHboTY3kRZezQ2fcxpHbhFI6/Nk5T9fQoYN3L+k6Al5/7b9ksP
Rxc42XiV/ScTaA1k6fyy+K611ej5Zx+RxCLJoEJXHyKbLHd8GjN/NdDypVidO9V5SDl0APcM9DLt
+dgDJ3jCgP3wt5ojXrxt1rzZsCX+zghPtWNKZbRERZX48ROw2fG7hsZHhz4DBzioeUHDmtNQk4d6
Iu3ehbNUz1okqNRoSuneTfu9Z0nK05x0CMYeeEdV8TwsOOfd+edlfpONumF4kwEg3IR4qpezHSnQ
EsBhZmCSK/TdeJudqMjqtDgomp/K6aV5FGegH8WSFN4tooAdTYC83kzxmN04qOV86BxPSJwhTWDv
4cd/ISBkkN6qVGZvYQzytvnVGUiAYllQCB07houvtFhynXKAjivdUHvqDqsvuY5nHf1OF/c69wim
fh/1WyBw/gax2Ilb/+MxCJDmlIdvQAdJVIjtXQWytG64i4HJ355fri5CUMlBF6wuZnn5WPXAkA7x
whlqbEQytBkb6yCzn0Ufqwcb30JoJXqJhCVMUfpplgKSNT0SL5ehGVBPRPH/N6mraTuTYhOClWT4
0NJpUZjIjD5Dxo+aAO9F8/tZpBknYexS7di/1+bSKP1GP9XV9HF4jV3zDBvWbpZQvtX7TP277GD5
YYWW7ahMWQU020yYX9nIxXlq8H/WTVrnKcuKXAWvpzAWRpcEhkvg8zdthDAz3ZP3R8EgzbLWRmpA
RCRFyF0b03YdcjZv1KF2YKF6gxYKBVWH7Vuongt/8Y1lBUAV4sG8alVBB+hTQIiybvb8V5W1piN+
P/twxMe9pXdNwMjRUIrYWRYUkOr5VQSGB2Nx3X0cbJTl0d7LXKvJ2CI/PMLrksWOyE3azR3XSdbC
pnrmMPluuzouS6q81wWjkxEEJ8zWJhRpUrcy24vvmvsimkxBKgg2Am4wpw+DOrwcs35l7kOM0mxS
9ELar5cN84KzXSZ9KkZEeWmi4xSx/D+7JXHADfZE4AYY8kSgsFasnBLpXO0fplZ+lzOqttO+VmaM
i0QTGCgy4dNqE4dw1admlnlw4fjlL00hcUC9t+Sy2toSvoF/IIFutiVcMMxH7nUaXO+82/c+xVkP
EoX31aw0Leo0kQWqB+uagpXA8K1MqsMRPQbIirBh4yAuvJYgSWirIsS5okZ/RZPSsCAwq0ft/LnZ
lvrFE88j5AJ/iJwnVOJ5jyK4CtmeaX/Q0SnG0BqI4dzpwYb5zV00htPlMFAhmKIXHUj6YPuxL6PT
PJt24qtjAkgfxUa3ibZEcnos6wEgabUNWKb7WVcSWObc9k57qFDho1cB/lcUgq9mL/cZACpbmgnm
P1YsDISZZ2gD1BuqGOYBEPH2Q+sVXQBnZC1p7WtMfZHVMRmmZFn5+530CozQYbPheWW+oHixLWZS
GNZEFnsdPZviq8rTHOk/w1yA1mKRpzKf4HiNQWRnNkUu/ao2GPeb71JKD6SIHo4nJOZpASXOXEbf
UrU4ZtQZRfwAKS7+Dnbyx+amT6MRbxCiIkDHALhZYhh3PM+bzeKIWbnEihPEBgv4XlWymTddjsR+
gUCwk4PJvEBHwuiqxblACk/OtYtNB0uxvRBxVcW/PW2jtNmGTldOmSMJsAGYPTZcTa97m/HR9ahl
MgYg1Y+buIVTIWXx+QbPvtvXdptQX6f+N3ehGLpTZUYdw0kFzZpA42uPcU+akXbGU+6ensLp/tmb
++PQ96IT4nE2Bn9z+Ee3P5gzs75eZPzDDDHJ+xdc6P4U4oOPjd5crJGL4fG8H70JFtAGTyHNer2v
u7USpMIXG1YA53m4R1PgvnYLu9IHUvqc4lceV4iFNiQu9oOfChwt0AQGw8k69KAemWE8CsY67xEI
4myhYjT0mMmse3iMDufvUjindxu86/TjRsUGxVdyRFZJ8X9opsEwcdLCV8ZmdW9frdS9+gJrBmSm
9uEYfNcOt85aRIDnC4wwWHuVhpdCsJogUizjy3yUy4zWXjUnBuMcnFXtLDPUCpL4YbCwqpDKN0Pu
XQ9RviY38pih6ifNxitwDtPtiJUXx/MpBF47wlJwMqNIhoC6HBBmeLdFG2R93J7skTMnZB+NcZRK
kGH055yv6Dv1jedz1ZOLe3V0lErYJ38uT1Any/8P3HGvVYgVLkg4bTrgrn1p+Sl4rCBiStPFtKDa
0UplClxdxj4ja9MRo9azm1PiQsZANbWeRfdI283v+VpZR5mYpR+1rsCLIHl8K7z0YyTYOfOzVuPM
xHcyN7YvzhnX7hRiadnDi8GztC9smH466s2CjppnC1Y7wvK9hHqfXIHCGZ7BobKIUNVHrXehgbPr
roFPNbHa94VxQwaaD9euPrP62UBljFHKa/BXylAMbbc7nMePKGmG5fAHW7/zV/k1JKCoKOkI/PCF
EIGq7p7bCYiy8KYDR25zdlgw5ZwLd8CeGGzJN6fA8ffOKxJVg30WmC7UzCkrE6XtMdHAHdjTnwNz
uGfU92lGkY+mMxoi3fiHNs1QEjPYvKthI2Sfm0HctEOTaisjh4mR1NlT3mPk6z9VZqK+Ik+OQ2TC
bvqixCPIGsg8y2KPfoH7oCr4jONAskYfXuRQ5tInYPdD5bJbzSrku9GmeGY6VUkdGC9Le6hy+SpL
C/HHVagllxaJQPwIVfGFlVBv2tbyjG2QOAfAzDheOXB5W9A80ZXTq0sFFrwHz+951qwbfL73SbIr
b1aNzEH6TLwLQ1zz5VUQ4ValeWeJ5Iwh31E3gLNj1m7XYrMFsojFdhQzkUTpM+JiFNcPnKWAq6UG
2Dj3DWfRei07dQUxOiM6baTGPjkxLVZpm+mubZIiyZySudqACVb7cL9HS597dPeNX+MyLUXB/K19
YALqHpFt+A/Gnz0a6VQa23Om3KM43fOPlYEDQu674gEcEaEBHU3t3eTPx5X3VYsa2xuX7KcdtPSK
2sL2dNLxThDvjA2nsAlCHMksN9XqPyTJJmH51KBTsEnD/Sger/RKKS+MZKEZC+N6aJEFyqPgScSk
onzUeyI408+fKFW7+FKtm4nzNm/M7YcsacjP6aFmVIYBPFLR9nt48W3WXf4LkX1uD2tDTgb1h0Lz
aYdnFCJD/Z5hvLfHTzykhVBDeSOI4LsiOK9csr/KL4e2JrSwThDEtScqmKN4tHUH6QeUndEci3//
1VNWF8eqa4o591uAeOgOEfP7JtPkVNmpP89qh6xh3o1tbjwy/rhBLERc+Mv/FaNTU0S/T5B2JoD/
FMQ7PwHb8boBsKOpsgd6n56EwCyBFOtdMEpurItc9KdTg3WHbQXk61qjbzADWXpanmIynXx7PX5W
c6znixmCboQO+YtjziBnjwp42D9/+GT3Dd2SE4tSffnUdcVvebeLW+F3z5nZaeZKIwJw23VNT1+k
4wWbXZVpxG1FX1rrm+H9IK9If6Um3T3JeudanFp3rqvnC/cJs3VgXl0lrHpfBaXISsrMWk2Gq8GF
F7wOG/TGfObkbDh9s0D4ruSIWWGhzC5/WoMwVmqM22funz1yx98Trzv7G1pmjPHCVYhQX2Y0bUAn
2XEecSGQsvVjzi1ritd5KVohcZqElaOIYu8wPeW+JaiHE5HyCpbtgzdArrC32AjDiAcvuwueRE9F
yeDlUFX5ub3rectIqzlDoagIWZ5YkCWsvN5xeKIRsxad9eCweGloalo2DyAJrj4FGNNgUjhLl+yw
uKJ+1++USz2DxS0cEiuflAmlOMEI6LdzS9ctl9xi5C+LjvzyvYG+Vh5BjwrpMEk+6FT6euOhUS8y
3NLLZUuDmh6/o9sT7L7gHR2/6B2qT0/2gkiZ+AqJ6nhSki3cy+JPZNhxW9GdaEv0W+J93ufHetoK
0YcT2Gl/t8KRYzxe4B2nMrkwqJOQUk+F2bCB7DTRlpD2DUntr+//9iOphurGlWAKqMLDD/B9zqlO
dM1ZP0EX6loeZTea+k1ZWW92/GtowIxhKYvrJ/LRwaNuZqs1sFY5Xk8DeVTlQ+bXeGOf+ExAj1xs
YeJNmNolH9ZrsILh5x0tWQnvAQtAITPb6GoFTyPKWJnDBcjn6Kf9V2sEG1sJ09QHdkwNIoeL/VKZ
GwdaXVtHePGbfpKULk1YJKdRLMWUQKP2GTROhQ/ihqgdVxSbCwnTO2JOus3NjFqoojlBqkKVSHoP
S4XtD6WItadEOGNmjOufOowz9IE5U0A7EJdtjEe/CLSUeRmBrJTYiNDIn/m/wnCHAqwhpGArE6D9
bCTF/w4T2jpcPauCh2+klWjJplFne8HTXa4SvwpfFB5cdaH3d9e4NCMARtgVrz4dsFsUh4ifeV8X
2gvd8mxBSoPkpyOaDJfntvld+r7lSXJh95rYvL5n2Ygw65QphZjaVQxy+aV5JSBkwrcyDLWIQZRM
VX298absxgneYkuTNAmEcP/ObLqXigvCeRQ7PTni+o9J+/KrShGa/qGE4lvRxy+X6lHpLLheWNtu
V5txZeBY8XTJI+IG/SDof/DRezSruFuGQ3fBkHxYeR9kmpxKNYS63SNSX0Bxdn/8Jp3uU9GvqaZk
9YMQwvOqDR5Tzu/0rbdMm/cPIY+GRuMzWxO0pUcrrH7qBjSkMXY8s2ucdB6e3fqsEoKwN7YL2oe8
FMP9/UecLaqLidnype/ijHvF9XbrylE0S3KjTad5r+qUL1QF3YvVw2WfN1o5kwuWew623q8pIFOt
AJr+zuXALu0Q7R12T2h06xytswGOhjeTgpkgC8kNcs4B9PizBpEcezS5sHYUS6bCFXi1kUrbfPfr
XBrl6Av6Z8UJ+B4XCamlNtz5I0gTFVz6J74As/SLz5hZR0xh6LPTVqx4ahk9WMQ6zPKX9NYeI/V/
w8RZgHv1C4x23wz3nAsccvmO33hZriNAcSffYAwNBgaCMKe0BhOKqf/Zo9oi3uXA5kjRcK993C2N
HUlvVZLV4A+rJVGGVFL1jj+KLU0+UANCNvN6H0bO/dfvRdXfyHVsQ6NyAzzxEcwh6w/aoC6vRYRG
594RrfOBD3nM6qGcKMQgL0A5GOgjiw8FlOmloXchh1V13L0G7+Ds4KfuJ9E5q8k+YaLdq4VKMZMS
tF5tQud7EVr6iCbMm25ld2MZOxjNmL2OR91SuURGiLugoUrI2Dclwaiy9SLmdgjCNjuS6sNLpej8
dA0P0Mt+D0z7OlP43MswXis0GBFHSW41Q4feYc5ST8R+ZB7Z7HMq2sTHZBPP8AjJKEfuiOVyw82R
G+PmWRVfU8otPRiUz1HR/83tKVN4R38zFoOJZixjCRoalVYKB62FD5FOSZKQZSU5T3YixXZwWmVT
w77Ln63+k5nIYPhpS5uRdrQeMnnxbaSHDkgmDEb4HACgbEG5zfeQK4DfBA8msPiAKkcaXdC5xChr
bEOreagCi8ixVyKP5KQSyVxIRsQQPYckIaC99Ag8rikF0v3+ha+aUqmCZa1FZEMxxKPM0ZoSCxVw
z3tmYmE6xwgysL5gwGc14JZjCJ9KL1qAM0Pzd2DgSra0aTri3B/UBZ7aDD+6wAL4Bf3LWbmeli5k
su29+9ZMWHNtkr7JFV4b/2GRGYL4Mj5g44iZW6UPJukn/nVPJGZ5tRFDXMUNVMFjkQsp65niOggK
2GYMsSVhbZBtF6lt0VSFYoxwylFZNgpBuGQqqU/sdj31Tbq/s06jhzEAl/tgiX6VprlYom4xGcwW
s9ZwSw2DzCYwcLF43Wqjtcih97pnoghymb4RjihYbJ1tC8mEShPep13VT/jlNYIZvhjYJnPQg7Mk
be++sbN48szig0DCOo4TEQ7LYqSs/9MBDWqwfbBcFvNx1iVpLtnp12uABkbNRMsVRVE0/TXHXTIW
/ogDz+3HWwj+ChY23Ybak9cYMED2beRqro9TMHgkhBE4TjGVayJezuwI127kfHH5CsOpE76NbkBs
D4zcOv+qry+vGBN3b3CLJOHKxWqTrAa5Gzoouo+qdtiO5RjeEN7CnQZc9DnfkBjsgYpGhp9qmZH4
SgfGObK318LJ+p1nQvjPwlw/fsKLxGN2WQhvJbzEizi1LDhoKOuXjO41dEmIpv6LfrwT26PlA2/S
E6fG2dXIeBXdFph/R8jvDvCA+MXvk/EL3aLdPDpn3JtL2bPfJKL2lHoq0qN300xBG2olccBok5Eb
H+r8ccRdWXGq2V/GH8Xa0HLHXUMqKkXf3C+nCygICNxc8VdZaWU+BUKyylmb8J+M9jc4KX3qLZ5l
Z0LRBllhQz0al+0cs77jKOCoDSfdB1m8F23oKLluM3VnBquj0IQE9P0tthoo09OiWV+a4ZBWn1hg
sB1cSitVozDCSZBwZvsLbOnc+5w2DuTQg1QaAjkJ/xmg+I0vaap93mwdJLw68g3L+5K8QuUvyWpW
xoE4R9WD9w4Bio4eEAEkvvC2BQgObJezg7T9YsdZzNoRW5LTxY/SqEd2B49iog1unz3ApxM0tdLU
+FVUeaWuiqq/cX53YLsNx/w4Lj4CrcHRymAkupJiiB++S6LwZ6fKS0Ee0xBDdt2UqLnQ/lQ88XNv
OflqiFpAx14esdELQuRZUOBX7Vbn2UVBavL3niPCbZ51e+821VsstFPPMYXvUuS+MPujyHCCBWGe
0cJVjX19G8dNaHSx3Y26Xi1DDI+SvciaKPOVnvcj1ydl3QQtvjWoVp3NWfmOA1Zzf2Ai55lvuIXD
J7MNYWQCeAWTXeMrP1oD90AyOMm9danNNiD4Yha+dLFRbx5Se57jV8AC8MsQlmDIZTqcudwRSxSA
OSoncbUoVbBUw+osFR4vETdvznF7Ujtv5rFhvvlaF0s6UN95RiP8RNsjqwhOwAhBXJJF4DkJL0si
mia0DoArxXpZe4XEXQ7QN7RxvnIzDoPJj39LQRh8/AMkIIKXSxIWJAsAGkhMXO8RKt7hw/yKYs5Q
1P6sRUH9t9g5RZLmhx+fB+ay1Ex7qZhyVh1qQU6o7nYde5V/ZvVbbBRcs+4MwIeHRBwYkCUFt9Ul
u295amcfwHYRl+LWWWYXJo+H/IWmJsdipAzJPCtHEFX/GyjbALlSZckf8KH20GzlDop7gSi+zvMf
kH8Oh5Bi4nhLm4VM3w+h2JC27Mw+YOd/oaZa3WBeVhHxb1oI2eX39bqrBi2qryirHAJAzbVzQnew
xUh3R4sIszkrT66Sb6DF6dZ6e0vPduf3cz1Kto6z/C1c/5FGI+QZCMmm1cUietOHOd1is+LaFKip
5AtoXfRWAcqTlqZhRVld2X2DtZIMTSUmoljdI7uXgbC/+Qa26SbU/KPkVdP5zre8LrhCHpkKB4Vf
89BVpXjaH9EMb4FWG50nbTp0dtsMYZctmkePSF/LR/T/BEe5x/7d8l/rn711LUhlQzZWapqRN+WZ
3MeFkkoHCLqPBpU+rQvtGlRbR7IxydlLZ5cfD9cXdP8UZ129QO8Q7D9Vut1ywms6A9oR1Ap3XdVK
+T3jat9uMgfIkwgu1x2BngSYZLMm0GAnihOYMhnLihtMtrVgFO2SjnZN9CGiTFvpT7Pm5gqF+0WB
0YntJcWV4a9KdFncYYc98nW1oxHYorR9iTdRjs0bqtGxBRgDyrcltnlqah/VLX8cbdgDai+xRe+t
QfF2QFwAhLFf1UwO3m2YUT+50838OoYBXpWj1prMNFag5rp4uul0ZGWHuZpJzmZ+jAb4MoJz5Uom
bIIwXZDVomsEpXop07EQTBtvK3AvWhgo0poAoXOnWwdNgQQ8h/3h+NBBSCvYbI/j9eZyvnfD+9/D
fLlfaVxIGZZN1ZaFzW6RtZvYtxJ+yu+fd1m7fU0vrke5HeedSulczG1VczQ6G5qRSBlY99WehQDR
NxvljBkSwUEjNpUJXgr46RkeBYRQ3PiLYGzapXbeeVsSpwN2/E3QifNsaejNzziOBgAs9sbwI9Eh
+DELFa6WUtfOsTov51bdGTww+3fQHR8dRo66h880jcLdXn/Zs2dPyHR91qNKveYoWmDXaAAxboij
ENFjwvgQCAi8c0NjkzNGoG6vggucM+QzGimoEp2PVcFPru7VZgsSeFoxzT/gMpG1Ux3lHcIFgfEl
PALlRReuyGI6RIisT6ZoXrX4uDEPr7YughqBXBSx3cCNWWU2Pp2Ft91bX5SQh8xyokTcoLQY+fET
3g8t4KIXABKo5u3DX6iqT9X7I5JMWrSRSxncsmdu3/t0sM2oEDgBXUGxTUdoYDwiqGaTdNtiudHp
x9wog4/yfv4yCd2dggdO2EwTFBkF0RwXiqpEJrVzijZ7TSAwrm1CdhAKb2CUorHKyflnA6U5Xk/l
U/s2TlDvF+f/BO2xfpm3CVBd63KL7Nvv+LFH43kekoVPyMyO1tqUhFvkFZDs0BPvsa/x6S1/xydH
A9wL1ZY94tGG29osqWSE8VE0G0vykLEWqXC8T9+oPfZRdHd1T05dWr0YzTOMFonEmgH/txCX4AfH
kxBN2sWjEXrHzdV5xHp1GlIKloTgNbNDPcRZ1nFNeYxo4i8Bm2qU7Bi3t9Qya178GAamai5DsEHU
RVaVmzdhcwoJyO/yFS58I3A2MGwOcpoZXNJ4pphwq7nQi+D7L3ZKu5ch/33IYvnJWg4Id4A+D+zG
3IPXX68TI11xBBfDvVX83qnWsojb2E2L6HtfhZFCLYezV6/QuQeYi1VGSE5yZXfMpENcoRxCJLEz
IUvOKigt8X6vysWl3cx4CTCf6ka5RUoMyrRTgujc0AigMdaPEFe7nA2y21kXK6ohcgtqFLMtFfyS
4hOa2cNL2NNtbc3B42Bz3JTS/NwPpItdXwTMxH+x3T0KVKFBKMR2YIYDNZzJYIJ3YVszSxZ/WLvt
Gh0KCKUIUWaO3TUR9XBMpC8YnsJSlYtnHDSVv0S+xfVoSwLfES7P8Q+OGkoI0F5EyjMp8F9qs80o
ZKDixy4c5ohayvVkHdcFI7btCOW3T/GE/obydzO301j+f4mD1eKR8AAqdAyKCHKPl4Fl3gUPVS1G
CNwU4vi8jgRCNTj49i5pYg+Z2zFiEe8hpk0+FbGcE4rXUw5AjvlIYKIZglyjYjSgq/MwS7w6uPNo
7ChC8a2ikF5lfTHg57GxOTSgmRkn2rw3Y0PsXmvRxMMuPFGrP/t0V0ozWHv6lXGgDwi7qdhEKpPw
kX/WPU+xM5uwinPZuTWH9Fm2cog3+LEWiWpCteGh4pR7nl4LzMX4L5/8iI4UvxxkR+ZcSpPHKJnA
G5ufivV2uAmZVxlwE2bSpIIYkaaWqDx7PzdMRWzPntGn2EJ2wKpUGyhHAfOq51Xj4W44nyT1mPV8
5UZeN6KLckE+L5Th6gH6Jg3HzyQmMu0x6wcea9ibXK8/tFe+H1lVPp0F8sPuUG0tLYIcUx6URSJu
lrbg05x+SjtkcP2F6gJ21e+VbDvmx6B4sb+a++g4J7TfAl8W8Hylb6aC4sgOZOD0OQdbLtVAz9wF
KfzihnY9zQpjwjs8SEZ/IxE/jyf+OFEPOVjGvkS6qw6Zz3uWzJ0yfRWEUdQRMPCNoZI4Lc+nAM16
wlv12nIDcuiilXUc4RjWLxZD3bmU1HBDK1EkJ9BTjuse8WCGMqmZmKeYTUbtS4wrD2ImaiDueO7J
y+UnRxkeVtTljtn7Vn1yxrvW5sLvQ8usXKGHMLL3xUUL82f3E6MPNG4xU6G8/kH9HSN6+mhgBxpC
hUT0rOF+y60yUapm6PoQZjhTmbziINJS6mCPZR3A33TlteyDiLiAlFrZ60knzTQvyNLVbBroMFfA
hP5RdjJojSg+RG720ZtfK4fvSvuUHXy2iYJ2YfyyxwN3FTjf8Lcqx222CpAkJxv11vEd1jdaVi19
4UXLGeEKPw9jXQSKFR1qQUU4N+KECRHkCh6WRJUTa0ng0lmdaYXCQz0BrX9YtE3AG+Y13cOBx+fJ
5IabsBzPYoOS1oOEw5/durP1zB1i6wABxz3hacdPC7VbnVyRAa4PiHbQByhbON6jNw9o7s8kOWZ5
CoTlBibznqmNNfmqTgZgws+41ui7FIeqr0Pp5GlXuEZov7YoiD2SRaSgvVJR2yEU1EIyO6QxDobZ
QfDnpuDgqb4ictABvgfdiFTXY1jSo7o5Dp/7VmUdNarJN6sXij8T9lDgUbXAVauNPWWCglifwnPl
qK6CH+DdsrhJNY+oihDcvvOeagg8asbUh/nyCIdHj86UQPGyMAXML45fJxH+FVP7Xb55wV1CSxHT
svnGqHegyVRsIm2w55qNzOO56B1HwmCvdtYAXbfGlzV4hskYXlUyQ9xYyR+xUl0hyusrfEHO7k3u
g+7PT7cBL1kfefy+pP1NUCddHt1uYBmaJSF6Xx2PmTsVRARMBy2r4FN9paPM1BYfuyRY+Klc4OZi
hOeB9/XV2qzu5mtvUmXVrftNi3d9mFZvzFTr/lN8T5pZdZRpMeqsGLZxyo85nu6scq/4dKJbf30Z
gCtc/ZrBkgMWi3Wi0mXqnGBhXqvAfT1zmS6fa3ysmc7XTpKuYog5niTcXGAFn1fcuf+AtiVmRK0o
TQDbE13AahbYHn13dd2gaMiwtLMeh6jWpnRT6SwEUeRKYtVuCTV3vALm/+ABEtHvY8/DURHb7fxJ
oi6PeTnL0ejbkbDeE/PeuqsCQ+gVVMxq6dwOYAkYZu7hamHx77GZqzfGgNGvhroWXdDrRugpsjZP
Nl9vebFRNSfqeIhCdfFCUgr/uA1C+jijb0ranaw0+b3IKEryZhhlmJmLZiWxXcH3dSS/LgXk395z
6yG8uoWry9lrYgM+iCIzUHkyeYm6FQ1NNtogk0/8dIe0Bs3XyHIdQfoHrrFOL+YRteowJzIo4tGE
TWAfbrDnumeJyVFzGae1GRqsgulktMfjPLU71Gnj5Mk4epTndqIz9Ef6KH/azPv/xSykpGrPNoBn
zNuZBzxlL6lD4xjhDdBKatgShBXLT5q09ScQ6J1E92mfoUs6fdEIDOz0nTOQS6IsahA67U7EuD7g
B+HqHAE3K2uWLMgahoOmV412luz+r6iq4h+d65BuUpfhZAW5gHqMK//pZ8Sw/kSuvm6mfhXQo62t
AjnjFK+iFVHCZgeKFXe+YqgUiXDZKdW08dfOzVw9gpH+eqowHFCAJ+wfDBcMBjRPREXE58Vj/kCJ
JKqh8vD7+CcnyRAVJe4U2PCTmZfnAn3P2n4jJ3MTzkTwfZNWrO5Pp1d/zn/4Co7FynRjsxJnSJK/
yxDtLvphPsa2j/D9Uvrv1mT90rZzkKjnxK4k390/sO4J3qwLX7lV/oLYrP0UHkElXX+oJVjv57Kl
ktNjCvGdgp7n/5/90T9IU/tazya8iD0bGcG4u6M3ecqXB76GlhOiDg35jUb8LNeoSarjNoQqQK81
8OudtpjXk91669lm+pW6Tghit3Eurah7NLfRDdhja1y5Uy65YwW1P5U85TRebtP5bAirmV3HG7Hb
E2p+390uCHhroByFwF3tp+6bZ1H5wkFGLfR8hqyIj4L1CPHtxpBGV/28sJHV8GqH3bVqZMOh+ezh
1Z3BUAdOthqX7rYvBh4exk7cros7HJGxRecsop8Viuh7VLF6zKetY5lL+UkgyDB4AijSsuScGXlK
gyJK8TOzqCgalgCQU8YWWmt/Q+PCTkMEf1HlOkwO6lAT6lTdjbHp2N7Wzwvn6iok4jtukJVKi0xl
3ZCX89PV13s1YuYm4Oqy7kVArzxRZLNfT1IXZ60YCsEaAleZ/b8wd2bKtoED4wkKLMz5P4vFT4Ux
WSJXdgVOPZh5DhLgNxFLrrF9OznDX3bGAG9ISeZgscQm8VG6G3sX6MFCnfSD3HtgBbd6aGSOYQP5
Hif9p5wo/F3FdIlNfRk/2fZDmdolDEHH2yJ0rHhg2Z9BgxTTOYgTp17wKF3loHH7fmOTuI0oibki
VWI3td8GAWDn2jmM8QN0djgBqBkRzAxZNqpVnpdaAx6zEtQ/X+FKraxYAnzpGksMFHJGbTHgMP+Z
tGGq9idj4d5xqd+yWMNsp74dys9OB5JC3oIK2RYwSNTqJ11D0lnc00zwUtnvh0DSRsJ6czj+ecrI
8A6harrME71BJDZIytBxbJRmUVDJBvSPTyv7oaLq7sFdkh4znBRss5sMyZQ/BgaMhrzBldFJ/UYA
AJolv4fGO98h4dbiTYfuWh9OKPwZgiKreCCi6Rkf85pRBtC5o9HTUqulfB1A67rLXtRaMifjxvEr
+/Ba74oMtE/g5lAhuUFilIY9ADMclobYfY6m6gWPfZ31O87uWEmLZtWxKij7lsIFxbeQkvdL7eZT
8d4uRvq2jGGmuTW8UVlKMXgxrrl10M2oxpr2fLwBdX+12aRDN3/boCtLEblypdPj1ZeYyoTSBlmT
vL3baxnXzt1t1d3XcZyDrVG/4aaM5qzuNPnSu8QtNUnNFNiGjDDMJKrCgPg+8zsjAcn4cWtX/eH4
l0uQyR65nv7H/eCA1Q6HypVZtXSLjhvQgEOu514ZOTEZ1Xn82XfuM+f1CFvGjJQWbTb0G6xLmrTS
/X3dCXLz/mykGxPYSMaj/ro1bY+tyfK7wAllef/6KJOlY3p62t1j+iV72o2k2vGHNSirpAbw9v2y
w07O3rFPlrje0g2XZdo60XZg6pSVxRvWI+HTfbLifo0b/f5eQucP3GWWNHYinehflyPVWOxl6lFW
xtuirRu9Z20EG8jPg5euiS16A2DMMknYF5z5cmyj/o1dPSh+JFIqZFbQg9iytcN4plvjMySR0Tl7
0GvPp6uYweXBGxJ2viz//8Qp3gAyOg21pZMf+IZG+xRFMZJyZRvYWQQzaL7xJ+Hv07LA8uW9iI8l
gSRjykLg7px5KIFMk6QLf12tXAPAJUI3jMCicSQauP7mfp2SqiWeojBZiKdGdfL4lk9Myyed2lwk
/tS7/aUBZoprpGqTWC/pIm1atMhGsyq24lLm0tGGgtNPrM9Sa92LMGyEvYXq0mgg5SqR/49wYN1N
Jxneflff4Uw7J5h3pwE8/B7U66rm/UnrgD07C1fOZehNF6Es0EnkYKZm2dWKfC4Poejerat9mwSE
PgP6ehOeovrrdw2BdZoxbPG838aDq7iNw0h2d015TKoMnpGAYh4hVydLA+Y4IDrTkF+FFb/GxFvg
wtaGowHqBReFWjeXAjX83dzQPv1ZqZP2HCCghaTo5K9Hv6ULcTzCzlQzt5xMQa9HUpzjHDdMyxhJ
HWEnu8pDedn+5MlFecVBdFZvB/B841ETW/yv5fJxWHGABOhzBP3ey95m1TmQwyAEKPCl6Hemfr7T
X0JrA4Wl5pa22JrmzGPQK8lx4XQBa3xAuDtd7+vThpO3w1U85CtMsrxdNE+LtctG5JoRIMt8UDIx
EjAIYQjUlHe1PwpdqLQLyZGWojltqQtiN19DEZBMYUM0OiqphcQLaoTKQA8DWOdQGjZB8/X3zpk9
IE2Vd3HBlJC8sR73dT+VEL4UfmGWRpZ8049PgxejGIqsY7FM+M3v28It0XoH5OXjYhAWyuWKkZUb
0Xg7eXLPraWPnFyQnXJpdQcXgMJlaYeuT7IAz/M34U0TIESLgeOlYPwoU/b4s3fcfUFBSRazp9Rs
H3PS85jofLXKmaMlYNs4Nh2ON60IGVEACblEDayqN+mZQxKGfQpFRvjYAEy24e+Yu6iVZ9TVLgWQ
/9W30FqnsAhmZsS9NM5OqTsEhFpYrJ1vMhpa03vlI+XkKwEQDQYP9rkEJo+CUYkvOjSJuRFuI2fb
YzMYf5druarrnkZySaY6hIT957v7cCHy2OR8Lb7v0ltCqZmV6uslGm0O9W8erz2RCMmV24JNmFt1
wuBL/e/sJGYjIFfEh7l34LcY8sOhQwpijYQO2P+SSGXRtMkwdqB9sNWcCy7GDlSMfHEiCgKUtyUI
GNyAUX7KX3TLUeU4/2OCWmIn+/6kf5fKGd5pY6wbQ4Qpbq2W4G6YyHK2j+gZJ1dowPwEAtNCgscN
dJ2eJPwzULUniTbe6XCDapk4Ph+9ZqbHJBvwi14G4LT0z0EWQwkp7LaqCbaroEpKrAX7MLXhMKMj
HQnH5QSKkZEAZNuhmps1tzmeYEYRP7WfGca/saKlHT2ihoT8M/ghLGtjY7sc2OoJ8WGtK5KEXxxi
mlcm7l9A0ziqUnZFzvEMx1H92UHvZYFBdff2pOvOBN9TZ6B/qUJnKUQQyGfHEvVHJFZTPBgaibP3
R1LX2t/NQzoKzuDiYUHltnVV4gT97no4OZ/UvIBQpoqnpQY5KK9VXtkOSn/HBvjL77ecO/mjcOOr
0DiPwUiBHHQuQrmXDSkG4yIBPeSIEIVcQ0jBspisX6HW4wuY0g0LH9P+RUFnXU0fX4yR7z0GCxFZ
Kzvr6vHyjmgY86AKTJnwGNX6aQsU81kNwWPF8CIHwlzBdH+atAK+3HGMoM/8wOg0zbFps5WFFHw5
nsUvpsi0tV3wV/JlSCLfp5JF1wGdVIYuD/WvnjaJdpqQfcWU01uXTJOMITq3ejoU3F90S1PjLL8E
DVNyz4MpuketXcEVM5aoOUwlEYCkA87rVUVyId7zjBWy/L1WCUNi4j/Yica+3mYnfd31WhvULYVV
y90xQ7QPejEItiYjBAt3pflITr5wcR9qzQ1oyDgYODytqkaVIXpv7w01+88+IqIGJvoIxvapPPdD
UTjjq/s1bebIDY9ZUi0+3kPsBiGjaOALeWIIOicv3yX9MhWoZ3PY9N0miEBkNMKDc2CfSDQ5wdKm
PbFN1hW0/o+hfPGTdHhzI4BjZnpDV3rhFFCl3Gj3WQM9nVFViqCr/NnVYLwxcqV0k2rw+rr53bw7
Uj9Be/99ty+47pv1/m2aW2jqFZv00UaeCq8zI1rxCKAaLHhkMIPGHe6hD1vlxRA68sCiGl5GiYxx
nYtQxn3NACaGmqu9wf1pkDzhkSmzKUK3nMwwvCECVr0//m5Sc5EAO2QKbaOGzSgu7+0oUwTsQk3y
K9+kkDh6SPTiPAZ/EGQgmoEWc2aiz/xOYyl9PqEQpSpYMuo0kTEEdLRJq2VBvKc2B9E47n9IBKp/
zf/kmqH/1UOFaSct+SUnEcgOm56avogjtamBq1/Ls77lWpTtLd1G5unVlG7J2v2advnxgO26LL5H
gGtSz56MubqY2MXmpk0TWKw04ERrnOZsYbXI9mUFrjDueUr53v7K8AYHHZa0RBslzn0gjjcf3oy4
mYSLNS0n8FlWey1/PlqqZRL/m2KkIrdOiWjLfIzYPsBoUy4GPySHjXiQJ/3Rcy6PdHCO7hVl1K5I
Zx37YUykaonGqZOf2rdzXEN4yi1kV7vf/C4X18cRVUPkXMFItcZBMuB2tAOzzwDXWLbqQMMR8uRg
/GjigxTTM6tkG3voWq4JAg2k+pvR2GbiXgqZsCCndBlNmA0A8INfwBu8UP0aeAj+wta6pgaUFmDE
vvwOiXNh2iOXpf4PR8G0s09Q8eDBZY6Lop8kHXQp/rV4xM8Nb1JjN7yOOXZ7d1VYRML+czy6qGT5
GvqE4p16Ce2lRgQr36efgpbTLEAxa289r+82//wKRoRc33WoeWeDmImm0YWGY2FBHn9KhS+7GEml
GPMjKLKC02eZIK+h+gnyzUb0Kkk1L3TyQPg/X/UVDXi7blFhIcps4P0stB+bOsG7Ahuk9ifRjHvD
qjjY6i2UhmdZDmdB/nQK6fxjDZV9uwcK6XLjoNtMxE1PpOsGSrc+mjUYT4rX5xwvBgGDxwMdNuSw
gpYlXk5jyLQYqXAWfn2J2hxgYNsrINR4udIs8zQXr/mEiD522EU+5yn/jTZWLGcM6vORJxJCU1LB
aO88qtNryyN4UkgtwbPNFdtmLu5IBZI7qx5NzI9H/iM03nTZ0HYyuFDEDM+kwJqcjqEFiF/f4fKR
t/HMwKTQjaTCYOVkcoBq0XbNmobUgwRW6yEMmtkCSLH9ngmYNCRCakey6uhkHvLdfQUx3Tg4d7lZ
oCvGDSuA89+MxTZ6zLPoCYyndVVSj3F7Dfq1GvKe525tPYxY62r6Et4WX3Sr8oEq/La2Gz8YmIRK
BXfVMOHmqFfxDDXbxIPBQm9EoHnzOXXfNNFL03sVq+IBRBJSQpHzFNdS154yZ1yKm/3W1dsp+TnN
bx+iNgmvfWJ1u72SIu7b3Q1UwvQSMJATOZ1FUYzTNYa739i2+GnhonePpb6aF+7QPpnw3znoPaTt
Q/6cdldR++WFAp54FA4gbzd4n5hHP9vW/vgFm9NLALgZTq2OiJhQuhMcbEMczH89LqdQbNpxZdJp
7HRWzVaC3vsZwjHKCuMR/n30BtnNXaRiYlhJSYl4pvCt8TLStwROJ1vtNiqeX25RyDCQ5jhrGNql
G36BKozqzCvoayu0lFH4D9C2vEriIk57HBQItjTrpZnTOR47hR0dcR5+zWQs29oBCmKSO/2Oda1S
JVxx5lJbHUCTV7RE4HUdN+t6FkHwf58YzJ/q2yTjq/XC2rsrl4Bf3C50C103HgDyeRqNvQL9S2uy
iY9i6JIitkgWy03RJEtjoCAtctxYEK9WEj2HwV/ldm/OF+06WOWPtQZdzCut1IZaVH4vBH2XoiCI
2qIEhF5UXBsiMlfuAelRPXTZygJ4kRhUR9LLRGp+M6TRLlv5zZnyR8XECjKSXusxi3RztazTVMCe
Jvfp9nViYJeXWhUGcpl60LhVlGsIWHAjF21pJI3g2anGaW99ObIwSUOVRaGdf0G6b24fzbBJH7zZ
fgblduwrZ+aPL6BzYLrM+JQlMuDbIZXG0LIcOQly1AsWsHJIrubNlSFdi5VKf3UzIpyoEIrsZSFv
vioNqdZZ66zCYqfwiE3rxqjVRG6g8Je80W7MhqcNzS70xRXdbwy8aivdhQlO9L1xrv+JTH2/ufLL
dZXfDcB0gGarr1dgkjTHKS5fMKUdlW/yakQHCMoXDMkDlLPjK9l53qU/a40uiRKHfi9lJnn/iLfd
/cc9lDAqHvD40AHYoebvqX9aeKWeUHv8XUbyCd4RbKeKXtDKwxxahJeYgU99tHQDua3SVzQbkEgf
vc/XDxRXhw5USv49cLC4RKR2rSPZJRvKrLeOmrkhg0eTOMiGzCMGT4L6TCyKvCMep1NwEVDPj6uo
xIu/CsuZq1brd6Oop6ZC0Hs1C9QlsYfb3Cd/jo82EpeUAg56K9VsT64Bizgm6QPUhuNgt4wYZEBT
Y8cQ1ontA6auN2DUW9Nf7utIvpwP7RV8M2dQ7V3DpvWFUBv6Zr4o3PJrHSuDam3FAO1S9oNZaxKO
HKOkqqqBJCh821Xjr5yp7OreM/g8bWny8ZBixJGS9DiJc2yzKiFJIoeO2mYFOTLYKgLkM6IiW7Sm
M4BdUj7gH9KIv1+4D/uVQNHbPd4xIGgV9AdTan2QZUPOCyui2Nhm+J2ldHdkfO+ztRB7ZwJo+vYi
ax2bYMsz+4gEQhByu4+97F1y8sgqHKSkyzGcG7XqQXtr86c4l9Tjdv7U3tzzNsAS3rGWIK80qr+n
YobLb5ew4ygu8ARbUvr/CU+oktCv3+F0c5o+ijDeofV13zKmH35YkiqHXYT42RusrrLU/ve0Vyey
NxmjJfam1W4eMfISgPT1fwS1os4TAWJyEwaT/k5BBH1dpnBM3c4IH+ELBkSu42qkeVR+GhFNOja0
fkQisxxJ1EighxycqApRx7sHtVBUM0O+5K6S6GvI5KkmelQH8woOJNvTltez5MAhfKKkUNQ+PMxL
tlE8WRCs9ZHsQrJKcp+H9dmxXcJZpDzria1GLDzwcVdJmO61XoSxEXXlrl01pCJBWVtDkP35QSYP
12L5bOaE1SxY7T8lZjjnV9bJ6QGapXZy4zEw5+UpSwwEmw88nYB/N9eL1RGhqwvyn9OJKZM4hyxk
0+5Y1NTydpvcilmkCk6B+4U0DKZe/c883wAsTRI/xLurZ5gbryeD7tJqt2eWUICYA7YT6TWyGG89
5oNTPb4sl8VPn8DlZGD6Qhz13tXRInqkB5SSLhJs07crcd+K5Gyp3pxxubK5hxZMNaqr9RMmvG5J
9Cfaxh127XgnVMUHkzRLoAijIuMKRr4Oc/txCc9t8/g7QFOJ+8WDFtcEwkJooO2//rBgLH5/4gQ7
2M86L1klPnvW5wmV+cRAgoJwQ6tPjOxqS9hV83BHivcsJWNuivi2IZxc5PU1yOUmbvS0yWfGi69P
PyaqtdVC0K1xGWZWM+IcH5A+5l7+WYzmvGqCzmaUqCC8xbfvGBQDBWp8GcsHXTmHv1nXa2wBcach
s+TLNcCoIoOtJOESttulp2K7GE+JDpUcqmCN/WR4jF1qAAVnTtNLxEmE54SWEU5alh9v0dbmGPYv
K7ULN6m+Ssgp4DH3yk2b3oHvfEm22rwVlORuZ9LR9JXeV4fq2eicuBlRYhUJsK2N7ho/8fjSapec
JRGxoujVBM2LG66Er5U89oIznNGZssopbSydoQMPF0+ubxzbRdCG+0MweA8AnjkOg7R70RiQNEd5
QQFM5LCyHGlGfA7/1XJe1m5wFVYBiTdVGXzdKme4zQTzVK7xjutqu1AwFMozmlGO9Z66hZWrhn6G
E3BpUNUM+VZtJ/N0LXM3CjrgT4gyim9iSmWmfArzQTPh+wKGDytTNlKWQAuBHXJ0QoMcHPA0hIRI
MO3eaIgV6CjDZz67x2+ZpcDRDO09vUCkjizg9LOzmsFCzbMfvi+0H/h+QmJGwFWwmDq0e4+Fibvq
pOB9Pcdi/uXXaemNmkYzyt6RFmXCLJxFmdK1CuIIHmdRiGz9s08LBbvC3wsM871PooAEqd45bfH9
BQRURsjn/NNSnRrlfoVKsH7YtbPuE5aUcly5ba5N1j4/yZY8LTi8LjKfmk2IWac6WdljHGA4TdwD
jaiGg/ms/2ZmaoFNImTtWCzvbu3+E2+qKqOgI0QKzy+2Udn8zWNOz7U5EWS9O4K+AKBflydORoB/
ZwNW6T/rwg/SrAsCDZGMaOTE7A3YlN7sBeoy1DMSSn0/0oXkbsJ6xtscOVbYWpYJEz8ICJQSsl4D
ozB0WfYnGDvQQDvfiyKNsfMVS7r0TPQRZ0o9uOlQi6tFTS5GA2oLhRvm0cJLq9kyhbWW4CH7z35c
ZnVI1VrfSER23x1f7TP+xzlblhd/njjQRJNXT7lnU+on4CFFyhisrxD8TLhAkQzXIuQZwt58miEp
2CfhYkQNfpBrRe9kBYm5Z1asXw70cYCx4JduaK02b0flA+y5j02Zcz9KYIVFaxtdoem8L5h9TBWo
SnGyPJyvlDtAWdo7SFX+p1rGXVAEZY6Vr6lnwLEf5EJonExMgdwidh05ASMU13gFWyGTEp49fXzO
gMgxyt1WXGot+a44oBNVkTVynD2umMZsmXD3+82WtRW0dtzNqL3fEmTeVeKQNQ2VpYPMqPJWNu4a
g3AKLR4vJZJfBG85QM4aThrsF30dH1JTO0x1Zi8nFqLFUtHe9cWjY/NMqnokzOaH8CfmaQRNjZBr
fb+LA77NzLP+aOAHfR4HBl4tkR7619oiqq+AnJi+KRICOSWBBb3PIEYuSWoZFi9R5EhUPcEqItzu
LpTbghtMFCe7XjrcL2z7pEdVFBha22PnTQBb+cmevg68Is1RMVBKEzCxONC9xTUUtwFX+Cd4l/ll
Uz0xscClUpqtGyN75IkNjR5xtqkhCldvm614QOIMrQa+lWK2ahjVRxzc7gZ+qVGbJrCtge32Gh3V
tnzVZpJPEK27Il76Xy4/EVeyj63KSfXVrraIVtxVm5zmNa2dVulyKUHGt8X5x78dli/4TLgCR902
HPL0hez2IMFSUN9S2k8jL3fuqbHTa6HApw9Ev2po0Bkc6B+qNgLxphqx/qBfOa3olNJKvU0sGdZh
KsD0GOrxrxqTwI7nmDfqV2JPBl4fQtu6t/7VoZfMoMZAwu9Fu0fBJPQr0CumHjK7rvxMfOsNQQha
bEIrmiY7UPaPV/1qbIp0Z8PN68NO1CNU5IayXslaAqPyWZqXKRK6YmKKMpW0AwxWJN0ywMzQ9zRv
ZGNuS1k8SJxcXdlTCdnf4YVx5Rn6HRtfgSoqCWLnuzX4k2Rhu/n+/SgO4WhX5yYzKzKXddUta5rF
kxQwoEV1tWoULdWxhQ+45gqJP8vd/Ah4Uvv0ea3eTMpS/7v4CrHXZ7ZLvc4bqGECJzzHwEN7VzPz
Hd33uuruaHyyTwUBg3QSmjCnEbmAcSz7QxEOYWwX1Mjog9iUzZxtmoC6Q7xK+CGcJWfQvR3tmrnT
2jOcqJ892VySygzVf2Bwp3Pv5ewwGDYAku/+d8Q6NX6440HTIB7Laq9zmxE0CmBPo87I4Y1DETOq
WdIm2+XzNXiWeIRKXIp+IaNLw51w39TWVSZutDy0KmlSm/Fdb/oKXQO+btihnXFqoUhe23cPNu4W
GqMb8Gm76NIsy1Xmj+uvxJ/QVnByzLL8FhDejHgfRdOp/rRGfaXSojJtUfID34aq4adRl97f+Fky
HQgXQwsa9Kyg/E9TW8CyaMwH4yLM+bseNOKXoPxcRAvmDsW7yPaPOrjxJW5sjw8RgkV1YtUuBkxS
YrV+Y08Y6i5aHAJPm7tO0BozInv2Rx9wzoNQImP/G5ZowCRU+Dk8wzqxUv5T74hDe/A7MImlmHbI
8yIp3VhhI5yWX0cFrz+jxeqDhuGOXx6JPrmehrxro3TU/BpTI4RpXcWsCcDmdMJuXDN3sqvrAlTO
mJRuHCB3DM2IBV5uAgFnFMSJMSZ7qPCGGm8Jk+vEV/mplFGF8c7ocLJmG8+PMltEJozZLAnF+zsO
2KemMf+iViEjxbjBtXr6wsB6T4T57/8sNOECo23cD1ilxprJQQfHLeN4Yuv3tfuuPejvZzOgFHaq
gku6230lm4FiXgttEBtCX2LpogPM4JEyFXCc1QG9HDhUySYKYmeMT7xRj/AD4z36ELw5eiAT1VEq
u///Js0+W2U55uvNRbE4IdqhZ/jhNz4urVDmiM6kgfH2ONC2zYriD3aDZuqeTlBpQVxOnj0SIAPH
ZVG18QpACFngSqFBR9doz5mP0hmPoUwnPwTILtEGCGf+8zTk+FU36NvKqZcGlUA05XzH+bmMYxsx
Ok+4tzG59tsjJQzsGcsTUbMRdOjMFr1zn0EbOSItvGrkwU2NrPffQoKpLIx5BUnGN9EEN6R9jDqD
O5A1PsxF9Pirzzx1t9qAJU8Fds5cngSaElwHpBJm1RpjUL8RVevQGaQfWEyRDj6t2j8jMZykdqX5
CWrMzb3/G4h0J7Pyk4YcAdR14KXz5NwXD9OAERtEbPvXtlaP5/7vCMiIXAoHkSgaD8YyQsLbYdHl
274LV10TyutEmtrWq2Zay0C5pXoxpQ16cvHFjLMI8IzSdnFblo04NtlVPrAberV8wH2jR9C5UwV1
wpNza5GW4uEk871ecbIjGdvGA4pGdJ11n0UFgOtEqs2lZpVAMKk4KZEuwTpR5zsVKToZImBmiSBi
BuxkfyKuNLOEYOmHkQ/bvmPXotFIry9d7Wl9UTVzX7whsq1df/MD62roV2RiEdO4e97YfKIoZceY
iMGsSDJ3KMBrASlA7gQTDFSPymnyQxoasLuHJS/+4EU9mRSaQrfeCNSlN+VwrcS/IGFbQzbpPpUM
18jFkEozHsNfgmKQAGgnnHZ0px9hmtdeZX53+wwu3RIcsCQD2TkvIec4nerEXyCy/wsySM/RKDzR
sholUpfWrCkpthU7cohBPV1OvTmRiCKL+CLMxBOsbmydfRl2jfWRV212H9Vn2RPMmeoiNfeqbYcS
g/IF1EVsdQww8yKPO587z7QKVJMyDqDe3L3opEPHA6MG0TZVbT4TkgEfhirTXzRFejZIQfA72kYz
JAvksbiBoQ2RhbDNoZSHSvbt1U9Pwe3lNpU8SjK8rEbzKAjaX4eTksnaQDWr1ALLXxwww4JHfjvy
hPMGDjmfdndeu3aejc9rcEbH1sHEDtCfOTwhe+TsKNCj359YceKVeqeFRXAiSEEYgMijB//Q+7nw
qA0t8lZqJ8GpVoK7bwNvBB2qJ3x8ocLcH7K45pNZNr5I2puKSl3nr9qZwIPyIqYklEwUSrnXZvBZ
ynRgXJXPLWAoZlrzl7IZy8nG1hdyd3KK32kpRwXMiwehnKp+yAbAzuWl6GS0CAVZ58OhQxvzYxYE
6pT49qmpOShb//9ME6k/zDINbidWElyRNKB47OLbw1w6JtCBFxVfiD7jviGDPWjUVV2Wxiv7sqSx
9kO3ifeWV+L89FnTzkqD0I+VjIoQIBCVG/oa71Di5kE2J/qC9B1kM/Fxru7ZVCM1rvbt8RWPFkRI
6kadSgX/jydKMj+wQvJLA5YExM/mJYuy/joSnULGxOE1+2yo1ZlgcglwaK7iqOqJhts7KGxihzhB
gFExJjGmSVkKbXcuKN4gPuOEZN96PYGA5mdDNpRTOcZBeuff75k/XsrAu/qJYfuTer28tcTiBqXx
sZKQWmrNv+6iyC9vbpWWLrUg7sGOqBD9/se8Tr7x6frXRySiabRJH9Xf7NLPYu3V06pRVUebtjYM
ZGKvLdUg1O9Or5MZl/M/WzJtdF5nHDQ4SbjLCzk/fGnx+J0Ke2QkswB/84Q4TMoaHORxjJ/z17SA
32X07QZ3hgrmVocEyceitE+FAktN0gBvTURq+y6izu4ip/CfkulELKaMqTyQF19RAaNN8z10EDQJ
lu6bqO6dmabZGGXbnYQsCJ8x8JAFq7rnm+rqy8kpOl/NqjYfs1qWgpru7+oZCehI4tgLUNbFcmzP
habNC6O5ihol02mPPlHJO2fw5H1re1TVG1v58tStJlUtOq2kLHwcS76lJsWB9wqLWshZ5gQcoXUR
Pnl2u/5gNxy+6oHKB/YCljWNekSyKgSm+p52xKYryKh8BrqHwYzgnxsl3vr/90rUDpD8ywBsVkKx
MirrnWtICAQ2BakKlj5vsa5ZxozgbUYv8DBDUU//xoyX1cokKrnQ1mmnewpoQy5fcpfTFFRqD67s
pkmZ7LTbCxXhCfwLUeY5Pe2cNdEQxYu0p9tDaMAdEk/0MtfWzpsyqsN27hfHGY60vriv0haCiwCn
Xtp+xs69cHBCWt05EQ291ezFxG8hchzp1Ah8wPAxt+IbNlQRjSjqJWltD0+875wJ4LKsP7wFJjI5
n3dF+uaYMYhB3/FgJwFUYiFjJN9n71R/rmVX9c1O4eMPxkEHs5nZ0dkGecLulmGrheavx6MMgXlS
C024RFYK+aoIDX9x2zxZwNxJTZMNLsOy7N6YM0noWYnhUwEaKLZ/qjLrntVnATFWZ2o+YBnBwdJq
VXSZvt3IjSl0Lv141QKuMz8uwRJZF308oh171IkXx/Gh7ZR2QfdrUOeAIPAWvtmYTy9V7t/rJFaz
eW/laorBZSKvPFgKj0vDRPB9WDXFEnLwP5ZtVpDlXHxvpFQxWuipcFJM9nacEyO8F8pzs7C9hiff
/Qg0KMkJj27Ao3eFm6kEHnQJeZvZViwhs207tDZ36bMFRSsDrBdVWBhGxpaj8Oq8HAtHdUCgvpVB
MILf+BbjGbwqPGtl7dh04weJwGEu45Bzbzx6UYo2ZSBoI3z0Ywv/r2jnkTicdAlJMld0xHcnASmT
JxNm3bea8oDZEghNajaFRSVENL4x6f97gqX1pQp6Wj3XZ0qh9Ay1ri3mg3NQO6XuuNbOBVjzWknm
zCcFZ0yYJMlzdLkTFrLigZXvDnIZ5wOl4oMWjrj925Z2e1oi/PF8IeoXd/VVg34DzPfsmIhqygfT
e3p9och/2VDHAGTskhkMZXCHmKpk1f37zo4ENkJaR3vROVfomOnePFbQER3wtp8hA/g6PPZzemkT
Cod92DXripwIoE41OYbry5YLWjmgSHyRPIPsdDK+//LK3Fo/R0LHiI3cUOM6bNdLwK7JsPXPqdgc
DfnNYNyofXrzA3GFNLgKwReZ9/4DaJXJFZhhrvtR6U3i0HHRrrFTexfbvwYnBNZNcSwWLnN1+yP1
2HcylgX1ocOoa9St9stgmBWhUqJ27DS7y3mNJIK+f0XYl+zeAqVZy1zoIB67YR7CxMjIF2FFBiMN
Qw/2PMHWI1/72RINcmwJPiXABHJ26Je1W0cuT1Asn4mphTqOv1xZC7m7rb9jylhBEClcYd2L31qN
tjnLVtdoq4588cOccvE30TNvzDTYgDs5WrXFAw67YUwcvId8WgYK7ZiDvGSUSbf5KxmntxgCdhWR
9z++OEwU8sSPvDXlSFHB4e8Qd52OMXyvpuXJK5xKYW963ix6ZjXY9ESy798GPFlsAs3tDRrMuNr/
+vzCAyET5z/1TBKB3+26bPUb5+IguMqL47d47pXzvoIGCSYBoOQ9WK4WHPH2xFi4iokDmKSgQ8sy
A6L/UpVZMxglUrK1Qvua6rF+KjAYGN/S4qOYf2Fx9FLmCGuDB/7ZLKR68WhRoyRR0IzkQXyQ5bik
J5C4KiUbdVrYa5bKfQ7QhxOtnrxJOjjQLfzEYVRSyWAbhptK21WFiBpEOrT4TlkjMBaCFdPiPYq8
QPOMClEO03QAZopJihJCA9UUriaavrUGCqf8bqLfIw3ilcLjJM/K7zWvO81K7deQV2hh9oHpPMgm
+jPXmvWEri9NScvEwQcMyvTcFpQ9JjiORZJ8S2as47G+AAeKNDvzv2QY9q4YFX5Hd3WMadtNRzO7
pjHq1Q2gKjlE+MeUEwWuXkBJOXohxNcyx2nPhxxuvqkaKENwbRGiRetUcQmQwpBhjiVza0D2Eg5X
PpXLIo+/yF6d7GvaBLFPAvwGCxfwqQ2PG9rtO7GKFtu1pd+zerBK7zUtBh8gktnISYd7qV3jmC5J
Vx+KMeG0/4bZiBtTXImgd2s2mhS6ezzx81wr5z5i9XprRrQ6BpFywhnLy5Gh5eBcLhChJCtEEW28
kx8Q6iAk5VzCEuoyCWEXxW9RT73e5aUBHIBkoejHd8WB9+c4EPr9A0E4pIwAmietKqy4Ar4ZA6fu
ZMCymIU4WZKnmdEIAm6pV5x88zU99z2LSOv5oXgoxliXctoK5o7I/t0ZTD6bIph3CmJgrq3pu3dh
PSHnVdfC5CGJhuaWnBgSw+vVPn1Lc+PEd24U16Ma3h6ovspps6cOpYS+rtaddPodnxaLMXPBFEU6
hjqsG0cBsUKVf30P/mEe2k8RU67zBKpbsv5H3YZVt9oq4mGo1PvEWbRPbb7XT1SYPjjKN7y46JWv
ilQeYtXs0i+u7F/PWjdPA7SEnpH6ONefWaiZE2FIh7UKjCwAqBuDABtItJktt8sh/n21VFL4+PBF
V2d6Fp41+xlNeYEhIoJOmRX9La9h21hbtud0SDhBE9cgfF/13ZaRB9K94qMJ5XRxYAVqqiq4MMsm
Hu9x3Z3+64pnGK7zSn01mz4Z1IoIih/pa1jdkp5dtN7Tkp/yfXxQceOdIzfOh8+2YmcvFJQ3BuE0
jbPDVhxw+PGuH7cxgBM464ZFcPYEcKfpa2F1rfOLXJ7hKoGkkSy25rVGqi5kg/1Q+0iLM7afVXLn
ZffTC1Im/SPClLwRYsKoTyAy7x+FG+p20XHjuqnCasW6ef6JtDJrvYeXFq0hCMw3wNECLQnrbAxX
mA2fUCzOAC/lnwIN2zz/lBtq2OMTbxLitPqmmjs6p1kSSIGk5OMLSVZJAj7qUw31enOJt2VnnOmw
5fsfeioZQ4lSMMwGRT+d7sMT0+K2o4A3iaXnOODPEgvkXeYi3btUxWzLxSgEKKg4zB7+YIAfyZx+
Dj1QH2PGzYx1hnWs9NbNR2YL3YpKQNVItomn0bOkI0nHnM6f2RDNlXWgL6Jx25RI2sFfCV/UVMDp
2OAcN+5S/W+vaj182k5c84xeYt7qyj/aJzIxP2qSq/eBTSAyrj/h4VS3ajD6O2Jq9tOgEFWWtpZ1
xhz2Yo+RuCcG6+6r4zZ3uN2bh7CGrpQpsG6T+BEn6lenCQkjWzVg6puWupXO55le38hQOTDCsbf4
8EWLqP74qNnOgXmGl6Qe1mU1pPaB3pkdGWr1Ny2wAg4eTysGYLsnKa5i2FI3XH5rYABtvaVZV4aT
HKcb7XIJgEdniI+D7gyogsIzut/iYeVak8MmPTLbFtWnwNrV1TBHOLFEx3uqbrSyEcDnVtt8P68e
2mkbO9C561mkrjviZGQBdfDz/i0PISh20RxeSaUVyNMArd3Tp+vhtot1PPJFWOzv6c1ic2NL2QGP
BzgkyV2y/WrnMs8qu+vTT8sBvJ7nzgGoOinpcrWDdJrb0rGrYcwnp5nTiX06Fzg1eefVrcXiQJ5B
HWsaQsX2nBKYVtrgjQWZDUOkefIDOCwKf5pDytYYeV5IiFjA11UROyeoRo2K40MEPGQJJADx9CMZ
DBR9VvpL/qeqCpeMtDrUgDWMcRQ4WRUhUtQkshWinv/6p9E2YLi11Tu+Hh+zLQm7YCi1FTA6YPFN
w/DDSxADYPd7w2ica97riONkZxZeQHE7nOohKl6KFT1FqVcdE61f8YbnD4s/RaIpyjIEBDZOW14K
CDp8DAweMnOLBc26D6b9ZHNfraNXopgcrugqjbX4Rqs4x+Q0OPLcfz/KVR9/jrHyBh9c1I++cnyj
n+EKUzYyNUi/SdOIX2rFcraYqPQ/yXgTMyn6U45o8SWo/R5OiTo31UwnkSrNFMG0psf4QqRKgIYq
vL8Taig+h8wXpZsXbcMN2TAQmkJ5TjZnEwmHSoRCVt75CutjCyGP8yKvt2cuNIR92mcNAk/MG57U
kJT81rmfvyWMf/ku3P+2KO75N61+i/m1AC4e0gII6ZcFqz/0Yujw1k0NN5EoDLG4ZyUHyzx+Y+AO
qKop3iXTaz1WZmGKDu21jmcjzIg5zQiX7qzOjGbIl+4B+rUfZrsGCFeIx6N/kZVuh4h7W5n1vGPQ
O/bdv5U3lLYL7IvRZ4BCy7aNTYk7XlGADHXGXU1Fqo0s0sCfEBUeMwLzMGwCs6Qi2fZHGGKFI4fb
LZKzSYrl5g3jsgWW2E3KDqIEA2kPQ0todPNcBOk0ceFcCWHvuoazDidJwIESGak/2Vmuu/TnN2Ag
DfR6SaLMjburwyaRS+rJNcAEFUzzU9gGQhAwDHAGsHTy+kKnK9sPGNjP2xHWKDymwQfhzCVvVdy4
NCxH9mIR+hS92UqfUqSoO5kt6+A76uXooiDKVEqV3IHnEdfYlCs9eOICcMYeBMGNSxf8cLRkUZ9P
nVncEESvDU8dmp7aKgwMQ9D8h27FgePZF8nDeipH7o2NBpo/dWcl1y+l//b/qJf00UYwWzpgZ+5u
7CtNvMyYCxVBZyxpVjFz4xfXRXm4eb7Os0TYL8lZblLhkeND3XlH3R32LUc+2e0tFzvgu+Nbcv1H
qTrGn7ACVsZvX8Vx9fhD7ohUNdfW5R4JIiRMOZB/eawSc4BVQDF2YfdBKix+zXFdeAkiU1KIRMMc
Yp5fCS1r1p3Bn7xWbd31WM0JALYpVTYESanvENce788kYRT+CMsSDX21DN6ikPzyBoZFiBN3ZHpj
KCLzdDoHSkxSxej1gkRAeeixahS6l8Pxq2ONlvSVGMOO7AGwB4bBwRNThXJFMb3nyOZy9MBLnTWD
oNyGf9bfg7IekCTPZHIHPU3tc7O36w6bUFnXWvSAmzOeWwVyvSMkSyzGS1DE9D+UBWbCJfgL6s4B
WfOZwsmfP0y/3/CYWl9E7D7GaZqINDP1CPoDd3klxIVFMAHI4amNI4KM4i1sKAKjh/bl+Ip7HHn3
RWRoXPqO2o2XOSB3yOuuRwRnQrcddZ4NgQFtZLtdjYVHy45Bow1Tw5MEWHro1IdF9w6uCtAD4zG1
G4qXPxlT0RmRLkC4qmGvrGa1PFh7qN/3Cn42qjBKW8pIHAOjvvYeNuTwvz/jXY00Y2/I+sjoI9Qq
7mnA6phPuupmFV5++QTx3Y6O9e6UtdwlboLwUpZWn+7OfFz5DrMpGZgNwHJaRbIJsO9C4X0zQsJX
grUjsZi1Yi0hTZTbSSNKF7xBF1wpoHcE0OaCDrsYtlt+VHOoNzrQaUamFIWLxrM5J3DKZsTsxf23
3puT41pP6g92JN08rK/JCJqIVEgRROQ6NfINg1rkYD9fEcE3geri5nxcONjvJ8N1+NqIW+dGEyov
dF7I/+CGbNBg+pelQNeedSh91LYNXx5YzoiVDndcw0yjxYW+VXQlx6GdVXewxxaJXHrCiXJptpBG
VA+pJFienztsMd6j0c1GfBxqjlsyifqTIo+H9itjRnyP6PebaBK8oN5c+WvI8Afs1V+2l0Zeuq0L
P0G59nBuzEzo8nLI5uDk6qVFTxRQqk8BmRmJ9pH84Zmch4IyqiXyE0+ThXE1SgcU9n0KQ7uYHeG1
HK5ctOHfnDVOmDftzEeyi7jc2z+A5zdphWs7in/SPy70gQXaRr8kYy5OdYgnc0BfXksjvWSX2b9E
F7icGKcFK1iv6CJpth5/1TW3aiCLXHCD+lOPcW6sKWHWOzTihFZokfH7oRx55lO/jT6L2MsZsiM2
vW+vswj44LHQZhK23tMVk0GX4KgFsm3KnYIW/KY3AOmeNMWuY95kSKKtlFZiX+aZnWQMHyMCVTla
vQ8wcy2tlLM1o4tjX5pzBBoeYAqMNFtxzc5ZFcoZJpcHy/JNPfAwEHOV+VD8o48cIaZVQ33JFCuU
xeUz4hC+YcjD+/jJ1Pub7aTx8RUDj6MSiw+1jfHrs4UzopQ7R0E6NyMI8sRjx1bYoKHmZ0XlT9+g
Dp3XPp4Hfjwyblm+6OHE4jYYjYGuZc4pfwB4e3Qqr5RgGc2H4Qq3h/iZiksNJ7+yYg+L80YNLf50
9ZSsF3UEh5RwinByBpPiGNyt4MeuM7cEx2vcIxAotR682cRQHXgAR17SWlIzxrzGDXaE3k0fpwmZ
HeTdEPVSefh9HOXTSVBrTQhMPWnANUYAF6PxbUqts/Q1NDvaGQecELRD/F6KyNCDSWgUKcdls8b6
b7Qv2ol3D338CHhsifuYq21ShmnhGvXPz1edlE079K97YWCjFWcYIXVMAYgmNK5BO5YsQvRnmn4U
LkTTv1+oKrSXsE54QJPArtzsg8dvYqPiJ8LkCm8slacKDjxqmInogfKIsUQTP0AqfrD5pYoRxOlf
H5HGN/U1YJtt2gLkYjfMV3B7GQkU+ZKO+iVntBh5XjzUBjxAVrBx8hWbwXX4sQlk6/rwms7dA2B8
zNWaMWrnFPxmHwQZhqSfO82pf561UcLVZCas1HNm+nhFwqaKFt5h46/gs7SWSfO57Ncjj9eVcBf1
3Gbs1fZM5qX0cJoBlghCue18/+84gv6XhD53IfWTNiAWVo6fzLn0+S8fkrQMGVWVdnly3BAOmWt1
/B8pSgRMkcyWTpzwE1NbIRvbcaYyNv4ACz2XCnZiSmt4YzW2H1mQrgeuEgw7gOHFtukly4+GrYAk
NE12qK5OrpZM98sn/4V2eD1S9pZhSK/4aeeRQ3HsKoZugZpP1e+a7ZYg/46FBw3DYN1jCuxKd9ig
/cbB33wHggSl0T0XU5ZHWznpnRSj45nfhk1FGNTQgShjckyatVoogbmuqBTrNhPoR768z2weUihM
REQ33RWkR3WN723P8GPgUfGkOCPwhYdAvJ2Ox9LUFw7bcrJ+HHCg2KcweHbVIKiRP8/cujozrxF2
n8csSLPYCAE96Hk3zlu9h30Lsf7ab8IKCbc8oRMGvL9ApEOihIK+xl0ljZd8jnpBH6xQw0Va7GlF
ITnMyC+HZdgOUasj/Hr1/ojjueVwqZWWYgaiq1NXG2ZT8HgR8Fue1v4abdhbCyzIIEqOZHWzxo9J
N3pnHfB+mKFWjfEHHI10S7t+PYfQcjaAVMTxHGW4GDfzIBVF25WyXfMyXyB6ng8FPh5FcC1nknBO
CoUE0skye5+0nxG+Z5hf9lpzQFNxlbuPEEupXB2943H/WFK4k4Fmh8AIwyL6nHYGWaon2x/E1Z4t
7UG0mjptOMoc90oA1GTQ8mO/oicZ0KfA14CH2OvedLVXtr9zSFltESE73eZ4nEwilD0evF8pYjhC
tDnRFF9xyOEemX7l+nl7aDxadaN9v4fcOPssaCxCfVaF+o6RXHvRD25c3OlL9nRH9IeQvl1V/eyU
M2m3rk9I8XPlykP5Xy1BjHHEmTrvLOeNmvF3/JcNOru9Ai9Tt7f594XzfW+0Gy2cLvxoWhUNUKXq
YDtBD8CoFjVP8pgOr6ei7bQYVsQIe79et8f+tAFIeB5Djm0Rka1w7g2zlelSPmaWlAMWqWa4SWC9
VK8P4yn369q6icS9SapLyCAEudJqF0SOVB/MPNI3T+no2Rm/dGUkRx4TECP7iEs7LqXaaqefGJEN
r6RBoQydnxoWtIpXICghl9hVSdpgcxhKXqBkAKuGrvktnfPCYfcRZd2RlhEOloVLcQeSjknQK54I
V/YqQQFRCvebwTKY2GY5bghzer4R3cLa2p11nYCd7HYf6djId31QdDw+lXFXH3cPr7tUdJ6wwNwV
0SYy5IeE15skYcPnOC/EpMd3UmIbtYhHjqnDiLz9dVme3HpruJZ1yMRur2jbIy56psRbHxbmWyBt
z9UQjex5qB8UTMk+Ms5dglSBVahbkLRkvyihS+ek+xH3oJO/i/xfnF/sgrHrzicRUDlbDElxgEb5
yCnzGzLvULSEBzBjP58KywQdARBvo2F2CSYp4b3tOXeUCiCykVXXmtVHRJ7iS7FxwF3lINn61DAA
LC0ohZv4tUefDx13SkqX2qJs8GLjVH+4whDeC300IP4nnCAAPEmjDSQcWmmulA/lOMSWCcwomYfe
raFq0ZdwZ/rwuBajn6WVC567a6WIC5dXnbkx9DHdkSVUNnWaiPweZdBmg3XQJoSy/aXKuSiMGHtL
BvocbTIT2swmCaRqyo9h0DiuTDMLw9a8SeBuBdIfGEFAp2y8EXKtMI6Vf0Qd8geKL2XfbnQsTaYN
/RgsHooWvXkV28IwfqBvZmyuyCoaZ/JSQ1Z1yT2rbweZgYP9ULv5EUAKXOBzhYclg+3hdLuqTlcB
GThM+ijCNrTRGQ0YbnyQEkkRrsxwnCLpbpE9wn7s2MAg+dEaE4E0lgaju3ulxlnXk3Ke0Vn+VdRE
sulwmWqBxb/tTf4XQrdre+hIEH431+7Fa4NsvpCvXouIT50v8bPQBe/x/LWpO5Mzxcw0JVJMYEvO
i9Rbs/lpQauAPXZAtXuP7DyzBfCo777LERxFwCw05kZ1mErBV16GjGmIcyU+jeYFMzAoyzbaykxX
DD+fdQbO1C/NhyUM4yI+IZZNlMZaL3TkiPcUbzgxx1bhfzgiufvo1mmTxUq+Zj9XZC3pxeIMvVSH
vg6VkBz0YfuK1+NXF0ZzNnYVAAbYIJiixP2scrItcRmYE+Nyy8aMzFS/8DnYw7mFcFzjRl2ncRrm
jiW3wKgz3r0jwZTA58dEBZ0FqmS1OhU7GAntVfrs4tgGaWAVhue8lkLO8aDMWDI6aud4YlPBD5I1
PP1Bp+tQCDSpdntGbW+01S2zKXqrhrNi1zM79WY1uGdD0D+JmyOvLPDaxE6GkVsgMu7hXVAXDC+U
qw41z1AmWSmMjVthZiNAlqg18KGwVn53QX9IVQ6EyPFnZtrchSbOMV60faoZCopXi5lpkV2YtXjq
shIlIANdQnkO+LTicFg9IEDEUEqEMjPhT4alLxUBg7mJWHceFL2KXurjjf1gDXTovMCi7Dpy5kZd
TcXradV2lZdV5nBAKxTbUBA8cQauarF9cQU23KG9VlQwHO39FX59S+8DKg21U4pxCrEPtEkhkzuS
zIOZA49SP1ivmsblttMkael4bGPl42T61HEs6WIRgQAcR19wKw1i/KxPNCecP/ftNiKndv3suqKI
gl0MsA5J5ts2RnNUlEYyGC6+9OPLOpOND3GC6yaN/2TI/y36PJ25StM8C3yRU90/8F0+TC95v+ql
Z+OzwuKA5q1bP5HnkbgqTutPY7EaeECIiDC9JFEKq/JuSxrEzjIdugDjvjYSTuO1SYSIC5nl504I
lup3dMeAtRGvCKrqPkXClPMgwGsFiMWkkoqPMaH3zBOFeqjYs1VL6BkRCGLwMzdJhJsXbrKG4PRe
X/9fy0o0F7n/OAYIg2L7uKPMBtVki1qu9lEzY8G1Bh40biACg/+ouVV2m1+4O2ZpBZkGE0jC+lqD
wlzo9nQqIVEosoEu9D8e//Dkmbr8zMNnApdZjpz2lbJKg1Xs+YgLocFMrzaYp3ECLnJvZMaZJBhH
hStSTRSgNEn+9bRLig+1yA0j4mFbeuyaNH42CU7fKqoLOEWorI8gM4WO/VwMBUxdqo/VaadKE6jZ
xb+wMpwTj+kHNi6C0LOEfH7VIUYr79pIloUgHKJ/x4C0VLnJMT8dMvNBzES8XCEdO7IQPI0VZosq
u0GFye+4VrXV2Hm3KvvgvyCcssSb9oo64PbOzxiNbiV6vnty8SXVV+JxwNRIrWmB5mozW2C0xg22
AwBbpsES1mb7o6L2mN+hbB+I7712zpPpJY+idLYpkApGNjgsjoF0Bs1iFb2miXnlBftejviWpyQC
htlQy20wl4E2aeIp/+WfAMlIVoqEJux5lpTUqIsfj+PiyRzuyz+XokFeD/y0ecG4FzRRkYgvm38E
ZqtiS9zfsaMa6QsCfzGF92AMeY7BxahgGFGm9I0Ap7frIOSHkUhoUi0XxmqYraIv08e4GGIl1upi
ubCuINDaPsSaZRiec5KW90cttlC1raEC6ZN9uOgQ+Vovyjc3BvmOstsF68fmAqh7up6ur5zXsFPV
j/I85P0PPL2swEJbWnbc9RQRrMUDFEysLa3ciqvNb/FPAPOqg98Nau9MxJNxkP3+wZEB8u3B0PMP
qQXU8igQIIYy+mVpMDPgXEZIB3dSrb33KXr5fArkYaG+IqkizHOPYRiCaZS/x7UHyUKnwr/7ELFl
9pa8WW9S6eL5yA1MkUNfLNqNW0NAlAei5XST3lTHtGLe5G3v4juWX7HJi4yWcOXV+JEAKR7RuXLP
T6lQlAf408tOHVW5BWblnTCdfK8j4lvSTdL0Wi582HZUTJKjyWQZmPnio1BUS2WR1/OQgkSsbf3K
Cs7Z7oHoKn1KDOvkIEE6BzV/Jl4/ZlD144fSjs+JZqn6H6iw+flGWGlmpYn0KZTq66eaNShIidvd
7OmbYoj8f2S0HgG863CkKvKFjdPdt09TOxldYBfrt1ESnZPGfMmmfmsYvldUW5VTeyUIRTftYTr4
AVexr1FJa/0lhpuYpfBOM5ukKBG5ApDtTPe2FNDlCTYDkREwT+8Qqbdzxpw1rHu7x6Hq3eIr9qLM
SV1H+8EWgMnjzbvfcOw1D8qVe87vKlnvbuIN3Qmvea4K0YUMJPJpe5+HgmBPryZh6CJQqhyd5N7o
nZ/TfeTRy5q0o/2zo31ytdMSEYvnuiWWpTISAVoKmA9qXYrL4NYAfN8to0FqTfQcHstDJa/O32Qa
fGiLowf1/wxifndEtY9iWKgLPvRHlvUuKF7ZOeIcBRuQH/Lj+8ssvFgApPHYB1bMSxcL7QYy5uKv
Bi1UFlw/Zk/+go8sC13vuRC9MawqM4V+vFYKBk7GzxIW/B4E9gdUX2MHeyNIL5K2+tYwHEqtfYgu
3Qse1hLMEIDBeBShgjOaa999cTBswS2/ME58/nlwojVr71Jf77Iq9bvNqE3mp1T3kOTkFIaXXya9
EvUrlAJcBfGz4OnTjFJDyyi/DkPomFFCZfr+cjrfskR6gl2BwkyTcmoYNtMldEcKhWfUV7IpGKkB
is9a+7uDt9HQEaVbG54Osbx8lwjiwVHAbxWm+zqhmolHx7pksMb7Uza+soaUK4KTLQjS1vdmUAYU
xbuwBbf97nQ37kjowEZdXZb//YcOrTc5vI7L4+2rMm7eIzUa9KqCswt6AaMKknYNg3bTacu1RlRS
6dTNZRAbqR9Iunq2k6TEC+AiXzxIgRD1BQLzkAfk15R/H9NyZuE3NkV/HmikJ4GYtG/QJ7NlXfYB
9tBBBgLtfWAB70a4A4c/GZP0uyKLQKZkVUonpFVFQ7WAzMLahSX394Ni+x+GTMfUwI3DdYq3Ou7+
zwbAguWxdw5CVH2QYHlCPjahDbd9Ag0KwPdqxeCFsKid4n1WbxiHDoYBhG//ehxfIcFBEHZ26kSD
BConkRha2ws2QYyVreao9wyU7x7dkU/5EBck9f9w2fc8AAhXcNjBLXP14RysO3oBoBKiN3tFE1uq
xCKUVGlNOe7E+Gmqe56WZ9oE/1Cz87nt2sUajex4Oa92JvtBMdSMBiA/lqyHO3vfPoZlUXvziP7J
mLq472ZHXP/VD0KKb7hGtbhkMIC3DnjagnmaYdwlf4zYkXfveZnaR9KuvUyZOdsnmdnltPADunrI
YTV/W62o73kH4OlXIQyg0Rr3qEsh+xI3KVckWdQkvEhlocF38IpJ/ONC+OIHKShWzCJ6mX96Mtt+
7hR2PuSLKoshNkVgiFkM27Df2ZyKYBg6p1Y+an9ZsB0zdxHG2wdhvK5nwriA1haLDMtQ9LSiZ9aC
qeRXKjsFQPqyoDBlxXnVQ2Ec83Txth9AP4p68zgtZj6xs/+c+w1N5j9KyVeNDtIwoUjCPEJAwz+g
pXTJPvOD+dkWvF2zcB/DCoycwgr13ddBQMT+wwiomkPLLKB6rhoPOBVwQmQhkc3Ue8+g8YFvIzzd
D99bQ/tjMUZhpKZlYiDcE6lxNuAYbGhI1nEhx33kjgRIGD2RgXzV743b+3Gz+pk2OgBmjpaIR2/o
KoMf68jpH4z7BAKv/l8Vj7Y54iL263AgU7nb+GXoGmOhuR3gU113RAsFC+nM36WN0xhnw6PRTyW8
tOc3XZO+fhJn0oWk7cwS+WnTbrbmfwjh80HOwtKMGgolcPjuXWQxUzSF/gAtDUChx0hvh1sNCVXt
xUToboq08cYs0iEGM47eUSdON1x3mV9S2OGpI09byv+jXPrp3xFDtN1l5RBRbtasDUrmSOUvZOHz
w9YoiJFwCGmviTV4JSJKvvfx00Ie5eZEd7Foe/8Iq1CrIM3aJc5MSt5Mmmf25CudO8n4GRTcAX/A
S1QCZVrFwzSAMGZOHnPu9i4kwfhMq4KQtD5UelBgNRvorMANgN/sxTq3tuVlVkUG/02cse6ujCs8
kklfIcgLR6mPmPJnWKFHIjYvL4jw9ZFGjKtjycRr8aR7L2L+mnRc0HWlPDdNyOc/vA3YA/AGk9N0
xU/e7I8TfvEdCfMjdWLB6RtVs1ALHou9V8+6vSOTcAyY/kW8vnK9S2dkTH3DunK/5kRdzqFD7Fa4
IGmSgrhQdrzTM4ZSWLvZfTPKPnjV8juSwVZpXjwjptHpbMkyW7rrrcLXn0Si1yL7UyccTS3Ds+sd
otccdPwOPIH1J/9zzcHQvsohHBAJMY8tmU6jmsE7piZJAAx4Xs63pp/CbdCjKEldbLJxU+xwj03l
Xayi50kFbp/Dy6Sbo2Elf4NUm/0oSDklKYgmB+8neUQCvOTIJddRdstEYyy//Tx37051gNTMOrDS
/K89mboxgKNBtd071EjomG3usPZaIPFB2l/Rg8h6RxfLtuo424N5vhdupyR+WZS96eBe38lHMPgu
nijQ99TbWxvQX5Vk4VVOL8//P8nFz8JBRf1n4pTXMz0gT28GyhG+OHh/2rDO8fgc0w5jXLEXCF8q
HMruRBBTOJY9EugGQC+wmbypgaM/bG5KFmLKOr0KhnuM2v3+E1QqMtitesrKb98KtMv7/J6gW/Nn
DM6zMmEXdvDdVhRW4ima2hgL2aCCKLZtzieh1NJsD3/HBjvYEty3VgNSC3+w77Ze0kw8m4pBhy99
Y6chUoWSFTj4uFiNl6KA985QniTTrgBCdlprVpt0liAU4Ue6aXI14vHyUKwgjqJ8QZZ5rteqXkbC
1jlSm2PwRzJoD0wCUhJsKqivxfxdm4Uad6tq56DLBUI3UjYYvoYPC9cu9IonxwJnVgz6MUTlUnyS
wzPH3HBY7c8sjBGtqjLRdHKpT1PhrZyaHDSgj+EayzWBNu3cVeMt75jGA/N1svrWt79DHKT+QIyM
U/gCGqOva/qa6AwPJf5ogWGzJJwdCfrsWgA5CVh2LFfGPGRqdrzoav9LBdVH7owoV+7zlvrMGDgg
Nju5cfZxg0rdPP9EGPJxwS0TMNQh4Bha0v7pbIhhZiuwQGtFpUUaPCN8TEGErtIPhJ/EZe8H3Osu
Y4BkHe1tWGsP1R39QMCFrkotpDYsF4o3xZrs8sywFAQkHeImrlP3oMaNf4X5SU5fep+N0pfQDNwT
T+ptBYQcP5oVNAE8WNHdTewsLoIPciku3CEp4TVaf7Kkg3/6oGWeLG95YyFd2SUhD2EnNjqVISz/
ZXDNxJs78bnII0hIRTPFgNmIad+3LHuVmHb7lYIbxvey6I3R8+mIzzHZLQk7+ZPuk/OtS4+TANy4
mxAYi6Qs4zGCHGENPKYTrQBvgNwE5QOSm8huXg1SxxECAzcsomgBAWXNzlGMwO4WC15oqnF6NA9b
5MEDk7QNqa+9kQRa196pEmgxzMOhwT4MInKwlr1+dK3QLhYADrfcgffgbqtbUCoP3SL1830ZA436
iC89RQc6w9DEhzGAeG7bloBDvxSOALbi6rKzycDCLz7MIT2/Gx15ITfJfCeNNf6cJWKVkHgGDkem
fDAPQjLAzm9hVe98BZmJsYWehjWzMw5dwJlXEMPG9vS4pJA7lQya+WqrILsPVt7SqHUZ7vG13yce
LBMoF61QbtmivhHdNL5nNB+wSUjYcY9W8HaKlonZhfEtRi+Wwr+DMupTIfO/7kMMlK/UDJk3zcvs
7uxL03gj4nD6q4LA2c9myCkUeSFoiyXJy1eKFe/mV79Mk8fhHs1Rpam0RDzK90F9ov5OalGtlmLR
XAC4yBkaPCWxKk6sgzSHJZwvsnOHenxK3TIjSSKJZXRn7+mjU7wHME/R9TlX2PCMahPxNtU/eq2z
yrqTnrOM9JhgrpRslItaVtOmA4dWNmaZ2Joe5CwqV3HsH0UeQ5bT+AAFZ3pUC2Hf7CNO4bi7z5A9
X9HZvxQOdJ8twwuCx707j8RqI1CcZU4nnpO/mT67mmWeZbDuCw5YQXFvig5xpBH4dGh0UDjUhOHa
0ZR8FswE+pkKOLBX5iSwAIZ/7sFGF7+Ym/NUKOquWbg48EIc6Ms4jchUZpTSzwMN48+9cs4KK0nj
QBxtY+DHFne71Q9pVypIKgNPdSCO0aUJFn8vt/fLGj6FM67QX+eigivuVbW8iimZ2iLsVxZdnlhX
x34qt32hJrtiV16xLSsoHTIAkq7bKE4JCUOrVFJwEpyF1fabC7ogb8C85jbhZKrs/vqK99VMEM9e
pFk3fyyEDKB32T3yRYwc5BYlx3Z44QdbvEnIOE1Q+H6toGVSMfFfMFR2Z21u+2N0GT7ZImRJG8Dl
V+Y44jUhC0qhrS/Rr3k//AHgx0ffhntuM18NmUciHtK61roEW5+0R9l3N8ppgbhIDu4LSIiaw+0+
7dmhdlCQCO+UH4KJdMLnGkfQJEwfWBAc9Zarr4OUOXb6HWtKfz92/jPSG4sSXuOY307Z1rbmKVtJ
tTqZ6JPM38VGJ7KD7WkHaOaZC5Wy6/2KPQuNnZCHraZKFSnm73c1nlYfYzMD9rof0mCph72JjU1G
cYPm2DdX/XwpHmXhXDBbkoUeu3G8lzBEI8SQKYhUIcP479px6b/IosJ1yaWo8gfRX/EtAbVu5fWV
3MPHAHR/ZS/iHNNzk1ZGwNluG/UCpsJrTXy1wWf2uCHa2C2FWIPmb1IPdcserD7TTqqSv3oO1axL
akuDyLcBsos8DSu5iDhM53JIZxrr5iQv//4PuNWMIsun9NPTTTiXo5n5j66URzVu7JgtRd+lY192
TTVE2FUm8Q1IzXkVcXk0AXFiyLJgxgf9YINGIF6UiFL1oxY3DpaIJE6ZwDCUDxc/pdiWS5Yf1P7t
XyZoFpGROxoZALxNHsu648XAnOl3E4ZzesPZExmLN7FAoWIa0mqkAXV3SVeWVq5sdb/to2qHODz1
x8lLXnK/C5ATmOHUOSfUlA5r3ZWWgBrLrFSeE50NtsL3dwwAsg0Fy0vJNK0R0NtxYG0Gj6PMP10b
S9tfECsRd07C5TPjXF+okbCk87czl8MszWhyctaADD608AImRsbXevPb6gZBBj6TbcMIE20hEQ0x
Df9QqEjrT9YQBlZ6Lm3LibC00bbxCeLuodrFzHXM/tv79+iYmuJh2gTiwlH32hS/BRgzlKrtWS2o
QR2oLQzrYbJY1YSJZlsZuBzPbljfSlLrfvHdz02/eiwbYLWI1Y2zZhn3jXProd83Mp/kvqCGCfXd
n8wBWyIbyfW8lAjHy6ccW5YoYSttFhemEkLPHESi+lr8vgrMSxDU073BxpjfYY7ybL2aUYBBXnlG
syXvXHONCx1xHYPEZTNyGbDhVU38mOgNfvzJA4B0w0y2HgLEumXTJp4xhmAJQE8gDE5tCKHSB3ZW
AjeeA50D+47UtALCdEywao+81smEMa9C4k+/OSwUOTjk06HvU524x3umhQjSo8hez/vPNkGq3I0G
KlmFgJ4L6mc4KckNJHZ7RJOcms++WGzR3P6T7pCW3laOJb6EpZ+NX77osicJsXHjnrNGN6MmnGMZ
sP9FBdjJambL9HkrGT6u5hdr57xFiGwigDUnzY316ETIq7GNaLPeXnlNHHC+tpKW6htxQ5T3bHk0
PLlE4yIxZBhoGiGiZk9C5yENW9e2BCuY2ZMGeYwJw/gwpDiGY9dU7J2og3mtZbQyNyKRmdGM/Pt3
L/gnN/HY0GiTGjVqR05AuFAfjdoK9DXCsawlBmswQ0VK2TUJH389N5tI4h3P376aTNhRaJ/lDKv6
CuMBftpMa8g532EePKMyMDx5xuKt5bPlP5NZAU5l6hXOiZH+vaa65rV2aKYF4krvYh5XwnpX81m5
E/ubKxl1cimFJQlgMcm3AuTGyQAt2Gs9sLyxs3rJBVa9/ZkMvR0Qe/wjenpHrVukVJRNM1qNx2xg
8Bg1j7fFkuAvA9QHzimwfUQjLsY14jMwIWJWKVhU8bykifdsfwRp7T3gIY+AJgOWYV2FHs2/dCoz
rQ3BNz/2qTCT5mtuhzcJi0+Jy8CFccSi5YMpw/gi3AZPwqqm63okMdMvdtYt1iG90ERaOgLL4OEz
kHe/uAymzxW2OawpFmCem/iUZeMm8wlrx9D/iow6lVPA3cy7LxJXqTzQwcMe9atPRleEQiuPvbxd
V/j0AjHcjMfWF5LVs9NjczqySxQWPTEc8SF75Jjj23/q3/X9gaCYteBDJUsH+bd96K9+hmP/ZMMY
8zFwb5xWLPvCs2lkum/xtT93eGXquHFuOD4DlVL6UUFxbrEsdlcbrWOJQLJYPsvlEoKc6ZWmYoZT
VOvkVvgj223BCXvVpt4PitMfVEf2RmW8lrRMs4AGUHDMH4YwaYDCIyO5n109x+VkGqVXnxS3kD0j
J4o7Nadiwk1MIvRhkK7Dy0Sl2I9bqKgAz9nBQ0NR2CaT4Uor5l+tOtywe2UMPfmrPeQFhnugnA8m
lcoey0yWrQJt0GdOdezfqaSUfMapuYoyIMIPwzDcS7gqssl/mmMnqyXArPUNKOCpjeD6ajctpgsc
VYnkvTmoJDqOOmSfLzgA17RdmNjz3MXK5KIMr/4VSjdLp15D8GYlBdB23OqENrMm1EuO2RkWwFAt
CYumS0wgMkOU+EwmFsU7i0ivmvaTU2L2SCuFn1ovU7Lz83OECEWYgb5yn1KsVwp1MgZF+uTcDdY6
BAdPpKQP3lYMuFb11z4JhzCKaO59aF+m7I3wPtUxiZlbH/1W1vfzmlWDCCWHyTaqOx7tJC1NHT94
X+sFPBLXMvhA3Ji6mZ5Dcs1JxO6SHoi/jsrGP/uEyesPRi+I7d6DzScAnQIWm13X4413fuMEFTpo
4tcb5OlrhXJ8ZBNCNeKUyRJDaluyRx5LszD2YCr3oRznzFdV0IX76zBfuxQY9xNP3NDd3xLg+ptp
3TCZ7mxqSIh8CptuTgwMDUDASkUc2Tct4l0FmQPc/RUPk8jmTGhEEQkpcnQZFFRpClEo/Qr3MgyZ
TmENUAdwS16p7jv1sYkn3JZh7qdJW1Msn49FHB7aNuQCiVJL42rqC/c46FdzjzoTDBKGUezXa6ca
bC1pSNQQFpQhoGBB20UG1MQV10tx4g9lEWpeSf0CZ2WlHU0U+MpTunHt+PL4NEucTIhWDjMUsL6Z
irXiY2VSzIuiua3SoKadxBlL4bwYTaI2XAbzQb8HU4N7va4iG2o4ZM/K5R+QTwCUrpUOUAa7KwPZ
+vgWT7gcjkPYEh7YPQvsPwK6lnXXiLuNR1NmpX+icrOGug89vMRyKMerZmMrrrYhJLiXq+9eu9KB
RTM54DvaAHzMl+WZ1Xd56p2Iuy5oT+8siePEmSTVUiMEZtstQa/nLwtnvx5/fUGbngqN65/SnhbD
8yU5hjxB5QVHqeRptamo/xxXRQrMhZx7UjaWIi19BdYbqfc4XHpEJh+CwqxVTNY09bCJ7FSjXi2N
V41r5c++j6gbYVZFRAt54Xkutt32rGpX4shL4SeydqP6DA7a3M/NX3GsvxlKmvzMQL8HbNCQkPG/
eqMEfJcJB/rbAAzKEBBohy6VpES0QgFmWQjSfRX4/LK+5EGwRZBqrrCwl4syEYtpdi9cO/uynO5p
UgM2g2lKny0PEtMjHMeRRLpadGgFA6Ownsi1sKDn4rGxJogcRWNepp0x4mCmcxq0al8bishNBci6
VTwHHpleHz7Nhbb6Ync5stFIVk6o1bPAb6HhvwVAm6aUOupOqVa049nVqmXmRX9hKFzZed934Sm5
V0elWrJkVnaTWzIRfk47pBwVASjlIArycST/9Os9HTI3ZBxkiSpwOdRU7SL97RlfzlWqtwP3w0pZ
bz7/Y7FtOpq+Fdy5zopFQL7LJ1LBa6fFEIafhxkxoixvBmzkd5ZdeCSk9PYsICe1CltBv1F1+l5B
oTuAQctk88PehOkLjDDLt7S5zE6kdE4JdCdNXTadJV+sOzJDctHpYTU3Nrr7PjXiOOVywM4ygVN7
uzsT1ilqrCmTZdqn1xNf53ogSBg7Ivla/1JWyko8/N/cRGCd8z2GKAhFBSEqdQ7ud7/XGQmxSRX2
90ba/3eNG6As2kfChr4SZoZKfFOOnueGXS63xSr2zxZDK8nYTVlHcqFFKTIVnsxgBQkIefj3kOud
EuGoGs2C7cbrtObd9dzI2nJJhrzrvc09u1Qqe2Zl0huANHUCM1A0lvaAdVKku3qKoHoOMMof7WqY
RJuCFRxML5KyktcCLg0GGI3AyNdxR2C7SiiFdgHdfGBH65r5kHfI+3Dw64dNX1IdAsk+mb2Oop4w
vr8w+0LCwIIAzI2ountpz2LSIKd+MKWq4Dl5VBsxEUu72oNoJBV8PINT+Zd78pgEqmtsln0J5gGx
7Jb0PGOYFVsHK5MEzjf3fZOjfoKmK6uX8/9C9WCvsI6KiMnTeFW2/+ncKtOA/OL9Xkdibc35JxL8
e8GEob+8mR56JFR0yiPPXYnlcsg/s7irCxf+fG/55KaNH2t/UVQj1zWZWknjyuyTuI5p1hH1fDaE
Hndtfct6EEaRDJJYKpxOOCZGymJl6RGckn44DgIN0P9hqoVqwmxeHH/kngleLvHaDsH29Y/l0rR6
wUszfi53HqQ8W39sqhDZ3wjQKwbdDapdZsLu82T8eff3EHNao6K+kgcxIHGuAUButC+P+xw8+YfA
MWHjqhF4PH+e3EXittfplcvQdvOIPG+fXZzbGWy5Jp8rqQEvwM714Smh+8h52pwc+uyHCnRWnmdD
OLuhtshtW9ooWt2lDRP9Ow6u+AhI0e1FanrizMr97zyqcWDM+qM5K0+Sim9RlWkNVLvx0PjO5jDC
FZG8V0XZXkghK1vr6rWwCH9xMQ2EfqHqhGPu21A0sHl6YYFulzQIgtgT+DdYcS/t5hs1VG5DjJyu
GYseYTO1bGohYmiF1bLfuyMGDe/pXjHNKl6A+SGEe1j69/w5REgSK4mZjmClRRLulZWeT+BXHi1o
OgWWfTQT5QyTi6CaxDMYimdI0laz4SxRmLQqtS75sWDXxYWSF923xLILmFZZu7RF7t5GWdNGcfxD
1Ucnp+gcKrJubYhASNL3L99FS6Hr5ltrGRXHuoqtRcVaWjpIRfZ779y7bClT41RA7nqt/mRPH8Bh
9YFcAKQWXm1bYku2MnbGdR8pa2U9CPbfeL/V+ImIb4UV1QbAicolcuNk7RzSEl978zb0iTmRpCT4
RnMBwNNUfUyFwKXTcEeF6LrjGxb52GvZhhn1QFr2dFVF5jIVnm25DMPM+NfR8gO3T4QI+rmxHorx
dyBXvBA5WwRMiuqr+o/BaBPN5Gxx0kQ9W0t4zV+gUff1aK7djRRSk+lCrCC3MERRBbukw25/v44w
ljIKv/aq+oNDlJVVyH+TCNetijIfCXQi8ibe4O8T7e/Reos3mCzsVFaj1GfFksi8HTR9gHOfgrYZ
eEHZRRgUAXCU3b+0z55uZAVdyOl0/nBxyZ4trqoW8OG3/uCBzSwwzIq3JwCGsm5GBsLeG8gd4q2T
3MTVfZtriKnMMHNB6Uao+4aEn+OJhyDvZX7a+Dzq4R6zs+RUeqsN+NMa5dQCXvy9BPQt/wdXIAFx
BGO6agFM5n13xEUxOQZY37yGdey0nO66eFkI0t8AtIoF5wO9xDzxUlTUnCnP3SPI9h/mmi9+fsch
q/zIE4mPhY95EbLxHNBknhVn2dFIPdXO4aZYdCpO2byw670vsuqcLA1QsjPMHUvZj+x4wmHe6IwM
x/NktOL1wf0kw80U3/1f6c7d2KU0u8/VHdkKX9XA2zryB7p+jslln3cuUGZxpP1E/OpQPt4GeDWD
6qWX6n8p6lYUClfBiZh8b00abJv0LnYxi7CPurlUnLMdfeSB6Itq1DxAgrAqc4GPSUjrzh0841/r
dGp8eiU7LmmbHVWmLYwM/fdbwqusRoTNwq82N4JNhfsSIy/BCgNK8i4b1wf/HUcJziHrgkojiVg4
u6LUP7MNoZ7cGX3JCZClkZCdxNbIQlKcJW3HLM1XpLeNe0I96DkClVZrMsgLpNq0IjrGR0NxBq7t
WJM2dC05JJf7PSJKrrzVW6QiP0/MFdPthZGShH6lOYNAkJrrzun8q+SQu8xFOgJgn3QCKLE1nJi/
azGJa04w8rg3K/z0INBmX8oos+ar6MyLdBBJhPMGCXNPCk1hILv48P0vH8GU8EUVkIfaLOl+mvZs
GZXK39VQIgzKm+gBg9bVe2p+brQL+v69+mmtkEFFtI6x1zWLisuI+Mf0pEZ/P0y+8LDUkQPrW4UU
RGgEggK8i1NQ4UQW8x/5HN8Fp9+y2JuKNSY9xrVimGZ58A+05Ls6iC4oQ6cZGmuiHuiE9RTF+QYW
gMS15CehTXN9rmstxl2CaS2J7V56p7wKDyLqL7hEMyJAcKSlGSQ/kghd00G8N3Jzo3VwN+Ks7U7Y
0hfBQhD1Z+lo1WoRd2IMLqBzH9tr4QVrF8B+3oE4dX6NUXu0glpcaOHYbbXi1vCjhJlO4CPz5aif
rb9kBXUtDqbVG7kjfA3swXenPcIBGTtTV2CGuUu/eE/EnxkI92q+X6TJcqX/LsmTZJRXaax/YTfr
HSfM0HFGTb6jAXnMYM/0Ue3oUHONXYa9IRtvP7z51+9l+G3kbOwiZ++AxzwA2EbwY7pxaBHr/GgD
bjwhk3vvGlpIEfBxNXT8ETXGllXWPSjC6aZz+OqxXTNjhFhAq8GycVf/6jG2nGADBDUsDSWwvJqh
9opZLM1FySOKnZKQU+fe3PH6WyIVEX0VFdd1bmLn2ZKIc9qOcCvm4cpVC1UdIcZ0IgumsJTO6Uoj
2VmW4SiIVCPDYCeBz/JhlY5lsH4jHhjvUkmBaMje9G+u2YMg20migxomWXpDCQj0G7Q/yD+I1vSS
pQ/9bZxgXux+/9yPuPHQxt0DP1RkZKBI7nhtG3jZvPVkBevpiMXoY4KS8uz7ep4acH4fP1x8DffS
q8SariyQWi1JXd+UMy3s33ldB3uolMf69+4FN+xJ5M85QmXz1xhGrbv80LJoodjs1PNwI+dXHlP+
KNy+UJKtTFAWQt1225nYa3cWOgU5rzi9+zXIrWrTbGGlqKQ/4g+q60PPTnCLGPYJlgJIj5iObcdD
Z/Y6MWgZ0Q8CCavZgiUamNzk9FXEZiogl5lNysjV5eegL9wzPk5fip9DQqNvDVd5GpCvpAg0I0HW
KO4gFVJPyNf0h8BA8+Lt7s5LS9EAH+UetSISDmxzQxsyFuUZLdQmu/A103r920ov19BxXLIeD0Kp
G7uLjuc2n9JinE4qlVgSTBMm3p/U7SYlp1kIZBDZMPfRU5fpDhCeZGO5S9W220qtsPbqm5jQvwgv
evclAYjXUjP+WWfFCgtPxx5gsdf7oCh249ojKUcRSlkJdWfAlslglc9dTFjBE8jDpU7jKBKSbnFZ
qEKbN1gblv3hONhDWp/aas64W48hzMQ85Sl+EQSsl3blxa2XXnJsjMtlcQklZ6AHBefHqEwehE2b
v4r9IhJTCEAdEUfb5qpY27t08J7wC1haSLjH5qNOxlCh2xh929ERX2yGAknkjnI/5rCzHSCbsubT
uosJX6+TSwEQ5pHb0spDnL+B6CLdR5Uniy1+9uwEFXxCTa60ku5IZsgLQ4FMNpG3pUVvxUKOLRGt
F8g6OhvA6NgUOFDp2ZtvBJeYp7GISJOIodKCwPnBfXusr4ByMAfLRlOSsqN/uWK061dfeWvDKqfb
Mdl70KzBg987Qk82B9Z0LASZrmYbjcaM2nXDcgoM0XezgJzH6/OY9O4AC0TJcqsoyWnu206UfZr8
pFTZgOFSdb4Q2gVT/cPvPgEbbJUA9tyxWk8i2W6Lsn6iBRbJLhHwuvK0S8+vkIj+UkCdu/UNqDGN
fdh4Ebamx72cBo9C+Zri8YChO4MP1K4/xRUoRVnk6k/zXzaRmO8Cq7MZ3WJ/OjfVLhiswuuNwFnk
bOYmgplaS454hoPgGFo1E/KKDs1EhmiSJ22I/q9G74iy0HpMhOD/NxvoMW+wWchr9rU4Gvq+XXjM
1WdFja8mvMV0q+nNzub80lwqpy+SjmVwxOT8cmrbwDLYQ6ihQAozMDzuPE52QH5PYEDdNe24i6DP
hPnl7CLceYuJ3BqphRqwsRvI9j4xWqyrU4y4vIFFYaqGmLBbTiHRhdrCl/4+Tzlz/FyOT286hVFr
tX+zN/IMkOTB+hzag0OcSxk3MQtcFwQ2WklhpTvxt2uXKeumvH5Xt62A/EIU95LT91+w4hr2MrBn
YzSeSqe1aJ5rnHUaDH22ylAJ2WB9Y1/Bpls7X4DtQoEpCX4aZa9NjiVqjLxzpEd4rzXiNfV0w5qX
uiyjquoYKlc67azC/N2sqSAfMa3pYy8olIPxSxoYrmiC/iWMnHh5kQwhSPrS5fHKwm7sZ8vx+ppe
HVAGW7zeEPtt3e15UXtCgAB8nNe7yi7ZdhmUL/dPDjDu38Dvih7zVepBL5q1apxQE/Y0DAWSRxI3
WEFL+WDxXq2kEvnLDZAsXTjJfx4DUHjmNrSufbUdWtl0eiYWenp8qua68VuIIkGYz/4DQKOgARLc
KU5EARdnAM21a3xZdMnY68Ryrs6epal74HQWpfPIU7BH3qWUnqmKzA7+k9VJE/K9OfjvjfXTETNe
wwUSqqvCoR6VHc5hiNe/xSbUK4ZJwNSvZTWZv45+nR3s3GT2R/+hsfeEhukQgXMipp8cAjzF67gm
J8d5YghhJCvtg7Pfk0sWqP5eBWpKi1mLCc/bgCJDRJ69yRugXNPINcD5q2d/HDmRnlJyqrSMmuCW
hlG3V2VPK/ML5iLueKraCHlY1LlZXjZEm4U7PCMi31VezKi7V7UA1yH/9IOhHuKZWOuXAq95YZ+r
LgbllExNYQAkzzsnTbbcsL3gg2IXvpPBVy7IF1WfwnQqGJHcl3CZBm6EeGv1QrHQMgogvV/6rrZL
nMPXdJOC3Demo3UgYFKb7cf2ZDgIPrajIfJ/3vhYEKY2UdG/3Swpltu08BHs3geNHkbHJqONUC9U
VB1594QIYOHv+xxUUswqj86nn22jJGYfAt9xohD0/ihL3mOWNsgeC34WONNRdRPHFc5a7coFShvp
wT803rsgBoKitaZmUUC26I9wkRy/USZUE7r8s03MxI46KfEEiifybyxhkViXL94OETfrT8pe488u
E0hdnRhLBIYatM583EAMylCmmsloIUHSgbaLKuTXGet7MkyryeGOGPV82hWhodaQmJGPKUaQHVFz
P1NYWZrxPk0LJ8U80s88xLw+H4Qy7p5Bvq9VnX8pDRkWqE2obXYYEVs75i+OHZ/IecxvcCq0LCiN
Z4zbPstzKhQbxaLzstZAhShiOfLjfyb8GVtMjMgR8A/I0a7tFb57CcrA0cMWd1QPXUTBdWCVOmqY
5Gw71/QAvCWYK81T5zT81gMr2YTcwLYWpBtaMKVpUbJfcNvqtGRSrNMekuAVkaKmJpb+S7iWTqgQ
uKdggf6cUQ1ncKIySyu/lo1dAV+VpaSNNnpItWsgX7R9f/sgDByc2+igg3hVjvgEfj2i4bVEi/q+
3rjdbjpvq1rMH7R55/gXNnywNrJSMqB+TUZ/Caei3o9CbdMRu8IFoRTeRSoZdT4B9N8HfJd2EGaW
6es+rx9ciHEeOYLBfEoV0pblVMltNOcn8hMx2F0vJEb+KuDWQDF51MJE9sTSuACtiufcNaB0r95z
6srBibvQALIWUh+U+/OL35kajflTadKnyvgcqE6xi70wjgQculBC6OsCJZ3RKiugCbNS6tzej1A3
FHi5L8zt1Hllynb64VnfuZFOLYnsfNoA11bxFOiO19Wx7hKdUqBCwP7HW4SG5QeI8oESLw3GMMIH
juUwfoFLFfRREpZEHXVNkFeo215Ap8gX4eOsCT6CHaqNKSHD4ULzNjylhcFEilOfF9ZuXjMzAvYN
W7tN40OwXQSFUXUK00eeIDQ+/XeKQKd3ea+6f9AWju1L+8Yizj4xw40cOdUGW7RqBPVUG9p6S304
53ALijp0SWJotPl7HAj82bfrpIA2SJlRK6EG3FPPUeC5Xya61/Qy8O5NbfDEHnANoqFFRaNCl8sz
DbTXwP3Ou5eU9RkCzhLW4YuEn7Jgmkn22euSA2PJkWOGKqu1+0IwajvRnhPCmd0Y7aHMBklaqyej
FofRJO2bu0Sd2fP/LAsWKHMWTltTtYQI2oZYsGxI2rrq/jTZHAnF4JktyQIuKzJV82HVGisPZaOT
41tuSM9KPxnZqUWFWuC2M2ZvUX3O9icxw/mUM/5t/lXJz1ctenv+yj37JYYlL/+BUdWsS2FviwOQ
39L+kt3MRwWZ0zDFIr+NKqVj+N2dF3FGK7+l2mIBoyoOeG39FUp4N3IJquUvJAMBSil77hy6sH4D
JTyDUSOUjAylgt5+Xn6I8LKxFahP3Grj0tM/ySvqsvm51FCshRFJpsP9dJiOkX16ztKNT3J2/Zcx
2RgZNvhAbRsDKgyvDYgXnIiutP9+u73s1ZMNV9Uoe8ZsqvrbK5pPXbJxjLZESJ5efKwQUfC+YUVd
x31JaEOaPBi29icsjdBntdWecnmFBFC2yl801jEe8xCiI4vx1g8lx/RWQDpP5Lk72Owg9tumilbo
0SXAPNl8PZ0BjhvKYaTeyhNtihNcQFa4sE3H3yWZx5u6Fltr8ljFttGSjaJ5LaK0U8SS0yUHJIsR
aTasmqaoSWIqrgtrqEQqYdo7ApY5xCUfcw2OZpn2qxwb6xyyVoZLQM1+K+dj/TZd5rq9VmoBmtg2
E9sNdrdht1gqU2mtO7khUiaEJCD73xpQp/Ff1LRJ4OTvqUW4P52BH5Zyg7IYqy3Go2HvifsjcGmd
qO6UMSwM904wwLrGdeC5eVTFgm44hD0Eqrg9TyTUEHj5y8//9VnSTDvtTizytyydYBh8jReMmeb7
DgjpVGrHrOKklXIckEbjDO1bVET2Ihm4TN3sKEyObtkGnNVvXzBy0Y24KlEJCMe5/C46nzY2ciZ0
7aWdEUyn7Qoy1i+NnSEHFQn6lv+Qk9sEo2hSd5iYlkXjf/POXwlq2/hPwK1CReyR3eARq4VyHJV1
11IuuB8Kgl/L349NS8U1kTwJ+2K+gHr6pctlUgnY6ZkVprPxU1kduSpivtqsDf61JBzBcFpSM/bh
mPXTZkKYOwczlw2J31EHBbxErujoq82sqJeOLMTv025YWVIJ+9ngLxjY6ttZ+xaj8aF6Wy1X5si4
UYiQlN2wpsBy35V0asbEotjG97JTEvhgVFwfbhiQvEpyJY/j4UXimkeIT9ZY2dWkmttibUFsCX7q
rdg6TNozK80RIrIJd/nZ1tOG+VHjgN6Ojbdn/ZuCHHJv7rgnNLsZYcuPXrwyfI0vd+wD3u0Nb0Q6
t9EPQBmI4Wy9F49e4dr7VeoVccF69wwB2/2cjQkBSowjva2C0MZdGl43lubObgVPKu51aj35xDRQ
4gugQQh6xWQY1JDddl3HU1pgfWTtsMOatHGAHdyrOC8LWtdxnR+JaN78gaVmyWyDNbilWBXUto9l
QzzGysjFKyHfLMLSOyvinZvVslhGW5QlmU+THPPzoYpzRz568Y0G7g/JrTEI4P2rLzNLYNoOhqfe
OBJvrANFPRH1SNt8Sq2cvbcW4ulm44qa9CyzXhlbaPWfwOD9sG7bWKPj95DL3R5Bl0t+UqQKA/p9
O3mTACxiDo0ZkzQkP6Z9LwEepUSMZci+qbqrrY60p/+ft3P1mMEjzHe038hjCfyRdRQ/LLhJukjP
zhwjKhtp0zpDaWzWzAWxiP19nJCSHnxpv5eK1z2t0Z6vWehUql7eqq8Pf7acG87kcXPSUYXZ5n5I
gcSy2Wjwk3r4BUIBdJiUZOzBKfPRdqXgs9hJYGvqnGBRc7L1gGxY4D0Iu1kZcw6dCbNZuf7+YJtn
vRON44d2nZHK3Hp7vuEMfoKbnkDBUk8LB4lau8XH5QQmy9cmBo61k/y3d3yQOgAwffMWFu7850cb
gLPQPey3L7R5Rp3xbHrAnn31hPOVtx28shhTTSJjGoMOBcgeJ2LCG/ejt91UzR48zXvO2BycbvzF
B+W4s96uMyKliSeYXb9V0sGtqEbEk/LaXiQGahu1r/wbHXrenedIwYOwgn7SM6mjQtOfldKnmQfE
DfWYJndc5ue/kDtJMj5j3FYG7ahYMQqzKx5gx2RGq+RqTAmOnww0pSHIFX8WnQM3dXTv1vbovHzu
8vtxKEtqq3vuii5Z9kebgMHda7u5EnNBsXpBz3YQOh2sXmd6FGWciGLtHp/nCRFLdi74Qqnm5zft
p3iy9NbJ4UtXbdVAb/a6hNqgNFZ+FJO66uVM0RyqBEMA6gP6tOgIOp639qpS4vR200kJulc0Ydg1
fzCSSMKZW4fSUqQm5cg1MFIX1RVJPyMk3NQSqzDvyfSawB7uZTBxftlmlC5DrGb9ga+suW0D96nS
qA2+uBsHBushWy3tOK/Nha+ZecPb8+pQmF2nJmX3do40GzCxeq7ziVO5Np+I1qdPSdl9v7sNOMkB
7u9LyvdNJS9JTyfDgXqjNzjUhnLJaYwatKtu+aJDneBOyxoSLNVQuvbMqRR5D+i/fsplM2PIHLAk
DCq1MSw19xgc3ZCWF+m1DRBa1f+tvmXjNrC2fbXNXAGNDkZC8rxuMH/9FILnD4GglrnmoTgcAEG2
QWmMUi5YI6pjEfaCI10efcq8nTGBa3ZPFJ62cnDKGQ/YSrRfZTkpG6IEdYEC80Qkzd7JXpviGB0a
kKiTj7cmhbkNUQLGnYeLYt/jdb4/MbFmIHH8w5vTbALvvjZNKvJsgZV+vs9qLrVbJPxQOKF228gu
Jt2N5BDrWKykOTrtY5ru8AWItX4L+8if6zBpR5AsrjSHG68VhqV0rlWMtmcXbxbIDj1x8bDPQ+92
eF0DkLR77Y2Th0diEAwA9QjO/LWbMPo/xDhG489pullQpP0mwGnqlDwZ1CTYC8fLvxHbqYbfm2J3
qRV6TiEXmPoGiBrdXSFzcvimoYEL44j0ZxPJBtCvplkUBoq9Fu7EatHpDfU8j9PnNIanJovYMnqq
HLeKutl45c3/fTUV8otwADCYW5ISoejh2uNq6A6MzjAMN4yC7XDklX0FgLciNEhme15FyClgyn1k
jZ0ZZd1g8gjFoZ97ZDWWwdLGjrVgXtF2F+GKiRayhJoIpMa+YMgwQ1A8vM0RKSApKMJzqdSr+7vT
JfXZALWck3B7RxpxCLfqakNfA54rnZ/DaPVQ0nbzEdsQQWvRHbieKxvPqn4O8YT9tzJmQ2L8f8se
KfdE54hU8wNtlKZz3lD5HnzFaRMwCyQZTsbcIGERCk69D0W1eMFynL8DfiO99POw4/eScGMw2F3N
/4mPleDrJbasHYbdO5dA8ibk8Ugh1HJKWodHvrYa5EY6kbI3KtUFYTz7jwmAigr0hTULyBN2qtkO
iIn/rBeeICvhV7MmHjpAyFc8nwPhWK+2aASKH+zgfb0FL1s7i6Z18iMnLt4enLLRr3//xM6Xde8Q
3/LkwZW1e1Fp2DChnqZNDYbngqF0q699fLPUgUiCsXuZhZsEtQ8G5q7QB2fEv3MjGfkrzBXQ8FnT
TjI+L9ys+Y0raRzvRg5jzNtZzsLAeN/0UhUidU9EvvOBzSAyZMUkgc1NdlOuLykkthYmRUubdvmQ
l7PbKHFtrYvX0A9TNeHeON4hOOtdvuS2Dl8/kro5YdO7J5Vsx+dj8s9Zk59QroV1o0qE2CJ7yUI6
8awq5n78gAyo6IfaPqGOAI4D//IndnaUpWoFArbb0+SFapusLP/+59SI+I0C0HdpAOkUlbLXEH09
IBcwmxtw9A/TDxzDjKq/g1xdbRXFGme03NU9HIA/yVtHqQ5BXRi2nStUmXXK8P3oeHG0cEi/18MQ
GZJ2ACILFIkv8+VNh0LpTwJttGURvYBFceyUXAbMKdScnkFgw3foF2BKjUbxCzyg9eeC6OvXi4fa
FDBgELwURNJ6yI1M4vonK0+63zZC6xfLqzFo8etke+u4gg8KOGc9iFHBb0yOPmC4vg5t9RksJHQq
SyBj5S+08dAdFOu2egwepJwp1zWBIK9e2aya9SLY4jM99Clj/RcDEkCyA4eXPrNJQKE3S4rOV2p1
GPtSGXbssrlw0npGN+bJ471zDSjSe0I6t38dgeG/XBnIAymiyOsQuTJAwM9Q+yJTTyvwzoR5KpJu
H6DamBRCBHUvupNEepeBKDV9Z4AMdGeJbp8QJPL4plLgcdrQPbc3Y1uldv4lnjhndNhiOVaqMnfq
P6MHkE3QD5QtnT4SaQz6CuJV1cOKs8JueowsHbgwqeaqLety0AJfLzIQnqTU+QgbqlfLZleDUl5q
JitL2pA2OmijaN38bxSRkaj2CjYLuDDFxTG22ec8rRO7qi0HacyQTfjW605033Khit9LR/INLAHD
24oHSGhGvJgTbkeF1ICYSkg1J/Dq+HS6aLv2XSOit7rzrWkiG05dgyBOo/uaMXs0Jfz2TMHg/a8g
MWLmlQf8+IWkgwYmQBKpmiWTekULZpR5oZaHONGP7f8G7iLgdPN6ExO6o8oieR+jB2Xi7BUw//Ri
eCB0s1Sahgmod9ZWt7cEcOaex6Yf0K2Pwv8h2Tr7P2KdAoptR/hxvCZ/KiV5OurJWqFUMH5driOw
+tvJMUx9cCJ9+r089SO992Wdpq8RgjVK2xL0gbULFAwiIGTNqntf/r7sBexc7JynyQgmEOpj+DUu
KV+tYAxJBvnSF89UMsEvH1gRkLIrgmNy998yJsII70KagHJnraLN5w36toaW+HiSpJCYkapKGFQu
3g3upvQXUKN+Htfi0widDpQ3sT3fPywTF+6n78fvFkSt7oRVhliriZ1x5ro5V7+BJMcMcVT0ebIG
1nwfXv3LeCRudTzgGe57tsuLr899emforjTXPGNoFmKf6EuX/0/XGiUlMXZnPunkqNwXbeVCDa6+
2zjho3jPfZ0KDe3XNvfZ+yKCrAUuzOFNHAoLBP+qlVeOasiBAH4strrg8i83XR0GUhGEkTXzlQA5
1cwU5Vrt+C6OnHIoFxVr/Z3fL8h418UN44E2O2vVcflNCL5jpItJKiJVEq4mFRsIWKAcnREmL12o
V2Xsb8TMLPULIAMWDf/IKi7V0nrBAq5go3+YV1Ri2NhEywIKQY0FiU8isH7Y4QkLAfTCUstAktsu
Y1m/8qoUjjO06vEGvOANaC/xH3poQ5Y8oI4OvgtJFHAAZLOH6vdptzjiaWpcrBLZdjiSKoUg4D7y
T87wsoSukNeQEaPqzQYaRhxl8HsMDi0vsUomnhKHNXWCmY7dLtP6C3AHH+Ehi6FX5VrwzBu+2r02
ogul0JFR8FjjU+IqbP+1uXp4cL+P0q+4eflzXQTsliwQzLwS6499zorwrkRIniXy5p/Cbw3X4reU
+QAHE07w9T1Tnkoh/Li9rx9J9nhu7tslq1WMj6KAjIboA61EzGEwaNskJIDMZhuD44zeHiTHGG/L
cYUGSFcHcS9qNcOlz8Tr+YNO8EHCjcqu5d983x3JOW5I97o6kPaeSzJd1hVDCt4yu63A4SL4Zqjt
IopkvLFWJLGZcy0QN6XJNmlyXGoG6GmAlIwp/Ae3apfLk3nSTzNJyFkwfOAHR96Eut7JxydKQwh5
Oc/T+IoMwuzerey3IBz8JOAzdpIJMK38UOCBQreC7O+VoFv5a3VWfDzbQHANnj/17y0l8g+PjNDN
nBibrGwDbbpuQ5WB8/IYqijlGVvQ03g5ZxVY5D0bLCzBK6iuxCDbcEvEwa3cHbG6RJsleRmVWvHz
gMfe+DiMUicv7Doa8y5iQAz3hv/jbYqJ2iCN3v2dDtW80Yy6e5aXfPq39TL7WoO0+VDkFyD/zNj9
C8GQUuaZ2ri80kpWYWspRQoKmt/kEJYjxw7jyDrZygZRXRQ2cidHHA5V9nnXqEgeStb0FQtcOrjX
twNd5nUYvJXB6hB1HmXQyLTMOmuvMdYIkYoIBOKt8U9w+KCy6/D52pQAN9HBRvV6Ajhacmg18A47
VdOu75PiZw0R9iN3Rtn/UL+6m0VamVEcHtjP+GNbZoDxOWJ5EEdK5r0KENtr378dUZ9foVdGsHaI
S0wkZ+GtWQGjdAk//yDs8vn4tK37RqI3H7AThf6qPCC5M4YnBY86yJMVqWF9vsR1E+kXEJhSmlMO
n5Za2/hRv0VHV22Uoa5U2gYchBjctK3ub5BnhSoGEZVzBAwHy6UwCWY9aNGS6816MevhfscI/32O
LIUUtCgitKHkVBLvSiQXGC5R5NewgmceJr705X0aKSXenR4xmoll1m8BAYttoqXHdr/RJfjdneoC
zehGWdnf6IVL1SGHB5haIAGyKNZjO2HnONhF85kRUH8xpWUKomKNAsEk+5bB06VHdaL+Sz1e7/0X
lzPvM27aUJVI6o2ehZhdxKPrG4vKNWlEBuQpxMJmQORtLaTRbAMAQJnItophxSCxt/lFrimSQrq6
Il7fF7z2hsKtKA8gOs0Kx/ID4BIMYi1e+9WmCbMpnhONeocMK+OSc7xb+Hm21H6YnQgehMzpfIkm
/Hu4Uov9TCVByuD2teD5eWkOdnstCA1R7arbaWSxWB1hdmz1K6iUuv+eitcP3hINJ4Az75GpT5pi
Digk0CzxjR29u8zpbgcWM0JduTRlEvlLdUNc55hCKlCNF6q/QM8wMH9jGfld5ka+ODHWPwIihnM+
n+53y8MxBLsk1eSZKMlpNUyxpdagbH//SMWTJUwhXPVFw5vr08QnM2C8AR7TZh46jOT3M3yJIefM
ZgGN79YN22Gnr32Oi91FxyiY3i9TlyWFKqnc0jS4JJNR4TRILInBbK2vwSV5xfHvR8YosA+tNcpy
kPRRcYsOJrmEwyE2Hqi9JrYwe3rJ4K4xSZtZQ8vxm2My8hYWAsERvo+F0sY9Zycn/ylAYHwkGjz/
Hzq+NCgKzxEQ1IX96m/gAVewRH81YHzz4qjUoo5qG3GAzzzwdcSXERs8LjlS1SD4ePRQBN6nSwaN
0vTowWU5fG4ofz6mdeDMWCYdaVjQbPa1XEzWqaI4GmFadhUiBHZmTPtVwTiV75FQMpqDLVvhgAn0
WI+bGZ5Jr51jrXo4cjAYINsjPRoPSDixweR0Q4aHHVykc1XYdQsQMJm36al+XKRAuLKM3yLn8gQN
B/LlDzIVIq9gAeOlsl3VpwcFOS4Av4ht/bjry5v6SVLZjr4WP3YxmBWqTcmx7Petr8cCPoL+ajdL
sq6lJKKoRhWkm5UsF5sAXIA5PsvCfyrWm7e5L/2kHYzrr6omTP6n0fJWEWbqJ6oPoTd0TCUv4XRz
gAmCPBl1gbxNMm1Dho+BPwSnim5I5l1EVXK0e7seKQLxwwjj2wtWa7B5Jsoq9wAq5cztYBHHtE55
3Mxem8K0RzMMdPkojFbs46QvTDTKQLKbcNV9GxLFLZpKaRaAtbdp+KzZmToT5EQbNdP4g1BlSpOe
ZpS/cV9NyR/EfPc+LE2c9oO0uiRz+XDcOBglfB20KzYbTi8yKuDpLBAmCdaGYKgOSJMMFbcc+LPx
ImYh2MudxzAQBl3qMzlardWTYrFBzJGQkzQ48Xp7n2sKXQ6v9RVqTicS2h9PwnykAoItbDgtxwNx
sUvF3LjoLpX9yimCw60UlrvtuuGKvDgGEkdCejrBifQ/UH1WyNPIYk0ixD+rcTePYFVpU/7T5zGH
vS2SuXJVj8B3mYzX6f0J/GNDTWxYIyi/sEVZSN7iO4nhJWbOH1CIYBvY9eQtvq4nhD2pWSAP089W
QZQo8aakHn6GZuWf0hDH1HOmgaEe5bkhWQTxbDHlQM+YYvzxeN9GQonXRv8Y36dYqXn5V30f06P6
x+Odc+gP/WDymrteo625DGRhhxFxiFlh42V9F4c3vCUPzGvf9DS6++fxknajqclZOkJl5GBPoMHM
o7AW9soug5teeqzE0KbLG5QKrHdcZXUV/qqmQyL53Aifq7QNJeTfmxs9sDBIpizYTKGXR3A6IPGn
K2/HODdX7jKxY01a3mmWJ3EoMXlKUSA1KPZvNSTFMFu6ebXLMQtnSSU4HsNeEirrZvFqJ+YmTxei
I9qeARBNnIpJvdv40cYF1UCkBP/gnXXhIHn9davnFFyiYP7Hn9KYTNYHqHkfCoKN7XBh5NN+xM0b
4Sw+GPGq1cgLa18Gbl9Y7QUCdyHxmP7BsK7HCN0Y4Cens5fEEcbHCgwTXEVgNStbzh7i+S5GlVEq
wzOujdPZ8PzYV8Rb6lRFUaTzzR5lbuBeDEGvkktTrt1FRf4iONDXDKdyvsoFikGWzKB935UyacWd
IKE84e7PycKgoUMQ0s0e+GPATcT8f/+oAIWtOgkA/uOr7tGMU+8l9P5MBsLsnZctB63OsRVG7ofd
q74y7PmOGCArWvZYD8coa/RbxqgFtwKaWwje9mpEZGSitMdUPnR145kSRN7I8TBolAhO4cjH2l7T
3fqyKuBsxLgHHFR+DyswBRjwVXR3b/pJBM6BiFt5gMamBwre6XhobLwAVUpHKHYfjcFastJCbGB0
r8wB/JMZlV0LLNScMqmSEtImGbIAHckrFbk4+qAVp4sKiW/uuhdJWYiDMTuP9LHGLwZ5eKz5wGpF
NvevE62+wu0gCQ9h3USYvJEDOVS3nVaIOuc0JZq2FXqvticVeQgRdCB+Igrvs8vQlLWKubMXd3UO
SvyFwa1fUWGSF2CcdjMdP94XsgRPStwB6ie9AmWuqnnyasEkKcPrQeC01Hy0lQvEAr1fyWeRMply
cM5u15EL7K2RSdDGG688ln9hTQc2hO841zE0ZK7FmA1xvYAGEWZAiVM8ZxiTq5Kgo/dGW3joXdrR
Tdq9VvItk80o+gA34a87FuOKwpK00wZLU2Q1DLhX50uvGh5SuPwOj/SZyJvFlIukOxOoENOh363n
O/O4G7Drl7Gw7+bAiPaLh2BB2tcZ+wEaR/iv+Dii5nJEduEOgBXa6/Cakgo/+6JH39YrtDQgcnpC
Pt+69YDZoN7eZZc1u7XHkU/q1QphqDzYKOZFnLuEafag1P8T6PqQbDBQ8cxRHW5zTYjh1yD5lxi6
/fBbpPJBGG/fgJc5fbff+GrYStkRI8J5BBnEmZJrW21g1cRtuWu+yHsW5tbdQunNugFcNwlsCRjm
8vnAczkpqQRMAjDCRaGAAIMQ+Xsy7840+VKmD1wLBHaovw0c4EbVUDralUdrxmmoIm0fg+ohqMQk
ZUFWtuv50wxShNmnZEr+pC6xLQ6n0fXGLISe5QhlGWMc1haB4HeO88vstTG6VcCAGWk/Bb55eTLR
o5ygA7YI7FGQK/3mJPKPtW8fxDju1jx7O2RMyyAtsJK8pfQ4HK7AXzKbRHVWpzU6Aiw675DKWCj9
K1BPaJLQM51zg7ebwzZnPu4zE0b1J2cpK2z54bpUVy9zDQE9XBXME5arpGIYVvD4FCqNQyYGfYAx
qxX0TYXV9R2m9P7wUc21BXOEGJ+pI4Qr0czWiANYczlSMxeTxX7v3A6Pip39xDl1Y0rCJuCsNZw9
ywkuG0s9gfFuxzJZt23XTKFHBfrFRg3MJA/cvq9WhQa3HYqVumG0u1TxOhzafYV4WFKi/M3Hut98
1PDNPYlGFVr37InSo+FPedAc7paHNCSDxTcQIP/8tcligsv7+CEkXOwGt4RjY2e7DuWB7yhpdW0s
LgI4fWHR3u9lwyGXtiJjgca9vNoWGOaxmSiM5kvXR+5FgaEQd2M3b0XmNSZfl10lQNNQoQHBUB7s
C2ER/ukwyO4r64HfWu33ZBciCoqmflq2zb4Ce2om74OJ8lbZoEjC20yfQi+eH6pHxPKr6NtN97ge
IwF38VjPSZ75QCjW+ZxTtA4RnwUdmkheZw+41f70gqLGbSCA1X4X9HmO4J9I3S1P99udBwECAzbF
+GVrfN+hdf4xXjC63Bvn1/DftyehVCGJ5TZ2sIHpiJDRt8QRtzj743lMmBdNiBij0LvDZ7zK+GTz
zD/GMK28J96wvHtnrpdl7viq+/ybDDgoVXfPHpdZoMNGYzokHKgF5J8lxEfKU/Nc8CyMR1Lm8Tta
X2NL6OpR0aFhew87/Gkj5V7fW87W1LstgtQMGRx8trGD0mfk0N1o2msra+VxBCcxRllHAn9/svDJ
TB9Bwp5gcVWdzsBUHMLw3yCVAnYcX0HjGpdW9Hl+E4grZ0i/gl/uORmUsSLG/x2p4n+nfTKVdtfo
f38FMJXGg6A7HgUoOnHJBo6rWuly7lhEl3FhypLm2T2W3u1l0pi/pniBMCzlHMNTA0Rd5w9UOwfU
8so7qAeufTLlvchfBCvO7v6p7hcrxrXFHQl5KgF5AJKsd/3Y+VDQZPfDmYRrJ4x33gpBgFwOlTSj
zLkEuJhuEqCKEKSY0pJjGPiYJlRDvX7Nog3oUSr6ycCoV5MkKVYa3n92TWCf/ErZuK3p4AmzcpN0
2IH1HL3mRbYkAlIMJMSlv/OsR+OQmWrxUacN90XmHFCpPxHupxgCktVzpuRYOAfKCmir4qBAZUAT
JSty4cY0rJ12oamGV2dmMxROHFdqTP+LtJiCyLveZ6FIKGmg7OaOnGZh6EyrlbODYOxewNtW7A1A
rJ+ksMWlvx8UT0Cbw4uo8QO+JEy1/yZzMNG+4SGp/vc3ZCKraVU+fXRiK54NUgghtfWc3yEPu+qW
vg9mEiaFpimQCBeCbZhl9mxCDoXZZ831MTv26EtM1+T5uEgLRvw4gkKwMsXay9YicBeoCQRLggQl
Sq6LaZXKxKDSaMYTkYOORJ8VMOGxUPJXSxTXJ8KKTLZJmtYoimT1gvc8llFGdmi3ApRKkgWrdjFF
ieBV4vgsqw+35AtXDr3HXHuYpAbZcmorzzQqnHKL2Zg5emdYgp3jmR+5qDfQdCIMTKU52CyWhPyY
XkoKeFwbSJsQPrmyOOhbIWIa45lRGsam59Mj6uh1lH+u3HW5wHSAqY3OjaL7J2b1eo3j8GJ6uNnP
F1ik2WalNsteXRggsxI3dIUumZ3ElPU2X3xw9OFoCpMhJFzAUO5n74EjptfO8RAJqaNTT1OGCmY0
sod+AXpgYwCExL9xt/+uiYtwXYWAILNijinCQ/P0DzQXCidIV3OgwrpC7u+fhA7KgbjmEQ5JGo4c
cY63WqhlGtIRtqEotfHUVNeKNvYtEPao/6TwwsCnq+FpufVabXauDLfO09chg4kazLgi+P8WWZdO
mG/i4+0VJ/lvxbZ1K/0eoLypXssY2CVCUeBG0THFNZWH52TL4NXOfLMRkVFGeTpPsnFXo13o23TQ
YiuCuo2ECyGzK+9gOZuPI+cOGgo79HVOlzdka0RlEeLTcnQ3TpF4XMnBhRElrcI4oGFkWugJ4J83
FOugUGEonua8B4wf9d6BwzMJQ0dkGhe6f6sduGNKDmaymHOEYiVJuHGUj7JFMdTxL5yaqNflkBT2
W3uLmouruNc/QJfgBB8n28MIFWfdHpkHeC9Mczx6OmO1e13ya7QMAbxcVZBcLWLOXNq6r/g2A8si
h4TARbg1Z743+n4nWkIkPPSdt8Lwi6kWlTSjDwf8w/1RgZ+Su8cshFbPE4dVlWFZaMluBfTScgx3
uXrjSDgmjINUhu4ocs7Fid4qaghRFrhJniVXdVeKWl5nx6+bF+CZ4e7DXpwQU+zAuzLVSeRYQcWT
/6qkWuLY+sLPHFWv2UpY8W9O8UOmuGhUxRQ+rSxZGgut2HbQs8rSKcITbexfaocpQ0jK5u31j0qn
MifISUCd6/Ey9w+ovNIlIOPxGy/jFAIhPw7Xt6mKTFfrK817Pxtcl4pvcq3Q2jdBtnI05+R/AKQ6
z7pohNJ/ZB641h0H/RYmbilPBrj1ntNtsNrKVG107HzfT5cYIvtjsD4hy+t8hIjKSkBFW7mXOQzZ
Ai8EGE+DvcfYEsZjGilES+8WFdSDNMmARLnOLiT8ktAY88DwWBa5m+i6/D7DCDvKcXcldP0v1EDt
2zXai5zWm61BqjtFNE7DSsvQfncJGAv1aguP8gFwPTjvvMJaWGwnl6ev7fhkK/ebySH4rj8ULU73
/uCmS1jYLtnHntDjmtTaMWp4wu7pF1z/pzsV8CX54PETBjOdLTfyBOAcsl9hgy0tpzxC+7Xjkff6
/TolGFgl9fsqCdHYp87/J3D2PLPvHLQ6ATL9gT7h99bTGd3sRes704l4jAgArwTcwZMEBx8Qp5xR
uWya1oDu6sp7+8BVsDNxT2hHKsPHWZA/VTEUdaJhlMb6mfSgymuxSX3BB9SRaA5n89Al043ZOqR8
g+J8NdX7X12NMjfWutZEC45GWcIfx38fKUhO1HuS7oW0bqGt+3bXA6JXNokStUITk7dia+xUDq+I
3bPnwhu6E0iXww6NeR/YzBwLhHvpW+DkH+kekJK626OkPDJ9rDdpccESfHsdx0d6PxHwUBCItifx
9qjcP47v1V5xUsCM1vIfAz0TcAZLciebemWWIgwjywzYCoJeE/rWRG5R56HuSmAmsFFKLRnXo33D
DBBBBHx38ilKhzbhFx0KkiTTBniTyO2ekf5G5TrSEKnAirpXXjcIOloX/CTd1xbM3HvTQ7CtmDeM
nC4CcOtnXA5nYbQb44b0qo+LcbAE97lbBy6A+Fel7beMkiUFhIDEsZJpnFGeT7QuPnSh/qG9uJuE
bPF0eqB29SwCHtulf/6BxHqSg4O6R5BfA/Gnmv5sjKdCmho5yjbRnzqdZZU2AIEV5ORK+6uJqA8I
m/PLUvr4LEdbIebOiJKrM7Ojka5fdsFNus4zNHxTARM1NJpEERMjmOW+xFoAmctuZDpFJTqzY7ho
Gd3CS2cuVrxWduY1ebgr6cr91Aal58gKoVXUlHub9mjVppKlpKJD/d8jP2rscjy575XgSIoByNBG
5Msz+ZghAtH2zvgnTIwV3qMqbShordfgDK26G6jaJcj207orz2KBsbMUqnLq7OS/I9jBlh1empmV
Ver0bWkGNj41e6JSgdAPbOWT3WvfO56LuOstGSNNLBV2/wdkdP3hNZISzrQvrMlYWBq55hboc92E
B9QTYNhrlRjMrsYo3Bh6O/KNtkRLYXDK3tNIXOhfxp1dOcFJXQEoPcQtO1bE8ED8YUKVjOtPUelx
X4sD3EVg0USeMPa73s40oOxeX4RwncYGqMuNzypoVwKe6xjXgNugMt2V326qRAvyIIlycZjulCaK
xpCrHUEJvjZWteg9Y0fo+3CWKzP5Whiwv+jQlgWOC4fCmEJ+4l9LHQEHCHfq3VowIYW/F9cbNo2b
G7+SMeLI2s/aYaX/1U/FKXnkYTX6m/297T59uc70DidTo9WcBWC1rhFEkn7dvlm9SPnHnBIHM0St
Z3OB9wFWEQHHfExTsiawM1+2ovWdijfUsATyUIyACSSoAx2H5z89Q77EzS4yBqNug+iq+XW02Wlm
i+tiNcBNNBjqV1xmf8W7xX80ApAAH3X4oSZ98RjkxWAhearOmZaO5aZVM+Ks7dz3FHjSBhRPRYWq
yBDxNUA4V8OcD2OCWHWdy/W/SP0hH87nSZAX8v0jAgNRbXPoaJ81B+DD6/TzDJIDXoJbpDcGBPwy
ksxWVYlkmuULZySCmIoH/WOwxR66Vm8Zw6UclbOMJuM7uNlQVK3gsSmS5CSVbvtwnkqc4Rjf/upH
3nSm+NjRnoTWe7EMeaoVtQC0Xl7orvF9XnndFMBqVRLeF0eyMKu8hJH3Ra/CVLqW5gQ9MRW5KlfK
0RNO5XjFiZ9KhotPcmIZqlvF6OgWhloqk5laMuxuTyOlLmxdLRpqurfNfANyfPbhDm474OUdALYw
lBQyJrjHifg9ghFdrNZNMyOxqnXPz/RUgCK66UHfMNvKa0L+bfE9x9BYqaNH5nt2swhcCBtr1iMP
I6p3dRpAuU7OPuIxuCr03+hG54sFeHb4O5x/0CXQVeg7NS3U+dSqDPvXQsJqUt2MRdoIUOtVozBF
VpgBARKgjKVir9F28afKedmrT1fh9X3JfstV4CcyA75f70aQFmlPB4U95hhGe75wZzrCkhROekhp
bCGvqaNco88q/R9bgkAPq8HIMM+Fnoc6BOh5IIPJt1gvTHjFlrmQGR3ud4syDKwdZ2iQVMwyDzZ6
5F57Uopb0qSAGbfkl9GLhXyuOxJVP7vBYifZL0+2zJfqiF7IV1QL8IX7jQxE56ElZOzybnoFlL2k
ACjELBcY4nWqK3AY9e9Tgf2yyiISUDPLVQBE+pUndtqYxOefLRiYYHwtC1Z/KxLA0E++/QSC1oCC
Eo0cAET8DnnndyFkauRsRa7dSIdNhvJ+l5Nq93siID+B2w9UHHe06w8UhVmVhNwx0z+gqdjcn1ef
/CB8VCyth5aiGCAUblstXA366m4JArQ+y6WFLuy5BQixiPHrVcMma7KNp0RpI+fwvzAPRoluIhRh
Hgzpq/Fkts3CdZ7jU2zcBHlX0EQL5k0fL9OVEwuNDgw1y/3IWsQz1FdXJSyBEJ7iEIRfrB7dGAx/
H5h5Sl2oohNO+BRHiXEbvrFtXpZYDrwsYRbd2RTVnMslkbGABIqE1N/YvsZ+ZLSd9rmxFAlHWgZ7
PuRlMezbFAtKkJdiRkfDioqQGFyra0eckO5GCOnpu4hkpsJcdw2cLaXLKkcFBg4dkKQRbWlMOm/i
gtK23ccNxLQiXLWRIEjmffOGkGnl3qSUiLFVhUjfd44Lpj/VEMnXe8+rqRhQqXvlq6lK+Q8qWjau
cAVbvB+OJKNkcu+vGWlacA+PVqcBwOv6/1eGYMKqnoepLFPXUTQvX4+zLyTnv0irnRLmbQnE+45M
mLkqtwpYQ2qXmYRPHUUQC8qu+GZ3CKa2WoluIp6Ye2LczR0b89uWpggY/1mdDgetDN7vSGy0RVlv
lZRmGFv3+VIqYeR7HlBoKaHlz4LUqkJ9Glu8ebUTatSbT1K/nSJ6WS2ih/l8jG7rOu1UWRarQzdP
eGlnQtNgYPCzsyE7oNowcG3coKiP6jLKvLHYjeB4zAG2DzTydljeJMnwsWLAdxd+HEZZ8zRijQGm
DBOPDPnt7JoP+CI21SkFO7qpY7osCppFhWuAc2IQZ9Ez0oIt0Ma88+V2/7b3NnGp6c6AHsq8YLYu
DZa3JTviIFzaIjUCsZi4XcttMyZWcNdftWoWAKE6r3WeeCZar48aVPNuCc5irbVdYfFfrrJDMegc
7IsbVYk3yUiODkvMX449YYdKtnShoEhcSxrz2CvDcJa4vZvXnAGOra/+q9yUDXfrxyi3aclk7hzo
oVxLlUwF8xNBx/7107eNKF8D6TkL8/inn5+IVZeCPAuA/eRdRqtcRgQ47M0WQqbh+X4sI24Kdnza
WgkjsyRgTmHfIyzzEnnf88/gZ5XHoyMEjmgFi7DjwjMBJBC0s0wBtrdz0keQQiBiYrSt3dySwWK7
JNOvRZay9QwvGapZa/YqGJWmMIDHJibHZ7+wye+KYFUI35YkkhiJsMdUEboAJUTN3Gl2Ywjgs6Kt
MRS2osIVeiDHevF4hRdrpx/iBjkJtjXVewF2xZSWmVM5ZA87RgUuT/AFiD3XbzHsdYJCIrjr0yZ3
xy3mx5tFnwo7IjQoejb2RSbJGSn/BrpztP7bGQ5a6tA+Kk4L3J94FIWFIM73yfP59sbZychm27a2
aJGJf2jBsHO3e93tLeUXbBc4V9D+FSn7FTnnwAEQ+ONJ/IeHkN1djgXHDpJn4mRZgcJ5XVzVuMGE
wyEqLpZgcqGTr5JcFFBdYnw1nO4pj805SyYitSaLX8NA3wYpu5WBfTL6fdTDJ90XF9INK6BB4gED
OcvSKHYNlk2eskX/l69bjWOYDlxbuA3uftUdrPTIYaTKX599fLMoWPV4iolAUnRxVTyIN9pKXBsN
OBSAHIDWGjiGJ6anr6yqm4OuNKlyIRqyvVaQxMFbCs6cH63yehCEdMdR7iyWc3mu+1jRB8y4QbT4
wFqYVX7YDLRs/PapHWdeGs+5bRKZZ6MqqeBP410KmJSsUHTv8YKiToRwoO3+rskGDmsTnSrerfWy
rIvaDYs9KH6TkhrTknTWxoDLrccZJt7Ze/e2jlW+/xvLhkSR3h8YxbOkuEcprHUD0aB/NpCNMG2n
318jnG4E049kH367Z+CmYegnirFElIpKAYMbsDOjnl6btrVnP4OvgywPt7c/Sj57smnQc607MmEu
NtvtIbFE1Fy6SyGEA2mrz93WF7E1skrzCan3gKWjMHUIBrDXXBy72NmkLdE5JX9mH62zMb8MUZ+g
AkfNAbbjifq9YaWBu2TyOzFMLCquo9crAiOxOrAN3UTNQPYS+EIANWUvqn9bOrR9KtyKWLw8RzbF
CZaibAitYF5cttmNEEiZ+qoKoiVLGQJR8VlPulUBEzC84NQo7t+V7TvQPryn0IiS2H1s8U08F0qH
rtxFhdFNV1m68xHC+iSlMkVbRB2PweJvDbJ2IEPgPwUe+XGXdROWcNIUlvcqV2UfMr9MbKC8UPy9
36mQ6gudF5B1RsZOQv7HbPe/9oxPzpPv6cJJyRTeCQzGudQUhRyH74Pz06QK0izqj70AeJlIhN0+
DC/NvpjRCRV4UnT6xFEHRkFk2B1roMPMreyFcE8nAT1f9Jaoqmc4Pt6Dzthr/i8D8NJFTQPrw2gZ
1t1M9uAl9ehZ3pqfQbOm4KnRt7BlZRjiTRqCsi+ZVeFKX7Zy4er1ISS3HNPJ9bYG1QxR/TVbSJeI
8JkyHWI8IK7g8KfO6BUYMbIYzAdFvRhA6Pyx0C/HIkGRD0xpgYZth2yZjC/+J0i9ij8/SUmP1Z2V
HegkiWMrMrloS2uLNf827mhyDnt1b8Dh5sOFNVCrDskPRzNgU8OxfG1GP/RwE+oJ7XephSvVudGr
suJgdHcWgihg3qmGQU+ZhWkM+MqQJiPqeg/YzNqjoxypV+54Ymo+cML9rOXtYaXoUIP0wxiC/5ND
XbtX0XpDFb4tTEP1/LZVEPXr8zuZrIod3v5bN9+dwWHUCZCgyiM/NxstN1CZIeoqhbl0W3RNu8vj
xgaxti4idFcr/jA4sqyp8b67ClxOtqsv8Mgm1bIAQz2rPNjzr9Mt5vNY7jib7sZVTqMbXypJMg30
pBcuHpmJU3xfdsQx9Mc+y4qvYnREZn/+YLDH+JktERPjH2uzjHCkSIgahQR6f2BKR3zEicK7idIh
CWojxcm+niSU6axzVpne+kYngyCroIb8IKbpaiDpwZ5UapwxAtHBtL5Qbr9hPdPSA3Qx8uELqaiV
G+DUhZ/xu3OY/c8Oytcwk9uB8x4nxnARsL6Tomsn1ln1vGf6FRJHnvscKFWb78AJRnpXBg/psTdt
vmtyPgUbdyh0GTDChAO+P2U+Al9e7Szi3+zpbsiXzWuK4LZcjukuWSRUV9TrLhRx5+GxHAWbTHZf
BSueGePQ9GxDNYIlwgwlG4a6j4tkpxiJP5mXP6bTvlkawKzGDVnSI8c5e8WqbF4bm11eQQSPVVzQ
KjSf8BSlvuPYwWLVmMZ0vRSmQQ4TInJFUV1npIme4G5A493NdRmM0c/7Cll5Tk1B+587rBw4Qo9R
O/VLa1W7C78gO2/Qt+JGkh/F94e84nm6donICRrdUkJ+gnYHf2LP/S0jBXNcMjoV2q9Zz9qr0wbE
Bv0yx3gD7aa0OV/0BWTotNFuxTuwBBbghIh2LbegFvS+qGa805+rWR5wgmvyAyUKtZHi+9KIU3h1
ev3cRbiU6tuxRBAAAvbugxqIjBhjGptvyoO+IDi4hDCYjXti/lP/gESN9q98nypG7KBS77dLq3SX
slB2TfyubLTNRfxTVTARmSL17sZxFVO20rN8+u7r6bU5mRUCuQdRK887n1sdgrDCF325ZZsfOxEN
wzc/UjUOc10oZ6lStC3/nGOppg0oEebNwS5saIWvmQgKYI9p716ZaOH0cQXMcpiaUCQXg6uKso2p
tO4Zc7x8RJicH96jaLat0ZPMksCFueQaExAubqcBxe2FicooJMbcuKckyVb8WsLFsEwA0zpr8QUq
d83i9dIox/W5GIkCMJizWMTKfPvfNP4+16Z4ClrYlfrH/Q+xULqPlRYHvfv9PuIYl076imgHhGe4
zdTlzfwqnDJR6Tl8HaiMT6l236S3jbT6GXHzlkIhT/7KgalQMmbet5U/Je+bPEBcEPTIhusYLQU0
iDuTwoLr9TgQWlr6/lr2XBAS7QuqjTICEnqVZeYDF5cGQWKkrMYTD0+TVoLncSJQXFt2yviE1Ti2
NPPO6Mg1P0xnuwk4w9MijnBbLXKjuAzsZG6Vmkm1ZIUYiicb/rJwxASb5JeI32NOvCIPExuhOdl5
tJ1eVDUfH5pHpq/SXO3PxQIIRyM4SVIPkz73Fe3vrCHlAvXYliKN8Vz+EjVNoGOWGjtikznJAZWV
t8bK38YCnK0GGO1GUESsVwFA1SWWuCm8KZCqHYLxWvge7HejLvDvfMjcrPBIdYHbvynnyYOCS+sJ
qFV1tFmxzR9j++vqiOZQBg3lzUfB3nOiZHca5ZrGN/4yoy6I35h1TO72tdSvfNg3wb3a7tB9duDc
aGdFQV2FjzNeBS/ogn0UAwMbN+gL6A10lb6+iIrFemx54Q0R/hweypKP/12+RzJ2cqg26ubKq1KC
XDDLWBthcxGr0EmIpaxHCZb7aQJX/co6F4NwFY7fvXMFXhICjP8H8514f14JI+KVTBscQ5NIuDNc
1sqCcgYQHCYUjnmQolye3h0PomvKxg9rAu2oVuEOYVS/L9VNw8PrU7TgUvqCvAmG9q2zMZ6Pzt5s
Yff9vZYitaPVYZ3a06W2hgxcfTm4Gk+eH2VqAGV9NR1rdHMDmDmv+20tBQ3M62sj10+1lbolXEVh
vywSPC7CehEhpAISS4b3OhxdW2UfcdH40xv8PmyNqQb7kWUudgUmNA2YqzpeoiTLVgdfsjHYKd0A
qU6iruucVytEvBTlQ0rb+WKEmFFmHwIOzq0W/YY7fQNMPZlmqIjWzaKnihpm0/8/3Z3MZ3d3BAZa
EW1QM2LJYc41RVuZT3/gUaMS8xhUlXS/vnrlYYqPc9HE1CnY1Pxt0rByNBxwujTw09IBXV7QWkW6
UlsZ73zKJ2sHCnVlKEa/ZL76UNUj6mfa18wzStV0A5gn55YzHLSIqf6BTIBuAT1DdwiE+EBDEgip
iEpklJzSAPvkPmJZnRUWaarCCSw80S+ZwA2gA/wu2ujxeWKfh6yhpri7uvfgI1YBn6PiKwcYfwY5
veFKVdkqCfFVLgMDO4vP3wrMI+qV7Z+HFphNKIujLUe6uy4w92JOpksUw6F/drLjLHHmx1poADOW
4sBqRFjjs81ZgJpVarlodKSgyaSoq6ROH26rRaGgCGrMoGI642FVwlGt3IeWfWRgYbBdaaSIoDjR
bJnxcQE8D4JY7Zu3rPtR4dmVdgnn9twoPvZEk9NY5dMOAcqsvwo0hi9Pi66WB57n5dXO4UrQGhe3
wjxbXtjK0roSIwjrrvlrMJcizs051BbByAKsQ7/Xo0k/NI0gDpnSyqRgRmYDhWWnKxwO0c0zJh3M
SyklNvsxwlXdAyb0zO+UgigDFAPJzj0WR2dsU9bLzPjQzws1euT+JmIjd3D8jjrHjHs3ZSXFwF+/
7klKBxwn3yFa/UUMXuSqvVelR7lAkoVshb0r5ZC4RUgmhCEuf1qjMG1BNZ2HLghL7bnSqnN7EQIv
aFq+U23ZjHvJUtGHs1vYLFyf+sMn5Vo+0lxCBii82ePUY0JuzZ1VAOfCKchgPGWhpAexHcLJPbIT
4AQYpZWBDGmDURtFBreNLvcJqJlYPPReCYWNbDIlV839aqrfwY/2LIiVpOjwEImzmqpkSRz+VuyA
ZvCoue1cy3UdIVpmuarGPQ304BbrBhNCSqz8Y1kL16HEEdz9j/CuPiLXV4KawmhF4X/l4jLuU4fG
8O4hXCiZvQpFYbS6GOKaQpc4JCCXiByPQ6DSTfgSmRojqWehGrN8rikuw1YhcesVHK3W6vWGyZeS
MqtBJYevH3/woJlSSlLnzRkeCskd4x8TS99IQP1g7Zfs/k5dNUsa0tQ8Q3WuQUwG0ibBhaW0ws5P
I846uGQK0n5kTVYWAWDSUtZ2u2k4JDxFYsDOpfTNDaT7bvLaaagrfZBPgHivnGh30cueSzGTkesH
ti62GHox1S+8ulO5Nz+dUPH20Ef1mqD929qwtTsYqkAtd5ZohAR0hKFMdyxqAI1YMCWjZhwP0Bn7
2lFupn2RGafABfG3O6eVvtdz0H+C6sH7EDI4rT1lDq+/1Ke52SE5nmUT34UBbiBIBeka3ukh40rV
0YzCQKHRceN4ZZcgJnNbBMELF1fxSoO964URkFSNCwacj8YceHBqATztNkFW/tKCXwCG/n35EBc/
4NxI+a0W0wOw1aUU67r1MDwVGiSrKq6fqkU+e7TjRbDuupVxnCqGuXlP+Vl4hmYnFCYMZbCMNBgz
zIP5lqhZ0jukQslTvB0imkiUmjJbP+Y8uMLsAqe2fQBjoxMJ3URCt0f4vKBnr7wUn/XvtgrbOmAd
NDcEm8ujCLFqu5H4k2JpVVoFyN8mEQDXAJGKKndTq61E4jbbpyZ96HxL3PDdYEcKbc+8AKSUgqZf
oe5FcBjwl5Gc7xjEcqGkkyuXzwi5/Nz4lQ1c+pqB9QkE/gmhPkI+9iNX5h7a+5UcYzOlc3m33cge
U3ZiKa6AS49ySwv/EArgcPiK79U6G3xh9JX8WnTVQOz7mThEA4ItuNMwJuIX0dDPOdxxExJbJeop
1qKQE1G4lGvtKz+FI4p4jQdIejyQj8ug2FDeBWfoYfi6vqGMXgAzxyxdMxQgHdNN7Cnc7/HZAhGu
/80LRKcsPdC3w0phNo/49M5ZlBr22kdD8PKExMmGYrBNq7stzFGWRIzvrjIZjH0lxWwdps93BQZd
CKhuc0QLiM5AY1hCUeC468IPc18jF/UqhFiMxeSSkVlb8nNzui+k4se0wJK8SWJuyrkjts+dv+j+
gL0G/ETAPrgrQ3zzCPCLJYlbJS7CKQ0VceKgBhLEdHF5J/poS0syGxn2r8dEOypyQG4LQMVZdiVR
0yV7+y5gQ6Ol3q2n5mqBOKmMs5w/yl1DKy5iWBh91hlNIFammUH0+EWtfSSxVGE54vm8MrqJsok4
py8dzVKEf/mpmXEJC1riQkGz1dAHN7LcmSE7asYuPa7s2hYN/NUmNmygvpqVkS6NWsbtLpR4HYAs
tj714fzuE8y5N+fnf8DOeTuGywRzCtc0+BHwsZbJ950R7m4QvbG/drA8esyDHcS2/mVx9CoOmoKM
MPdlBFDGwayUmDwOnPIvlbJYR+SnKcsMhicU+v+m0006dfFhpHal2ZuooTrf2b4i7LAl6Zpogx6T
iAsdF7o8Vzhg1rDH1tGg6bnEbxU+JWFj6x0TQBQsYkbt192XwjFq6ohoU7xLO/puXMv5Lrhs9y7o
56J7pgBkoK/z4TFX0MeMZcd2F9CPqyxRBIJpmBlhf+MfYc7+AZJQBe0/htRyclMjppB9WTYMHVVT
HPl92lomNsxAy75mLrQQ4lXvqdIY0FKliRzO2bT7rOwL5wcvEttOvngtIgPGnmlhHEQ9hzuSJrZ/
5rB51iIejyrjozNFlvNoHXgiC5oV/49Wca5pTHuBro9Rr4Qc32Y8JDxpe4pjoFbHpdi3UI2IQoqx
79Kwt5sTz/X8MPcZLZQUczJC5wMHGOIu4IMji0TLpJOQgopnODRgzflpTZU13kWV20adz2Q9I3Za
N0wUYGIX0j1oWu49JEHjKofJ8/PvfOIBUCxkAma+K46rxluSfgLg27Vhha8vIxG8yD+54Iwh5uA2
j6xAUds48yCMWyot20v9McUnImTbiiA8yizlXHDnCqknjUhz8rBwb2Fay5fgocqrBiMA8Vn2zLd5
DkaypFbLiHmpv/RIXCc/dKpsotqOvZnXotlY/B/iwI2U12c4U1HhQQxGPz/QfPx8XJ/RL0qTILsC
0Xek8z4KbmZUj2UouVDeZfYMGnE8UiWBcL1SRRYG8ggbOM3fusqE5vWd7aVrFVjkzupUo1jM+yyn
r/iBX9kzw2K37FaqlWqW2NwULU4Izi3L2zx/9G48Q232JPlzhyZ6o3iPKsPUHmOOMcEoaiApU4o/
7IlMgW81QFek6SkNT+h6FCQvcmxuJrN5YFWMuDHGysI3at3WSfpAc9nbwI5OLBK/s8bhI/8EHQGS
XlaSrWqt3escZrhoMbXHFQotvpJBpnEbxJEA1HwxqN2fR/unh00DTqFgBYAy7fASP3WTzErHMtt0
qcMIu3OAgjMl1B+xHpCtceSmWTy/0NPUe7WQQR1rDQv/+T+PtGinIvsKBHGgdgto/EpOBqS1ldxF
+pNpfhHiyjiQAOPFKWS5T40vmjse2U+9mfrcRo9YlpVuLzHaxAVzwIWdGaQYclkAqt917OAufDMm
LkBIZ2SwGmsyE7CSY4lRkgIZKmpoxjKtpuwlwPNHMs0Z+btb5kdkrJzMB6W6H8hkWhX/4hR1Zey+
Cspcax63UeIETATsHhSCsIHjNBcBOKhe/zS4mHCC9YLZ1IVmmCHZneuf36nHOx5Mqkym/+0ti8vJ
lnYDMsE/qS6pb25FM4tPpaJP+XZnhojRqb5tw0Bkk3XudGEVerwJZMTrwnuDEnc8O1cmDe5agij8
O4aOguSc5sDvKIRs96ZkXe+9fv1oJw5XFG7S1qrHGxSiyA+JUzUQcOJL5SqEQh3wN37DXrndkAHA
01hzFVjp4QLjXWtnG6JBfishBhyBfTOWH60ZULux5krC7zxjfYjrvBjGFmtVCbieuCkoVUg1i9hZ
eQ5vwdAsqkwWREmx1zSEmItGEFZ2YF8/f/sVrsNUxJ2bJHS+IPJf+G4D6NHC+R9Z1pYUCx4PWbeR
DOIf5lvo+H1t3o8/VUTUgNVk0y6zAuwQSqBPcHZ50BVZ4vDg6ro/LIx0STLRjugOzBzThJzcNELl
PoOR/GjKpVqaSVuAqWIL+fZNk22htGU8nCO5zkzO4embjWj7+Fm3nrsA+taHXh2m6C3Gl15Yh0D1
NosOVdjhp+Cg8VK0qaL9u6lEKcjLTkR7Pe5aK/dHoyhzf3ePP7ZMhqvOYctPe51iNyNRcs5WUIg3
kIY9snkFoCIuvytXQ3+w7s7LoL8Ma+0kihUhhUsEW1ctIP62eF7jXr84j2gjpOez/a0EAhqssFJX
pYDBkUejWUpC/sspCvdkcwe6XTsPeHN4s7vH29gnvHpVuDqEVr0Nw4fXMrxmBqF6RRL5V6OIzGWq
49I5rPElolp/LLbXiw4EkECM+1KSONaviWPsZeIQKEdmuXWZwQRqdKWsDMWnfAvvWTiC94U7w8+Q
fFn9BA4+QFoiKMPuPW6CqBPx1WIp0j/cNGmGJd5zYAwwaAFrwhxDF7ck2aA7LC5qZikyhx2+Mcue
JXwkWz/3lJayxXMGtDO8uaGrIECNd1LIRqL+1BLhxYp8BS5+OhsXIH6Ek1AYW7grCinX7UfN7u8/
879D7ajM3t56AHnMWKC7BraIW30EWie7T/QJAFSYk9N+RCjh9w9GwjI97EFDPwre10P1sM/wiK8o
9UoirMXDhVjjZ+efKNBBgbc43LKA2fWre7zzO3LQh7pwyi+eXDBTATWhgcpqF0BXqtx44IqPSjeQ
rbCYap7FP11lSFsELW2JlyoViFXuTPs9l3E7L2pELpS2QpiWkh/8EuT3oNgbt6+g8yn4Pd5uw6rG
FzHfR26j4XhwH/FaiY5rIZqzN8XzMiTdpnLUjoPPnHLxuu3j1f/zxSiXYxzTso7T8rqHN/V5luXr
OSTt5HGP8g3Jwq/oaXd7slRyKblr8WVwUQnL3LXqpjqcF75PGrcUEOwckgLQS3lJgyOe+DilrYQy
OIqiG3wIj8n/c1Rx35LaHvOmYbsrcVgGswcKcXbstALMlhyFN4zfwbOzwJVx1rsK10Gm2dNZFUb9
+cx5qRONSm8lszXW/Iay+NjSgnW+IPJkQPFNWlPi29J6WFpmhiny9z6oU0k2ereaET/4/0S+s+KL
0Dhi7IK1EyjyyXr3dxWh7GpIUn5BtKm7qvCfC54DhUGB0Lvzx5p3M6bhiVTcNmzN2pie5d4VZ2q0
s4wdc9EwY6CVo0EzC1GiZ1QVowDdpsWR7jV0KjVYThthpDEtNBJUtNztQ/QS+JKuFgAvvDoYErTF
0KZqZnYs0dHne6+cNy9dsOy01o5prgPWvuLZjaCu+azU3QUTU1MiXOD/arbJ5MrRjhFAtL4COHhG
WSif1uMT5MBjlOnJk6ngvHBaYytxRSXV4Vw07+PIIcMn2o1lcZT9UUxj9rKTHFGqbxpt2Wc6Tnwh
ByQgcOVYAEwAPJICfLUJEGbfI9yGOoAGrofP76f5wNxwmHmEEeZwv0Z9Pcdf+2EtMlfMymQcUQA0
AVVLr3LTDvz0QhOn/Wo4GFG0+dyDotd4rNMwlBe0Iukyq09z7jwojdQgEaSeL+cALskfMsCyeRdr
L+s1SbEf1HVDEzshy4FTSaG/5bf3+QW5Qh6RQd+WTnfIVv5ZMB4OCSku3Oyof8uMytEjNo5rXuxf
MeayvGe4+kq7J6ZDyLNIhxWHk3FFkrcnaDvhTIZ/i36UF2lupWHYpBoZYoVN5U9iH40ntY2zRj1h
CdrWO0Os1doL58X73RvjvKATNDZC7eJIfTFNy+PvlMhfw69YBPKkCdaAtlQsnKBTcZLg2MgmEmoF
qc01rWOnmT7lN8nbCpMe6hLPqf3ZqJ+2Pv3yeObxGRMv0BHZM9BLxeuDxq11jdf/81d58hZNu7Mz
Dy7Q3bxPF7uSi925hs6kcVI98vvrVt54smJhIPQ05wnSsmH3CtU+76KBgdIyZZENZvTyCGofVPGI
TA7C7BAcKAz7y6kb+aaBmBhoKkJMT0F3bqYGe1KhLZsYIY1YREEiiFgpbcNUEfHyQGdkoXUUQ+64
yzcecPJn+O4DFOXAX1ztNyCN5pNRfX9EqLAlwmwE1zdLvuQnHzTvrqCQzzw09QCvGiGKk/8Cv3VJ
y5n/QF5VMMw4lx70+KWz3+wTm1QKDDphrpSrJ+kEBrNvtFTXaMZBPH9JpWnlt0XrxHo/kfLUgozl
rSdAuiwAauGB6CIo/+G5Pgt8uhyd21yruB5MgOWxsE+kRoyAIbJmHwbLzXFrZ4B/PkCgclYPQIz3
msl4ZDYdU+8W0cT6VSYpGzULsbyVOjvg+tUSkCCaSrEI9IdqWyPkGDFR2oP3fvzZSoPsFup5EVus
Xxml7ya+uAnh+ZXWCoe7zifOhVMiXgBJjvXIiXX0N58MaPBigGBszAS4tCQYxiGh59p8/iffsQk0
8J5nrJc8Lv67f5Y/XaZ5NzJIoU578OZgs3JKxmq//dabTBg0pN4U1rrlJ//5MMyiCGbW1UD0Egjf
HylLVU6LaII5t44K8gDsCX8KEtTfyGtUYidAjY0NSEC2e6ySU0JKZpeiOx7X90P2zwrRj3tgMM/l
HPCHK0N4A5MsZXxupayJQZUCfhVZAiwK9T5L2/8ER2MTsQVcr82PEJAC5KsinI3oGJAJIXckoHBe
zxfp3p4gLIA28Dng4gPPf76FnG7hvng1nyIVTr024d9j2kySubKuY9SeqYVpwU4X6Kdx+t9mMSZp
BVjYU5MAb2+59ue/WDmMFh24olYdIVJNOca4OgKjwhXLB6CXxvL+RtfjZxMvwhZD4jYV1IWppCt9
AZTcvTFNFBtR5DS5Ymb7uegASPSamYzO1fEHG7VWYXWg+PxEheCk7YKjw5JAqR1GcuwFc+2kx1C5
9rXN99bAdhrGJkVoUJBPvlGBjyqR4zend2n6aRpUzEgLcfoQvTirnJtR0cmZqP6xM4KmqKjp47it
WZ6qr0a82zPnzZR1h/s5AOqIjcZpuXqwgHvC2y/JLLW8ka/G3c/JHuJRtbfkqDZaYhHaqUp4/5Cq
4X14IQ5RFvopTxaNvWzJ5+h9AEy2dePYeTijbHi+BtQjeuNam8p3bGu93HxYWVzkV5ryQImyEUaK
XNMorW4Tyfgt/YtirKgkCzV/j0sZPoDftA0QTY0WCr0phkSqIhTzGTP1oRYhguTSv84+YDzlrzOV
V6YHe+DXPM0P08GyeFaudS5amgHvLLQOzlgJWyXjFBnHrBM9FzpiJwqgzpC0Ki8NyrzACNmdSSMe
4ux7JuFC1zYUT3bNn+kt/CHAv8wmDxpL952M/LzyvFt7e1X4Gv4WVaMzYHg6SoMLuAPFGQ5CtPia
9KjUDz6VVtg+BUELBNrOhHhEa2o+6dPnt63dKFOPfIjE0IKeq6y+F054/7pwITs0a236fhQ1hl9Q
OUXcgVAHM5qfhs5C05B8JSHH+QPUaf/cmg59qcV/EUEM3rSxO+6NvtIJ5udkcHWaXOEdk9KSnylf
12UngNrbNlb5cbffnwX8YDLu8oH9a80RakwFVG1HtaSrG720/U0xw4TuENeFQU4AXS3uROY7stZE
MUX5GGo7kPXpiHLythFTGwM+Nscf6er0cvZ057Ia7C6xGu5R8rZZeim4kpf2o6rbnekTbRnxY9U+
LYk4E+aoBLDHpRu445ZC1k8ryskJIr4f/+SoLlH3fzeAKAGxkoJ9dQB4i1vlo7fQk3gNp6xAduhe
0lXCv16rR9ni7yuDwO9tnk+EJu2pQXqhDkG4pB587aYF7ipxQC7r7ZxyQLbpDQRnflXDe9T0rSPX
XmbbfKOyFsFOgBeYPTV3JdIxFOwIRs8anyBFfbRQAKJTLPnI0J1m+E5Ic1aFXqLDGA/Va7rIzvM5
PY+XIXaOYJXtQiSR7namaziToM8pC3JZkProUePlYU8bnuIT9GhAWT9/0GQsng3AXZgAPrbgtreh
l6ALOpn3tZDhvG4CHRWHcU4UoDAsW/xmSxq9HJOsi9q/DKseFtWvwgDuvuidJAGhw7mxHjRrjDPq
7xSGrZlzmqHQZydzfQxaN5iG/1S6xp4ZwXdYg1/oS6t64dMxGbhfi3XXTK5YfXI+z8pkMCiTPPqb
cuDczpR1xeFNfyAAc1LFAcuBl0aGP7eI1u+Wi03kDoTKBvNXDkX56BI5lEKDTlFRQQQyeewJwdqP
t6FPMB13uz2bqyPTUsXA4Ou+oKi/0MUTBF5zTm78RdepyuOfYA+Zfr7eUNTO4fTKOx0nR7XGjDcm
R1qhPKfRXFlfLXMJT86Y+9UbHtllMrPr/A0abcbefupz4/AbXozub0Uuq6D0C3DsgxZzKGKqzrgu
TeP7UYhvscFtDzQLJfa8nXHwPwDhA+0HCLZNoyyeV5YiiF7qhXnTGKv5+yLYfzzBEA6uacWfgrGr
nBZ/IyO7CdZcCMYLY8nwH/m/cokZWxUnP725vMtUg9u3wWEUMBv3zR2/bcnjawJ98HpgQuYEzNGT
r4EgXhqxHxfCHbURQn2UJTk1sgW+r0T1rdmKtcVv2NJbuYMa3SB2NNIZZFRODsZsX5Ht9dm3OMFH
9pZftopalLfZgNUfvmaflZl7J2GDG7e4yXRsTx9MZiOhsvVvDHNqQsqXZp5q7Qg9I/z0lZJoJCFy
hLYzwTi2noAKz2qxr7IDXL5/DYT8K+puDw7MjjdPTiynHlPu2KgCL3cX0Bx5CCsaR1Jp6eo9HJUR
glcXII/mgSpISAvh2kX9mOAq/54wWZrYHCxkt/EsrCgctG9L3XdcbotN4sKlnHHQOZfanv2eeXEQ
JteXIJknOJqsptNu63QI3rHtOq0b9rEknroMTH6aoxgyLHfuEfEg2Eqe6RzqfirHJ/uSyQcBWLcf
I87distJpMUbapN+qsl/NfN8uvAEPVZH1UETcn07JqHgoOEvPxtqLcmgp1yirhVK86zcPSJrOXoF
lOVVTjXWymP3fdAv/BzgeKEosBGkGPKpcfteVeAxG0IBIRZ4ZAmDRjXkCgbljBJVWKpBZ3nk2nGn
+kCgBSqeCxIRPSkjaLl4iBeyqXJIUaoVsBOHyx7D1p8wCWDyZlMijt3AoQP2syMOpaN1rfnUw3cg
bvL/1+oS513jLvEf9AvsgzTU+XLY+ZKfmgb9L7jehv5g63Av3gKKyftkRLadxY3XljB8U6/6uEKO
TEUtKM8fFUj9OEvsrwDkEQ2ebJ1x48vsg6G761PgoTCbpZU0ZuFnnU8n87vgwRKKhFog2uTF3h/5
U5T45tmdtr6vav0joJ8S57KKIO+bCG3zHsebP4CFvc9RNAO2qZEnptz3W+zNDw077cA0v9urxkIG
J1LbUFhjC2goyfKobO18ifxaYWLix0XP7a+ucR7TGcqiLcRt/4xhHPmLzFrBuJ3MvJBFOr3LM3oh
KheE/WU/GVRCRpApdiLDfDCwx3Y1zCxYB1mqDIa3BE/B3OMIBrfv91oIBZnYjG61DYUOmRO5Wk0Y
jaMHSS0qTDquTdQfzckRM2srNv/CIoUb+tzKiZ5oi+iopsjjuWxNJB4HLBv3iP3i7HQEFOVpeBe1
pXs19THzQoD5KGXpgLVUuJppytthRXI6G3n5lGl/Ev49l0eS3S92O+FgqZjnW4sNWsK17PDfOHIR
N9WZDtjpM0LNSEaEpjqDrSZ7K3g/0DyeSRtxYM/3S3kSZEuwY8Z8IuphR5f1NbU1ezCPjr2U8ClH
AdrONFr0/VAEwzqaSU8OkyjGCqsefkxX/LotFrfJTq6+LXadwAaMtZRijhdeCcnRmLLAyV8l8GSk
SMhEebmpNVGr8n+ygm/oZUnrR58G2r/V3w91xUrYwMjGvbH5ByTD6VEU47WTI1WUPk2iNEA9twOV
i+v34lQIqBVXIFjhPonqcvDWszT91u99qyTw+AR9yFRLE75KRRlDBO+SL8xL0dNvqrTA4zAX3k75
dia5dKeBIyJz+SrfIiiAigkwb2Beda3KmO/1bpF0cZoOEVc0UWmjQOYE0lIFnMkeLqZYhwtwlxwH
I69tkYmx8RNxh9xRe2VV3ogp80qJOCY3+ClczhoVkD2Vknxc7+1eTZKTPIQq30iUrPs/uBCgOiip
feNoECzOh7wO92r26MuXnXlpSJri0b7jdOVO0Qtg8zUHmMFD7KrB0MtKe+yb0KMYxu6Lm5Jhs6zs
d/PqYioDhFRtG5iVwZ78vJu0NYt61VLlg+AfDNF0Q4+4oPH8iOI/NW4VjxxyIqjZk2JNHMspmo1V
Wi6+IgT8uni2bVX617YXchaRSk2E62GIzXMUSSsOhLyXHFHBUY9xp2Yfq+6zRB7VpJsh4pa4cPbu
E3afq5aNSkIEf2MXVx2FtTPp/JE2Ty3GlA/lkqedRNSPCW/RaMnqefzEfOnpHOH14NrNGXE77WN9
ZA/Z/yKQiyed7MtlYmwcUkKtKYhWBY95w+xDWqwpG/gN0OuBKMWX08lFvZ/usvM8yz7ZysCc7i3n
Fk81ljf3KH1zWullC37bUax8fjyNaQJtTZVsNR/XhSI41Jr9G4HmEfNpx+WKC0GaCCuxRX7nxvxm
zHzxxTsYf5NpDXuCOz66kSNJgnwTd/YZEe3KCc5rtiROh9h0j89ZYrrUILeoUltzsV2QLLsdTtFD
SCh4sasUDglJU/NDjKiK6dpUbZxopRWKA+aQBSq1ZXNxnQLGbDQ1tXSBcUs3tWsJ6JHts/NOf77s
MjavH3na0RIG5/wis6t6hQDIz9jxleWv+XxLrcKBIhfnU1iPE2IZCcbLkVnTGZrZvIKTTyU3PaX/
KWNWsB1JKiorLEt3ZvS6vUkFPAS2GBQnCBz8IRxFvEez4Mq7RMZm5S17DdplRR5B7zQl6FbbB5OV
kX7D7J5awP9aMZm1OdHc0KgMg3j40naJMVpsKYLqw5HtPkjj41erduCEPPFe0shd2XhJSC5D5XkD
ueYySZPsoPKVuajnf/Gs5lCwsDMfY2mvkByH957ByaSsqcw6jVOC94riU3zyrkjAZDqOQczVPvBe
8HNhsYXKc/8B9LIeE4jQ1z3Zfj+3dFpGOWvHAL/w2NsMt1/HEC0C8oHShQ0FbHvJuKNQhI9AgjEq
DPDsh1s+31wN+xominm8wfBF3TvXpAB6PC5AOQDcVi6v83Ns6pBup4jJJhFQkHGuJ05lSYGmZ+VQ
mDhFrbrP9p5NS+SICVKzFhe1HO1CB0g8d4sPtziNQ+oCE2olnZroZhpxJmkJJl8WGmoMYbhrMo0r
GmWIxkqubJ0HQlEHiJFH3KWqvvuJd2hiE2uyk+6/pxXtvY86X4NlvNGlTgqlih9qVWCREQCGBbsK
oieTvvScYolu9TPCkG8nAFdI0AzTgzeHhhpcK2n2ZCbZUtgvnyIlcWxaGJ4GT0TMn/wVygyhYq8F
eG06Qv8eNBD7mQwuqKMqzxsvBjSksVxt7jFQM90PgrOuAU2C87V9UP4eK8OHk19OX5ApPRHZBQVX
vn3X3Jjnb6onnjfi5V/hlI2HIlwhi5Z7DklEXK1XaAdqEfQHwffpRRH0255RSq5MfcmjNr56bJu5
+i7rfmkJFlAW8RFcxNncuEv5LkK0SWn0CKFTBVW7GLvUyoAjPnjbfZ1t2eM139N+XH0ZXks9UF7K
RqNyA96jKpQf+NbJm5aBmlzqW7oEOGSyWEqfyBxYhswnkQrOOB4sUdzMDqhcOgvpL4AGRLk90t+p
zCG/hG6WRwSdOAHCPWS1iB1IaolS2hqKUnXwVvu1FQ/eKHC9GHXXryt9HhF2LLEmxebWxmHsGpaP
t5UrGGp9ayCYYBadqh6X9nqKwtbRHDXDm/yTDd9lguY6Ipee95djl+fxi0eQxUp7FsZUlOKYFMjt
0mNlLjOwzJJPLerrV10a+1R0LVHWCyur741R3WOCkDfR2JdrZPaV4vMviMZmyoxu00jNG7vseK4T
i+H5mVq/Tx56cOlcD21VI56QRqZ/zUYyDbecixQs/xQhY1kPgFKwp7U0kURfa8Bp1sir707exX0V
AZXjNv8nSEwvnukvfuoHLdFuThzDIGSfNpZvqDBgtP1N58uoKpX/9w+uuo+Hh6I8JCTry0nw5iwv
cHexOWAMgUGEnxzwlwKpXeb+I6hWlKTW3QHpVW/pEz1oycU8S5gJEhlMCD8IEt3JgrRF3hh8IJca
QPKSKXdxooHAq42+sWiPrZaJ2mnzvIOBcizrRmLus0AFc2/pSWh4qwDKHKzPJnr6Ej9lxjIz9/19
sZ4TjYoM1cdnTLgln4g74QYHtGZ/xJMLdqS92PNM1PNbf9gKvW3BoHHeSJirDE8P5VFn86xoJ2n5
j+Vw5YUXdRdl2Xw5edU73U8hc0QkRCTyYHFILGrVB7QhzfplRLm5d0HB+BjX3XUppi22h/WsfYss
9CwNWk5qpTcrPzIupZmj0PQuu+DXKzhjMrFl8jjfZee0JHlsns5XWmS+33ynyAxXysWzz8YKfLKZ
2XmUGo9IH5yNz0Glhg7Pp0ysaeBm4AAUzRA+cOaDm24BY/pu2V51B8eiaiJ2y7iIh3kRXa0R8gC1
bglAa/qUJMoc3SvqCLVbEeIyJY7nu+rIMQXAYWKp+L0BSzy+hrivZq1hDlpay+zRD0s20wqLPWe3
xmFl6lrqUdW2FIyyND+eZRdkUL5+9T6H
`protect end_protected
