-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
HfPiOgRIwhLfCyWMt8Yd5G9bib75s1VKbkfRaoxArZiYc6DU1Y+8W1Y/ros/GvM1
NKdIWE9R0w3HU8rggXN/95Y6/GsSXhcRhIt/UQWEBg1rFJzHOYkTJIe9OXCvXgte
KD+iou3cqpB3vaB5Hu74by3Cr69X9KQNEE9tPJQ2xecN3PRk+vIPXA==
--pragma protect end_key_block
--pragma protect digest_block
KrOu++C2kHVINobaa0eAJ56mSjo=
--pragma protect end_digest_block
--pragma protect data_block
O7cRHIJasm5q45vc+UKQoOJ31FaD7oZgs3ldaHBS1xDJ5h1iw+63ljKXY/kt7Yja
n/0x2E2YDIbDjSzplEJ9/4dTwVTktJVwZ3Ut2L1jbgOg4OE3dG9yH5doS72lHIN+
c0CAfi4ca9etD6EIHvQ0m3hO8JOLgqalr2Wjqqhs/WsN7Q72RoKGJZVtXSRLfk1+
K5adg0NPz12fvjgMqYzyRtT3lISdMd/E7O8/j7LbEyFoXO3p2mqNzPA3ZvzWMUOv
S8nfRmgtLOxZ4jbqVFwAs8RuCN5M8m8TfGIHLSWT0M3IBq5oTjuhroQ6fJdU4hQc
Gqe9Km3580PCAk5AmuDNED7EDYAmNBH95peqndP288V8vUXE/kK0ja22xNSVnFq7
OZ4R+VN4NyMRHucC97Q8BChmjridWPOLklqJnWO2AtLjEHTA0qqHzrI/f1DlEv5P
KZeF2Jjxhv/qmqFlGw3s5vHq9MStN8Z/r67R7QlLaxJGLXJvpfmc1+EoeODyPg5I
jbcl5Q9TPSTvYYCY6Md4NhUU1Gvn+ftzPhS8F1QNTfAQB4H6ob7ClBJjEdx8ZrF2
bhb00/SIuXcrPVmOTB1WcUZQYhjzRUw7u+/5a6+BVxWJ8FBBylbuHmSc4863/ASi
fTKLgc5e/TfZf/TtdzvEV0pM4rWkv7c8WMopS0FLec+5zc1MAsLPajLnM0i72RmD
PcasagYOtv9loN52Zr2JClyCebnuQZ2c/aJXInMmQlR5pcQcsP6tq2yb64Ws7KEH
3JgMdn2V0m+KBC8ZfVoh1EyXbD8vdSTHPLck5RJlIdOcf4WDQCH9yiHTjn6+yPh9
5tVz/QUpNTTMCJCKNPCImIZ6dXppn0QBryrAG0Qko6UHs3zfdOtdf5FGbzsrB+YT
m16tp68NigQ1W7TxQgb6JcNzhmWtXuzVMIQcRYqOAmnZVZ3CuzCih2G2gSDc+sAd
Dvo/RlOglYFxe84T77V2KglYYYWDImkfjb89ZNG8DQDFM2keIR4rNMBc2r/UfRym
nMDrsz3a+watkN7rY6m+5o5WQl32uYwb5RytqL+sCTAEIcX2J5SuL7/v2SsM99c8
tr0rZeAlBdpIgriIlrefmSaCpZiRRnLfMa1YABqvCWuStx0akApzet8Q4Ofx5SZd
esBOHO2rMXAVMC2aNshdjdPut4lSPn1xUssiAEx0HU8RrAeB2broJBu7mgXVzmRy
LQIU2VrsSqBLsFDH0rQ17PlvcaUIEy8sn8/OxH7eoN8KI/JC8bV7uELCuGXX+sph
sneCdAQ8aIpsIp+jTgxC8PV8ZzCeMTr5FJOxmbteBQ1a0lXe9b1sjXqPVv+gSkay
Y7oiafam2o/njYsjxMA5GsNJbMwm+pv79yf3AdB561fs6n6YhiRVN5HxAOWy3Xvx
u/iiuMkwtvLfiXwHoF26uRuczAn4bFGB+i7+ooT8AF5r7J9obuDMa0zzlcJ/8tDa
r2YQoZhpQt+uotS8T01ilOQHv7MJyuy7pHrtxa1QE73Pnz/ht7lwdeADSxKIIXPy
M3vvwgameLTKr2aiYyezUvmUhibJP/6GLq4eLkDTpm4uOjKzVpHF8+3HSGFOmXiK
NjZlwjqAJVN8OlT//NVrNlY0sUvrM+kxbQ3TnOHOuS1FnOKQqBmourT6NQEBpimF
oD+EfFd5br+6MGSvCjmMFaiEW82jwm4JC6rchFPautlqm8lrFuEIKyxxHWa4X9X0
aOn0uIzyu6Kw2BtUkCei+r+FUnQQaFmWom8DjML2xjZfFatx060DTos/1e8/40SN
d5Hooz5uxUCKlloa8WcHd9wNw8aJ7D+kV2raaTh3eNlAoMRI8k4/hJhj4MusEwe6
Sthh5+jhvAEuAfZpq29vMkb+l4V7hXIp4Bqi+51YCkXV4BCtnecs2b4WOjiHespK
hW2U7wz34Hlwmp0KFWsHMNUZwUH+n3fZkQNUWueGw9m73XKsjCcCuFFdyj5ZCoxG
COX0mOF0tKGUkqrWMlO4AOZyfaUcsRH/DoRlj1CkVoor4Ya4apSbFtj7CkJFJhRs
x0mU9LD0p0VdA4bOq7dbqqBe7fxTmlD0g3LNvkMF+Dr0jZbVMUs0q0xxmwrn7DFC
HbQYY55t5jtBOACbp/Td3HCy4MdxLS11UABlnPnqqbIiIaRrp7NOfvgAeXaAlKIC
ksoUaOHo5lZhf3lqdS48SzcpMLNDXgO6jWufclx1irlDBL0GB9Xx9m4Cqlhbb/nT
y+n0lqQJeDwJIfrkrVmSiT9UvBUNrQiJSRcD4Qbz634weD+MsK5njLl5veWJn9Pf
G06CW0VPjdr6dgteadUuKKLaP3XWFY+sGp+BBOhArhC63qsXnECRBkudXWjp5YuZ
Hu+ho9dgxLJnD0Ac1RAj0JYu1Ul+suCQk24/PGRyBCv9kf7nzIEw+LgTmdlz39qE
8VwBt0rouabbVeBv+AL9q/d3IT6xCOEnClaTonyIhsywBx7GZQmPybrMkCC5s/yC
3bkduS+yXG5P2V8IKFORWYelMudvvtOh8ZYMZxztst7Ex0L85Pk5NFfvauhyKyyB
LhM5fzQXbmP+aQFeAJlim1e0DP36fI0vvJuWHNbUXCOOpYKhBhMbypNceXiu/zHk
Qt0I/G3VelYkp5FtEB/CLkM8Ni1Ia/SO/waJ7q7huYlAWWQPQxRpx5G12w1sbI3v
R7BS/NyveVrWf7I/LAxF0ug5YzEnvx1oYA5lRC5l6RTdHBJPwaYU4w7RcdFkyATr
kpjt0Wfh/rjSJv4c/4pll2H0THYm5L/mSJWWSlUXtEhNH9Fe2R5lvHIK0ySCuA/X
DC7Dij3wfsVMlOe4dfK6RkxPQG4WZCNwBlxYk9FW5+Trx5gus4NS4AtMINRGUiYv
QGkJqFPg0Wyo1s1mDXWQzFVEq8lRU0FLKcfgh7RdBlbldFQntA349fD+qihyKZPn
yH6t26QbKRp1RJ0aqS/PtEYpEgSpOMvEISrdPwMQB2KUgyYAdGPzDxM+/0QVAG2Z
vvOV/2JDj9NI3A8Pgk8SwdjI8lY3zE9dkFO7yhphszvJYDY6VgDj0B9HQNVITmRW
fBOpSkGNOabSxelY7Ws5UAzVatw2EJI33JJeRNKo3aP9jB497eJn+AJpGObmphpT
A/3JySYiB6I7D2IStS07FuSqgnnna1Lm5It8Z4kWEpOYvv+skNpi71JwhIS6M+s5
j4wXhd86IAPkmndAomhUEE2MRczsVtvMIGCHtgHVv1StlbYsHLFeTRb/jnsCn/oI
Fj8np2JfX8Z4T2aPvbPddMpMpOxxWL92h1ZEGhQmQWH3RGGzsjYZdBZLOgijLpZd
VuPhZ2PyXw5w3EdRTawxjzTwtEH0Oi+8ST4IpUXZaKaaAYr+9zfhtq9BH/9GkpNi
O79+zWvLQ1XmvTFWZkFWQW/8Iw1QubqkviTfZyNlMaq1bo/0Ewrksz82YIp1lcI/
qbYZ9IVbmOPM7OlU/P02+mpdRuWGg3ofFuLot+nK2U6EkS2xHWaDRNx168Adlyh/
tTciLsjBMy5fU5OvAltz3izKeuYvk4HmLDPVoUAK7Mb236UG/XYsF0lMqdixSwyj
LM3DLeHTi+5VnwqmgQCxWUWUvzjF3UlT4l3/biKkJDkMEdDOZHLubI/w5J5JycNR
s2vESBCUWgwujuHn39PaXKACzM+/WOHuyfi4MFpsryK7Pn8sekpzBN9NFe1qhGjy
1aM3glHjo2kV+sYtlNBVWys1FzRi3V6Jvye8FxAtzt523Kt5xw/gyyQDcaWkaFE9
nuYXjbyWqVheEHMqDIwfnczFLPGj3I0v3FHEgKElHbHbu13VRVtczocdU25VL2SK
xcbXVxpES/VnuUIgvaP8ag5hkO+xjFDpQZT8OxTBw9LrOmNAYUTxWathkPriN++w
4bQ+HHan8CJ3d1QLvGmoLVEXVj25NXmvVWH8TXnz0Vh0R9ya5y/6okm7oehVTWyI
Xo1BBcJKq5isJa+M+ykLlWr4E9690+4hGixC+wgY6tl39ivrJ3dn8fZHuHNnpkYY
BUu+faQGiPi7rGa/68qYte6Goj7M/GLX1W0uKofgjAypfrtwTNRT10nu4arDyWWA
XXCmnq9LVipuW0SbmU2zt7Xq7Xq/jhHXBrHxaZqGFfaHvDFVR7b7mV9URki+bpAX
B3V3FWKB7uHGgN/bO136LXCOOmJnWU0JxBsdlTKt7XLtvEqAMNyR+LshW5Dgi0gs
u/L7Lkg0NCxx5XJho07jDhp+LdLysjXbaoKNWvUyOpYPYNNNBQMtelusF9cagozk
+BsieOnpulR9mOnjaYTXc9dkyCIQacQZfceLo0GD3DPSn/eSZOXPEO4e14daOBTy
tHUe2F38+7ryb8p+vkoFNe8CR4Hg0qafI40l6ra950Flj6xAL8ufPqxiY1tma0NH
rtoxTsmcP2ANk4akDKrTRaeTJmuveTibsqe7M0Abp/9GkKUAMo2BMX/l0Ab1/wfd
e7Od/4PG1HfGVlcHiXt8zd/ceZntqZngage4a068eBvL9hIqBoQg1ZDpnocI5u0g
9ueaoDl90lDqakSzQLW6U9trcqnU35n8pD45fkvF3parvYuh+Epgzl2wsxYaOc97
wa0LjiStCbxH7txRlKmqc8aYFK4XFJja65a/doSu0UBFZs7d9f0CkhuaLebaYq2M
qFSGIOtbG5FGgit2S/F71UryNftQXrAj6t2xoIvB90Bp5nGKAgjB5uT+/HwOhKeb
36SkNyHL+0etFoM6mrZFJZ4y9vtuVlMdF4aOzS1LnXT2zsO+J5KCNryEm7FVHwGn
Vzm6qOyfpk25gy5ii1Z8rRRwAGDwaYFkZSZdCkPqEMgIAubq3cfjybsOjN1k6HOc
Qipvhw46cGMzVZpDlo8JzZqzbHsbjcqxSyerK9Cx4FJAgrUXzOOLdmEJCg1B4iHn
G1Pn3qtxoG4z4kMb+fwTOknY5dO/waU+OsA48XI1uD2amekvU2bxRj8oBwCBrZHg
D4aGkrbiagFAsMvhUIjTeB5vI+NiAOSimA7QFQwhc2bLsDNOfCdPJprb7d0nKH0C
6TAAM/5YhdlXLAkevcocOvkyzmNJEkYMshEuIS4k/DJthhrQpuP3cQCuooHU4AtS
K3OqsRNO0Sr+lJEkoDjWr3Q/a7erP7vst031TPTBwy4TRLylnHl5i2UJyn/1sCch
APE2HsA+l0UKspiyXGUYLT7+g93CVaK6um60b77MIXsOelSLUAs96R/2NJfJMFgy
4iN9lfGGQUkvUccBgAjpUJxJP6ebSiTIoTEswSJn4keBftAqPayidvP1hAbGEWvL
+6Ry2rG3KUeHPQmTfcQkAXnYYg4Cm+trqQP6nw4EmAvtKnnBNOeALHTgRKj94ka3
L6N/GiZAJUQ50BNEy98dQC2Qs05fjIX+lNgO1ANoMaHK0ALqU6iX29tcwtq04RFl
VWoFqq9imnXy2y1RFM4uiDoqDfV6un7ycPW/wxYQo2lwlneP1HVO+ERwILPMkJDO
yBAgsUVzr23Xik+82H8pFiZZoClRLaYdJeRjcVCVj109NRiIF42JseudNLoM8L9H
WI+tRc19anbbJDB+nQlkIGreSbddCBiMUBvPRl9suTh2xxqbSQsXOFelTvKbkCCb
ybo+WBh2lhyaULUQNxC6Ub/OHoK0PNkhGPaQIDkFEPVPEpT5hXJzE/Jsuuou11GU
rVcSYVtrn28iPw4zEA/ZSMSPh6tHBIDzepOtDFPGmw7yBEt+EbOY90PQz7a0eTmN
W2wVyROghROB5V3bQ3zOVU0ZJSqW/WXvwvTGaxA1xij1vlorCvu7K4sM76h6MvQx
Xns3SRhmh4th4kegmoSTndU/hc21SxuJiZ1pspklUKHDKwk8eOHqrclmcuvVOtL5
ToxMCaP1VIon5Z04hH+FL7EvtwXOvKl340iJ4ZlAG9yCku3CEDzeT+elOIaY6ZJO
5wY4iUqfXr83OcJTPnKJSj6poR4zWZY+jZ7nIjIl4EdehNxvrGxGFUEeucR8XpcT
EiN/GvYOVXR9uDfCiAvtvUVKeWwWPAZDi0ySUL6hcBWfnvaNJ/ht+FjhL8kVxIlP
l21OA4JJXDCn0Q3tkla/EhBJK3UgGhbo4lvHdK58vI3WNOL0bRvFlVOxILuGGFhr
DvTDiJD7m+XyWD38jZyXk2qNhMvCrcusyFzv6xYPQHRw0knMFRliVzx/WiJ0VqSI
a8jQfNFd1Gcg9847zzWBVUgrEET/IGFQa1mVX/2TsroZGXYLNneR6UmtRt8Mq8xp
1ckxhUXgVfXVpGsVbvEbR265Co+e3QOuQzrc4i3LC1KscgUffoLhOuNEmlB4PHgs
ZWLUxiiw6+8A897AptsxrK12/BIYOcIRnGwEceutm9w0w56RpOFZ2+Nn6vKk9S7B
Zd6lC6WpljXE/XPlZHpbBaY7z7UxUDfqNM/8UQ17racmMs5oScdjIrmYIxURJoCG
wQgWLvgYdzJRwYvyypuvYAb/3g3KmWdyNeLoLMG6e3YRilyjRMJLfxyecvd3Wt5J
WHK3lTaarMQqDyYqig2MA08Kofrvs5WVx4pCwJ3Sz+g2WFE9lEoHGVUx2J3L8ZM/
gaCEdjoM/jn8ePbHJvEpLVs2Egx/1lGDwhMzecHVgvCJw4TMz7lpWIdr9gyoKZmv
LmSFeGzUIwB9tsZnfkzml+m1Fp9hs8U8Hda2K71yiTSScCSlGz+Ul5BGmTl3o5ZY
Lvl9F7/BYTDPBC3vX2YzDFzSaVYqW4mCrag2c3UaGYGJfqszKh17b5Enh/wFV8TY
j5849evcskdZi7LDMENoLozcKhEPUBg9ZnpWI7v2x7anKgPbXvwaRKDJn6ADlS/k
Xd3aO6b5mw0iS1G6gr/j0aeoIpnpxAQFhlocBAYmgadf6eFE2HNWmXrTZ9EBCJUL
5UrX6itqaAEOCpSD7q1w+aPx8TFF+7ulJ6p8S+kSl+uTYUt5aR9lDP1xFzj3GdLR
AZ33tRTN0rn8PgSlPjYzHG8t0nsZjdYD8a8mHFzNxbkNpN4EEvH4lqxzRVywtb8i
Lny3Xeu/uJeoPhSOjVNPiozCjViW5O47VsZunxrkniNWZ3CMUc/nwz4R13NSimRg
Te9uGO1cawJbdb26xNQUE1iF4uPIy0fzM51MYUJoz1dXQ1aMaJZNf+1NoQdbxZAV
H24nORpPHdd4jl/485c2dXzEvSgbOXuTed1PewDg6kSsyFMmUGK530PwHQbA3CpY
X4wdNXY10Q1diwHRsBM6IrEgoOWUY3aV2N8VzrVytrq957jahxWT03Mrb+7q/Rm5
Wxw2gch6MUl40ya2c6VAps9Ano8KSihqatlZKmxmeMyZyNwVZKzQXekGiZjtd+YP
apHWFMKhyk0hWk50np+JdzPb6+4bTaBKPczkcI7ptxwPSGzZLlNTRnbWgjyfwhm5
Lu+1qozuNjBHc4ijh7XuNwlw5FGt949EudGZ8q8IIFxxv7gnYPOQTa/FNlmOjdXm
O6175lmvGC1VoalxJ6XZ5Uy05z/wn4rBfCNcoRr4xj06KunRyZ6+hElb1m25LX8O
Gp5wZP66WOrrxYiW0dvI77xY74aQwHxyLRsBQ+F/KhUzpOyvnP3u1jknPi/BD/54
EhRqm67gKFmJ4MBtAJ2TOhkh3K/aROwRNtz2EVIzTH1AgCMzEYMO99tWdU1ICta6
FdpYy0YXpbC2tg3KwKsYKOME4U9w0VNv0WR/gLN3pCBb/fJNmbyAnKdGT7vfWXRM
LE2tXdc2HlvjO/RAfHj8cOh/VqYRuDD0oNDItiVjITCkQq+GLrk3Jo8Zoj6auOso
dNkZlETG4BYqCPsT9IIwpbGHs24NO7V+oJH9OAI66//X+14QMf2du5rtfC/ofKfo
74NS3wloGY/c69XzXcKWmGKKE+NdZfVYQs+/mMO9nfQn9q79qKn941Lel/3Ojn83
9nSc+X3DjneIJb3SQWAtroAg0Q6qcTTT8ySM6Pv/6ScCbfY3ilbNofEVE9/Af3lO
je+LXgIdAl3eE9Xr21fz1pZbv9bsyApmG037Q57RRTFwH3C0iKdAWMoBtCiks7UZ
8kXCtBxIzt8zjF5k7oQIF1Vi7Q8fI0Z2SiuJHVu2KY/j/q1spMV8rDTk0kZ99Swo
u4ir/WDB0VdjapJ7Eoy7iAlzPGq/BoIXugo52xOwVEEyIJo8Nt+JOmANQ2wAQWtC
5qIztPBcXVsRkiTw32g5QXyCXuJU/oZkIYAZ361MyBZeRpg9QmK5i2qpmV3LGCpY
wQGciJ29MIZVi7lo8LM9Akohum8fbsBMvtoyqXCqYvZ88+4VCqYKSUQtiEhFtBKh
DWDK/D/6RYuQj5p6HlN4QuZm//dMqY6tjFbNpLQUlZsF9g0CUU6c3XKoa1l57M4W
C3DmcIyto4U9S2R5dwCeXvgPUlHbH7ua5AAbK0585IAKKBy+1uSpxKNC9/xte9iZ
cXINk6oqRafByPDScngoafJegPtZGOwCnc9ZmF/7IvvOmjMduhHVGC7wqfjnwFNN
wLAqVt28Q2LhpQ2lYkfK7y3QJ/Up0/iz4TfGeIiomZgVEuCZlNydSCTQMinXKpIO
b92+DFm4NFSvcMCoAmoKr5YfcUTmlwzzHKonRxZ3lklqDfi6lLTgVI6JgWYgx1Lo
Uk60/nWUZOqj/UiJFAaGl8uFgZOXsXPg9AJZRCwTT4ygDbfWLg3Y5yQqDPmtQ02x
pYgWpkUxdIgtG9mVSJPYsD1L26NOwNUW+zkwSpgzcAgjLEf/jn83NAyV8xSF2BYp
auXfDdASymOp2pkMpxJapaRgB8uehz1o1Hv2Tck2bu6eyR+7LNLxU4U2/cmL95MJ
h7DvVTqOVi9KEndgYXShrUwVshkGfkNU6bx65YSeqooZmAW3cA2E6hd8FyuRZKne
uxoawkVppqhwG9bdr2Wh6nDSoTMpagK9X+wfh0CKM0H6oaY4T5xdihLzM1J7+7nS
oIA04Cs2XR9A1SPY59AN4bArP6+BdzE7SkmIai48qmi5DsLBxUryNV9VS/hnJl5J
e+D0F0SKPCQoYFCpyDNIqG72vtfJ+djs5hcxL1SjnQVDtWGI3XJakSf+j60uA5vp
qr+Pkn3lx0nUwwxVJEhdfjdewRC5M60VlQ0dGRqArJj/Oo5HODVacTi9sF5dQfOa
lpETvHHMbXa6tRI66u4nDf+mPkV8Dq93+yBpR9V2jzYSYd/b67pzUvrbbWiLQFFp
z6P5ac9hnDOU7ePRTvPP+n68vKvwZC+FPcR1aLJmWw0keMzTcTjzINbbRSF8bPHZ
d6xeaI4iAiPF+u9afdtunAuygKMvMyt942ZH39nisJuJ5Wd/Lub4RsVUJMdZwMal
Z4JR8p+fwXn5DSWCg+MFWONJgmRaK7jOxvQ8LHV5q10GZCtYWAVKamuDyK3qsj8V
NElGH/ISj/XSHGQNzXupC8Vi574GIQKFLIt5JqdsbYDrmY7/99YJquDN0osldCUE
6Uh9JAtFwkzChpqJ0ziX4PdNH3pvDrOeFp8Ce1jjpp9TOcYDTfWTu5u81frcnq2Q
kQ0CGecPsNYFc42pdL6XvrSdjAl+Euos99Ad/FIyzfgNRCuKdVzbiLUyOlIoHmtJ
Q5BFR4NPAyWAurUqvVsIRX6AkL8sYXT9AqtOTwznHw0yZbPvzWFNDWAPgwd7n/w7
V1QlwWNnjZ/hOhu6o9nTQElxDoESjYSFMnDSgUytiEk4tU/3fCG3ZhhOMfB05Zxo
fEIkpbAQetmzmaV46utmvv1cbHkgoBIWf74PM6HQTGd3e/fszhKlyp5LaUflW9G0
Jj/RAuYRzs460A0IXW7jXmbYVT+mD3tBQT9pgSY8C9ugcXYm6B3FAf19ZgKkbYKk
rGqwdm4krZVXLRG6hlNTHih22oB2XaYD4GOnPPYJGUpkYpOPwgu4G0eKauxytE8m
JUZtwy0beyBmodJxdZx4wjqH3o1qIVf6gWTD51aWKbviAmntPhM11mpcozDCtiHt
RjUHssBo4ZiIDlxMnoMkA8hKj/hqrn6AH4lil4eIKGRSlxUX42qEoIzDXwwHUE8o
W2vh665btYPc5mD+nmeAYWnJomnm73p2XlPs15HmERkzfDPAGtggMU54ZURpOMVp
UC5HY7vY1+R8GikNlccqrGPZHYbH2sRe+HSkHFyHlWGR1PPnyOAC32gzNEMv6m8u
1LtsCVb+xm0nlZsqPfWGCIyDg2lh/JBrh0H7vYfPvhRtLalZYUJIl2MqctPkTvqs
Qb9FerSSuEnBOWtY/C+fIesb5Qar0h5bKBUTnR9k3gkxLjA6jqibvVhtGKgSj5T+
OIAcwqT2shedg0C05iFz7H/Qr4vCsXF5rWblbGepEuZBYejpTJkPf+DDOZUC99nP
QZmRlDFfL+o+/2r/mvXhobv/tQhJIFgjl1zUUYcUkx13aXyhctCc5aOTeCvaBoNG
vqdz8ywWPKizt+h9Hq+1fr+j727MeLGKj2fRLRYKja7m6E5ESWJz1XMYr0PnaCsv
XOlAwvaCWvq5svDdQNSX3/DxzDPPqbj1uzShnDI0hfrLkZOEI4Uc3brehG6QLXpt
qLT081yEjOVXNddO6Hs4CNwCWjCPAKZnxkmwyjCLDiHn5VUmR80YsxcOTxK3H/nN
aOhKf80HxkyGisvK7vEXTYV0bAC/CHn96E0F/QUqTZzQOYhmbf+cfppEdrGnG0rK
cwOFZtn49nU1B6v8UgbkZJXYrJ83CM9jnWTFz+i/dvcrOnw7igVtofzDjgR0MhkZ
oPUMMlpbe1SBihnKhP28uOKrT3VhZE/696vjb3NPv3LMdlNvdHJBs5dx1yyAER6f
fvzVZb3F8URMNDZolGD53snpZ23KPSdNgwBChZOMmHlDz2W9h4XtymgLxBCFDJSi
2GYeNIx1tpMIMlK+G7DmdZ1eV8QJcxjzvPi6wdvRt8ACEjpYyvod5W5GIGjOJapd
bD7XGoZsUaVldRtSa8t3s7rxAfzm8ojvX7nFPwOTHJbtrWI0ph5l4HVoKSyx97e3
+XE8gzU4+MJWO6uhxz5qcdbVU1rhzQJgFlAy4yfOuKfp4lB3QolFsaDVWH1wrkRb
xPk3iGdd3GYkqGTubsX3M1plXor/Li85qwefwQhAc02cit04jXsA+YCv6Rq8ttgY
NXt7ohAHlp8WN3/dZ2Y3G0qAJbY1IexGl9MrA/Mfo4gVRl2FBmmvhecQlLqS8zpI
w0wjSJBxmNWUmUmrx6mHNX6/Fk7CH1dW5bcqo6zPobMt7a9p6i8Cuqp15Pm73Cpo
Ub3m6irLSWomEtef6HNMsPNiDv2sv9KlgXt0ruYsGvbh2SWgI0ykyw26p0rNEMlx
9C+9H7MdPQsceqMERJP7088oH9DNUYuA+2WvJQnuSyu3mbzM/o/ob+q9XJvUbfEr
6yIqXaiAd3V7G8SzgR1BvARut4n86MunPOTZHTqecDmgnYaJPEw3e2mmfn1dzZlK
N3+LpwjysXTfxBcmMn5z9dFnG9JmY7KFeEIMbd1PmhjWSZZUKVS8o7UPFc4Z2ZSF
PR92aK8XNNLzBPxOylKrZpWkv4jdPndzKvJO6LxBNqvl2/cfyR/PbiaXFFF3gZWB
a4YChBsiNeARK4VbyvpmZs7h9JV+D1/R2SRbyvSHjILrXVlENFP2y87Z4JwOBCG4
QcP5z7/qCri6MwSgj1Uyf95UadgAmGO2d8VsTv2v+g71GYKw4rBqtv1KprsH6ERi
gDRyrDJ77DRnHmadqml8mfxu8yZOw2cmZmFqD94KkfBVWoqjsY6zup67m7kSwR9l
ZGG1vWw9y1e2C6seU23EQtKXpdmeyyN7IjSGyylsWHOHiFcWYlYET7zuV81KDuNr
fo34ITzFlmiw5x+cXkMEwLYyaQ8FE+Sf/K72q25VX5mpr4ZizWdEmptWFO6J7vmK
PmSMDvkadbapQkbnysYYt+TgfWeHGB3Guk7Ar/QCkUVvJxm2G6yuYSPXhO0gZBp9
Hdl1N94ojKcWEmSs3f8Ta44wEUZITuIUSlGvhOkRhayJaMFaObc4JImtkdKj5R+f
+gPbyXAdGiuojq5PhMVmjuApYKNXfAZhOw1ZRUuviJcOrLYvSf+vC04zUEsozReq
6P35NiePFSRSwSkYwVRKy1WK9FkrCgaR2Sh03FJF7aNr76IbOQsEPavvE+n7wPek
yBG9m2mb+ftrGcll6lESV5kTJObGJTFdEM823OUqSOspgW2k6VQoDIC3nkQ2Ejw0
JRbX1p+mJJt9zRZHmWFiVn/HpAQWf44GbVqkGBgt8T1dcAntqfENB8cQxTEPjDkX
vvYhbVqXgfFvQ3N1QxZP8tFGeUPsyTMGWMUItk+BMO1SAkIAam8FdZkgbLYsBpBV
H9nnx0Ld6shaZF2DPIalMUwrvapZw54aq95ZKMgUJeyzGlOyLyMziMkknAXlKOdW
0sZ5zmWtLLeUUJOk7pMnOswT0xwFu+GEw1VD4RzVv0DEB1sNcJek2Y6h2dT3Mr4C
vJxg7fCSIDkpLFMy+bXXZB1rGs2/haRSehDzmJNjxJr05mEc9Mlyjn0kUVpg7z0M
+o6oaK5Y7jn6gGNHMpK5kVDN75jKHcln4hW9SbyeJOMD/HrMz28cMIudpjj7+QPb
UMQhQjPRprlXmh9yulMifJe23t5Ok/FXMj5oMHvQgSpLYEFMTtIeE6h6MWYOPIqD
WCXXT+3DkU+zHoKnL3yhRrVZLzufRkA+vLVMGHdqaP7X2+g3sqFPToUCSiVWr9Lh
BXr/IgtdRLbSj1ckot1v1wX9tc5NLJzKtRkw7VhDHTz4hUryE17I+3I8+xU6uMZy
tX/A/kmAEDueQXBvlgHfipcFv13O5Sc6cJMyA1mPGXzDVtQpR5vXB4RECDzBzDsP
dqVVf54t9PwzPkeLUnopz2aiRLnOCa1D8uykUS8etuQj80fMHPS/r8Knof6jCyY9
yB4G/dwWRW9FGyrgr9uEvnMF9Vm7iBS/UvHU0MEWDI5JzS6Z+JC0QOR1IxfH4Cp+
I/7KtIEWiKvJENA4TMTgPuxjLUjRlDA6dgA7vRDRybI2/vY5tGiDctWJBmzpUJAZ
7GdBzDEZSOvtHeui+8AjXlczx3nqdOJQEZ6oq7gBIKoptHBQO1uskqFNhjYJanJX
VcahF5w3J1h1aq+9WJ0mP11bVA1uJRh2VRa1mXCRToY/1Rv8Pmt+dMUoT7/OUioR
x/Mr7lsQZN/StS4ZY9uax71jah1/XQXKmktY2Ha0Ltbcf81OGIvq4K22bBDgmiit
RWtr4ZKLCwvYc1Mky81+DOMSvGRhRH0wxUK7t3bWEnIyQIYDlsPTjm7fi6cX+JnQ
+9+0GKQsG5jH5IbDG1hr1p1RMVb8U2jO31IB1UZ86+spI1RbxLUPZ2hbJ1ZYEHOf
PCzzajb1DvPrVl0zMTG2Vm8BkuqxECtPGWX5wvuYFu3z6rFMkD85YlhOg7U5u7DY
t7Tp5txt3Njd0pdv1TZ72jIb3CTq7eXZN0rpOJxa7sDenRRw9VyGTE+qzixc5l47
73yM5mEVVJ0KCWlZCzHj57MTKkE+S+iGUoTEyVlBuNKza94zdA8jL5I+TA82cxTc
Y61PXi6cVXTb5lC7IV1QZqHLst2I7ESOrcUVUefpRlIAtL97ZsokDAv8zs10Bot5
zFUR785GNX7Nv+4rbThnDBYjdKU9hjr3VlMIDnhTFP3OaukL2+Oj0K5MVLRpfUjR
l/zx3W1qhzchUqtBsT4PINyOpWv37X/QmJrU6SIdTr3ZAjtkCkFdlInIywkMSNIj
fsR7IIXmAF2f4zkxOAI8vifkzMBKvv0gVeDxCuGWfU922icUbYGEtyQN0Ady0uxq
wzagVcJ3vGKvrWvcfB72gseXCvGG7f152FO7A+ZAxvxPEHEi/8HM98gUcUgZAfgn
9Bktxivrn3Aw6piXdCFiqKIMF0dcJ5ID4txcYljnZeCe6szz4+X1a1l8KQUFmN0J
n1u+iafBQ8ho2RFPQbxIyp79aA6z7Rgtlt7TK2TSV/b3LjIYabJ6HJ039gSh/UmB
v6KLSdf7cnCEmY9Ab1j2IweTZzvIJimnwzq87nY3aNss4MKjLYIuqD4GVANQqEP3
qtw3a0hGUVh/TB7pfoSwLd3QRuAsq9TfDkL+a22H/ewth4GqrfjTod1qnevOU84Z
jQkEBM2gemKlwAaJX1jFTEij3VXL8OLZAfceAjBY9NT6HxZ2lA7LSekep9sj3zCj
pR8+vRPhHi5kt+qkRebMhDz/ChF8mX0z78HENto21wfzNuQw/pciWUYh1+pLAdI9
1qIFvdeH1+2ssQ/Qr+0DpfrSSmzLgTlHlCsyKBQvVdmRIhJwxZ0RbR+jW/KEXzQA
m9kGFQjO5d/t2bYmn11ZirLsQHF92PAufQHjrH6KnnkYA3GIXTqvgoZGTLMHDzZe
Z1AJ3ye9BEG2UHg9pLQkTrMGCmNGvNugiyAttHC8hW6s5WUsDm1Nono8vrXYik6r
sPxqqJekvWYahll0nJpUTaoZMX0thKSFD2SnWpxOV3iVKkXur6vfGITZV6+nAgSI
jgEBJdJND56r1mZo3hzT96xsNSVHuOHJndRiCzrkc1kXPxREsIqQDYfgMVAd3B64
3DgpVwb6LcPCem9pSTNkhB8lvsUF6Wd2k7m899UwABuMkgd+LFnjI5Su1nRik6WH
NYSr2175W4QF1ikaiilIJt/R5WjXLX6Ww3Fzlkpx2D9vdh8LEnQs8HmLm19iKHOw
EYPZ1+VulLNaRiYrset/bhiRYtrwFS9UnHIHwmQmBew85Hmj7myJd8sXBbIfoGpX
x5YHCZrb5vLTSRdoxObZNjB03Mv5VefurmniWDyRRcCM7Rv4z1pgVzPS53gdRwAi
oS2FxH6owBRaQrncseUg5BeDWlK85R3M6wnXbgWYwjkMpQF0gdCEVmTNU7Vxwmnj
IkCoDXS/HjuLRZhw0BqAmwiXnkvtmzQU4Jx2vZKEyLLuI8zK0a0OThZjpID8T2VP
Pvfq5KeS/6NeheFC6qLr+a6pifnFpGejH6gmIvigWRaAGNKz3BxnJukxbAHJMIsc
gifOhAN3aTQsg1lmivs9aZhJkf3tt+mDhJhr7nO5TtPYNbMnJmPk9AmdHhPbW1fe
QkOxjiYn2Ru0lCr3oHqd7O9lg7nmYkeYf+l8I0EeNhMQoBHpkL0A2dbpRCNLGOsb
5MP/uV4k2pAGX7LLr7sHcbxoWOoBIvJJB+HzZJWnAVO1ph0amHL6P3v4eySDSlj3
fD2qOQz5PWh9/jDWNX9IDM0RwZrlzi6CIKqljVo3YknQ/yUcoUNn400NqjVzkNo0
m1YTAaCXmA5j2diQMHRvTJS94/IVsjt+Zp1+0jSE1tPD4es7hY9OXPIJFJXTTVIJ
5vYQx5VBzX3ql3/AN6EgiVOa6jdKO/RIYNIXehUA6OkCAQVvnwGMmOIWBdTSF4uX
3Gokp058HkpNDQUboSWhHYeF2Q1ob2aQXW8qj+HcurbCCrAcfQZV8MBwJQaXkTQh
zI+eg73npNmOE2LZ1RjZBUjU/MZymwCAa0mUy/O8Tk69Cr78qZ5EGcoyyfoWaMHE
qldCuEzlfv9BPqwBVCPfHNC1pgpJx6HjFjws5/gAkD0zRqQH/BYlP52LQMqXa7w2
PMbvE/dVZsdAtQNrMjn0njJGlKyLZAut970GOPYUipvZkWBXUJ/Xc3NSwe1GU7Bj
fWDEEcpdxyhe3lw5sM6wPww51FnzikWqXoh36kylt+OwI3lglqwsKqbF6pfwwnPS
LBoom1Tb2GZXissOeHMrhgFM+R2CLtZiEXv5Bq3D5lzV/1f+B0flzo5CGNV/aogU
mjYmI4/UNuqSOAKFRfNEGSpbtke42Y0mogfdbxggu8VupNfG7LhsZHA8M8Odt5PD
iP3V37JiHiPkTSkHKPyx2sVqhEGWTtw4IJqh7zDbLJPTHEYuj0ambyf70fnomyR8
e8jZQyTSQKtUmrNGwcDHJijyxGTwLxMTGDtq+dR5zmFqKoWChyefXAfvgDcfM6R7
JkOU37eIFD4uOumOYh9hqnXbedjtgMpNJAOtfZtEp2+R7g42qltLQ2A4DurdJwJW
MmaKEUM4OOeZQiNCCJRp+cDUzLfv1600Guu/CoR4FqcJ8xGLzJpcn8NJTsezBc4A
WWm3JnB+Y1TWBMsxrsm19Jy9JeAD1kn2VLqGhp6t7S1EteTtYiUk8St8rK2a/W7N
oy0b8l/9YK2hA/AU1tNgrqRXhbQ2/h93E9CBFnqLXWs+trh052eFCJernzb2/60p
9U7icQGBtFG7zDKbbkjgz+5nwps6/T0iFg8ri55nkbE=
--pragma protect end_data_block
--pragma protect digest_block
lrsZTuQZLTOGtx/8Cvu9Dpr5TZI=
--pragma protect end_digest_block
--pragma protect end_protected
