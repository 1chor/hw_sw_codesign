-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
JFk9SLXkFxwFKgI5yKC1giR4IW1L+becaajhdOn8DHnOStNa623avxzciUA8Iv/m
UxAq0ijxnAmgzPWDL8VO8ieqDzO0+b+UKPRDNvbyAEKH3ludmippSFU+4rAQZO9C
g1lWxH/cAbvHnYT/hn0HC/ODZ/nv2Kx4l0Cr8rkV4Mg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 88416)
`protect data_block
aChdQp4j78NIOvJB/8fWMfj2xHOSsklN655HwEPPrkZaS+LEnPIkJXUshim0kw+h
bCzb141fLsYe+4Sd4SBCLDQn8tbvTYPTznLO3xjfukWLpDOiQQcNnJaMC1KC90uc
LO4tYTUcOKJD6lvlBGE3pIew89i1XC/gxWyFrfqj8uIO58SLAeJk+zivnL7FdmaM
OR87lTiIkhftOIEO5wDCw4RV1hQ6ao2s1Kx1AHUZ+uwmgQb7StSabzGW/hcRRfDd
Ufu/KYqqtlHugw9ZivDNGQ+w70llAe6k4GpR2qtRucNym7CLqCjpN7S0AH6L5qce
VpKq5EGujRc5sHtad1J4FPp1GL1ussUMylwzOhgzDbHGYlzeYEFw9ACc5p3EP0KT
g1sDZVdIu3q/U4bG3lnLDOW7eWhhIho9zqs6a3OzbDYGYpaOPwAO2QBL0aURkr81
DEk/ENb27JdXYg1HwtVNwdlBcNZ2w/d1hYhUZpcdTfiNUcMopo0RM/T3gOR7v1vE
xiEFQvH7iZ9onmuEvF4YbnszgkpG0vQzFRTOUwVQkcqNoWaup5o8DkkzytqGW+ck
nOJTpn83N0gAp5x+4cjkCnz0L0EZPWNwEBl1pyt5GGrXS7C7uK4Zl8F6Ld1K1TL2
1l9n271WxQOWFT3plumAzTSQUAxaZO11o/VkTU74FmNt+nq6K/k/rVbBQS18wpru
au3F/PydTR4U1DK9ex8f2ESoNO0ze1OWgdu/l5EGPpnBtiJf0CHmSpMlI8E0rdCw
t8n6BD6PhFLyt7PWEabn5PQrVLB93FiwCP6fSqv9vhLxlOle4+yl4m5QhXnWdZx6
mjx1CWQu13OH5NBZz1s/G5xyCfeoMDDLEomx9EWyy3xXWAy4BiI72mKeG60mqPtP
at6UF6WYoSCuNKzOdHmlBfnZN00iDZaWZTWn0GlWG55csnPgNTBeNmKfDkaLCJSW
thkOYuSn+dsmtpW4jPI1YxLFdpU9chywZP05UPSqx5bzF/j5uwKALlqG7y+uzQjd
x/YANUZzyVN4AE4OH4AIt5lvZGGDSCGCSWJeDMMe5tnPXBWYs+mKZmtFEo7AiLd9
BuICoYmgSDUVZZzsRAKDy1YE1qkVxRs5e4hC5rYdmsEfWcPexYShyqQEgpDhrbI6
qD6Jsbbz5nOWknukA+FnaVInj9k7E633F54rrlqSjYsG0h/GSojunNvyw7KX6Zyg
MvX27zoAL0nK6C2zaEtrV88qRYEWoNNBRZxCmR8a6LofacMXTRNn362ipeYvnxlT
DC0AnSqrNeh49/tVEf8Z6sU7EGpvk3MzMHzU4O7mjhrukmQ7HgTW3yvitrstV/f3
dF1vNZv6TktjDGDeviIRHjnYAG3MxcVKNRBqhBIggCEpRF+vvBr/8n5WyPyBGN2D
A+gNb7nfPfzbLwVp/1oU15wGIalMpVaWQiVcjBLhNfh/4jB+nwcbCt24rGrFNwjj
XRoRfu4+A9D1VKrq1s7GYZ6N+s4Egtt1OspPGrj0db/xgRlnIyQz0180aszftTeB
POyTcxQ72/dZDNIwBnAaq0ttvJITi5SxFhH4LmE/x6xUG9R+xibi1VtsltdPe0qQ
bwWnpa3Ql4s4iwoqXVs0wtoymQyUCHen7f4MOGZ1w2ZQEhM0OsK5QTT0VwbWzOGP
UrwvgdebkxYuCa9dr++tvlhGzwAJnrfe4tsipqR3Y+RiuOjG7zX4RD0jfN9CROWr
zfyW1kh0+VqmypM88I7GTKlO4spkDRgKuArdHx9H14UA/Kf73gd/pd8QrBsOXr+i
oMakS5kPmG3txZv2X4Ufk5IDXV2XdKtNJA5t6o8vqqAQD2W7tYeDWEhGXbxFWSvd
wwHUXh61QctZYeYQtuASOu4fcPFo9fqGLSXIhv8zRFKuKYEVn071/FBnkxTSiv5J
0q76RGfZBvy6Uic1nyfdeRXL7T69k0CiuVWamt6pr3M4+Wrok8iRidM6X8jCNsMe
E5FrfbfazhDlkcLqwNurEKJUsncu1OhsQ4iaGWEzgLAe1U6+tJdMLN9QyH1IxB1a
42jszrTKux+dN4fkIcE4psLbdQAyBL/Tt+quJF5TsOM5d96JPa2KiDp75D3lQwd4
vmuRSROFnwsbj3whltnBtkcjs7YZA/MuwtjvAhh1xpkdiholeeigWQQ35qVxV3Ee
JBaZCzX8P4q7KRY/PprbnDEtHdmyNKPuXkRkag5RfmGQxbJ8UVeiJ/LxxdmARCNV
tcFiiu8+Oc0/l9cUPRYOxxbm9eIXMFPYlGu2jHsxnLrbojmebaCr3XtcEtI5F8CB
mpbhiy1HMk0Ar74mrqHE3p9J2nk5BKbWLTCtvAeIHw73qbjTDGY3tRaALVaPk9nl
VUyb43Ehoawh4610RgEkNlBc873cwOUtqZHDxCmvi6vtmoGI9qaVH3JpIRg6Ivnw
kY7UI65HnWsrEi6wJcQZtgp/OGxZW2WdPrwxyEZzV1d/sM1b917FQ0o8/aa5JBDD
M+l3PzPjjFmEhHvbQ41ycCnNjXq0IyU+y/sMfhebg8DBXQV8qLzj/uM4Micq9k1m
jGScT86KYjV2rw5ncKnIo0uLNGuhEZy2HQBlh0/XhYG6nVaTiZJ5fS6OO3JbSXTw
lss8rRPKffe5CHXHKw9WYIyswnUX8I2Hptt0jTcwHporp2n8tI5X/OiyJDldR9co
2Eb8C747L8guWSLzSpOWfi9nMtfvsxLUez0B4hfG5NFnZoGgQei8y/rNnDhR0bzP
pyqwvEe7e8gz4Eiyv8YnaLCmc5pvG32sW2WEhfarzjAVQF0+I5odnUtRIUk2mp/9
nHuR6eyIu6lOVYt0ROmS+kJVuTktARwhVvFsIh+ZJhM7Eo/dVAf6CIGxeYtvQ/ZU
VGnYQRqcfOyOBO39n435Fx0ltB3POL0K5CqBud4mYhSq+A4rnrlSBlY0opbCTulA
xeYEQ9DJP4E0N2BTm96foyxFAqYKnP4ln6f3jzibvuVDBievn+SAnap9KV+nzyQf
ZmEiDgVPzW1SXw4TLFHyikZ2z2hu5bGtyaf+2iOR/s0uWJFNplHWFucDRKBriWNu
XbSpMxq5lQ5eql+/JxGzDFz24mksiQoWz1pZJ2hYsR1iLG501zvB63hGuJUrHAwy
rwTprRXHOrI4hC6LBtUDWGE3lp/jlNs3Z7Nl+kVPIETq5K9THG4f6Ichvtrg205Y
jHF12CyNqz5qn02f/JHH+rkrjHD/h7EDDKFRnjGVZJq8hECNeMwynPbTS71BnOYk
zc8zkyGzExG9TQIxadQ3d5GJYoEGUN/olUQIs+Qq50JX3yV7QuGj2notT9fptdQh
Zl3Yh1ZQLRgfCbddKd8lByLGMVAcSH/SeqgYITJHBa2m5K48dtI8QMR2x6nqZwFH
4WfbvDWQrLdQv9z5dixVlhFXExhm7dBTndV9s0wZMs2mvv8/1QdPPoypZRTTeAQg
pPb7QVUNe3rukFJwtDfNfpNHz89Dl2LgyqHRh+WgJypgHqKMhFqMiBctb+lC0gee
TDkcDJjG2Ru5rZlQ46FM7U2vyhvuAD83/rQ6P2Lx9J6InDyOkx81n8//XIoxsmGj
7wA8gxOd26ugnkghNQJ+qgAszc97fKxV9/mnn3NcivarDu4zYPnsGFblGhkOdN6/
F1SUVmolQkmHZWsrPwtjCei/XjBgrg36WCHCHFlJI96bzctkgopE5ie1hcja44Np
yxYqs/lRf1xuHmlSXqXBewYl7c3tI5DKxgozcW96Sc1HDjPWGintfmi31m9IDKqC
Y6Uaw8rE4FYmd5RIzxsnDEZjH0C3Os0JHyy++cg3WRIz7oY2bF985l8LG0fYyw5F
ccm2IoK861R+5kPYGirDEkO9VRxTrTVUdkgIRNzs8iFR7Dsroa47NiHAQr9nAkxL
4IxGHIJZHIrommCxX3Wko/Mj+oeTGIpzsyYVGVvVGeBjVQoVXM9ZKeAkEc5J4mN5
BdlQJ4o7bq/cl5IBYQ4ZUspeqNOGz0jIOL00uw5rrawuKg7HJky3eCZcYiNHoeJo
bXOQNixwB+FLJ7gv/LTg/ln8aMp5fg5cEH1fUVZrBNh/6nagLcF0UOQIbLPtK/Ft
Q6BTy1BNKvy/UUJg2Acoq33h92v7XVvIUkQsidrJ2ywMvbzctuC5wro1V9gSb8Lq
ZbeD4BBDKlzwYQJ08ESeetovBnKd0qDfgFvZsERcfRdisS1vy6XvPOEZmxAEhCN+
nOT0T9h/O/AIXYEBfMY3lruZa1+LwSRxMqyaKP424AFSmhSbuMXJEWMAgcsYPKW3
qJKYUc2kJr7pIaKQnMPDJuiGBk8o+O1VKPj++cTm/esS9egIU926GWtAw7MvVZH+
Tb7XVf4pDqOoXoaGisiu4fOzOBX/+rCoJTOIdrjq+T3Sc412UIORmHO4WW+YfTNk
c1NKySAijiWDRTnMWVa5IHzeEBEt9hLbfsbFgVQXWSpnlZ0220eumgnxVHU4aoNv
cPRfWuL3u7QQHeqNGxmygFeWFkhzpRdo2338iOonlfoHG06Bqgzar4DM0+YHs3Yz
kMrC/m529EOXtQgpwj17DNqkggS50mqx7+ZS0oVCYx1Q+TM6xLYO2ojGm/jCShGU
0d7wn/FVPBy7+OXFvgoc6tFGOrbOWVxFlZ8mIRVcbh69zDzwT4zUAOBH28hiJnne
yRz02vY7NTDZhg/rNQl8jGhW5taTIxvuK/URdEASBLTrrBo8yOOz38MrHtw2E+dA
zz55AMB4zMvmez74LoAfxuwwigsL3REjn+kjOy5EtQeXYJSjwwQuSeng7LpWHjau
zK+liWJsHTwBDX/5R6u2c3PM5VC13Wyvr0jNZRK9CgvKQ8mL05NWitlDoWEh6mJ+
tcgFPpKb1T+DyIbU0oCCW0KAUFWYpkqCxUKMwVNIqUlV12BX6ew0LfnMgPNGEaN4
2/ac3xZXfY8PyrxwzCHPFTalL16CGPKsmkS7G/XGOvqLeHFMYska2WnQFTMyLa8w
h66oCSqxGOiy9BSnuDq4hKFqFFi9h0cPf5ZVewwBKaOuC35xcMG9+0HpWjHRfigN
6z7l3FF2TNoy6pyLS2z7pqXFL/WEy47txdwHPcRxNVtl1BCXknqlBQg5VLx9xArH
DwjmiaX0qyMSAlxmEPs8zIbHbrzNEemtNrbIMrfU1/ed4w40g14u+87iMVLl5vCt
ThpgDitUGNu/p5zk3Ppzi3z4fzUwnDA9o/DdRBcDkjRA5Qx1/N6f4Ej9pTzmsDDs
vd5ecrwjCZh4iZBY6pbHOldSDNC5gxk0V6X11ZIMZx/By1E481hp/H6ATHfVIzKB
t3zg38JOCM/PlCHdkxgUOhpP8q4e+iw89Zi/bB3kQVl3+QzGeB4UHHPA6wnrbfRo
Cv1SIl51Qd9+/XeiC65t9iAZhMv3oWDFBDLBRo7twVjERbAZPW68nvgdeYUMZBRm
Ew3DhhyNZPDGqqZ8hAY3U8/TX67nGoDwNk/BHiXexsf75I+4WOJZeE3SFs/azdQI
eGZm0H60yQcY05I4NG1UKFNqTZFdtbf6Jaooh16XPXPZDvrj+W3ImQ0bRpoTJ2Iu
5Q6z6crOSQHCygMzc0RfPpGI8HhMQD9i/4+Hc8/agxPh2OHs7LOJZzFyRdxPK5wX
j1WWqzOU+ZDULFnODTyuqcrHwiI1G7GrPsAV2H2Mno2UudxXHOVE+J2IpO7lB/3e
k9ibw/Qb8hjhFkFjwF2tgNrvbpzdL1/xxzYuJALro7/UIByKScXHm8IaPIF7tetY
o6KYC3ALQumF7Q9uJ1XjhHuqsqENNfyuLQbM6OQNkUhyS8KR/s6oQyB0oTDAIkuQ
6diQQjdK1TEYpJzzCS2oJJ9w7KmJOf0PjPeCH0+ZhVXYoRplYHkqwIt/lVtYgruF
keO8btKePyuFRpxJG6c00IHWWP8c3Bt7mENl3uS1+DCKaL4XDrUgOZYkz9+HEqL1
wtkHvyeJ/kekC88F5Ullql5LB6B7BGmtCV8fM3KcozL0qQ6HprnI7nG1iwZw/fBI
RFQfAyeE0Tl6dXrjyjEYPiNugjogtFd0tMxyM+StujLwL6nR9tmPXuVY6DK7Z5/U
Sx8xx7jEKs1younYFYEFrZUGaexow9dGAl2N4sA+dxIP4i1jfBYZu9GnxQQivWpI
+y5YbzhjCuvE5t4g8tvuTKguSm6ay2j16jsiwEla9AC/f9cxPVBdD7yxseYW/IRT
6DnrTwd2BZeuD0uGWV8WcRI3Zi6CrtciHOIZdpR0+9EqOSRA8xQRhsIozGNKwpSM
sy7LInMR0+MsROGRd0T4z2GinEDPAM9yAu10vP5qvjsIPgljvIyU5H6mJsfu9c/0
QO5GlI6g5ZJBHg5la6xr1l9TBrUGM0e0rmMVvF9kOfCOSioPl3/TJSLvY7/GWS4h
SeqGYtV7U5RWUJAzKuBDCeqkZIToRz/Qspem2Ls9WcgoCYQblOCI52+j5xwlDWrB
5puPdFhdwBdLVW7Y5tWSMt2zZd3Zqc7IO6vpNlLks1HofPZ0mW69lMuu0IQNPeqm
XiIz6wLTfUPVD0urE3KA2Ld2CnkTS9zxk5eMUGWHytmUUx3F6SEVKyGcTBh6R3wp
0UMn+gpTyguoypHZQXPgrh/Fl+tBvwmlhzDjgpVVyTm+aTuQKj91pYfsOjltBSli
yPfm9KAMV72McW1XELuBfm2i1esuYMe3LYUP9MyrXfMhoFATyXcc1WO+dtqyguyr
jBiz3zJCwA02hJHom3DhY5g5q86kLU42NyO7w8H0QaEyI/puA0HbtaypJqfqzlXV
g7B0N+tsk8vtJt94wfWR2aPrhBQspR68Rp2pBIu2BTZY2st049eDtH/k99hBFZQi
C19UYYLk0WMYY+WQ5iP/s+HqxyGuo6/0PYSpVw66xMN9sBtkHmUUGlH4p9yBY56p
AGPSJbBSR2xALhH/zyEPHVT+Spym6ctThS95CUIDi/fcGbK6Gn5+0VtYrJlou3i4
ZdjpRr/5R7aoRYbHmqQNNZDTaEcRhaoOqWKiT0aHm5IzLLdAZL7cPbiwQklIpjhy
0XskI/a0gkucp9+Din7DVtSDw1zMnPw+dJMn71AINbV6q7FELmKiyPqGpQtyZAxc
yodNx6fP+ciHBPxXGivn/X6cHbsiFJQgcLv7NduxTfNnyI1hUuzcoNgDBGDvJYpj
0Zu5YIt5V3pxek0MK2mskuMYIKEl2ID6qK7amnLtjrN5EHAkff1fC8DQjK9nH+lM
DTvR4zYhdrJakPMswJBsFcthJ/Q4aY+TgmFUsULUY0NXOu9KhG/BDVAkG1Vk7yr7
HAd9jkc/MKuI3niiWJ9lhbix2Qxyc476Z3KrVJVrqUOyIeVgN8RzWPLEd6MTfoQT
7jcx4+Co4y21SBRNUBBc2GrSbPvIVyxTkYTNih2VVy+5rnfSbhDKpx4bOqCBBeSC
KQRuMFIm9IOLi0EJBMfHIV2VLs+4GgazHWnMW68mS0v2JHg+2crTfB7H9SS1NQKy
Cpitq/MedeVrfgwUxUVlZPDSn5jDE1/Tf9ZzQExVktNNN7BEQ3d5fRSRhwcj7720
a8YTvCTIAokTzHbVBLQbzI8Af7kY9dy3zLcwOFksebZ9u0yapcl4XFs9b7UACi2e
VTTTqMyMRFdci3tkO7l5o2dPcnCrK3lcUzXnWi0aU42+/Ntuc/6iSc8WxUxt0ShS
ycI6PbCmNECv2vJqM9xmwcpTub+rzdQZ9BZ1KlMy7bKQEO7pG5D7BTT3xsgspcZW
UJViI4rqfCBoCPhwyWKSzJOc1dKX8CMIDm3mAUEOi7PkWXwsr+QkeNaQlyxsdRN9
WXH4ib7UqrakQljMuHqy5PsIyuB1SWFiGzO829XXEXXIp9ogKdNYvaFX19tCNYkO
2VuCIUcoTPO+OZsIImSlmjYI6TkQdIHyCTRjN4b/pPI9ONfguUXRQggiKY2OYnfN
bZ1nWh7ddAKqlb6it0IkRz4AQc2cMcjQe8D72SU8BJ4EPlxsyUDmUESoLHj3pzGB
anMf5Je/tkZYgXNhcOr8TJOKIzlY93Ksg/dkC9yUcJwgzwGjBkBW4OSoyHEnBO/Y
jMXclDojLzK3qdih6VgnBMfkZaI/WMvZFP1zBzwWhZ8b5LTUVsYuWIrPHWX7zrv2
jbseEw/bswXfpR7h8ouVIBppQP+klkANR0CJI8RIC8bsdtv5uIVlKKO9EsfznmkZ
NSz+kXclWkCQ3VxBPhLOTaEWPiVjgptdyAdF/PzvnnyYhkJXwnQzI3JybMFun0k8
NvViXlYBtPccoLTit91MiPnQRvDn7p0RscAWE01fNINst3v7wQ+TN4ksQzkp+xGr
TM/4L7AR6+cMmao0dOFPwrbUZTes34brBHLWp73oYZfd4Lp5p79crIKGw1VZ+mv9
Uw0K21niXyeoyWU1OzhjqzuXpzuYTbozuo6lzdqIiGiXjYk6YDd71rOLfM9XGTb1
nxqHfp7vcJe1otjslQltQs/biDEap+NoR7cLOSyup3Lh6kny0Be/tJtO5acacNvZ
uYpLi/6CK4Q/SuTNiHGyJ25AmmPjwqzU5j079MAyR/rtyqphoigWjujgt6NaDzbl
mszMyUMdEqcL2mtgcvD4/DMd5ZOvkDicTmCxGaphiJuoAzlbGzUDwCrxRmHzMugs
LWy235GUYVeY/5H071bWGa/dt96f3enyO6KHX+yqZF8mHNNEtkIwpuz/+fJhIL1o
Y79Yy5Iu/r3fnMh8nwe71NOB1TLg/AE8rartl/vgj46FeZnBEGzY8Z51ESviA4r1
aHasJvUQjlmRonhG5cTIVb6j4KDpLaqnZhyrT+jynmw+/16sJKNG/gL/+aHB9xf5
hY9u8/CyooTghnnKkmwufZbW6VOUnYM7cE9wfd7cjwzze3+Yu7X/bS9ymVIjpuE0
5GxeNTmcofkpEgdYmUdd9j1hZnkfILBK+ns2lTq+BGQDnnC8iVYXQ2GRSI6KgoDe
DoFIusD0S/gV9zSAgAOk+f5VC3S7C1aYVUaq+Y+Hu/o7atxKT8a9jpq1Ax8zD+2O
JGPtuq5WbRIoSxX7/ybFlzA56qTDPnVeRu+zEITTxzrbvyF6iC+vXVuOFtj1cazv
GfD0yF2gW/T9IvLgLHDdBlHirtEwjNzvOok2f1TMyfF3n1JP0Q40ozsgCXtCQYRP
4GFXGpr7FiRE77dTiwA/izHvaaWXm4M28RnSLWKhhdIrBnJOU3bj/dQNSXXNEGz7
frb5ULFqgZH3gkRQELQodROSiRCuV0HptScu3vskajWfv1YkqUuWzvfOk40s9pku
2EdcsZmGcOX4fDUx0LU9ucIBaP5C+QDQOldlPtlW68vFpWyqxZRkrpHuOFLxEDNO
TJHSnFjELzHs3taO4i6tMeZVs/zvAkvtYfD4Foy9EMcFd23EIgrUe9nzgij5IJv3
Aibd6VzjM3pMU/Xz/6QSt0Rd86RRvbhUDUmVRVSkuVHu3OPkpZcmwtEfuzNiDV1S
+wgn5UoThB7mdPx9/18SAz+AIDQSO/QmkQdrsS9o2bbszbQ+z143PKIV1w3VdVRM
annZeCUAnU3RKvwDDCS1WFyq3JMk4gROlwv+BLDhjM2LNnCFde4C4YOXYpXAmEl6
dWM/tm+ri48Q4CGw01+Se7N4QCo0l/7JMX2KQjJPLh21THgAU6g56IrJbrj5z8Ku
aiBbKimhoL2OapB93FIM28ZWwBaZCZfIKNlVsCAt31/qK8UIbQVWjVJm2RDuowde
p0uG58ec++akc7FqbzH/r4ShjEU9trcLnA+MWHC0btMR2vi1SZREEPYYXFG4NBde
H8OFpfFHmz080a2eHA3j/F2NCPDIzPIxFi3y42M0mTc+o6ZhuGlD+2aNFw/xSWah
4q0go55mHCYT+Ci1UuisUZJyH3I4uuN6u0PhVh0XUuAKrMVW5qQuOi2YFZfn8z+O
NLY3i6d5FnWLeOgT/R72ChZxmt1omIRnJLHRVkZCN61MOFKQBPCr/5ptpqcBqjEG
gmhNb5qw45vxafkN+QCDRoum4oJ4AiJ4R8ppcePnQUVd9ttZbKfv5l/Zo6OJLZ5g
cvleRr/8Guqv10GNCJBlouy1djM1QDY6IV1JSEYmo/5oRB0Wxgc6QlfWNKXmMM/Q
9Nwf62f8e4V6t/NGHoKYvTBe6yOk/oSTN9oWcn9KnsauiJ1eFP+AAUhPy8kuBNaB
JGcwcQAX9ruaA7Vz7HPQUT1ejYD0yu7ocCjMNJTxeJkcw/kfmuzx/YyzQ5t7kaBV
eJMSkK35XhWOJacQDRs5/IMY6C8Cf+d08FMkoQ8x+JtMSj6OcvtHXkziQe9XCCjo
l4p5FprQxXisIItW/vlEwFyouenEkB8aMPJeCGFzqpTQWEMBpNYEPUS6qixhnaCO
HF1zChRWonQFw0pPZpUVzRkBMWOgz+l4KDAlxm3PwsKLwQK1A/PqDksaNu5HMm8c
FRcOzgxK75RS1JJM2qZRig7AzJ27TbxGEyWCA/9IqFZwWNLAEwfrgG2SqQf/+r1l
pAGs2xYdeMVbmI+jgqkJnZe9JFyZpQnSg70xHq14xeEMvP1UZK4oH9SClLM+7T3M
XLL6xgUHiqBFyg51gDMT0tjkWmZW+ufPEUsDWBw9LrWu63m6SI9f9wWhNKJ0F4/j
dRu5YamTTVy71E7kXgrL+fIj9THfL5FgKrVQwP4IElawW6P3ja2qC/8Wi4i1KZAF
kHK2qyNgC7UKA/SBa/6A2Cm/z8ADbWOIy8Q4MxVHvLi6zPVmMYjBtcsSSgywkcm2
SaX+DbPFp6Zxw1pxLTtrxZVOzgG3Wxnrhfn4vycYGeqaRv28h/h3NffT+CdztgRM
5hJJRQY9hucwVOrwqscwb5w+6gJ7cf+4HkSwjgShqTfj/n3613vX3Vq3+/6OIe0c
k8lgSqyNz+CsYMzH/foM9aXHl0jbwdU0Kv9Dhu3evsGOpCormxMETMqL3QQXhrCg
hVGLMxtrPRiTYH1Vi51PYPQB9mf5XwXRuc80alGqc8uexwDWJvnh2IFHxsN5kxT9
I+RCSSs8UA+o4Ft+id0aMi1j2axd8Q4uvD6rQErRxtwjHMlFE4PuXILJUvkE5s9W
NEVeNUWa8q0hvHsZBmkl5GW9FNogdH1ZHd3+E0hA1CqOUopARXTWLJzlb6bjYriJ
Urq2dqTi2VB5A3g6DqrsfFrkmC6eyKW2+w/v2Om5IFKW1LTQxqymV8oJunHAjxaI
n6q4GCGhzNAzRbyFhhpovfisYctHDOx9bNbvHPsQovHw1Tbm2VE6sv540zZee6YQ
Zi5m9AFaQymaY5i/cQ1OJLbxU8UFNRIotVWRw5t7tJCOn5VlektTe5c5HOM/7qpY
iuzlO9gNW0+1QBkJ+d4MDgclDGwI2o0AM8YTERzxMnsqM6biX9dBjTtdAsuQj/5S
slJiARZ+dvNioXsX1XSoG+ze21TUJfdZNI/wJOiRnQE9+QHtsJODuqYKjlAK/GuH
OdK+zZ+lZKc6C29iTZ/TqLxeaugCwV806clOdco9Bxjf5z2LM9PT2Jo+Kcg/Isii
elCSEh62wbooSAjC8OX1/cabuG6li0aneC7sJcC5yYHm8jXE8zIzIPYSfyPnBq7T
q3wMIyOdQky+lMZryuULFU+NXzG5111WSeTXaPIPLitiyUGWPIxqLNtZbCdc5ovL
5dJmp1/8USDhokoeWzBx035Y4zKsoTIwDQFOUsQmplgIyzjh5KWYWdK89DLW3H7Q
MbiJcfAfRczbkU/ola3tB7AJldQ6uO0G3GzOOYO2fiOkr02tnyobqFsd76VMNt2F
pKUvv4XcrkQ9Mg5xUsp444Zn/CTDRxutaap4o3xw3v0zeCPfbVEX85SD7IPebJNu
wXFE20yvII4sfMy38pkzc+XmO426IPr1BSoPx8IitGXKpZwh+8m1kreh10eEXuyW
oVRRWyH96jdknJSN1KINDJ8P81wkFinEoeHVCwiXj14u2xRZhKw5gyz24v6Gz7jL
cITbN3SYZqhhldrkvlL76nRCwqUzerUaCseiM/R/II01ZVEp2jhnxPAyzYzZJidS
ma+O+8yBxoKdJp/WxBiSkrpePrDKKIL5naOTzmh2UI2kCo7nJq+IACYieJFCnAem
+crCz620cY6m6tMO93RqHoJC+YD873zddrLM6AwFTEsSLG2kzxpN2OlLI1GesLel
geUG1T75O/qJtHwNaDVJat7DcpzDwha1as87VZ77rI/MjNib0XXmqicOZYZVSczM
8Ty6fpvHT+ePR/HILnQA18QvaZmvfVnLkL88+bFMarDV8vKoUfxnn6ldG+FBaei4
Ugyrk27wKCCOXmpyvcJP20zMyrnuOBDfSAazM2Qob3TXunEH5SOKZnt9E9YmF9ks
S8QA6CXHMFftLs8E1IWAd/uBFHd8O7dtUgIF6Q+sCWEKmZcPUeAMsCpCRR1VY7Rj
mUvrl+ksGc9Ma4jJdoxe7CiKqP9tEOkKx4Eq7BTFuD/FheCJv51nomQNRwLpuO4l
Jn0QleQjAl5oOiCfj103GMHNXD1+9o5oEFzBNW01XAbAzHktZYLeDlFDE8r4hnXO
DZwEoPDK7oxCRPAjukmAHkAKqFTjQ2tQX8krM1PtsHi1n/QQUEiQoFnSJTewMdqo
lkr8VbDU7TKBwlaQ7Fg7kfwOZnPmvNvL1CxStKotLogzi6NormHcgV2di9jsap2H
whPHbuImWw6Ft8arg847PrLV2/6DqAyNTRy+tMNhOkCudBH+13s0Rq6hnDGd9xvO
JujcePmWxLetiPQDhYMCRPFwO7w/BwjqPk+Z0fauheqiDD2u/bTs+H4pWWJL1qxr
1SqfI0/X81z+gag5lfFps7uBRZEjVNyVrP7r5Vhn+l6PWBWcWAnn20XPoS8kJ5Go
coBEMGjtqGYS+tZvxGz8wt53SPdG9stGpqkEOkoDt3qgXNvSq5u1II6Vrne2TC6R
Ji4+3slKu8kH2gWibSLMeSI2fLkG5Kh6lwvg4NUr3xJqWf4NlUKe3BVOsU2nqaJK
yyADLIY1rqyyFgzh0zgGz56wnfEPNOSFUufSpvfs4txe3gQhttKZBDdggC4ftx3t
YgDaUcFPvGeRdfTO9S4b3Lq8p7Jnzuxwu/oOx9me5d0l2jnE6fo6+NQgj10hRdV4
KjzUP7DsSVi8MI4HTtLvOka0PQId+KklDPW+ktnpoefNBfsJoSW+KPUEMc6ri2BS
6RrQcTbW84RxWFzOpJajW6zuXTineCxjvrFjqLc02vvJ3uWI9MV9wSKD5V/+qcpO
uDJ67sYSQgjbxn6DtUBIBqBmmVcV/6Isibt9K8HCZHXTp5fUZqawJGsKuDJQ5tTv
Pz9DFoY6u/c8N/uhyijR707RZAWeU+uNGfeTYSLCuPNrDw0V+NUoBamylGKdCtKU
f7sjH6JQcfuv2QKPrZJ9M1LK0RLULZIYa9eESPieGlqJg3VIhtCpNryON5Hy3orP
ON7vR8Wm9Q09ZxgQW3F1DXhxTkuGuR5iZBNtI1nukHxFl3HIDVEFxjIOs3xWip/f
9qPGXwUyNvsuiKYMU8SmGF3lZG6YFS1iIk2DOTsIDA71WjTGG5EWfyyBAc25nKn0
hEUkyIuRjK0HZanuc3XBjXgNoBhrUo0lGW2t9WGdAtNJisleijQuve2MeyfXCrY8
dfrpsuOKO38W/rpYpQqsXN+FbNaqNdg1hLOhqbZicqaLMjvKRczc/5oL+Be9yQRF
+MP5EAmLYAv9G/4EAx3cGQmFAYZaChKGpctGjUvtHtA2WvLGa+N+BMiUM8r689Sx
tmfsYh00egmNK6tmn8aUAAv5jYlEU5Od4IJVQdmJC9sKOLzIVzj6l+dokzgDthDa
wIxGG/muGK++NdOOXxgaPZH/DWCCnN7GTl7Z/h7aOxhG5y7YwHuX2E+7tVJPqrtP
PP4Q0HnG6FYzrCVEtgAKamzwcFiuTwuOf/vfMw+VDzSDwuqwJ1lpjFEh0QhBWLXM
2FTFnUfp1/wf5Kaqs0TUjFi1h1jnF2nBPO+nED1foUoNnthusiJ9cPu6kf1fNGzd
LgbT6Ee2atyOHNg5KSdzrTyy3S5J1GQ8QUpCZ+6eKcNpYlJp34Cn2u7o+wI2YDbT
KsnT+lK6Z8W0pZblMn8Beh9/dJxsy73+h0wYae9F906Rva5N/Jy3LFUyHZfvVkRq
0Ebt9XWDbMtBFHAXp2mmGDlyT3f7SUX499fHSC/fjHakpyxf24AsJruc+Hka+PiY
MjUlc5hs0sHm3PJSeVEmLnBt0cPHaI1coqUqsAi0GpXhhT1tv96rzF1cofdKNTWV
uuCzyPhwO3OYqzsG592SPDFjFCEUsTA3PVLmeAf7Flov+HpuvhS/gBE6rWsd4/1Q
reRefeRQ0e6t01NnN4ErHHAauKqwKnAYkICNFkFH33t8qYzSp647fnLH7NC7+pqP
cSZBe036M1NE1oC/+Q+Qd9BFD1mI2Zr7m8M+9IVnyGcy8h+QTVoMKDUJcMNrjtx1
u1kTE9VcpBhY633/iS8jwUEoqLJGzk/UO1/LsfJCQusfzxgqHMNRmuNZtr4ENWUn
CWFxEbLnphlxdK6cOLH64AK+NxYmAkAU33plTAvsj+WKtRJnrGXqEjAA5Iiln5Mx
VPDxL22XwFfNg+Opn88iEwl2StWTZyBKLwRtv8TAJISpA6pZCN61PVxo/0jYwohu
YHbe6jaY+Gqu6coupWrzaiv7BaX/NR4UILSmwA3Iv6eMthgbW1s3GG0BoTxP3TWB
Tej08WZqxu/YZU8AkctQIniJ1UtLYz/B0+mKr7AzKUC8QbcQb1q00cu3xuaGBwV9
F3T1UetBtB9V16uTLkuMFqP23fH8UW4qFBL73NyoMIXjuWDTM8d48Dikwu62r/Ue
yVTDoZB3KXxMmN5AhN1zIxs8gpahmC4ZIggx6ofTZWTTkYF5MgOVQj996wSv/en8
MwI6KY2LZoJhUnUjffEw7kpRu4Fkyqf9mUlyYfCqbJJdYryf+Z6ljBnD4zGl5hqh
2xq/lshIK8WSm2spUyiRJwxq2JxDXgb5wybQpXZ9aRBTtsxuzM1vE1OyZaSMYqg5
kkR11ilw0d7XgQMzg0hjSFh6eMxcRs7aNCcCo6/wtE87KZAS/h0JNmSiJ7yrJA/l
xQzYd8IG7UJDvLB1NXboLxl1FwnmOGwGpCM38OTFMAqudAgkZdzLmVBd8Efy/Rub
o8SOhBQPiS44kPGCCACmfPKsiloq8WgRyhMR9oE2zZ9ntjtjymrmm9a8/W09ZOoM
YtSaxYVgOxa1l2NB6RKLQbyyWxhNQug5fkdUfiwV0O6lJzXsJJXGZzebapYtOvzP
Ch+KYoTgEQnX8ET6D2kWxX5sPBoABgiiu8sHPB4VlRY8B+JTEdWJCsscyhEHkZEv
Glz4ojP0Ia9hiAalGkCZttHKnf1mZanUUXZxLTAS1vR4BS2JSEDnOeIFz4OBt95n
EfD3fkllDFxXIVqoMxCpaXAqY01z1uMWrEjcJUVWbsDl24cSljQbPdQQOrhjbWoL
GxEs+xbEQj+aiCU/CMMeYKEw97DmfqHa6c4nLgu9fB7Jow339RftYYcbuQe4rfm7
Y8ESr9AZ/S0gtRPqRrC/EZBpE3VN3uZJ3uAX7Tq7bXQ5jL1NXSapMdYmmGlhRB8n
qAu8zxpQ7K70uEQpiqIdjgfjckLZeParUTB4Tg8uHDZlIazGSPfyJastSn7/RGch
oTBu99MlI9NYODFbVQNbBi4i7a1zaJR1FEw/4lU3up9cEqXwI9VTQY1ZtkVf0lEH
9jjjBU5aFtaEbgwpsuGB5iefM7Q24mQEYDbveLPXLWjSQai9JrE9IUQWpuiD7Zao
RfVoG+LZD4foCGK0nbSEWVnhlM59w/skNOaG1M9TxJunict1OCzH4p18lUE6iopI
aDKKtj+ei3q6hIqavj5/WFjIRXDvVac/ts2exM6u+eOZoswebgSDMOwZpxGqfuNo
oGluWD1SQm4VME4duyA/sU8g14jMKGaeMJtyHLD7/5IKE5Q1PDSbrNGCjENOq7iW
/WPpO8Wrj3FR7INQvLK7ngmM44cvvNE0FOGzMa6Z622JAw0qWYnxMAZPQ0mU/OVR
dOprHwJvhEwRmQ+UBQiAmDmot1g3dun/GpMs9Wh6DfDdQzSoJFuUIKxcPfgD4uAb
tWB6EZtgW/EuxOCEf4DQLLEFzoI38/GfehJWhADmkos/TTgfcGrizc9aSyijX+M1
jbRFFQTN8DK+8YP8XqEDeEUj7HCcyNxNJ3nMf6BKV6FRP7CYJsC6iBeNFOHS5Pzm
vtN+OL8SghOIWjeG+Pnu046cl0CvM4qzbPxz4Cc6kJZNXGsZnLwy+TFgXr3ZP9n4
voDkuC+fTqoO2STyCJXMU6SY70Xn4QBSJovXA+CrSgvPs/wPnP6uKFYOjldXpBzA
LTTmSpUdXWmAr48RwWiP2GzsJziE3738bEfMO1/q/j1f2i9tZ3obeIE/nxkk3YTP
zuwOyiPP5sOsDDTthFbF5mepEaHAlO5a8/F6xtyXI8seC+7C7kpv37o/gsbcdGtX
S2lag4gLQRRMRakiofW+MsGYo2kNgx3GBm3xYqvC/RDxkG+vtGUZeYGLNcV+w1GI
gm6DA1vx0jZsZ9WR3FXCCuOcULuCymWM0+XtRIdvXOMYBXma1xnpz81eZoec8i+L
swRxCe9HVtPoGOBhRw4LppdH3pdEVedYWpfUg3pS6xadD8OND8WsfMcNi5V6xIkg
WLvA0X8t27fBLDBztvRYZZuo2udDXoC3s33YLkTANANJ1TWKVh2ldRMw1wcMWJUe
6BfKmCnKEmgxitB8rjtNl9z6p08it9SV/1meKD2OdzoJk5UtmNuCQXDHKpx31tsq
D4N7ySveWNzShaux9DwcnlQi8LGNoNhV5honh8TMKDjt+x23JFc6vdMOK5MKwQ6Z
Wnt8rB5hCuYTek82t7sHGfKjot+OEQEfxTkMWnNkkopIOHyAaAks4z7RiMIYdStz
DGNL55dPJCFq+nkqMGsMdBrhK2X9ymhHbzi+yQ0DpkK7nJRi+S/kbNZ/XNMgpGeq
qrb3Bj+jvLK1FaltMJcSlXHCF1aO1DwBNJi1vc7CReyBHnVDX+FyqIBGR5/GmtBq
0cY/oO21P/5nYt8cRJWhYThXbdKVlhY/75DIXFJOFef3TrKfisIdu9pvC33vpE7u
I//ZH4y21mngTn5EcON7CfKaLsjhaiF6ekYuROQqiMTqM3tLpz8GIPGY8iXiFAB7
PzEaanlxlDgG41VSUkr+q3XqAjTJoP2N7q9yJo242ZrHUq74gK0wzzQvLwgTMY1A
xXH/4dMQxvLcNUw9LXAMNhgvWZLYZhqEyAQ2FYfXkqhhBo0E36QYqQoTvbo9V5WJ
y1cgo0AwENCERXxb7icxSPH4+agY4tyEsVm4z/F9buYHzC2LNE9fcY7tn+RNJj5g
y4gnG5+7EEuK9zWObknTsiKBVuIhovZwLdhhtTTwLzrCLc/5pZ162jjqPBjEH4DL
H2sA0EjaLNbyQC419uLas4WggjruN+uF/dyH566ZKEUQmMRofkSQeiZleKVaFXfu
yw0Hknpjplcdc4gfxz0TaRky7MgApvnXZIQJ0ioNi6ZIp+caJ/J8tIfSjVMmg6hY
Bs9EHNOSHSNmxudMLXvDtGq87sL/x7dgOWUxd8+VFaVnXj0XvyjZ8aUPXEoJPUMD
LX1a9ougTOuN/meH99liJvMdj9/TgAJiBoRqrah75eEojTzZJsDMUHnTD+uFxhhR
rRbJ+woY5OyYQXhppI+AkMYb4+JHUQ+zob5Bg6UcLzXtDrzNDAtcCCw3ALv7W0Yj
nEqIv28hprm+q7z2MjWoxLMPtEDbbkWwpLP2AsrpgMirApdzG6Auu2Od5FSjRwjW
PzL3Pd6JkYxRUDMQU8Yyktn2GVigmt5xHsfJk/T6hgeIHHQw2MqoNqWO4h39qnBF
i2gUqVGFZi0eyywPwAOLRiDWxg+IPdq6ocPSwVcc1jny93YciCstMBSDWNVhe57u
Px2Pn4RF/vekgB6PHEElxgyZPW+lLkbK7Mq8OXlBJbStFF0E0hUUw7y7uI1XEHeW
BBGZoythoJBjYQorJJN8ZKg/ZleYMVo78NPTH6SE0on+SajEe6OFLx84rATng81H
GJ7pVfYfixg2IN6NI+FYUOW4Bw/QWUDVFsLxgk+/AuKXZMcu81XuNSeahuy0+9Yg
0W2WXCETZs/5G0pnUde5MqFudlwl/G2CB/zwAdUP8/vHfEYhqK+kowE12XpmJ4cm
1qpbrsKQQmQ6Y2ogbqLoyFOR+7XsL/bWbdpVA8uKZGPSJE2LDDu55Q0JJCqnYblV
ybQGh4w33iigh1NhkGI/J4VHeXjZp4p0xeDny/NJ6JiDsT8GW7AFqIADpcgBMy0F
pbxei1vX7R6IOo52eBjavklVJWvInV7k3tAobEIyFiziQB07CYmKQk5gMIONi7iQ
VkQCQzREtr5d6Aq3C3ZkuunEWfeU2+ap/HDQ7tbR3CKBb42PYLpXOpZm67s1EbRG
EekcXVJwOdIGLHE0NT5IiolPRVs9ZgwsQmRuuemKbLrEhJcbNk3m8h5ufi09zE2e
Z0VEexrS2aqeB5HaClNFIcCz1RMxyQvMXCU44QtxE0x5BRI9/brzz9qatYoxTSck
B8p8zd5hLXHL1zjPrKn3mWRtlIb2tEtBKWo+tzkeruVaeXqZ/NGFxBKtDntzAEHy
ebaa3qz8QNLvaas/SU1j3P3RGuZ5gsRmZt1GuyFRm+p/oD63dSHbzFRdHdh8uEUe
L7Qwj67R5kf/KaJHMQIou5Rs1G3WmZKQ+B4CQ/h/X6lGfPL2I9MO2hOlevTy8e3F
tH2vRgqFzHCp1UeGRXhJgVeIjKC+QYWBPCfGauhOLfxB4vVszAhJSLPY91GPqklk
qcGyK8rYyzwqvvUpYgakHCIgpCQNPFt33THtlEWGM36fWQTHRwD/sH4OFs4N2WOA
3O3TW/8xtMnuxyc5OmTB/mP1GRzupZGMKLXiAGun+ZEI2RYMUFk6fsaXLM4e70aO
8b5vRhsT2c5q5f53xfxsQUbGa8hmornhmD8xDC+9MGnmocHh1MuYl14YCgAuuPwX
cMzPFcmRNYn48zYmV0PipwaxY5PsZ6z2hMVYDhF4SVJ6uVtnbkc2m2OeMqZ5Pg92
GTkFcJaEF9pFqT10rUeHfDkXM6YtwMEKdYi1pfU/FtzzrC6D7NOOxwZKQds9C45s
CtRaNYXFGfmTkFsITPZHbfcWSdn1OABkG+BmvBa7h6IYSJas/On4JyGvTOrVyeTS
6dhKOwScy8Wl5RBHs0erzu8gB+EMur8UN8ZS1Vw5huyf1vOvxLQbs1JR+egUJ5nw
+tfm++011WwS5sg85w2S+Og4dDuunzuZ/Af3dFnU7LEGtwJzR9bQ5PtEdNG17a7y
YuU5zp0/1FDVoHd7xhRCPhDs+Zl7juojptHWMjma40HRK3abELufo4qHWhWQnshY
82hayiAxIbZ6TqOG0Ins/eU70merugJjC4pJgrQfszoQh3S02BVE+NDEShup/hGG
sZW0HNPlft2HFkosNp4urc7aUJPm4+RplwVVnVdxrVGMtttcaTUscWGGdXb/wC2M
nM/ouG2XZUi+I6Eb8mArpbQtce7CtRxg5KTnrlaIqREJ/YjOJMKT3pdYjxmuf7Th
q0v9HfDQQe41TXWBDxRrBn/sOxeeVlDsa+d6DWGEsBcLFFXJ+8HSl1kcxiCrGrlP
WTN2kxL6B0muVYRfNCpD71GVCUXCf270225QjIX8fnolx9j95KGYEkKNCtJCKqkV
pBzaId7ftSW0XFmHUUaITOiqSy5aCqzEljZdfHV/+TvcMJkcs+hYsRDivUNUi9tB
hlTEJU+43HyRfFNGMtRCSlqU28qtdoCfAK+Zt/ZyVYWSe5HCmA6ouHDI2wJ8EjCf
FDFiEmiyGybFyXNwPRykq6S1H+EaHgQITS2YpK6xNiWLyy/fdnvaekEgi11Gwgvw
x9H2SZtYcAFspN9WEsGk6zdM/HkhHleHVOKCIZq3c3cVxJs4GZ6M0a+BU+JuSM2c
mPAr9PJejvJEYP9lTE03cVGaOOZNLfVvX0ZfejvVD4OPXwZeAxdhjRDAE8MUDmfD
e+dYeIVLHcqRxG3WHGN+EpILkxn/pejaak2TqtmEGisoCp6qrT+PYbJfoWrrhJTj
2v4RFs7dXDZElaC8AnAunvPV1uJ4OjhXW48ICvJ8p58SEVTdG3QT2y+1qjivY01d
gk8YHFKa0ORjZU4j6xlGehVtLrWt1Pg4cJOEf/uvC9PlXKtGmkea1CIPUiFDXLuj
UZCCHT8mqKQ1UsRhqVihRGOiIibbQCEJ22rPNb3wk2/73eQeAyH+XoGGcg2RHqtM
z6ezd1QUIo1u2brGkzFx44cL5e8jjdbm59PsjBB2Z7pklXzUtmacspa9Z0MLqlEs
3rWPMcK6PtoSa/EFucQgpUI5rC/+TOdOaZxajYn/hlLcalXkYHc4HhyonC2Ab5MA
5jgMcSfrkya0Sh6cANerirGzg13rzdq+zukFG9eZkexw6podCtMMwaaZWs6V4fnZ
9G2+F/lyD1fXyGZMdwiVUMG9hZAFVW+o+oeUR8X66ZEO24HGuJ/Qoro28Z2IYMwj
1IkEVvQFU0d/1juq3LooG68gzdSNjR1CpB6HsyZ4ItbHZmnhUerZ2X1CIlCLlMy4
vqWxcGTFFX/TfEfhHetHNrwNM6o6Fax5TasOS7gCVwhAWhF3SceM11VRqM9yOmK1
ouYkcSuG0dA8xFwLfySI4nVOcO3GOckI/7IpSOAOpN8nZ8M+5lAzgbOT8Oi42Elx
Y5LwsY+92hkyxR296Y+5ik+kNiwHYPJfu8+cZa60RVCXv9Lb3cNI3GxlTm6nWeWu
GBt+3IdyTvaQHvzOXuT73EgvdVu4HWMmjTWCipradLcLaikL772Y2u21jMNnn/qX
yWIAp5xxy5xOezOSHBIdJtulmeHnHW7/qrCoUHr5VxUFgH0pINIUUD1GliGwSmaL
M8tVeemxx02uvW5KzM56oxexlDURnLiCqnX8DSfyzCIMFQu5WhYuSdjFlpVG60yf
VFhmTC7icJC0TK7cF+hfMH/uwynJMsfSRvd/Nsp+sdikMTVkPFnMKQjHNg049qYr
Z9RSyj55v0eMxKy4iuWhDXkx5JhtC1kEV8bqG8HOkeQBs+8A8syOHzgOe151ABpG
aPFu5ULVXSIBfrCrJJXqLwYt7PWvQeby/5L9zAg8pT1vrYlRBBe97OysQ8IMqIh7
BFnxmBR9JuwpBJYocHz0LcahWl3QIpHQAAimsPuPrgEGO4utZFBBUN14eB6gy8Jm
J3OUyJAwqRuVHXGnRGZC9kBji1957Nk8ssEXDgrTYTU+ReF3osIM/WOfr4j3rOYs
p/CsKkaIgoKkyDob/nII2LXQQ9U7YkwlH4VY+YRUoX/3a6rvXSemVr1oZFiqJQXQ
p1/4L8h0eOW0trakwp2AL9aKXberJWaifc0/HnTwk3+CS+xX8dqEHr8/25K8Dokz
ExAPl3trQ37KOZRWZvwpF9w3jSOrh3cRn/mNP0xkyBI9KtQYxDocrEivRgVRlJ8U
JIisHqXi7Ut//x6aq5vrAwu7iJsWIqfy+5rjt09nUDp6x5hguzY32y/GfQfk0UNq
/LDDmHQisp+MRxkUT2swpM5jQAdVNK6dR0cjUT+TLRWH7fyDt/CGnqd0+gayPG5x
nCAkFVbf2nB5Dsum3MGB7eXdc6o4f2Jv2fuF+Rz9cKG42YZzCPPWcIA1nhoM44Tw
Q2vO1zxqT6D3qw6XR/gGH5WLHwXD4KRb99fdqOvPfLHAq2KXxvnwaohwCZrKPFls
bapZvFBbIGkNKlGVK8ZK/4CBGuRJBEo2kL4wf8doooLccCzZ80l3NBZUWQx1WcNQ
TbLUcZYaft3dPi2z/fRbgBF2I3bHjkQwNnlCQFE9QQ0IslQdsbm5pdeWJxskKIy7
DvzDdETIcst20+KzXI++8eoR62bKD6GJdppYuUmdSqTygN/sgGERZ8qr1gsbMDSS
V7Qe5rMx/xWPzKxeEXIQhbgPD5gPJR21n6StdNg2uH2jFO4BvJzV0BiRYIVvpR6y
npV0bQF70dhNLz/a1GVR7D4ScK108ZiFn/N6sCGSyXekTVjMBn6RVXEyJiWthq7c
wmn3klhCvGdoosaGtyAxLprnp6YNk0n0DTK+6Im+sZS6bGdmuStA2Z3B8bjI1dm3
p/39gXSeLtFhMjWeI16iCZWL/NB+GqYMXfS3UwmDJ+bkdA1tqy6eeIRbhfVBLWh+
dZ71Ey8yDG/of62soYwN/PETN61BAjj4w/4ViLHY+DuH/K2HRA4y9LXRBMgh+2/4
/N4IodWSiKXlLSkB2EHSHwKk4Os5evxuiZOshEWhQcqEM5AgGrK3hafUg9g57mkQ
Wzq8ZKuuJHKAtFZfuyJcpBVljHDyvRdYYTFXQybjSB/q2fnpjgjVsK2oe4hGruzG
mpHDmlSF6OuMBoSO3xESu2huvhTxgRD4zGZcf9Z4uL23K/434d9yMJPWLG2dM20c
QHLR9Rqb9j2GqzpFEh5Tjwu7DvKl4DoOuxnZCx8775zX5dgqRDzBs4kyW4bA4mjY
2jGUejGfMCamopBzJxrs/sGH/LJx1cwrJhOXgNcQGKChAh9L6M9NKDChlG+8r2hR
M4fJsReTJDBc8dK1LOGGp7d5EZ5S0XVzAvXE3LpzDVm4RSHuGDsKuYR/Y+4qNorF
3DUJ1hWAtAr9JbgV9Q0pwBLA2KIHPJUTVrkydP5KHz12Xkk72dbzYfglCNlw/RVm
vz5rr9I5QtzzjFyw61KTtX+kLo0vjKek9LaLnfmMltITRq89Y+aABdlRAqkmqCxA
5ztsRFJRTsLM9ws4YI3b8gbAGN/5PCOENRlePLrFzeY+IXDf2JZklJDN74WCqRfi
Nl/1foxOGedHX+7nxLhCWws7JyN3VpFLjSzjwOjFP5tNKqfYXUAf2YiArMBb1vpX
yQQMgeGikrQSOhIBoJp5UIJiX4tf1B6H27i0TPQDCer0UK54JcexyFKAnMv2oMo/
G4cBh4xMEpvbjuMMhuTxgw1+zE2rriBcdphHi63LbRCbQwxNVW9Z1aFiuq37QAc8
raaB9f4dVCn1gMSsNG3i9K8HhWXvZSfw/Oo1vDThpZEt6WwFhm2IKuME/8vXib/s
AM0gbMK6IqgR3Ag8TKNADIgJL03HVTy2apbLp1ifMW9rJ+vdmCrYwQmFDS3wuAaF
pMdBudlC2oRNr/IScC5jRQuC425umrVJnZDXEeF8FKD5kfH71ySYapJWGTsJf5Jb
YDeqkYvp7+6/FsvqCS7ivJs/bQXEEe5RSw2AgaCxRU+wiyNyAwBksIpFeORXz1hx
bJL2OZEnpsjcLgvwhObAsjQvW5jYq4jubB9QufqNCkCElTN/+p6kY/Lys4s5Fm9z
JK1th0MDzX9zH4ZeR5NlMonVAeTfjAW7N5SvqjJ03XIKov8iqCAyqrFvr/j7lg02
wg+XK8Bsbbj2sEIhsfqSI9GtxBtm1A8YL8BCHIYsLmtYiJ40K3TkNzLmhQwZ2r4C
EQSa8AFXaMOCYTpUxscnBI1e5RgMrwwaSUI9LXAqVOW0v9hwedZ/qfsxNep7kt53
AOG7PNSbnoWeZD807WmVspcvWVXvW1GNM3lsH7WeHUCXtZXPMiTfI5xfC79Y7Hyt
qcASkCgzKrtfdWtbUvKucO0BLdR3gtAKagA3viAi/2edAB3zOejxn3kChBRnN24S
pk7QE5b+lWJ73yn7rIJYJh+egXO0o676yPmAaGDe0+2/Qd5tGDC/numgWKvLkCgl
YVPWF9eAZFxxBon+1rKrNQ/23S65P9KA1sr8T6nvxxVNieCKrksZqUq+N2ZCneMq
pOd5PlqwI0EJmzb3J0YGt1CZkJVtWN2r76wU1JUDoVczPNXMGWmOm8YIZWOKGKOz
t6+Cgpp0mvFWcB4OTK/TdfDTyaRTYeBzXg/mBT2x0sLvSX3N/d5i0BWsaXER+qrq
K22zBJCpSq1UM4oum9YPFlFb8dxK+M1ybXtXGzw1XhLvKv+pszwJFRRIxW0kLuGj
lgQi5O7QeaXBP91lWpwWwTwQHUdTklGQ8vFgv+VFT2H/TP3YyHN1EmZy0rjR0kW/
omBLzugrVntYtlqpXf6u6RY1njUbj1D6SXna0zLP3quvrrDryZBt84az8OSh1TRL
lNl7UFX0nqfdFgFwhdL7f1x+Xvq8FWpXQXTDx+6h+O68NhmTNa3NfouZ1xHekDmo
yqzbdv4oG3uHfsodNdf9/JepK4OFpbFpghlEmrzd9F9b33lrOPvd19MplIRqPG+g
PM1LT74rQGA9CB/U36o9yNYj4hgN/t0Y6VT+6yhlmnN4mDYcQK/9vgz5HkKqo5q1
IWlgJVuPCJLt0iWGk+tPzqY8FWLuyKmfaUHZXtQjEL4zMRFshYoiL+kG72vTLbFj
jyguTtVCQAVjVkJS7mM9o9ZoatFkv4Dihcjx7i6dYHJ721YXTcPfR++2wpNMuVmh
gbZ+go2Vh2MiQC2Y8BMcXmCkYurojqTCJteqnbOfiypT1MVZI0s9EiKVjyvEVZ70
UK2XPfY4ptccerddnAqwRh/+yLWn4OcQTarP1InEa6BmTQF4jYrxyiPrlaaFtuCW
BI4SrbSGJh/ebTf4CjbV32CmHToN4N+s7sFL/8ixXsJG2xQiwVe6wwlJdK8fx6kF
E6rWlhz9bdFW2B3iQPicVfNH4z0zw8W9R9nUfa4bgi+H/YTNR9g/9RrxsVT/k7AO
8AhaqrDOAVEitPvcMpg7upcNEF3o5GxIqhCbZfq8od5pCBcd58I11K6z8nMyr2WQ
0L9B13l/BQsX4Ei4Sh2IvT6lnm4Qaru/TR2EohRPfJt1g9hqh2BkPrmrryPvfczW
qW60VjrxpwaWxJ5qP53ZDlYmxZbEaTXvEPEoPt0P9Yhbxn2Kjz8bVGCPUUMXQB6u
RJR/UFryKwZz0yS866FRxhJGIjWiEQh+ecAz7ImS+uj/fgDBqDRNSpSKjorfGc+P
0CKgYqMwgzo5wTZgXV3xJWGz/whRCg8NFioO02HaVge5nphfvybNg5MzqYqYE09i
fCMOYZLSs8zkvVopUqH4MM7c/Doh4z7b8cUOyKgs2LrDZEZzVSSqp6oNzzvJD97b
iVAxJF+RDD4yLGy6AVfD320AMYB6hcHgv1t8Hpmnh3ASq6e0MYKTIDameDjSONsH
vBRtXgiqX4W4zeyVTcwbWwKrBgx0bp55ATqC7InzUTuhHeBWbErU8omHLnkOgmGC
B+sxl7eAaO5VPaUQ7M4JBkJ1yylE7RgXmFRYIu4oxmaJVp3M24ZYMHMnmY/LDj6p
CvtlLjmXMj4y92yCpJQ3coV8AIcmW+fT3/bdelAavHp6a8qkGsds50qCspmLaEhM
yGIiU5oxn9IP5fsFUnxuJpcZYk+1QBPfNMM52tRrnIhdcGQlwcWZCIwICfY3OdYE
DhhBSHm7aVUHU10HPDgio9WurWPo6k02lIURKqq1TLQlkGUebAO4HOOKthiHnYDW
MbygsbYIOFlyNpsPuoIkG9zouq1dUEt0yuH/bLrLew7IM1/aoBMcCmOKsEiAJ8Za
PtWnrjbCmb2fGjBqS2wQ+EupTsvJdsXw8W7pSsd4Qe4MeqXXdwshWJ5ayp+t+NZ2
wX47vgAWsxDO2LQU7Qk7EJoxt5F7F/XRakXBjqzrwkveBxU3tMO+/vP97Uw6l2A1
bGH0H6DbUymJtC8zvqpGjQlZl371U/61j0N/ewmshgKLzASpWq2tZo/JkUhvaBH3
6RVve/u0NYiCTu1aE2iFIl6ponuoLF6Ci/3TyN253BfvsMFOVWfo5lEQiqDsfb1a
yM+2BdX8Rb5S2WlxILBKEybBBnkGlQTNWLnnIMoG3Yviuw72oll5qbfPZ44srpYI
SHL/+MUVifsKzVtrr7mCWtBF6Kacu2PESayP6LbM/jzsZGjQGRNMJMYJcRWUd7x9
sK43jd4ZzKl8yTVmPNvjrz+o59J5d7l7vJNAAmV6QD0BosqCkyWgkQripKLUk22E
DOMWi098FaWuTVxVqEdbp3BpOJ4TohKKfPEF3tJZ34Dqlwf/3fNQKGKJ/AV41T/q
V4NvHCyE90qWy1YoQv+08MxpLekauYknKi4q/8vBS41m0amQVvnIb7QFV7J18bGY
unMFm5CI4SlOU41ROd5DkijEtBaRBselPSpUxPiDmlWgM9VBg+EiaX1tDETJnEEl
36KsBiPayqZRwWLYV+Kc74m5w/6EdlaW5O9yESHp/oGOVac02teTzB84B6FrM3HX
x/twWVQDD3RwxiwqdCVZYoTQFDh/vAYUWeRW7ORnsL5C0zjPqv8mscfWzRsyW/Za
WGRBfpwiZADKEOwRQ1ZhrK68CgYuFnp7ywtBH6LEPhH/641trOXjfvhU+m+57hJY
Fj67p2PnXyiYVmwNSlIzuz7TydygsIEr/yR4HZgGwn1W728EwVW5JIX/Ay6L6P5x
kkI88YcPTey4ayo12/9Ks6wcgyVik7xZT/LY5y76nlWKfQDl58Q28IM7pkucBBZ7
HacsJw+kZpZhb1Yp9H3rBhGZG0E/yC2y0jJ6WyW4BhQDUgIAZX++fHyPWeXROlf1
F/8WTFB/fMlfk779hxIKMWNfk7goHk/5QzMccQED/4/QNxmQu17OMFGph2xuzJQi
F3Wgw/ndWPGJoqcO/xwuUYWEclhFU9Xurr+ZIIq4W/9f43ZakdSTWN1MKaC3F2wq
hASHNW7JmXnt3Z6pYjKYm3Qk18I7E6KT9Pb/ZngHjlHvZimiXuMxsqs8GkL1LNfz
XZpMGGFVpPYkfDaqNSF87NR+ETU7TWknBi5qaahJRDneaaC/beKGPnTKfagrsBWG
daVRL0AL+KiX7Y0539I+QIB1F652eJLbTpqg6PX4VOS/QVjlwHlTkkZQw0QJkG4B
PgN/MSr8ibqxoyVUm2XBgrkKIWuheunz6Bbe2lvHGpI5fxA00O3qQzGgtlom5Me/
LWLk2lCryLt+uzAEr4/KSCM1GJR1iN7bfZ8RyQq8ii35PvItNYdsTc/D3oJ19oPo
JyZOamuPGXNMmpDLtw17/Ot8m4pAPdQfOYo9tQ77EQoGCspdPfXaBr+FWg4lURo9
KN3hZwnvDv8PK7LPBfmnma+lbM90YdmrpOkH9gzuVOOH/KNbVIez+YhwogP6PZmF
GxQc+s1RROcrk1c+OuYqT4AS1ZI050OhC1qetEmIfKhYRA4MVEdeqYD9MfPkipw9
Z3UyKJGeGQ158l/+BINk4cgI8wKrAt3mYIFrK35HYl2aEtlzpI8E9bL7v+H6sUVY
lPFOFmg5IMBBgoBvlo49pW1aMDgbqyiWwv8L2rKK91oOeTN8Yg2SywsVCKaghr9w
Wdyuxw5kdMobWFXFLk5DXgOAS/I0gSl4doCzeQUr/F/O1riD4V7h80fGp6dAO4ou
OQk/9l8OjORh7z5Qu2dAVdpAEYgPF85riau7FeGJFke4r4nF4YWdlxLjRvZrlnOF
bkRIRV7AkN/5bPLCxXC7dY+Q/YvnoOVYRk/CrYAyMC1nSrdcyHYuKa/FfNlCN/5h
zTCYzexUIWoPsLDe0qd3WItjzm2zTgmdFs/ndUpTPeOrUBINcy7FD7QD5yXVIyZq
rm7g9VWPQ6mLhKO0i/CyDZaOlSMWzwO/xTAM0+oLDmRVYQPy2nwQ+O95WqHi9+kY
ttzwimgJxnry+8viv7sUA99R+gDaJtg7ciSQnNlISpY4GnOWCQVnJFcV6msWPKmA
SD5PjxjZ+e4ZU3kXDFKMfXRs5Sv1K5KvgD316ZKZorqwiffcBAFKB5IfyQeAxCOC
AC2Nh32oBUQkKZkUUs6qY7OH74RoMKdJ3Za4bi9A1yqYTUmNjXvlkpA/ZCgj00/a
MCzUV/OGDjxVG/C3HaLJvYPRYRpyvFumU0VcNkdH1LbQZyqbd9DlzUNrcvK/HwI4
bNbxjVGm44IZE4U5RnfK3Z6FcabgP9bBnXIbPHm3aAMY9ZEQdfDigbsVjtbKxsSd
NotPTmtKeGKFbX1BoI4kpOqzfeGZAhmEmfciSPpgbQqIW2a3xKDRuDpXBxMd5Wbw
E8nmU+TrTds1F2PAslgt+zWgi6kajtqfpsUWdN0Xf77CvvqW+iJ0QvfPyDXgZsup
HxMXfjBEfjUi3lwvBfl2EJpTcZElqqFo8ZhSletQxRMAxqT6uspQ4CQq0nosIxyC
aZVE45K/JUYZajrsMvpPGvgmpb6QPIDe0n+0Pv7y6MSAdTGH232DRPQr1jS9FYbr
/viVH1vLbcgacvuJVIzMmMdnHD+dZaidtcDC9yu0sHYGKJFI2OlIYYB6zWahwbe4
DFGjc2xTCTCOfVnIBmMuPYRkKfbanDRz6YFtt39ujB1G4V1Suaps3AQ+oy6ZJPdm
VgibU+sEnB/lt/81SB8mAon/chvvlJ9uVsYVU8ZMGtw3gCYugJQ2R0a/Q1KbAPVy
f74FI2qwo6cK3g4QZXkK3ytYPxnDpkR6XQMs86VTX4QY5U3ru0JfPUQmeay0RK82
1Rxmdu5QvWWPDltKHBkQlZnxGC6N/n6qsMtfdoI8mKGpX8eMUKc+XszMFdmFcvqu
ctkf1ZPeKi0PDDI6md0oTFGl9LXiVdcZCvG3lGKySNS7e/p/x0huOX+wVW/48IiT
cBtRYqu7uBEgSiZ75jCE4MlQPyrOBbeM1xdpcOPUB5EvhtFzZdeuX8OuST7KMnYW
vraK/1WHFfC8z17jcwRPI1x8Gb540053V0AP9YOFuDqL19vda+/+X1/7y5U5Ic0d
s2Xd2l+m5Z7x0NInH1jiBbQxNzXmyWyn4+9dWECC3IEEyfQ6+5+WH93NMnT9qGKT
TygzTVd4CX0dM9RlgnF/qQ7YcpGITcxzCfpCbah2B/An6Q5JgCfOX4ynO+i6Dwkl
BYiGYmHuE0NaqqE+KLzpT0VjVFXj4dLhIs5EhgRaPa5MGRq6+/nCeyiD2eK/m1I4
uNGD68GFkOe9vjh5xPv4N3GMqun5tcpQ0mmo9qQ+dzqXodWjFKUdq3giORxCBS2j
2+1B8QFFx0Iy/x83AHQaGcaqrZfdP3qttskD+qxLgr6NhXPFQY3yLIMXK6T9WA4h
qURl3CtnS02th9vGBFOHcOyYoAna8f+GS4cHVZRUCHqlSATz6xL37nbIkUtf29WS
oOP/vDtkpgmQEWruLEIulYOo5eAH4aSoE6lofYpG6ZwiETqrIgtax8mKZ7/cSasQ
whr2ki+EyvjB0WpomD9gz5RDz4Of7hUi+cBd736GPEDxjuUHs37nmSrfkrut7vQT
sC04L+DOWbNNkZUC15c1huBoKmCHFSPbmE8tNbSbIKZwxI8tWIK1eS+beg0gVnzX
2WmiTEyLuFvR3+gsowGe7kIqBYjrlGZG099X7FthWvY0XzsdOxd5p4xoBmWuu0PP
u7ipwbN+YtFNoxONNe1byD5LHcWZ2BJY+Mz2USoAKT8+BQWuBlZ3wCk8C+ELirP0
X/lF+px6TNJz1IWzFPVLUFHx4DEsAtXkBX4eDF/N7xBpShtgGdQQ6v/6hCdjWNls
8QlOeBYJQHud+82bxkY6am23ZUYd6LJMdqd/hXzWRGSerJBolqQnw1+x3Wi4agnT
jxZVjDeq+Wen871naiTI5vZtTA5T+PC9rUKpJIC36B0fh7e5hv0eX6yUQIoJaYs2
ou8YNPacA0Om1ko5zlvMGaCz+Hm1cUA1perH2/uGlo2al0wFGEg6JEV0S3OOfovx
nhh/ICTvQoDFkdK+yZCagptN/lCeypndMrjVsK1/uGH/MHaMeqxk9Jym5UfiCk1N
3NhMvGWFMapDi2kJZN8aVfftIo0Um7O8Wn3rYZqgC3Xkx+g5x32dJZP/IZOvuDk2
wUbAOf8erTNPcIpEXXUUMTn0LFQHxQNbdbgEH7nCiRA/4shK0lIZXLBruNhmtX74
ag17PIvuH3ih3L8NHodwOAl6b+jHwDEUkQ8igMrLYS/IwOozDL93Iq2mObD6VrNs
AnyQ5DnF0ZDEQrcmJ+qjCx0ngUw8f8aWWF6h4X5uoEaPn/Vn0mpJMDtwMDqigYau
wLLRa9cK+KCtwBUnPk1RaWE/Mn0dpXuP8SUoKhCf1NSSENVE7k7EV2p1c24VMa0c
jJe9iaw3AkTP0h9fkPCe+sjaXZWkq52oiG1MQJ4SOq3ZMNdoXtg0mBtEYg9hMgQW
jIZ9gqvMNpiUzv9rIUSG/9B5ye02mw+sxLGgrJbv9OF0RSWnxw7x3Kcd6FbwRHrz
DpcOgHR4fH5gqFV5r0l6vc3fnTv4MNdj4P0oqMm6Y4ZsFBv9WGfrw5VaIlF6OrwX
pnJb8/kVmHY+p0baVeeoSmfdVeRxop2YTjK7veZ6LOGbhJ5q9315uO1RA6px/aeW
aSjCXrAuHyaR/NEroOMFnFC2i+AJ04u52wfW9gcHLZuR6aKK0PPP9Z7FFisVHzqW
JZfOZzyZDL6rlQqlmdx+KPCwFxlQtc1c4c+D/uby4NDg2atepZp7W2Ldxpt3V/0/
BVvycYe+eUSTSjCO5X5idWhmZv6m1moM1arF9R4yMJxS02F6WvGbzeynYf3TL/5U
XMsIihubwFALN2qoqUgh/mLrN8eiex6/3DasTROXSxsKhYJ0Ua4/JRZPPPFQQAMn
8uh0cPHHGZwyXPTBEO9tfjUawz7wjgTnL068inNsi1g6QbhZ1+XEshne1yKhMouy
IkCLocT3gr/KGfmsXAy/qvfDYvtNYgcEb5ZeUVvU+kWqrBUqTVtf+UCRXP9OKMsm
G7H76P6nzUkLhprNEfDAvI7gwQLUNOOTvwPDHhK/H21tAX0HyJQOZHMNgT98P+xL
rdgSsMub4Ljqop0YltqJG1u/1ZzoQPUEX1hvCk/zaagh+Bbezgpwnz1S8WXMzcDW
buTdqbKmuJiZEC5RKJe+97HxYoINPvjNNVV4qQ8km8Mqozj/NFDlFZCLwiwXtVDh
kffZdg+rag2P25pcn5KsArbyIqfrAGvOeOndrqYXyQhPbu6XICrVNOxVd3gd29Y1
w9/sudkR9fuGJNQQb+8dGtrODe2HS0NGL8Xt1DQN78ia46GASM76+JP8katy7Alc
bpkAj5mdk2+WpZc9yyizJkm6QRcxKLqNFWyX/RZObJ5FBcLvbAHsAlPienJMD38Z
GJkUjj9cSI2dnXTtx0UqulIZ0Lnd0aWjVB/boT2OqUy9MiYwmCqDIlQe3zXUksSj
40yAg11im7cuLw979sSkR3LiV6oiJEbVL4h3Kn86kko0nLD0Z1ar4uskMHytmOvO
VJOLck4aHzqk/Osaaa9PEk352fCsE3bbB6V2BUHuXRe1ERcx6aMab2GryOE+ZxHV
a2mCQJRICieTmfk9WpnQow3D/tWdiEAhmuzDLrPBFzmPrzGIHoYStkf/pR9G00/8
qoS7Elqsrr0HFa868E/jQvwQReZnfj69mEaeZ0YzphyTpE2KnBIszOpGQIDY+ftG
4j32rsSSx77cEOFsE3gW/70SUghBTsC1tIecchsfwvt1qUOpz6cdxF8n+kLiDw5t
ob8vE2BnSzWKswpscXBsiThmKtbE0ZY1NhC9vI07FksWU2v9wUSG7jK6vUBWLAqX
ZoGGi7rZ5ppUr7lYYRQsR0o3sVtPjNuGez4pB6hiSLtaIrH/zVMETyBt5iELovtH
HSuHwG8H5m7bIkNDxo7MRMuwiiLANRMiQosRqMHmkC/2F+HbiwXy9XFVfMvdyvv1
QvDcG4tf9rH885Khd/4ns/EZp9tuK1MleB1SibTfl/V9b0CaFwQ2vXV85hlhg6Du
mvdtqC6ABWE6a1uxut0K5BPrqiZ50bIE/TdfAwCN4G7racwLMbSuhEBhzl91+LDW
Ck154acMA2JComdPRrGclofpoNJdv9kBz4EzP1nhXqXpztqeaZZloAlHz7AF7Ie0
DNxbdAK85fWGSJRzdPJOE2/DOR0hdamBAo8CXw2FyJRY6XmWfzTPoyOTvISw1KAf
P7vqkDkUNWDcRB0BVnBGWnldYqM5mTtK9bc9AOm+nw8KkzWqjyRTQiUvllXpHtcV
svfukXbWp1PALxiGFme1qpRwqEjgTzwHQ4kT+MDWlJyEaBoZNx6L0zY3byGdi/Ln
dpEDU0WiJn3QbYReqbCJO37yeygCFJPfFPmO2XW/tRPIuU6fiJjkHu0UV9EFaBSf
70LKbkPVG3M5TmUt2Spt+2Rv/yVgJaQK8HzDLsMbviPhc3iu3gt+OUn/Ur2pw2zR
kd9ZjKZbNKpEbmXYbAejF51JQo+y9rxPVkwsJViuxdyYltiLqWu2rWgLP26dCp7G
ILwljyU4UBSOHLjo5GSF9gscT2vJnmz8FlN8GCPzq5rBxZM+rmPLn+fADBydCduj
EXhi0QOQDWDK3tHLT6+QRyJIp2SIpSVhIJp1FA41kNGMd1sZL/6doOmYxbgFdEnR
JrMqY7PwQHtMrWVmyjvsKHiYDyJtXAWYQvkMGN7YBhWKd8nCh339LwB2imHgl6vp
z27Zs3OdAN+WQRkoAvVwaRsTmmHgoxB5/V9RC8T2VIP47v+Mrvh1v+daSFuSOLXi
cDXUxfRGn8Jzfuup3y59ecgCVgWkwrGQuJkpFui+KRuMXjD6X3Oy7Mh9KOO6ZqTw
e3VMlbcpm4BRWQq85r5mZJcw4td04cQk7vn4LJdJuOEAI5FAjvy2sG+2HuwxgSSM
Aj/mvKIncjF16n+88dzGq9QCi1p2FEsA5MYZywJ9wtEhcg88D7YmGF4PVdXoZUSL
RBrfX6Hz2GA7h0teXS5L1yygi5cMeLYph4csZWRSv/B97xD9WfKYziHGF3y+chyC
48jGTiXTfxBtAhoOv70enK4nCjOL2ZMCKMkYVRIzZjxaniQ2MrKyaWSTJb65M/Ee
Nb/jOJ6GGZzR01yQZb98UAbkWUNnK2bVjY7TtFIKmXAF0C2MCIBQ0XKihU/tq3fd
FnqdA/rgf0Ai/lemF9rp1GOjSj6uaXJZkTDL7nq1rEATwC1dm7qOvcA+5+TS0YD7
cqZeIRld1o3wSWLO/v5gUwsMua8M+0uIquoVqmS/vVUF7hiVAwlVFRvuVWtrSrYk
tdA49FW4Alj/DmVSc4Ag6AboUOTjjBzS0ZIYOVkTLq4jdCGc/wiqOqoHwkPEhCyA
a7TShnn5g9E0LAMGsrZ8VuX6uFcvgpT+eE+g58Cp7n+VeFDEfAZR1NEq+ezval5K
MDf4n7SF7p22o7Bs4uobHGT/tPYD85j+Tz5EaQVKIDrlozQSolaSgYEH6yQ61ZQ4
ez/DzBOU5LuXid5i43sGKhmMnHoG+BtxWIolhqHY8BWdrOYr26pLm6ig9MHDavJu
PQ7wwVe03YeoNCOUb31FJhJ3xiCJ9BL/1Hx2MgMGSIW4A1QEezOSUrQ1avhr3Jqo
bgw8OP1kS3sVH8wQoqR8LbNk//4KgkP7v/AQmrC9BUY93L6XlbKW2PWZjFePEDAB
H2cTFXw/3UNK2itsOJWfSZiQL7bRKf55Rtu3ESq82Ubf4nVwRrmQUbvjoDEs373J
XA53R3n09AfkQhwF3+gCE6IwK+NwxGBUKob2IPy1mX2FbxoeCxrkSlrMDy3Rdbo4
WNojqRZsXNN0u6OKg+apJN9BDDzNYHpP+VkdQQWJ9zWzIMIbOwew/2T/18KlOc1v
3dDcs2KCvx8HkYYKCZQRqraMFa1eXvKcw1zgfR6aYqGiK5wAyImYsuNaQS8M+Roi
a+5r5w1Z+OHdAvidHgO2cCpLKaAnjgzJve4HF2bCGEosZxoqUBStYMTY40ie0ksT
kMxe0xIjJM19T9/cWaHp7wyiNFoCyIfjLpDQlGQZ+qthuQj1Kg9++S9OOcS5r/xr
o+4tXU6wF2l/w7hjCt5zlZRF0EO9gZfm+34IBxgLIDtU9JNq12uD+u7tG+zLE4JH
FT5GeKnJPytvFvLiZomzfaZmTImalZgsqfQ8uun0raGgw290x6eI6Opq5w458tHI
gPNGLQq5kM6ELOpa6hV2q9FfsKlz2BObMqzh0bgfi+EfUB1dpgNgi7bbGKRSsF6j
S9ICuCK8f5FJSP0iXAzHxgn3YqGYcnwv2UoCOzxczxwNSZ1hfkWWAqu4tmXwbJjH
Tg5J8QI87+sceXOKRSa7KuAuY3INlVm5o1yq7lx9amDZzqCqEqraxfqN4ZO9wmd6
tJr+B9bzdjAsOIf6nkfWFaVdstiwiI0RH6gfXW5kx/Ny8UipM7uUvm05TsEkt+tK
WbSEHxY4RImBuzEmQamAiDb31FRuhRQSGfS6ZJEA+kQQ6mkOtU3tfrMk2ySh/Pn6
eVZXLfOhaP2UbG3erKRfbhAlJvOntK6kDKeJeVtW1zpEbuUBEOi1nQixlFa7x+wV
EZHLR3kQu5J/VRyrCULnEbCx1F+1CKfqABYccD0Iq7XFar1wYXmaqFtve9j6MCQg
AgUUaendttsH36wtJyXyLTWvmEFRaU/KEuV/BPAdNOfaOJc5juY2TM70W72Lv6pa
xUKOYPRvrYgN1BKKNIB9ZmxEgohLoIiNGDGkPLfwdqnMjv0GchWMorOOH9B/yhaH
IXE1Yx3bH6N7GthWX6eI881yIi9Kjpz5txZ6tZ/b51X1z07zfce06sylFvAWD1U4
f/GpV9dmvMVvrB/s2UodPeIaD15EJsDMt30Wwx9AsuPsNHmCr3TTckbW7cJfPdYC
bYYddKTC1SdVDvToAbM5STHRj4CPkYRyePCvakL4+HUXYqHyPbTPbTIQbUW+YD/p
AMHqCrJA/ydpyPRdi8kGknQbOGCuXKRDGEl7p0M/ZOdAl+d3qp/DCjW6mUnwIW3s
WxaOYcdn3O7lInlJXsw4GSkD0b0zI2UvV8IJgHylAKAy1t4UUsEF2Ldc9h/XxcHe
aNpqVASWok1rIpfRV7E+nDX1yFY6OTUYfpN4LBrYvMNsHCpL/RBd6BBVH2O6jWIn
LKBi7OJzbZ172YkIgEqgHOyHHbZ0ER7wEHcnxnnJOyYrBu2pGaxdJVijvmaCr8W6
40Rd5oFprr57j4KzwYGbMPqClyWq8jVc1Y2mox1nyJcG67n3I33jO2faxSR1tfGg
vKt89x9D5+fek2YUwLdI4tZrXmPFs8HZhGznYyizeK0Esh6VNqEzS/NJ8qnw7jKD
psoD2Xcp2CyUsqbs/U/AKHHZyP4jI/OZccxZnkcHxqF5dp5ufKNv8fE0KtEKMfB9
2h+fK95qcykZv6rt8iqbuc12IcHmQOZRtvPdAKQcZnSbHygYv2JHfe7jTjIphGaL
YtIlsbprHeUXCt+UlzsjZnIlVzhwKHsgYQp5o3lugpRPcZwqEp2+hgjmcWrHCqC3
KyZNko1oB5Wj2K+PDo6jpYiM/yYo9mVT0gDGAXa9xuzy+yGPPZFuz8txbJSCEVr0
pBJvgl2g5W8yqVQxebDDxAIJRR85TM4mbt7p2oBSqLD2VgOl6afGrPeQK8yNG2hz
Q3UW1vWDaZI/PifrnSaXbmMbGXNSe+XMgFdI4zu7wjcjsYQAvLRJ65LtKbxc4Gqj
kpASbj5kABOVi8VZ8UuX8JUFgthk/EDng+n+jTWExZgbAKd5a6mN+0Y1CtOGv12a
ukUKDYjOcPPTcfBkT9D7pnMBO+JAlqqzxFdzOBz35UHKYoDz/k5e2Dv3wslTFnjo
qpxs4rX2PyiTfv2A2PPrOgFGt6WNwISz7SCK7YuK33csjNrF2q2GBDwSxqJxfKxu
ng56NPonsimtz/PORTBz+g4zHNNPl7rVaPjnQz35SH3MOfMX9v+Em3eCth2YxdHR
xdvAwtP3nrOEiKDpaLfm9cpPeyMmVltZSy8siEYaMgNnfEq4+Hcqyp0NXF4Kl2TN
CKCTY8J4zGMdPLxSYjV5caOKfp9i54UBDvASplEwf0IODEIXJzwJLAhwde10AMkb
GFZrH1t4PyRL15Bl6JF7fKQMTyzmxM2jIqNLlTSNKNrgKP8hemEdfHVrCq0+KNY7
nxD1Ckqg8h5o+zNEIsCup6QTBfD+sN6nxxCqPmX9UI3YWtLQGpCOqeuXKkz5pWix
jkdNb54d5xMxXAMZanv9sYCOn13G7dLFf0ZSJUn0Cve6m+WWDeotjyV74E9kk4sY
UPEo7QsdLOf3KkLPnWM2xnP6PMq7aTf4YDWpx0enzpfcgk/pvIZ7p21I5f6firFm
m5rbqfXPbpW52iQ3/Wzgn8I8VNhoHlYw6/XGZmONJSt6DoATi4Y3AeQm9gw1IVpV
a7zTs9XjC8K3eFCY1CsCQj9n6WUccKHTYZ9z+aAvP8wpNjigslOvDgAwldnHw6P2
louftiBNEi5WIXbhOzrAWbjhUQx1WfbqKU5l0GorN0CQnN2nCUKBQDITitsrrvHG
+XBpQrICf6hOVBbQUg8oRQXAMDo/RrKpGN3W+2fqKNnyasyUyw4ygrvlusGBwBOQ
MaJdjd+Z5Ey/4rMAbvBoIyHiecso/gkhJC/4i7l9fGCSJ+vsBGeKOjKF6y3R14Pd
3RsY0/4ak4GnaFLuG51eZkDACmF+bQd9d1tu/NV6Jr4FWuaKQAct5kLkEGhVVzE5
PQhNnjeVRwWxjpJznilRZeCZBcctCKdJ4rMHWtnkzKJ/shEZR3fDK+m2bxDcAjXg
cu5XQfWgn15zOZgl+szqa9WJtjVJhlxZ3+kYzTgs/HXPyRhIjtIjKQdowcuC5793
XxU7NoDdoYB+wrPvl2dJYKVRx+5Nqhd4sNpMb1c9GD7Wgem+xWdDSCC5hIasKlBO
kaOtx9bewbyHfkUKNFJ9JazsPBr3fQgqkctpTrTwyTsVepzdOnFfkN2h+081/P2Z
cjU3oIjkyGJfL7HVHXPpnjFJoDCkfI5MrSpia8rD3iEEtoZh2dSt57TXFkrc8vQB
W/oXMGqLVRgUIX7sNJhCCTbUs4bXgIgrlDeFzjF32D7QwwwuvZht2WCGZ5K+lmy1
XR3aeiLUtuma3jrBG0XZrDAvrBrES2A61/Ga6o2ewVUUMT3eGGZDAFLgrxILORkd
w0I8RIw1a3AvHRcwiq0lMvWe5THM0VRRn8iIEC1IgZHEquU0Be/tittlX6zuG1EM
AKG7XNEiFtc5K6xgCXdQO/vBvM5ChpA9oaXyhSwEEZmyyeDr+jWkFcvbVm6xjvzB
7zGwUvTt0hm560hzcx2Ub3iQxATQnzHD6X9nDocOThSK7eimmNgmEZxjlCB2VsiE
zThWAaV6CV1gxA1CUBdFpler1oGzVe7kOwT5LXAt+iu+aF2zQHgR2E2qDpVD9CKH
Ruyoh+3kwfRTu2NkM57079dJT9642A3iPLvGaAukXPm6abW6g12a/V7+EghmAvoT
n7AIwgds02F95Xo2dWDl+J5BsE7Hlb6SDasHVpH97fZBtAR1iTUJbR3nSb7d7HYf
+hBDcWvcnhcGiysu5c8+XtJB/U1OJp/T55/UdQw79+Ca+iaZZnbsiNZ9vQcn1Cd2
b4FPp3fYLAeIsTYSQ/SKe8bgOg/7qRBgI3GXM3BtCFnEuuOmkzlZF4wORfQawj9p
pE2GcLVb5/xAD3f5YDjo9F4TEb38QAu9U+AwLcFx/eDOonGgJYbm6foWydUtQa6/
6IPEFVSEOMbs28IQCYnWlxgFFI/OBsNL9Vo+cNuAhAfkzZWj9y9Dr6XG5nP0sRN+
vqZKagvC8bXXgX62TySu8tKR2NBLhzTin3JKBmquQMhelaLQFIritDLPKv1DBWNF
WWvgJcJhC+4rQq+uSTvD5yP2DdgwBIqjbQISr7vk/p8ofS/iuj/ENR2kldvliSC4
afvWQA/Z5sh1uYxL5QEVHHpFpjEyjBbBbpVcDWcHw1iF6RCxYDDV0ZhqpbchvHuJ
zyPqOg/rBBz+c87CNNahPanYDsRz9Rndom3eoWgPBI7BKNW5jOjKOwvR+xFw4BXX
ggKin8B3Ei+wdO8aO0pvhXPZ99ZZOAmUw4bsVjveiMI4QNJSAYB7swJ3CEeNx936
JCfsWcnEw9qzoDvw1S9l1JJTqDEIKj03xSiMuKlgFIjtleUIW99b48y6QXtG1rNM
Hfs6YyPFjcxFpoaWIMCZ9E+x5IiSpfsqAyD8NWiJf0i9cgzSXsAsKRhkM/w+Ebq0
AC2wRJQeIT8D/rbUCPukfLlTHIM6go8qh4kjv3ctscWO81Xp81SLINn3O5qLHfeC
GkVDNomfgFX5Y7tK36W80AcOCiSgFtfHEqBtmcc4a5H93vC3zVnUV7bV/lWpUlqr
iQSLHoq1xikbOL0O5dKcGCK8nRxxHvOo+6Mq6Xc2yJffeP7Nukv6PqYa/8QdG0L0
0TrNU+9kOFWj7xm5LjfK2TxKt6JnZwlgz3q9rGFLFt46sYp4ubrbyxIDm2nWI8vJ
ho86iJEMkHBfYCI8671DYdXbGH7PbZfaiXps9F7tFf4kuLCFodOROJLBeqTfN5IF
xgvEq9f8TT12Twx3B6NZCMjiXyPVVMHvKHmjOABhnZhH/0jdSFHY9DVeRnAHdFWp
5ZpybcdXa2uMB93loxvxnSuGa3nBTofYtzyV9WEKiXtpSwluKjCVY0gGZRirKrj7
/Ajsla3oGJPh5l7jsEENXWLqUUxh4vOaiS9xJ13W3dPJg2y0EwLmAkwquj2P/i3J
D7GoHBbwmgdVd4WNFofUSNfM5ujjdUVDq0aTex79KI2MILK5wH/60hpcU7OoNOp9
ZuTLxreXVBEKAJFTPPc7IOCa5Z31rCPDRkR8aq0JTz4RVgvn2ys6wKYY6QZguqN9
EVTu7XIABLOF64l2V8iyriGjWl89/8/lpnZ4lRbBKzbZBPwrW7i1Y8ozcZXPt0JC
HgpPZltieqX1m3z19ejs1Ysobx126nHoitNwAx0IToAI3L2dytyyQ96a25i1PSbI
BfC2SLKVZhEfGHAVWz8TIzMXCmroWCSNALh4MIbFr2I/8mn04zMemu/emsNuH+Do
NhEN9kn+arBNgaZSYAS3GA1neKfLUOTXJm5L9qo3aKmB00H60XMak3QGHfFWLqag
VeIlZimctJt5VpjeTPWTFtOI8cXPTDDtWC7bhg3TJYp6ghvNentrMTVF9TM3EA4Q
E95s75hFCDsDcX5Nq1oG7LBSzt7kmrdkJQ8Az3uKUfeRPhztZlwa091+8yoxBLIY
C+wN7kysrqzMFd/RhRStS0yIyeIMyH/UxrhuGdHG5MANvBlPuWMwFzFXyHiSeB9o
KcslL/UBAKgfZdH9y9zx9KjvPbRI4hwm1JjDz5DRRcjDyZ+ldB+QUd3C4BbUNSiE
w2ytUbEZ9wkTpGY07fDHxYmr7zU9fpu9w+2t4DQqabh6V1gbJmsnKoLHYgF6MKD4
VJY9bX1T2qZs9gGXqO2el/cCW1CZ71HZ1nVcfXjz0k+E1CrwO/4JPT21kjOniv5Q
E+X5DyMmeUDRjndL/9nSETvQU3umdpJ7KTjF8VdPKXrirFQBoqql+MUSF/GNes1V
zn2FzZz13GbIDlmQuvYr2V77qAyE3TMNfm7KT3Qj4kVIckfSgZ6IO34Hrx/Y71T+
t5RPz3WN9XAGLxNiMWV88CcP0n9Bywwq9MDRBVArkVj3FJqkqlR3BgibgH0qgG/L
U5Xsuxb6RH3l8I26c+0+VNX3poi1lFVzk+J5Ucej2DM68Vl040LWSOBJZ85eVunk
+wieSYt3tzpfDtsay2GEZrKvHEOB19ouKFt+jddINJExSHBPU918m2/Bahj+DTcs
byp7JkA9/TPe+4io3Jo1R0P5Zy03w2GE6BKUoL1DkyC2LNBpLeX1yD7aIgpwYf3E
au2OKMkiIA3CqGxS+Uvrd7odIm81Ndzy16Oe4ZQphkBEwrPP5n804RF9xm6gxRug
BL0M/Fh/Sh/RWYSmQU2Z15flZMEvxmDTwsOlKv2twCKAZLQzFCVPzJMr7Nfw6uPb
o8PI96rT26jhyJxJ+6kEqADjjxAZxwV4b6Sz7ZxbMXSdqjDpeTTOtt82UFuVk+rB
Ke5w6PJWeBBFjXx65uQpHbvV/0gcVBNG9fY9Vrz4UcyRFHGy8sN7I7P/EWMB8Wqw
h7D9MCMmifawsMlNmPGA0zUH2YZ2J66a77EzrGk2AUZA1fx7cY8cMznugxIu85SB
jO3DTtgoX93DdiOX9pvm1oEv3YQ5WMJ1Z2cMlDNKtKkzlGfr5GuZcdtT/5ltSf/K
M0qsAi0Sl2PGKCQrknkuTUmSiPENu00nfhqedTjCFtDxDhTbUwJ9xbzxGmUz88vA
aDk28TT0sBeXqwq20gD9SmftvKS8VLz4KQstZa6BDn0KN25gIel04w1hLwHvfma0
Ao9sOYj7T+y5RfnnrM31zSYBeQ3NK4FcMbgTJsZZVViNPHXAk4yZHqe1uf+ZcLaX
9NFSN6RyuOmmiwqkUrdJkND6uq45txWgzFephif9lG8lhHHUshWqz4zXyG12fgt9
sjSdf2Y6jKvV6z0lGFRmRucOOZqViUgrY2FN9uWOYSZScBdczeNiDgA0w5Pt4m7K
JWYaPCISXpJdibbBUEjRfgD/YdMgY3iLkZBDqMjHMiOo9ClyznFHbYHYXzsd4qRk
tsnhglrWJexYFbP2exSU9E4OlsJzduhCd2YPXCduuiBDRfHxQ/J6tjBtTzTrI0WH
h6/lJMKuTl+vd4f2WyVmZzsD4w4xgOvw6LQwVTm8m4JE4sEE688amj1vLhjwTbQ/
8pcJEfAJqoWAavznRq0tSz7OZi5+32xVUs6J57RomWNFHWCxM3UsmlnHaTwvVz4j
C/y28x1g5NfwXd8jcO99M+JxoB/c9cPzDhrEMt2inISD7QxDqlulo38b21wT7d3S
AWQQPE6XPKExLsvRRmEt/FjlahvQ/oRFMrH6t0qpNSOJsdyxjNf9cNuOWCcqNUYE
Gpu3p/b9/lmi0AaWyUo1+O/ThY94afs5zfK9o4QNQsHE8iGrMiefEJ/HaLZ+pCod
wwj0Mj0Lya84XbZ77JYQd/5zRmDyKA3Ol0RtAqAM1pxMLvUuNU7+AHZVigcUVkDQ
WcsKCPMa1JBJIlgRuzVHkPlxpo2uMzlIQoqEBG2V088rUS4RQjO14vV826L/3153
AEfoJXG6dNJ9Qmd+JspOj9Ao5IQas9IloOo0myW7J4fehjSqKyTuHx2G+1KOJ0j1
Io9vjv0Tvcj4tzTOfPAOr5Ji2rpwmDSyfuKw8oF4SYGI9UbswX2eF7ZC8d77CDUH
HZJPzQTOUp06sRJa9S8171bzHIM1xu7c6qFwLIQfdktrTQRQySeSLKvbIRIMJ8Lh
Z1tmUiM8JReJF+GV8svEEgvRdBNFIR8I7BwQchzCrwTfuiKzB0C8qUmc3shpBJ2x
o1LfKrsLHPO5BuyrhIXT4l8mk5atGQVTn/jz9ZI/fq1aisIGl/QeJqJWcckL2nHf
h6hzGf69t1ycHM80toOrsPIfIAcsCNZRrvq6ckkCuQk/DPBX+kFeMGu3t9jsonBd
VbhWyQreszFzgFSTDAcKW1yulh8AWR8HaVCKa+edf9/NCIXpnlmiN9FeRNGlEp1a
QGOtbPy7MtwIfMLYPo1JH8I3JkwZ3U9DzMra/Wenf+tuKLdCtO4Vi996NpiSmIv8
Sz6D/w/2XlJImATroFvGMMlS45S4khaG3KuG63FYvvvHq+hlaTD3tt76pyiGMk5w
Mt0d21ER43lSa8Tk/GsJFcUcIYvy8zSeylLSSziIKvhG1MDqSj+O7VniZOrtNRnM
A7UC6N/m3Twq68cPKWiNuQ3chAaZL0JTuYVsbLBnJMQXxXVqfGykE+jh0fdN3SmP
nGhVkKqxIH6x0/6tK5TuaU/jyG15zEnna5PlIk7gdpLYWA/OyicbAKLOiu+DKB7F
N1Y2FVraYOlmRUh4bJ/S+//x0UsWDOSDxS8Xhhv5uWSamxFCuOHA7rxgXn8v+sDg
E2blzTmPqfIqg5dEURexxhHeNVNfZVay/pG/X9cxhxib8KOIRveLGBsTHmlbN0pE
M/mf67gdiSkDFxYVQ9GuQ5ScnVUlngMh7TzABHEAGtsavGk1WCt7I4wF2TjYoNI9
4AnMIJt3FwfbwnWHy3CNgL4ZQKFZPCwGueFmfLHCoQsKSTL7gBGraCogaBc1VKi1
7RXka4PTm463VzfrRMYcch9y50c6KBW5fIA4xBJBIIIFNukrazPXrViSIayM61DE
0+f2QoZHLHpSXnALXzrhAPa8sWWIUnm5Gp7pcCyCggZn3/bXfDcPrLmYYjB+aUQ8
ClHDD4mFRARYMUVW8HVw3BZ74XWeJRpKi3yWOz8DOkLW0aSpAeqHs/HVValsCIQN
xjIyB5/mZiTXDlpEvyqxUoSb5cIyQPeWtftQNvFt0Lvs/OHivF3nlrVno7NUB51e
RY3az7qTlM0zdJqeDLmBEW71WkpT65dLfshl2GkqFRoeuzEDJ0cRLlZCZoXUn0gk
6i9qH3KLoNga7Niqr2ikNNiK551hI/f+qxQs57az0aEgS2zJSci7i5HDWLUAyCnO
GAW1Dno1BiXttgkft2Gtvs2RorL3rXQcxmt+FvatdC0MUp/vLjIqoSn1isIEbM28
o0m4+dFTA9sZciCfi9M0IRxkQ7EA90pHD38TENNN6arWuO7mT7GEjw/KKrV6hvn7
k9RgLyR3rYQQQDWKMRQfguTEZ29iZCqvUGYisgfWXzYx1rPSCs5RoG3gL7TqLAkj
jug81cZNDskp9WP1mmuIuFAwjQU30VIfmM+Rq69oSVc1FVhV+i3ILCdGhh2YLBot
eHtsZG1agpi4sbjzrEe+G4R8qtWg72tX3H+42iqHntkGvAVjQVUpisi+VFhUmVla
3jBJTewnGlvolptegk20kLmQqY6KQeXV17hy5bfmPrtm7cj6erNUDWOHx9YOVrt9
06j5x6VSjQnxd6sWdOGhdVKXemuDYwa/v9MV2yM8iN9JKHobX37w2r62xiP/HkW8
c/WlUolQOpywEYsE5ATX7sbPV5RQGqOHO7C60DgpOpFjO4fqWcjRGM00y/zeOuLE
aQh4d+Wp5mvGj7IMDYIZb4n4sHAx+xwUk1I0y4WgIkkXFS9ly0yYuYd9VEjFD/hS
fPW8VZVI4icZxurom2z755r6HE+5RzsriR7Nv3FgJYKR5e6yCTqPQ5iBNxxILCT1
eoDMbm6HM1UmRjR5lG88GJZ7XZFXz9jyxL3RjD9b60PEsT6g76vURN6Ek3E3kx2T
ZeQQdjOfUKYGLOj0wfn1yUzYok+9h9YEW8cCl3Hb6guKlXJ9SmFDUSBSaKITpNe2
Qf3AcCCR0pk3Pie9oFxT/AumIvjY72fIG61i9XLPb3lQMzZccMUjglJSzmnfP3Tq
HdOE0RW+m9ThS4HVTAyqQZCvYxaoucxzWsJrZYNAO9f+Vxakcbq50o0giyoW4Wy5
K6mSjj0IWifGKLm5wlu2AX/AyMTtiSl6gZUUO/kOJbts3SGDy+W61RnicDvyJiw3
okwysTNnJH7LGq9k9IrHNoOhptOWq93ZVnSeOqmzQg6kOtrzScw/kxk7IbQKxa+J
0qfvCAyfB1bPiCTjwZCtIOQZ55Dyc15kOvQlQHnaHnPOETMb4VHRtS+5vmnV0o/L
OFjuJTz7U1StmyqD5sv6fVoBioyVRplS0xA/R9cjM6JeDJfSUk/AIPMVvG+I56ZJ
BxsZgFIQJmY6NArFjU34uPVhXmdyjneCtxkO+Nwr0vau8LDReXmwx2efFKAzXxyt
gvEUMQAMU/AXG4/+V1i+DyiPONVbOkX4HDYedzZrDTdsXK3RlkfgfC2cWnSkRLsB
AWsaFG/HCdf3OsNawWKkItejC9XSX8JzAOYxUe3q/VbxOB5ZBGHYhlUZLwxMKV1G
14UI9a/itjbWhXD5xaeK3tW0Q8k4F77USdVNaUlpiGmQSXTPkgOT3kCVMKPsr81O
9lhOXTHcxYoRHEUDBt9lbEH/ktXn/u40nr/ptJQUfhK1xtyVEE1Wxpp1P1dt1fEU
LMKVPVlXBnpwQTr1duU52HtMoSK+RICEXex8/5ARl5L8c/9FLhcTGP7vCv+WGHF0
C0hjtFkgeW5sfAtetzQWEdi+oPbKiPSV5rZTUVqSZ3qZ8NuyiMfCqt3Fh+NwZqmM
TBl8Enb6i8gruRnlq8lkGkVrnfVruw/oh9hkLpK41ai2xQ3j4kkp/7khyLP2UheM
ggLKuyU9yijXnCImm1wP+Bho6Z4UdB3UQN9NeUgp3EnNs9gZ1C90Uno5Lut8yUUe
8/pOrv2JMwN3pFLBtqQzbIH6fLfR/WWA5ZLykd4uo5/eCTWyugABT7XbyHLuTX56
AfFsBo+hZajvSEx/EDMugFoVWmzXvQTvD02Q1Dsnpfz0Wk6Szqq/M3p5GO2pcdVO
UJP/KW1QvyX2Lf608Ov64qwmVVeh6JCzPJZggonucmP0a88mSxaV0hTtXwCTf3Qt
EAHDX8fo7n5YjcLIUyNsLrYOSX63lp+ProExgmonV4MNoGN0w2XGLa/KnugucECu
kMVHCjo6ggWj9d3hxZO/8t9JZ7gr0wIsZkg1XhAvyAeOlTED/X5WbOQ8X9HSi8Cl
vox1NRtHQRZBZL6NkOCylxEoe7O+aRmJfcLlUoBKVbP792oOh7DspeBPh+8zKbEb
YujmwLd/bySIdzwv7kYdegfZ2XPLx82oAciKndNQmExw3GB1fcyrtVG5KBKAghKw
hUCelywIfXZfc/CjUCRMRTUMPbPy3KhlQ8x0gaFZaCZ2Tbni/kcuxNxMRskj6fg7
fRWrcEoT5tJ+/lRQbb+eNpilr5IvsdYaP9xnqcaqHi6OzAHEXPpnTG5xI3Y+hgS7
Y8JUCN9vRffh1+AunB4dR1eq3yR/bo6B6KV+kIp2b5DDKOGWRTvhxGyhqP7WCaaD
Cz+hpRlyquFGHl1cJwO8WXH8ygJ2NDKMnNytbV/Yddj5V2THI3BpQMVYBSTDlLC2
y2EOlMTb9QMaGbs2vkheYF93QzBACuaEqo1NtcP07F6uXof5FAd2cclUOLrDSFfW
ZSk5sJ7bmncvxHHHqGCSi949FYzhNE/DJWoa2b8r0MK5CfmE+Oqs8RjEpi+V33k+
5KRQPuz24Vtl9tSGTwOD4VvDFSR+vvzB72Wml3y7hTAIQFdFWIGCpbxOM4hdRaJV
07kLuiG++P6AHtRoaW9FQinVyqZsvc4vNVpJ6c5ApvBJXNJcrV1YgnR8O3o8ZBRK
KEkxZwGS1/yM96r/VqgK1AX7TL/X/Xp71QYLbQDTV3zlnubgJf83x5BJL51xcd64
cPoKeApWJYX4d4sz2rtMYJQtHYYWUilt4MRy1XEIR78TpvBD+PJX1eB7dO97mV07
+GD32UB+FWTZ5tP88bQqg5K/sLe7DzO118lKN4iSSt7Jr0O0IMSg8lpt9RDU6l0d
H+4uVc4pykb0g2V2wO8jCDSxbUvlrMHlvtgrWhqtyxRaBuRFMqOfDbL1cxMVQit7
k7HgwXjf4bPzzbbJ9KLl1VsO7Lo2jRjneL9mx/Ee3EQ8Mo2TQVx/hsmrxxKwWTtk
F0g0+2CWKwLArRJlDkcYYsOYkYwUOZC4hd//6C2RqrLmcjZVZwAApCgmIV13GEuK
lMM+sDqgPcPbJE2OvRsZtp9KTRfEFowPFwdDpc3+9S/MJqD8b2meEMsJH8muKQ+L
7PHNORBGp4pBC6+KhTxFNphSoipUkmU7IdCO7GmCmvK7/EQrnw+X9kiFyfArZvty
YyNISkp15dsxAz+XoSw3TkJ/gT3UD9BZOFPcTAAIQaErh01J6nEqZFhd9oPk5pe7
2OLBgILvPL3ltXu96c9woYhTD/4wmWYIuyVoEQu1+EZasEXCh8ERwB4F5NcQAVxE
VEV9Sf/akXl9DYy7GVLkVTQGdBkk2e48rydLBzmPP1AzlUOWpN832wJP5vTmF99f
T2joDC2OoOSpr9GgtH/8BIOxTxvYkz+qNsdNy/P94cJ2XhGhPa62sdw4U/dsYsj1
XEoNQ6Pyu2eIGK7Ibmf63v3D9w8LhjuQLegLgvLznXe4lrOqE8q/xWmzYF1w6FIh
py4h1FOv30c9PVZ8DnxV85ZFeJV9WjARLezUJmEZvIlF03XbQf0EGkpb9ELZuMzg
JfX1phVqUR5dSbEQyHgl90f8AMjZEEQuczuITuw1ISuKPbz1d0iC8PXgJHXlb83g
7IezUcp9gsJ3x2v7DjCu9sFc4x90dnfzsBmyrbePxiHAYJ3hWqdcE9THW6JDCKgz
qFXmkz4NndGtaUY93IDkIHRuSsVjxAEu6pjMl5UcF6T0ajea/oQxr2MXalupJ+Y4
WzMCFuHGqT19aRnguRC44V4ino2pkY8IiPCyxnSdW+AshKy+dyRGRNhSQ/16YbDj
0b1fbtcL2Qum8ojcPkfElJ+pmWoYgEdpaINHmPTALHeAiM6XnhSUDlqRIkkmCtDx
3skR06fqQewv79CHvpIDS0A1j2AGzpwt8AJF0ssnM/9TVSJB33z73kuiVXQugq2B
Pli/bwAx6YKnYI9MEmT3BL/cgl9xOfInb894JMCp42Hcq7ZzxlPazFJuh40q+9Tr
g9HLJhF7RWWha8GPqKE9oRhTnhLOyaHs9UeLEndEdpb7Du4g967KR43beoCfdurZ
VOxFvHYhKS0zkZexvUTyRcXPm9zv7JYHAYsP9q8DPKa/yMFz8sCf2LFLoaLTjMC0
4Py2cy28kH0Wnsw8K89Q2RTVS12CuizQrUJZ7K0wP6t8qzjHZLk4Pn5002YOkFzm
Qyofk78jplzlR6VQ7FcH/SfIA/u6dW2V7fu/7nMzZufnH72ymzk/khAp0f+BGdiI
UNj3PlFzTZlRlYAhYyf6cMBmn0PpcIljdwk3hhbqgNeZ1RjooOYKRdyKhvza8qOn
CLXHO7hZPxkkdSoSUoYMb8cdNj2plEakjhKoOVKq4tR+qg1ICfPlyhLwMtmXvDso
6H3Oz0H+pw6UfEMzjph7TGBfXHK42A7R8gFmWE79Mc/6IK9rObZ44G8gqkH9Hrkc
h+7E5rOiUOdusFhapxXcrMzilm2FqWDs9g4w9zmzOvlcPyGvlnyo+oe/DnBDzrxv
19DDLDBuis4eyLcrA28snoxEetI9MCLq5sN52mUAUHx5gJFITW2UiVQWw9NschkA
xykwG9R1+aPEjpg1J00GIhXes72krkEbBX8iVa4/4haq8puDkG++r+Ad0IzTzlsr
kKCObZSUTN1Z0uVnIGDOrJTtXYMBS9IxSj99iwBoRLT0S8MOdU11HkfLeDrW+qjk
9qQ8STz0BxkPfJ9VLSb8U+Z9u6MXPjJ81mRfW8qQ4gXX07ryECknpdWPbUF03ety
ulHh5gJxP8jNlHtpdJAZmInMCKdeXkVli6WJMGg0jjyAGL9sHp9Es3Tk6uOLy3Qo
DcUBFRjqzFpO6KxRjBOqZsF2xLd0KTl0rXa/CyUxoVF8CUcxFlv8l2mJh1jBDvEU
fYtAcxVFD5WoS50yBQQw9c0sjLx1TprsmKlK+0elbCqiOa6WQNAv6Q9P3F3QXzVO
Zf0fhTqW+84fUMdip4jY2sjtjjC95OTwxUJSBtwlR9MuEb2Bad4mtQbWTCagZ60Y
UWaMgJvDpI9g1ml4ZnuG1y8d+ph+TGgeDIZYjcXwxonDpXnxL/4KWPgzJUXBnJhK
hbfgdtHhSZrLj29EtisnKIyWVUEHEl7slfZh3O1PMuj5CdM9VtQKselXJk/gfCjh
0zKkw8B31h/lWw1XS2RcbMwWVQhQK5k7ddqVUeb51QMFtZCOpbFD7CDv4/+5PsvU
r0ERcQKPboDHAV6j2PE69/i33YzLum1NQz2WVTO+Yo7XpD77XRNSMemTukiNRPfk
f5nlslEejaMsEe4FZa8b8XGiUrqad+PcCIgQQP3XwjK55yKRDcm5TFll73W+13Kl
b/qctjAhzkLpChQ3Hxyw2R8u/qA9VrBiEowtBn6ZW67YAfW8c6ZwZNgUwnqfdBCB
ne8GiuyeOdo1ZQ6toGZDZePIj4z6hRQ8Op4ZC3gL84DsxXVu4LKLjTAwfihs2eGd
Pn5barMlM+WReEjldVJjxkOxzVuqGXEilAxWMR9Wy5AH3gv2JE4cfXxdoHF8XsVH
2ne1UgyNzB+KP9MhIv2raCFA/fDQ7wNvavyRNia7y7EIqjECu2M0QUXYl2hIwMQh
niG4wK06DzUsiXKbXzNEH3/lPoYywFLE0SgiqRU4WTgjDRzE/zfw3Y++xCzclPdg
zJB7lk+cyaJZ6lzWjp34Oe29ETt/blRWOjF1hfOToOqIvGvJdJtpDuVUJTLkJVun
5DsU/Ote7jEj9PttWSxp/lA48leQSIMaN8ggWDUs8QiG+v0pi3YwvSiwWAJDnZLi
djhdcM5JJQOnpYw1CpekaNGmPBNCcC/i8bJ1Uzr3kUqgFYkgRMOKwrxQ0wP5P4uu
jF6PABpSzeNpdhnsK/gSghrZ+ltZ2kjNMAk7POeNIo75v+VreCbf80h+KnLEGHF5
e6tBPe6bbVozu+hddHKq7uxrAJL6GwBBzE8zpYWJbg0j9Yo3z7q3HjnjL5++nOf0
48DO6Ns8ZuoZAhhy6+BIC4kRR8OgP5w+zSvxNIfLJfN+kGU+uHLtL3haXUvkB9Js
xdBQGLJRBzhkACf3e+Pm3o/+qqtP/Gpsd3QRsOjxr51grz7LMltdlHKBTs5M6MGG
45DZlRP+5FmzLk/AJzVfvqox6uwoHH+IyIeAT7rEEQyggn6GNByE+UfBYlZn+YPx
TDfps46MFci02aaLqkPccUBQEIEQPx5QrW/ZrjYTL83Qx+G4GNfMNYf8efGR6FW3
xcVRxdjt1uv60rtSEs89DviAQbRrEBO60JY51RNfkoT3HyNl3dNY0uoFRAYudRb9
zn3fu01Us5Lf2LXeymVL9dcXfw692nIA+4B0eXoPczY3kuc+eUFBFKkhjGKN57ss
VVCKQ/+Qp2SGYZ9SxOSp6VNppDobeSMNXXyy+nOEIjoR8VswxSkUtDLf0whg3oYI
rGKvtyCFXpgb/FR3in6MZWgWEAM05oZPOSKrn51Eo3VALuaG73Iz5LxTp+qDNckJ
MSynuKWNh6XQryb9wtvBnfWjUlU63XovV//UX3wkPHB1XZP1inhfVu722hOoWgB3
VU/NmeoftT1RviqW2N1xnG03At2UPH7I+FHJYUn0vwUJ5NbTPkQ+t/MEHUOe050r
d9HCmzxKmMi3wkMTVGjhmA/SYqrlZcA0YPE/VvfP5EWyASe37vB5iMxXJGJ3rWkg
1N8lOPamxa3KVO5TLIBgFVHMYmXFjB6jDzWqxmWTWSncIfMQkYYE4wVgQ9jumjMI
LbGdhIvIDBokwAGUlAu7qkOg13vpWoH1gS48DlVyDVKgnxMYreZ8Ssh/Og5IF8gE
V9ESvg3YIzwVrlagTBvIE1h6FteW9F7aG3k1Xk0sOlWMOZoX9xu3uvkvPjbqV9WU
5K+bDp3hW5T6TAE+T9mSMNprdnT6QDERlxsIs17zQyeZfTDMRbmdNowb0UcW0K8o
AeeHrNUokkXRBnJXlcQVwmSlpt38QRUy2f3MxPB6okIGQQYntcMpuj2SPH6Mo4xC
9PU9/XARKTV+BHJsUrdGCpU4Oc8FYPCS/2Y0MWX/+ixRu1Kx4gz/L8y4fiGvU8IX
/g8kEUSpCmI1Y0avhtDBGEuJOlupdoqaVSVD0UFZRk3dv4XCy97w9i1xUydWYBJ4
ho9kKI8WbXSljNzglL9u4ZoAI+DI8LzVXwfwu6NB1L+6tQtXruuDxR4E52P4A8OC
f3kD3aUOKqCPWC+sfys3wAxVc08infv9ie9vbqcu9qKDoTKnzjK86En913Y/GUrv
0OpbgmXItjQY0X5l3h8eJ6uS8Dbnu3onCbxCPWv4UFDI2qqITDNZjXPN7BVbvfBJ
39MO2rGI7GdcYAfFgdfMLg0C3qMtEJwpJ6iyfe9cw8qMU2D6aFmVhYBlTCe0bQ2o
nexhvO1BfZje8Pg5zEu/OgxhSRX2kDR/TgPtz/YUQXcDv37ypiongAuhcfzASpnq
c1/5Fw0y7ZVk2+UStTsHIKGW16LkT7gXE/h47WtP06QC5E9o9pplhb37J3Z49a5t
daFQ6gcbDsE2a2OLABX6BKaxQ4/kct8ufly1pdp+czgEi4vkJFi/iVvr2ljB+Q63
my20Mn72bihFzZNxAUcjJ/QqqaHjNosOfYDMYBCCJyVWDFzzVXZItZzD4nt5YdEP
JvGzJyZIaotxI1/z6YpHMca3CZ14l4fPoOA2g8p2JVgfXjhDuMa0ysMHHfbbgjey
5cg8DYqqLjWSeaR5cJ8j6E6I1gfO069DcDAvMbnIr8XnjJNWVhhD404yXq1Z4ztj
XYaFk80w7BOQQg0jrWhrF45M6yNUibNlFfjomlc7WyU1FcMDcIgwpNC88YCd4uoq
da9AIsqVkZwWt1EobRTSRu8o+LrRiEoqY67E+VXlrOmlEBJyZSIPOtpwtzV8Ncr5
sSoZqjkbyFdClT8N3nzeT3rURUhX+YVZZet2AnNa+EAedLprZZbXi1Ytjvbj7udN
HJ+XpfKptKIckcHbXkJmEW7qV/7UwvVI+tDh2I55jgMhMFVucdbcNNkpuJCnL5jm
tG0b1eU/xRjpUefPuGXpw/M03oVm9KNtzinA++J+1dRAQnHNhF49zaVjbsCcmyRm
/mE9iY39ASSzf2yPaNbDi4Y4aPVBZcwz7XEQhImWAYmMnrC8ubMyZKb7fNzKJ+NT
X9v6Q6F2SFiIWqE9GvTpYrUwzQ57Ie9hZmvnU8ltM6Mp1UtORkAxbiCnrLmmjFbd
J/DDLfSvqR2g2L93gxfIsM6ZearSKN5jhqI2Ys2IHj3ZxqOEY22ztqqPBuZruLnC
h3qtLn1fjVP8lP54fvH+KJ3Oi0Xxyt/lidplMgkw7cHcPxclkIxSvkmw5C3PvDwm
eAaHCZZMLHTx6/u6hSlS5Tja3DUDNhO6uScnlr+CiXEfwv7x/SzDw3ZRNonZm4Ki
o477PR/rJC/7Dy/yHp8WAdSxlbp+9d5ow/BtkVgZcLPsN4KXvPSnOQfasHZ8L1bl
0anr9aUk8IKnG0RWSxgW3vrwOSjAD/nTzGEb+26/5YFi8SQ9lCXYSKipohvzj2wi
UkYmwk20GxmaUekXJCIoxGpiMrc4OvLb3ZxX9PQc6aow8RlKwLCCEZ4W/graf+98
//o5Ns3hMCMUqe5wRTWuw3kE9eg43pybAH6c9XW3ttGjPLXkM9+iCfCW6s6qdOmB
6frS9UwwcOVY+AL18z6OZEuFSlo/QTRRV9aPKeH3+McufqO0kwz86qo+vzCnyjR2
sh9B/O3yf9HXMb4OzayAyFgtiJMfBVcPy4y7l3fOid4tzVZPs7IW2q8D+gwGxRRn
DAiwtNCcV3DZyzQfnrd3C7tK5wAr3c2colTEzpaWKNXHNQgEv/uhK0w+IhZ/ZhDB
TLvr9yuna0TG+J6J+Th7Jiba8P5Ry16LJ8xTa8ObvpT8LDdzxQ1AL4Ek3FJuASJg
5Rxn6rL2kT6hz+PnABDDx4mXVwKalgRpvVf8jh2jcqB0WWMwe8djWKHFFXcoEvPz
U6rIBvErTjxIpxFI6HROfK/OrWtFMuJ9RxAE5mTYB1oadmMhLavtsJb0QBRUNmAd
Yf2tpQMyAoP7PgnshqaUKbJYXo4N0++LtODxWomCWTU0Jg3FWsIfv5G1VpAklrjp
T2+sZRBMukjK1s4ADzy/SZaV0zdsZG6oDCIw7yWH2oJFmPQZlJnRSY5VjIz++KLE
1e2xb9e1AlMVOudEzPgJrMId762Rb37Z9gzzJs+dF3AE4LdDj7GO0WHkKEi2RhQ6
4T21Bd+pXKIkGqB9fNS7YI2a0ypIFFPzZbM91U4YtBPwU8y11LWEJyNDEBmzoeGT
f6brDJgYIUy9u8pmKJ3yzn/XVwaWubEH/4kvznMyOAai/xydPUtSmHR3ajcXAFQH
B8QNz/F4XM9oyIZwjKlGS2EnkSR2QAs6CyR9sqiygDMSBfZjBhlpF2vizpynLf+V
cm82BqaYJAw9Vc6PQpNLB7VezRMMajKM3U2Q1CUUTeBGzdr1Ee1uhz9tRFPYu8o9
NUaFs8n35Huaws++lUKxGkLGnTEKCYqir0JudxifTRTbJNEiJhLTZab6o5lQZopk
eksWi5WXJQy8DnZAyZbfnndH1rf2uEjGGEUBVU51o/3uPWD48eopg7JBUmPlxKDK
q9b6xRBtDspBMwFO8Xc9cBcCAU0styvs/DI86x0Zz7y+Qh+NL8l+OyzwVaHEKXm2
6Qzc/d9xXvdBf4kdCVIGxge4IQDXDPu2KouE5Gbwb8zDpXtnOufM+YIMgruuLf68
1NRydTYLB/ZUcda2V4R3saFG4GNef/KLV5axpEe8CrR6dW3Hax2iccK1aqdlDvcp
b2RqzNhlYBFT6mtybSnofaXK/PZm3xQRAjF7eaoKours305s6MbQkE6zsWtb2hCx
Vpna7WW1njdeRnF4ZNKzDddBdqWpqiIqjQFZdKE+mmstLgZPel9VilUY+wrvu5BU
I/Vreeivmyo/c4GAyY3IGTCKyFKiHtWKv9i6ouQNkf2051TYXxtYgezTUWW8JLmX
W3TgrOUpP599IYbMIhokoQU9MtHTkEG/KPc1fdNKCTLPcfW3DYiheMigsfm/olNC
pQCZ7jrqI8hgy36FT0Ioq+1qHMPc53a3GZHpP6CccTgnEeJsZf7yzmE+9OwHvj8c
aSVA71nGhQljaDx59gJEkQ/c5Eo3IXGQS+N8KdPtvrfPw+064EKq6A8XFtVffRYL
j5GWwRWW71FJpelB3bqbG2xa4od7n5BPk2zEynFdX22aTzms9VY/HGtzBvERkbzX
ekmldaE+OMQFfqh2xIAf5DIaUvbq6OLNtL/y77tvjoGbzqTa3gWnq+vwK3O7JNcD
RzOYe8dXgloeNFDXp9HrR7nyhX4YQ2MmpxRd92Yd/+T65w1rL7NsA5H3UxINs261
WuxJnRKBW7LUyKn/kIuGAhJRzVHTXH+YlUWicHoY70UgZm+6yehwz/RxiNe9+V8b
3sqcT8wv2OUuyXh44NDnutJvWIvU0cHpfrqQYl70H6ry0NcC2KcKSRZV+mUbYm4O
WKXSUWFK3jVRY2oGrx57XROsBNks8evCijrg2NBAxLpORrcqzIeuWisjrEaTaHSb
r/bM2OthGSFN/asudnY9THtsKk3xhimS8f7xU9eaqaJvLn2pj5ShKEFWaYuiqXL0
2YaoUOzQ9CsyDZHxym/ZpHpnzFrRm1xKatTp65lUuQIz/xVair2/RBAasAXwjcZ6
eweGlpD/yK8BF5rGR+7i1E16x33L1KgKir7l3tWe6RxcnDFX6Ds18KOmaD+F8JV8
ilkWzv8sS33mXj5We6gFWZvdqeBZDZhz5Sbce8gMtVWPbpstaVn7NvqQk8XsQ22G
vBnqf/uarqA0oKPydKJVlTceOJulqo2/QtOOAk+vR5lT5s8No+9I/du7vzloxab7
Rcbmp7ilcW1jFB24r2Xj1GP5vAOOj7gXdgiezCRhryc0OOKAEKpXY9o2CPZ2kazg
rwj6lpE8nUTg634aF9UGJzauuCUqSVVowznMeiP/tJUFXiZWUMUlQhIrVQm976wL
EwFC4plNoN5viNyqWs1caLSpsmPcoOZr6dzo7msac/zFAJ2qLpuMSD0vk9bHItYV
w3rizQmuSVBciwSh0Y1yHd8LA+xAxwMX/vqWGX7jwrswrUHHTOBBLWCfgYj9XoAF
keBYMDpAvyCAVd/hbME46BFptLY7EQC0cmKWtu9PDo52zQawjBxLp4hKqsph8Cwq
Zh8xmhRk2FG5LZshLDBkYEQRoGEwRUIgZEOlkkg+3UiqGwQHzX88EJFXhWcPvaXo
YxYHWyu7pyYQ3xWYkaOHwMbVuPV+iKtRbHMCbgpw53h+us/qI5Y5sIEm/9vugN8D
8SaXbVc+orF1Zuul+BJLOSAAQI5aWN/Nv7Lw92KwmszUHtd5Sw8cMejeENu/LQVx
WPCnfjJ6Awk26RWIpP9OlYo81l4i3Nj1UPSFLbdbdQdbuf2vsd9YOmONGVxkDEJH
wMuOLM9tCfW+Owkrb+IsJEhmRVv7PByUkTadOVA7IpiabpHMv1l/FwPw1K2+YiC1
+cfDTk/ybF+ne5m5TclVxxhGNmoheq9wsmcr9TVie1XNZb3u5qCTkkQYiDvTq+iP
Zu8Dtsjl+mvwJjN52p1ykzeqtMvFB9WrfEujt84SM3wufOPIzgi//fZsW4hVplp1
4u/67YHbbCoNcSna+w71pTAQrRMxdx7jdCk6q3VtSoiixUB+9WwyqAEpTlTO4WVw
+Fq+OvgaPtNavpiLvp5D+wTM6t96yqg0zBLinnw12E6xnLZhzHc4v89zOWrKfKAJ
C2zzxgMdj6vJJJ6+OkHIYzaYaO3bqKvnXUFDeMEUnpD8UPJBIsxWIofRC2Gw+Pe/
I077skRx1rmZok9sJBtn3nt/kndPohWW4m3ZgtUCCCybjZhVvecxF61q9nsWcyTv
UyAP75we/zGY+RckvynqpyxwAd+Ld3lUUG5fjB7iM/0xEWVF+DeSgh+pqFSQ+n+A
+B26czx4jEUzW/4ucdwladip5AD/A3A6/UMf+2MwDUSYtZnbmtIujsO2bs+cyG8a
Fq3YradqvTAtODJfQB6fbKOQbZ4Dk0LbGfNaLK5WsOWv4uZTjUet5wXWypiFjGTQ
7oE6QhgvlVBOJu1YcCbsoRIyMt2cGQqvdjv3OzzsqJ+1hHZVwkVycFEq06OGLNHm
vuC8Xb34ayD72ZJgb9lDa76pX2PZW4K8oRttbb03uUjRpA2DHnygJgoPBKDG/oCe
pswsBpuddMJsxuQ00TxS20xzIWy0jeH32Vwgs+CfxQMzX3Lr0IHdWpoi3IsFvgRe
5gK1PjNIKv/xfWxYlx6NTHXlQFDgkj82ceMuD8CQ2Y8q8lveQeAg5h6CVkE4aQQs
57bdkizxByK3vc2Pf0Q75EiVJhi/7SssboTBy83VSd1B+Zk6fzHO9CJDQYSsVcBz
e8GO5wKvHaPXEMXKSljK1F48O3gh2mY2eG0NmTYi5cFn5CqeUl56xvOip/27BmFS
JkgqakVTrsEdEIUP5NnSG4G5qLot8R2GuSPrJ8Bvg1/B0KdMptyHZjF8mrK7jAMb
FAx7Y8Rr/EBtmZSUQBOZ+696SPsFKr+zkMOhMfJCmOFYlrlplUqN0iuoGR1T4RkB
3s+eCxiF/+WMHVTzy4+dxmzxiVkiRpaTXTRcqMw397E17rbzrPKdj/nqLgPjWEQo
5MMBmMiVwsn5uyP9tQKMXqvIaMeF8byC4sZxINJSEebVE/mdI2s/4+WcY2BLBslz
ovLPSq9R/XfuQI5A0VzrRZeMKUaiBIwKBpwcmbBsAQEOoBVyP92cSVAIoorxOYFa
faEM+k9tQjBLUXve7y5vNE45u4hi9wemnL2W9FNoxoBI6pLfZDrhh6PfUVuoPCKs
jToZmUaE4n/Ff5jl5itU/eK1AArH7gYy/VOtxw21YcfNIZo3seNdeEQpDjcTrt4m
VlUoAW9EEV81l/iuywkhkTtQ3av/W1yF+4e2pCEpWAAXbeQxbJ5nqbfFDcsEUbvJ
RMnxhDMjFXgzSgjTWnYawhGFT5y5pfw/cyCGn9AgReGswvWZr6Rtt635mhzW6G5z
gwwRaSRphul8/7iGNn0Qdu2X1HRPAgup+6xwmRFc9lzN0bXiWroI98Z3hdxQUTCb
PscDoL/qbCsufH/tEd2tl8JpDeucUAE2uX4oNdVeRJT1qp9VUWPHs2Py4huVmNIU
gAsS4vykpnkqpxer79O/50EeFLnIH/idPkF9l7kXz3OQU0LK9pXQrG5kRstquktB
eMyp0NWLaKr23kjWzeJAKrIUdemirBGNvddOO2IcPofrYjH/WzaoAQziaqBAinIh
XtjBDazBMq1GbtR2sJ1gCklD43RImaJQrJkO/Zu+fvvDA+u0jACCLuc0V4Rp3kVk
iEyvKU228jCnDaCtBquELskqtdMj1XDx38FiLkVfNRIrfuvLroCVTzNtvfWJKpQ+
alQwjDFT/Q6Ym8kmNsSPcepIT68wC8OZsdXWf4bLRBewZW+DKOJTsSsY3LQcL3zZ
TqBNf6frob7iC7XfIuTTOu8tlDspsQFRV+y5fwy8Dme1nsXSWRfXDm0EUcuOFNJp
c82RPU6Ogibbr4r+gbCJY/UAGPrdF9NJmEwRmbsN7+CE0IMnmghwGAb40jbPNe3L
0LF5Jt0VKJxvkzefay5RZRvcRZv6kFBZRP9MYpK8qdUqrrXpvURnHFFjMZCVODXv
wBpadiCkxxVhUx7f2wo6X8ydOfczsbNKr6OJszZMxi5k0srb+Y3/4E6a/ry3/Ci/
3hwARKumP5bS1w9Ug/sBOzU7BLkwHvYRmZWEv0x6Vb5eIVbewFPWcpIFaZDA5m63
hDnP40or1qIoIwqJpLwVAq7jfrOOWksP4h+ciJrgeEiR6HY1t4/IUIRSuldZSlKx
y7xA3S216iLJZINcBZAljikerfY+GaOpyA21JCdSxPNS3YghLj/L4+lStYmfxnzn
h0TqLiLZsJ9v7O4dwEzNmyxGGgi2tingZb4wKqIpF19AFX5Vcc2IZJKHiYUBt/Ic
CqkbqA0fcegLesTF6W90mOj05eVzUxNFKAkv7IPa1w3rMENc2SGHKL8K4ntzVziG
kBmOlHFUmIYfsf/a4weUl/ZPY9JPxuMMDSNzRboj1hbSMmejMj0bEQAYivY7Wmxx
eukxsLlmaOI1KkTme2yQNWTte0mrRFpaBANtD+vEP7/W+M4B5DZebm6qSfln4Pr2
VTFgqmJTFZlPM3EU0uG8bARBktRFOK5EpobRD7rJLcq2R5VPefzTL9scLlAAyDKr
5FzkriOPHTla7B5tVdZuBQ3Ruf/r9k02GjHOZX5BVY65NDaeVxwL8wa+Kqjx6oFE
Gp8aKZSjokw+Dc3NJJTpc/GKR8UBV/fWFdvGdDgg1lRJsrQN154cz2GHxRUOV0r8
XdnxjdhUm3Z1DI4SUhYVbNj92GPbiRxu5dDZU2ELipZcy+BTZ73G1HVIER0hWIAS
G0f0dtJ5DoAZUal8xop8VklS2qFTqmPhw9qwkW9DknrzRmnslXIZOt9jOdFPYFGM
9uRiKooj9oiDel+JS5b+lveL7AnDCPVmRegxdWiBmzO16arQiK1lFISLCQeWatVZ
Cg3Mb18R9KTtSzEA8BErqy/sxDs7GY4eAG3zcDD6nhb8aVzYLglqHEgqwHNIMgFV
IwVJrBMe3Ce8AZa89C9w5hjJr5KKdQ5UtLxZRVxugUcjarP/NVi8OS/YxxmiiVm4
hyQbhRdNS7nQVrZYX6jeh6f57VGTiveH5vDPxV9VxT27J6oqGgW4aMdPCYma02bH
+ast9gQS5/Q0fTbGhwYmrtLEtPOJF7iPO7Of7EPPCTVhIHKo8+d1F+Ec3CptjY4Y
ogvihhc4lYO71n+eDDV4nwryxoi3Z+Xpv1Oe8Aia3pCmY/v7Uxm1iq6nPP1hGWe3
HJ0XYrbPhtYBYOofc6Hy4yTIHIBgKFmKsDUZ5tCFUNu5s1DzarqdolNfWFf30lXK
4VblBSU0TeHj55emxTyifKMHM7Bz3AQv6EZGbgxYHoEGoYtYuGZZOfLVHCDKbSnF
m8pSAL4IxR51XbPO86zcgEHA9WQT8qyCKR3wppZDr4zqIlDZsAScvS9O8MSdw28g
tY2XVL5PHmS8/yq5CZOpwWbI2u+wfCmLTS8QrcWhF1OO2igwvtanj4PS1fVYXUWw
n2aLVasmc+TQVMjJsbf1fJo9chxbOcBNd8L/mGEX9fVoUnbmTo6yaJMdFGRjSRjz
oT9U5mzyBDsNVyLEdshXehPiJxnRTn+bi4KX2/UI9G1ZV2kv8wT3cdwPtQgLX5nY
6bYjzxs5yQUvmXjL6Br8zyCKEJI1QQbaXzkOAPTRe23MeqT+T8/SuBcx4Sxmb7a8
0RHoixUU6azhpeSSjtvB7DLzWD/jOO8t1x55SNi4NemZWU2UkuAOiPETHHFcstI6
y3CHx5WHmBQd3irYxEwuA5iA4sZv5s0bSAgT5kpB92Srb45uBgogP7ouSGiVXVYA
gZGI+4nlE8Fpos8MMAT67z9T4oG6PPe/6SuSoiVrqfnyZRVpmVhdkFFxfVO4vNbb
PF7I3Z5+Hzduq7LRYuSMFnaL9a6hd4giNJ27UHSHOXiy4N6JDavP0XpQr3VSdhHp
uijAgjl4EZaVZm3ARNFcJALj9MDd0yJUbDRsDBewJ2yF2GDkdSIjTSvmpym4XZJ/
mDQxZSpp2ujnwFZ+8SBULuf6S7ts2USOHm/s1m4W/bvnheP0no3PhvVgm0HIj/Hz
LpTUi7UhaHNcqGtNA6Bk9Nj0KqjAzcCOB+zOIXfZe2WYsJHlLdsMUOuK43KYzfFD
Tc69aGKRpFIC247SHKGFnm//1gd9WieqDGFHxkMGBufTrHagls5QaHlImqMO8PAX
Hgcq4RHld8XS+3dzc6k4DeTjoF6oESKv8TQQgioIrTa3EGALaHIUp6xVCGq5FCF6
3Sg91cBl23GnQ9mSVxaWwZ7hR6vccPmeNUNqUGO5uW36BfMV+ghmMYJgAGZqjIe6
Q2WlzhUbcny/jyERIRqBjw4ce7/ALmV+ZByu27cWSqGeFicDfUun7I/6ulCIR7P3
EuY5KZ1nrcl8+aYulaMw2al/DsYRVGrbPdFZgz2WTau9kZoxGS9GXI5v0DaBXrvg
9ytseiq0rDT9JnGD9l6/ktA1WfJj2ySUew6vtyZzwdFmqcxISC/WemHiUayM7px2
2WK1NTIyK4UfCJeDrNbjSDbERcp8Ke42Zkt/0Hk9ODRAzHDtC+q9omr/d03f5cib
+h7vCM7SbCO5mDt8su+uN0xkupMlV6gXGrM10E1EBTIxlIJoU8BsoEAYSXj/ALAQ
nIBrgvnChgZJAeWRKHjA0GQz0kBDTXRWhrMxxX5B7fxnMJ5djwiDAPEdg1/RKJCI
hPQQM4dqLjw7xbALcKfC9wZug/qcaVc/oVdgJ+JL+IpZ4Sqt2mR/rq05T2TEjYTy
ihdR8kPK2hd/dD1DW1wDW1ifwCyvtpw/nWLDwLaxGL06uggAyKrOWyCdVseHraGb
8HIlZB6FqfQUYCR9wgmQXdAy2Nl6xNsU9QuBc3AYodJNix3kymstEd0DsxmQeQuO
hLCGR9rPTsHEfnCuV+WqseQbaz0ki0a8Wjck/xIkO3+tb3t04873GZ7GAVVIEVw8
6zq0/Ksd+IAhmhKsEgCDmZdSEgumkF6f2COlfvyTtWY1njMIFIKu1jwvhhVeZG8/
S8QALMMOPodigjEgC6JeeoW+jBQ4VSy8CCfXk94nbAP7l2CpB7izg78/wCcWQkLf
XzDWzkKpaz+VYVzsIoLjFMIl/4kqyBA4jcKpu3Bg+hRlwGHaxCi62iEK5jNwiTDx
LPsjMSoyRv2TZ5WpCAMCMwa5Oc0dybax0ozuZzHyKfn57w4hVdINm0HSEyiRL2sV
pCGw+TMq55/2xLRaSdn5hVbuX+IVjgnQEgHyfl3Ra1YGtpFJILCRU2CAJRNkAxb/
1AAImM5vreiQ5OlleVtbUU4qEkpGDXanWZMursc8qPB65J4o9KUUsmr+ySQFBxqG
zW184dX0rytPkplLlcuBInwpjghSAz6VZIEXteugoQCZiPeTPYQ6RCndSSPtIDFf
bijf/Oc5UylKl9Fo7HVTIyCVel30/VH7knZRVy0kiTGw2piVSpfxwoM9uz0pQ9rq
fqH/beCRRn//vn1W56JUvxZDVvbq5y/yMixSscK79yajTesXCtppyt5I9XDZ5D+u
d9lt3rXy9DKjSeIPPRwUzO47I74+lBiTtHZvh23N78EJyTOFEqXJ71JDYPGTQs3w
lq7YH9um3D6A9Wk1+xRiAaM0OQ2q08GeqUZsIyk3w5qU629y28BwScyLjfuVf8zW
74rxvQ0VpkVKxRvsdBZiihJpIDNwGo7W8HyPdfJnPPB09lsz6Y+BttukaWbyG8kk
67lqGljkTnwfrb4XogTSBtUa/sxq1CF+xG+uxWiUghJJPs5AueUF+eQkfEJnBOVm
km0epVCt07nsE0SrSuEebPzHWaPYL+8IOUKuz/KZhFWVTcg8d731xjXfKo3Zfima
S/e7vHAPcIGej3S5zls5VMnDxymknWX3mBjP4dPrLtYAphbmVC8ZEgU3NubxHy6h
qIUPM5/zbhHn4KlFd4jlR7mYLQPBw7DJ57rRNHuNgpf8uH6hyjGvQCrzm5NrXeNM
dvfy3+JWkZEgvdU+tlZyphhM9GcORQ1caKWOwHBTR9X52il3ui41V5/IDLlIH2QB
M/T45z4xQgjCxysslDT9dR1+/zHMITpfy6MVi+73ph33PISh7vh4X4W5kQJb6/6s
cfQUI76u41w2ZKYXmgKkn51gGVpvh96QFbd8Wk8F9UqNc+FTR/L8OU3cspeetKFB
1jKjQibvD7jtl2IaF6nGnUEfqS87ez6SX48lCETlvdJoeSa3YihUhFSOMRxqAsko
PngDksAduQsupMLitr4L+1UgtB9qIlKAofvA/UDCGTliAHpl/v+xOezLQrfIxGpP
Jsu7rvDy8SWNH0q7PmidHCjh30l846x3Hd+1Y754o8gvsPfyrC0ONTS3AEczEEMo
eqQ6VeQcaV+FamP/X38Qw+yWYRgvTWXiwKbzs9eO/0Bk7avxkaokCF1uPZOPIbW7
4wA2ZrGn7mZWtEl72fvy1V43Wwoy2n4jIIj0/QQKlVcHecXsI5T7HwfkKQf+Nkcz
7JUk5aLFir4wRCQxuced3txZI7TS2d8utT2AS6ygcgdflAnuUiTLQRmnJvIy1c80
PbrhUoV07GqrpGGR7nhoZn3BffkeX6RUnD+MlsDybxLg7ZQfwlwAFfbqnFKaiDvm
m1wWaweUv5ZcWS1SM9Qxxy3KcBajV5X/o6pMbZWew7Ckp8FsULG81EqVW5sSOD3w
JkxtL4P3HNRGDPwb2rXI7jnhNJRIPBZKgWvCX8G6bcWTmXV3tHtShmjwMTznIpzn
HalgIp3Y7Mf8RxD/Wu/Ef2m9FnE5c+xxDsIJYclNlJDrCk9EX0g5/sFQHIo/NrTs
cfpQjpZ6E5VgoObGP7KOXf+dB2J6Euv9g7JZZiOyytIp92ev9F7jruYcDQdXH3Kg
wfE007dX/U/Qf/Go8kW/djTiX4vOehGMEaLK45sHne8pFKmD1drOQI2IibjwHYAV
x4n05or6j1c7cNGWNWoBcYd3iERWhDABeo7i/5XUl1TRhjz+Nt+F2YIWDJT9aaoT
Zp91rvjysK4qpeJ3qywNLSoXkdcYtbhMABGgvcwHJeq8ZUECvBrMZJFzIM69MHX7
o2CKxIOtfde1LkYYLTjeKARAH9axe8At+udkC69q0xwR44zu2fjMFXpcXZ86uv3M
bTzqYDZTR0+SNcOfRBM9L/S151PxhKPQrWUVAKGRPqm17sU4/seMuWI0JX4WZojz
9PFhKH6mjLuooy7uTjdjrRT4fchbu43V9CRsCGxagZI63XFD0hjlEvI9vxa99NGm
PY8hJlEoQhDG1OHxhyWyVK6t3sS8IMYRQMlR1J/vzKQZ8RyOVhYOvdRb83FMCjY7
ZR8cBFXfKzNvjYz4+Da7sutMF7lVHenpCRWm+436yp/vgiWTmcbWTzC3iIY18fnW
zOE4xohQX116Rz2wWsm6OoZmP3mM+j2a65OuxkCW8zBpzDBcy6ICuUNVYDgEu/Su
W77VOwnqmbBKmV0cz2i9/yz5dZA2YFXKakozMJLZ1B2lOQ7xWUjrvSO15g96w8/5
/hJgVuGyP66/EPT/Elpu2L5NbA+RvloYgE4czcJBrKbQqp5xD7WvOqUgxn9dhrKS
5kPBoedVJDft0yrcXO+5Qy6wCJSjkkuns7quOCcEaPxRXOyYXDMVuSudyRUiFyDy
AVYkQ1mMHD6oSWnE2aac5MxC5Pl3227klSNsxfnfCopoJVhTAZIQpL41TQWBU7Fr
/ggfpfchqG1D6R1ycLcWPNWwYfMgiQ8e8wMjN0iOhXk6nNuhxEJm/9szxakdfjUm
7pHRoCHMZzt8rPBvEandWK40ouFePAI5N9sDh4eIQu7KtYR0r6e1PvclwsE2v4ir
uW1ChLueObWWtM3fLqlQ44Lc0vsMfeYG1tE/H9vLmLuxeM0AWLDZJmIJka2rBZhJ
FH67kNaxIgdTkvGi5XemZgt4sMKpqOwXWRtUOSBSLM8k8/CN247n/JPWvuig+Wq4
p8KyuFeHwGP9131dYyCbFwsoOSCEBgYlrw+2rr12zbOlkS96u4APO7SmyBE84Pvn
xpYnlMqKbb8EZtxAOUcMbQ52cqtRhaGw3ad9Usem7bbnvVQiHyUF/IDEEo6R3DBM
MzlC10afO8DkEkifguYmNqsmTAMmIHCNRhakfu+f6W05j3yul+3ZuXixxuo2yEUG
i/rN3zZYfWfjpxCmyjWYgoG8NBDfvnmqzU6O8nxueIL7rzBRi5DhQ53UJCzXYxTf
NDxqFS8FH1KTtgEHhe8qkK1vIcVYIPFrSqHMPfao4OlCZ4O/B0wFI+hw2/LJ9/NW
/tl31yEdo/JS/ZEjP/JC8Tk4fR8PtErhPahf2w9WZ8P0AWnijtVBkW9OFlSMmGfJ
IcxTIjTvFDMLn9ZuUdXwOrzUsDv+3yJ6S1DKOS9DQVeiUAfghL1mpBu8JBJR451M
/k8qeT2mKRXXK38FGQ3GEAfvCpVWmiXNqeXAZCyQXexEO8tWT3OO7Gsm/vLXMMAJ
FE8onClrpTmuBsiJgQcrDTpXJQBnmpNVS49VlWkbXI4XNU5t/xTTtksbC8dWpEdN
8cA/nSrkranwRDDj3W4qiGvmJE5wC1GFk5dWyVq+MwHfnetCCpguOdl9V3TI1GFu
SJhORU+jUJekj16fp6gTWGU+CbjilETErAGbLV9AK9D+E33XZd1biO3fUpVl70Gk
E+dPurM8o2vF/NkAzsvp0VIOug+vQ7BKDOdNlRbU7SAYFdI/Ar3cZ+rTv597I7wM
fd9EwURPgF/pdv48kkaE1aobdlej8cI6270k1um/gY5aZP4v/bUJpDt/uyR7qiPz
kc73qc6wwFpTO+X0ny0GQ9gehOOus9PdMlOtGbzekTS2j+CzZ29c5/1hV7QxxO6S
UmCr9Nq4L6OhC2mY/5DwRSGIsy25yRUPBrJKk2Hbbx1fQmKE+QDGcY6hpHP2DxjU
Cb5YEmNQ5z6deeX5fUKxnV4K97EyGaxE6ieRnqLjgcqG9z/uThPPWU5lMnet25dQ
O420XkMUVeQI8qqp4zaoHaQ4ail5chbmUl9qfeunQa4XBj7/YdiJK7IXvnNaG+hs
vqVDqwpQZjnX5gdcJsdjbT26olMsuAwN1orFlE6IgVWty/JhcnTnAxZbVJtbVe+D
G6vDLtg6C+3HF7NWE/WN/DVOL+R4KvDw7QWX/87v+Vk5Jcx9KLtIBV+kux18mJUC
4FLSFpxE2j5Olj1aTkEwYR54Ee9grMfJ+SOcJKhz5cJC9EK00MimWw/+1XGdGX37
ApNc5Xw8kZCy6ie7PLT4se/2UngM+ryz9caZC5OmeJlkm0OYjkklqzzL6BV6IYTT
FuE3Eou7Ufo/OFsahOLpETQrmAJhrigboQ3zUkjODknwbiU9QeYAvy3AuBzllvxd
bOw3OK6OWMeLueGaIQISClPpDYeDvB+Jvn07pasdZHcfEfAEOq80pPXJphNLGzT1
CafbJ9GHICEgjua8O+wvvb2TB+IzNs4/U0T7+VZXmA5p/2PA1PDb//K2kLMaUH2F
LDabYxB6E687bE3vBcMtI3MVTwxHd5ZWw+kfBTkw7M0wFsWD59kHgigIwQuDc6F9
2poeB4gEcUHX8H680vLYm46TQWj99AlSWfgZ5L8s4yGVPZXj8JlrY7+r+vGcVLjg
Im/slxG6t6eNXgKfMH7Kq2Mv0eWcniqSYsBKE5n8jdwsDj6TcNIOrvg4cHI0jNQm
GHjwnqIM52s1DdGLdvIjwd8jf+RImYpzPacLJYPUIHIcl28CqP2JO5RKIg+/Xuoq
GOezMqXpmQALp5N4bi8qFl1d20BwhNIqyiTePexRfCp4D7r7Ud11QupoI52Qpvgf
ySyUx+VKgoJ6216ToLfSD2wXV1ogaoU6pgoh+32lYJ2zQH3KOoVsLDxci1Y8l27n
81bGFASW6mL0E2pqafx75yi1bR29nQnHD3hRQ9AmWNRQhZPypHoAomxjYbLq7nDa
7DVqhEXIGhCcl46jiP1gou9GnQJQu8VQUkSrZ23esa3DQs9JLRLvci5MiP7h9yRE
CwIU0LBRePHsIp8vc8q/zY8Y4mEbXQdiJ4PBZIWlI8+cUbZjMk20CeSVL8tW27c/
e+ivvce+4/GHhcxpBJdFqzolbe0e/rtmWM+JoO0sAlvIymudaf/eDvlzo295cFHL
Y2FokZxFQ+ef3IO8L+eWcgh1666d0KZhCRlzXzL0o0RKOuAS1zVAmlahuYCQv7EC
h4b4Xk5kkAirq7GXBwHb6WTF6fFMMiB6Kr3M3QWjeysezco6cV9Wk5mk7C3BpgRT
lWw4zgISMVmduxzOgIhTok2KUTXOoRBufYxXflnX5kSKte9Pnbw/jS4Q+sggex0g
ClHBdZmxxS2V5xrGy2MeSwbh+w4gKtdVj8c9WUgtO3YctcCrP2HnuCzKRHcIFf1o
VAaBEwtW9hSZwFYFB8wGYazf/Q9xDpUM+lhlgbqMCczfMGgqOENu/liuY6NhdBxf
Z7ksCeh03f8wDB4o9qINL7dHtydMwyept+5aj4BC6ZJlJzuOOibKyrE4oOBgpoTj
6NQ33W6uU5K7mTMSJr1o/4ZbHQ8KQ3uA+X4zMoxqbNTbWzVxtvDx2zdtg6drL5Ue
+PuiNdm7jGCtMOXdduLr3frusoucMd/HV/Ozi83W9vbShvtvtfaGUYFsFszw4gqt
9FaqQ4fokI8tS3XDULOA3CGGlYdqiQJ1SAbjltVO8W/M+YkO8iNfhuyJpbDNg/za
ktbe5GOj5CILVWz0l6mj1DCxeDASlGmzZyWSekVNsmHprpQPGlxFm5QDfyZIUX57
iE8vTUJV6+USTiUz4oQ0ZHUcKTiMzt16j8l4jwKskiw6QrQhX+/pp5ru0LraNIQt
B13b5T2YuLNp5Xfg96CXlPuNzUxxPINM60x0/3T7EkeTOCEQcIaJzVhIjcp6UTAV
x3EPw1Hrn1XnXo2YOvn04XDUOXyu5BECEubpp55bFW214r3kXXoRiI0bjfBV5Tkq
j2TnKeVgGWM4fCqgA8wjzheHzx1xXG4RqStdF7D3ltDBeejlXnv+kCHH1vXhB1Qi
MT9SQdL1RZlWlasMpWGM59F9JcA1jGBCA6EmbooCQRcQlrsIXeBegd6o7DOmPU5y
RKfYHXdsQ7OXRZzfPuEZGZU2kWjcwxg60/jSsg6jDo7fXHKrqqcs3o6cGfC5trqb
1fpKVqqCHjG6K7zMwY7RGj70zq0LEPWrcbR/lmV7Rz7UGOEYyitMH2W2PpoHSf43
kntF92E3MOWff8OUW6WEa/4mzSJaMMmz1pUyLPBAe6EMri0Nf8ge/YmEZlLKMr7u
lvn+J1lWM2Y/LdqClDDyY67Ul9OrA1EWDiYMybi+wuB+E4kb+r/Ulq5ATIZrlG6y
j8kuo02z0GT5fOYIQRnVUITgQN6ly/BRmP+iCIMAaoK01/rjDzWM6GapJvQtcJW4
8cFlWHmSbVZK7ZJXOwfLzGWVa3agIZJ8+UNnZ7Izo/J/vrR9Ly8pC6bHxwMsE6GU
3XBHWhrJ+AKnnZaucu5ZT4nJtPBS2QSlyhOJHR/0iF85As79uU+GQPT/iZeMPYFC
3GdvFGyb2wUPT0cG39o3dMWgn3tzwAENpr667yVilkgGsu95XE/iQWdIchY0Z014
69d5LHmH/sXQeV2cKkaPgF5H/GgsaM+wjl/6zzz51o8sDvEIdcAh11vy+LaDaccX
n2bjC+QXxLp1zzXfMDLmyvCCn3W0x6n/WNlL1DzTOTxgdThIwCEc6QhhUTCI/pgG
sGbUyPpOAF5gJGSr502DIX+OW/9tQQzgPPavKpmuCKMHp+wS5VNs2b+H4i8kIOh3
Xm+4crlQW2s8caPqiZTk2DqUU5CRFujsY0y0J9IZ8lWDlwJDwOhqmLvYo5Mq0Z7b
JNa7RVZdghC+6cQZyTh0TuFSvphWoeyyhpe/ZGokZOqT76GFutVp+a8H5z8tQj+F
776WrkthajIMzXhJmJeUFhCKrpw61XoqnJIl46UXPYSFpnNx3GqWqeo7PKlpRYxN
e5jz0HZPvExi3sJc5tsc3fzH44Smlh3BPUKXEmYbuGERC+Z7x+WGF3AzJhPMsTNl
JD7V4q2h4kBb2sisD30wmAbYjSRHSeVNQZnUJNJBYcJNvcgyBUASqRu02xaz5Uh7
WAImst7KCUMj3O8shZpP9oeLVazRaMW9i5tgCulN3Id38Z8gj/LD/gzVddVvU+2k
+wpDOEvzW00sswkZKYWTaclDAUuExLRE2PeCFSTkBh+NeDMnVc4/APIyOJ7U9y4u
G81hZB/wRDJdXwITXZ6oRAKHOhUlvd3hNSniaw8ae1Q3TjdNMG/tIS9+EYwPAESS
km8FHXTuIJx3iLgE/8iBtrEDQFJy08g9TDG+xwDCDZaNOdOnt0a4+gyQLYB46leR
FWPSz9W8PB5WCO+I2Xfwo7nyO7trniteMoCWqU1AZPFjC5yGSWpRcT1HFajrsSHn
mKHa9vMW9m1cJcJSQU4CQgIOjRaPP42D6X7UInHOoLAY+Ap+QDXHnZjFYCl3DCu3
oCQunito+hEZuzbPe6fVGfsviIj4Cm0qHule7OJA8+3cURa9B0n+0tMKoZXf4u5O
IClLsrYzif+0PxFoqZMvSLg6RDrnM61Miyiz1q7R7E0/slnHjS6XjysNiBSPS4hF
aApsxiiJPAJEiR5/aJrM7nY+bpqkB+0v8f2p8V2pwKzAp7qFgCVBM50BHEAX0UsK
D9uF/xHlzod6r3GPZqnPJxPlxDEZvT69WlwNkc+P9RUThSI/4LVrFmFHrRXTSXks
SiBowH5oOorHbqvsEDRbnzucRYt2kPVUFiu973YjnMtV870cRhVr2Ox5Zh9l08S8
B76h+P5BHeUlq7NIOxFIoNlt7mX8FHhlLu8CLitPDRTp9oEOLzVG9sxGyqQzZbhX
W8T1mXVNE5WKUU8Rc0ExfQ4FICSiSCdqJsfydbF/4slS4lkmFC+wbkW7Yn0Ne1gB
w06nS+ABGOF15Oj8Sv/ogJZLtFHJasCGY7E6SgR0/LxQfe9x2B6cs7HD/Ddxtoms
0tvydsgEKLJplb8D9gfU5ux68fHuWbK5MkZc8+L79r9NEX8FBxpQmX/olyDBXmE+
oja4CA6Z0zxceReYANPCnxrEcJbKsEdv8+/qh0zmbZJfaASB7vaSJUxMIH/xlTrs
pZdNgPm2NqT0IyTaxyms0aE2j24Adgu4s7fZEgTpcuImLOaC8+/H6P5KZAfIlzm4
zZPpaz43tO44ebDqp/GKJS/gSaOKj7c9nJ0JpMS4rYxJgBhx1/h8nQpqsb1/f694
wdM7t/la027xXiblVRO6chGJP72Md383/mX/KMA/pyHeDacBBXR2m0AmKPupcUfJ
+KX4Prw3ceoTodPUGhMvJDt2/dFzHY5Lf/kcILTV3oz9aBzw005Qh08OXwC67MhR
ohyI8Lgn7bdeWvUiO3hCwj3wc7Huy/pC8ifIcXiCyOVVoXZR7Srq/h+JyWEna8+2
rWohhC0j/yQWFb0QY0wF4A0kkuD17LDJ5gLsb3aEW5tWB65bXqCJIJepSs3KzJyS
yh2aYivniKIOZH1fhLRon2rNCFujOrM4IDxUCOcXlXNIFSB2wSk6sPZXEM+kOJPp
Momi53Syz7fJ6SNak1ok7+8hRWBNCx0hOdipjVmVKonyEKapMqZQ/getSYheXMIh
jdpXMoyjTgqP0dQRsLnOHwJCERqY2q9oePAMtOJaWQwHOaAf+LDe+3uRNR4tyJq8
RMzVQqhaqQT1AMYPv5eHEhOYiTNjAsBNK6VfB3QZl3nuahBXoMCV5URmYfgfRZqX
6wbL1qMgqh7sy8Xi6I75gzPqbcfLFKeXeRH0J+8b1J0WU0w2TNME8J3IrXY7bssl
xMQAfgV2zuiGzzF7MQ17yG2Irm9DsivqETpl0u2vCzZJQ+odWFywR6kr+cSHs6Ap
KDoPDuiHKEWGR5h+PC8hexaqgXK2VMQbiMZP6kjviQ2l8knXaDSIJB5uq04QQ4FY
XyRxM/U2B89RhoDm2QphJsWvpM0kz7vTmdR6cHgu7YLZKFGDGntUvzFGIoDJIhz8
i6RyKIjR1GgG9K7i7z5llJeozQUhaBUni55doRfXgkzs8Rz0cU/zrTnLBj7pqDoI
60fi8pDtMB6MZzPfoJXJnAWq9ikqwC/P5xwgbKg2pKDyoosbRLaaviMni9BEOBk4
rBdEAy32OxhUx9po7tOyK9hHGBb26aI91SHp6beb7fsENKC94HgAFl6dH4k5cTL+
KJ7NFDqxQFKneRF6e/mspwOfbuySkxIBxmE4rwnJ0x7+6GF/Fvbm3AcnuI2puz1Z
klOrtwzjgCyZtpiLdQ8+UHvPC+wxqLH8cbphtINNuZ+WT2bsYax6bact1Tq1fab5
PrkOOt/o6hmrfU0L8/JU7zyPY0byJvFLKJqBEHwFZ2fhh433X6woEDlTuXnAZwpR
QTxEWZGApMQoi1myYRNxTLSGKIj58/uqbfs/nqzNB6TO879TuQAU6DFQh3ZHXnfz
PGnBywgDzWMlDb8LpjRl6uk0e9+xic1NDnysQB+dqJHjKAfuiX2dG2P2imgU7+/a
js72wEr4Jq6+T/KRAGrAbxWW25F6tqWKd3K0mLXWHSBNdNZev5bqvMTGmIoQPmrN
EJzqwWOyIiLYNBFqXUpdJdQYWYtxFw9m/TSqJiHPCjX+D2RzepFQmRBGfOzg3gyq
bkbUXGU4+kbI4MbIOK2+CrjIxaaMfTtd3W8jl7zm021Q2FKhlaSqXJliudrPs4BK
8RUal8Mzh9I3Uzr+z+a1unhA1bnIjh5bdbOCIUFSCHFOxzXHEkHG8C7L4svjAUbv
/+79WKNMJfG3EG0BwUKc/5UUMNCHPPuts3jXyXsdppgN73FXP8p/OZJ/kLbhFeaK
uFUGKncW6lGd1NQn89JvVHFzN1ZXuxsjglvZrpviwbkhVwMlEr5XG9o2y0asfHIZ
GHy6bvmCByz4GdSvYUZSDE5PhrqpwapIkQma5vDobi/dZGyugQmaVN0PXPvkNyMf
Ll86T1KniVmDgKXEZKryf3/GW3JXll6Vjk/RUHY4i+3pdTuh79FQkjEKutUbgn1d
4uqT2VCOltclAUDuQzx8cbxK1IreOJBdfnCT8JNzSGvT+i77jnlA1G1RccySLyJn
V+VkFdtvtK87IkJS8sVtSEOrsa5M+Rz5k6KhVhsCSm0hWntpQauaa3T+w23Fg7k8
ZHwbHabcPkZTj1ioOuCSjs6yCXFjF5tD/gqNY6PPHpcKEkTRU/NpBe4G18bYOEI7
mhkNCQfxPfQnAp2sW8aNReMYDUR15TVSvbrFIKz25rNhA2L4d2qpi9D0krbZhqbz
pveVHRaWyCO9wG3WOin8JMS3F2ZeTTe7tC6gL86FjOzHl7DrdVP5DRbN5GgslyWi
a4jFcNLLCT0E2jUpf2FE7tJebb0Tm7K1TlmpUAmDDQl9LrddwJlWHtcQVMUxw9h7
Y43Hlm/fjz2v73rSQevI0Bm0Sl+75AFZxVmfgD8GGyNzbeWIlegwJuN+38KhSM7B
YMskhEj6kakpd8SKYngyBwe93XAFUXCaHLJluLclZBHlb8C1JsK9aPIo+jn1TOxn
BmcAr7ScO6wLid9nEpjiGV+c+eOLgQUwn5AFcCzSaFAOxZ6wx9aYHhUZjwcx4Gqp
VAfOiir56KoEWu1xKWZbo6l7AKroOWNf9qjGHhC5/G8bcUlc8/uEAGv6GKw7bZSX
JWLYg9UY8IsNxG4icbHYwe6UW937PVt1HAxIRFHwTYVg4ZwZcmViV/ndxAlcNauw
sh92Ff9pOsgXP4De48GYNO/00DH3AnIJ4Yj/4f0BepSc+428B/C8srNZj7+I8oqm
QPEBLiIZmxfqGMa4nsopnpmmJvuivVlqBtHy0FdQYbKf0RSgAzBaTq/FjR1QVY8H
kNjDItLZeazr0d82SDpIvHUl8B+IUuHE/ohfDYcinPkXCcUQ2OB8Qc5Jll+TMM6o
fT3hGpNiuK3VGfXVQfPtYYJgV1wwGe6TM3CnDp/2rQcZmLrDzjKIDotBrsTKEdiu
Ps/d8N/+ZY+X7Jxo4OcpR19F995w9mm8nUnMMa65BQynpNoDOg7DGezb4BiacElU
wp9NmEE8qLs0KK9cdd+I/wLc7eZXCQsRDQOwOdTbIx1bQeJ4IVZDudyHbLg7itRW
QsjV2TAdD6/BO+VF+HzmVP0AT/efrz7/0crYpgD1H6glG/tN3rAy2pHnLBSXFwFf
seAbIAZTMnTffcHgFa8MdyhA/QQesDhuLaTzLqBby58/ffTbAu1376XOm1rBgQQV
UNOld6edc80t6T+u+iec/f3Vc4+Yh2kDJVuEOmAy9vR+Wy1UNeC6na/gxipiVMY9
313O9ky68HGIj5uYBivc6GeOu8SetNY/D+Cg3Vlz16MYQ0Dz/ft8sCcufBbKuwCp
kdMaRjRd7Ma7qv/6i11uYlaX1DDQFoyTyJnbKtTZ1tjeUcyQFUzY/vvFEVy/Ylmy
wRSgJJ9dSZaZa2qZn44CQVSsSyVUqkC8sRAlaeP+5II3sx78xPwh+Ntp40e8stfF
VSJv8g8XmBcu+R2lIgrYLZ0RrNyL/LZH6YmdVo/URMNXA/8+yiDQ+U9NkEIXcIIQ
04hs/e7gUmf88qSarpC4ts31swpovxsSTH9EKLOPOSmu8elqY9I4GIrspeTrOnC0
0r30bLawqKTvw7oLZnGLySCzTTh24A57EKoTP20+Qo4OMX0CqqXoTwXtlmMxwWcg
14uVSqCwA9sOUYhLpsHSbELASe2gVgLpbF6bkESt4d77dAL9XoYS0ccHKHH0Br9E
szQ5CpughvcVbPDYPn/vd4YigKF62qrFucd1OsOVbcl52lldH8NF8TH2AM4buPiO
7XP/3IUZGgzDCjLkPNNlLChO4GUInnLFhBfwqm92+rz18tMmuqcPaaLgzAxZx49/
Yq3SVg7tJ6Qe1jTUpVRvIavUyr0xlBwbrN4gpjasfIFUVrjfXfRag/RleO3Ewuep
FO3rFwol9aZ2ELwfFUyp1ArEkr+JGuzgV+2puFd11I+k8VBska0vXDqd7uY21L6H
7Oatg6XxNKKskGHuj5I3BYvcI+N9iR4Uh6Ml7+qa0v77QNxEOAZU6+Xvf+VtKG0d
0CIFcfv8iGr41MPMzEvfbxIVNWRNrds4F7pTORQyev08qu7KFDBPQwlF0aWM8Eaw
YPB6LZzjK7l6ZhNOUuLMENdcfx+cTdd0LcOGy6YUbLTT/cnT3djCpp7O3Eqne3/Q
PVmbBeV+ijkIGX4wtHwOrYO/fW6IWtrpPDqPOAhzqgI8OqmoFvoAuyyTefGhSnJf
FwYgCGp+nrnC/67dzlUgGApjR0r6+6FZKhZbkXdtN7V95hVbMWzEl3jLn2DGYlcH
cwTlrFvp06/WG3Q7zJhDYUiklkok5B2bcLnbsR5jk2+NBoAWxziX1kA9MnlFvbTH
W4hUmU60gNtUP5yYW9DfvXIJ1P2zJEHC7fAY6fWgHD1xNy2PX+qq7sdUV2OqzWjl
fTeZrV/IXDUC6ykpQyFZuKlTmXVW94eXNePfOux/gMJ6nos8f7VuY8jtvjMvAiBX
F0yMv+4wEbCACopdvvpjfCG+BQDD62cCKppb4ClOAr3yiqB+a7iVMtqBVaf8Xnnb
fE2KnVFzQVtnQATzJoj5q+x/Ic3U3nMpm5ipTQwxRpaj1cfR+lvt61LTRmdBtugE
bz78LNuXXVRvkN8wE30007Bjs9avw/R1o1KUBW1PRRjhQH0lMKNNPaPegnf0sASS
SrPWV3j12fRFOENOMdYCXDsZfI2Teb5s9BOWzubm3mvhQU49Lr3gEEXowJPP9X73
VQN1iiFPH6SET9tP90YDn1IERfQsr1mH04sqYn1G6HofX/BqMUWBecbF60JyuvYL
5SiMJVBp2ojzldv482sd+T4PlBf3nRbazMIL2MUDy9A14BAffsJSM9IyiPVMrcCP
SOWbBQVXbayEDsorppFpczZ1eLls8kCY/Z9j2mJyzjfZacuuT4YWQ1G/Txd2g27C
vzFvBx5ReSjHJy6IIONRwWWbHP+E2Xv/jsSircZ+mrNMcKDk+H/rmqpqRr5KhE07
zChC2e36YPNF29Eph9ZIsjqo+oUDdhCljSaCh+hcUvTyWXmLCJXXtaDA9ekXEJrE
jYgw0ySKj0PU7/d6WvlFTS4PJKnUQVIGu9ZkiZiJMMAK7NOdkTyPF1ftL77zegXZ
gDe5aroprBkxlFOb1vWRFUApdhJpyWrJD2fPuo0tw0I9cs3cqaefruC2dqKS+Qrp
OtDu2Oi3I0sBRTplJd/QhUTncE/+b9bXKA6N+9Bm3IkU4lKnA6FLUHp/lPGqbZEc
YSmndjjFZGbJIJtHlc2Ya3uhqBtYh9NRCId3SEUENejB0GKu9NuBdLd65PzDTWd5
wY6804C3sIPNS5tEe26mLt//EBZRFYm3ROmN+eBiNf4OFWTt6ZLW6g/6sw/h20iz
lT+48qKSpkK5qIjjiQmBP159SGNNtfZ0q2ROjtc8j56SQwAaV8gPy9n7CmyB7IET
cs+ovPGJx+uJdClucJwA5HT8L7+TODaafD2i+/iE8Uj13uYzys4vK0efeXi7sqNW
dpq4ArRXuMcLd6Z7X4MCW5kIpnGgYRZgcbfMe4X5DeUnJig3zzi2RESAN2avlCS3
YLwzWvNx3cOluO+tWy+DowsKlwGxifE5uXDKQd25xUiGcDGeFUjC1nqLncUcuJT3
0lIzl06BvlopDREf5ZnmtjfQo55xN+ssFXREG8XQvvLyFzC9m+kiA0j8UVzjAbyf
qOCD9rNGzDPOB5Oe2XTuL8KDSYV6cgGePobvCOWJgThGkZAUxmap9P3d+0RN/Ahf
O+js9l8qWu5wG3ezqrForeulVAOlEa/kFziwkNBq7ABnb4M4XyQCjmv0bdMv5pdf
Te93o8wq+oPaI75QLo9a0atdYN52P7OwSdGyeQPeaoDd38+/CQzCKxABvzfWEyCR
iGNW7i1E18QqbFGbITnVC2+n91J2MUPU6licjCT5sPgC+TDR8/wKmcTXCg3oH3kc
XK4A7XMSb2Ka150rnme6979CRAeZv2FO57+PmOPHA6XFtVxq4YxqSd9csfzGpT6k
5lxQ48D1R2aDlPbzoP4KlpOWoPLjbCUCFT341E1mnImaMoDXmp3jQyegzhI4ky59
+HXCAgDoGVbSQqzwW+syYy9/fU6oIEm6MSXJxvRwgtufvlSJRWqF2da3Oby0n1A0
H7YXe0jwtGHY/A/JQ4H5BlsgIs75WZ6TgLTQi28nM1ZsBgs17h0oegkQWx2zm9z3
MPttsALS1RpeS3fDk6OKpcE/oPgqZXPoCguefqPOBM6taVXIBIvaAv+iKCkTALju
3KCpo8a9Evs0+p7R7xTvruHwku+E5ZaQFrwWwT993MOouVdq+5ByXrIGJ6w/mELT
WwfOfUd0RmJNX4ewEW1nPHqIOaUFYlaABtJWQYw6lr72i3tPPmI28qS96MdzBf45
HJqxYcVCK9IM8JX7eccR7GQ1M9/x5NA2WuDLMi/zdpmYMNwd5I3QsLJJF9GpkseG
X30k4c4u3iqtlZeGDuTU616SDS3ybkFHxE1fH54dWE5K8xQSAjcitXF+NzzRd7VT
zDOT28tY+J4/mzMIXCKZNbPQ/VUzuuITHHzUriSGtzmbiKRTfTdSkarYl0qr4IyD
dRQ7Y3bDIlVoXOuEe5uZbyZgRoF4JFY4oXTSXe2wMPX8eEddu0xxpQS3IsWw3RS4
rtmeZrZE+y2liZNVSDLGp+2jCkVSRkqM690u2tlvaFyVMeXl0HGeRUDgcGO6u1ek
AeV57EoDa4C4IMbTNUC3mjaKDC+YaFcKSi86M/ST+BlSM18q8XZ0touCS/7fGQO0
5MXfvVALc0TYGSAtCQ0O5Gl3/Pp/DZsqeCVwA16fbKT5wB8wwxHLHWUHmzmQzOaX
2e/RGrrc44Y2+OUqeQXTgJTJUvXzuLMJiaLVKmwdCQcFv8tACU1o8CV7CxhEdmgg
cOTymIp2whhQKcynctiQLkQaU5J5Xs/uOxW3sOjQgC199E9tlXOrsabUTt1A/8jz
xqL5F7I4yMpWfgHHvwwdMalF7RQpermR0sp8fVckkMQpCT21KDjBV748LRl1eOap
C0GqB4MXaVCIE71I5g0UVJ+ij5jtphjX/JfNTKe/hnUN77LPWn87hjxA7JxZMUK3
Xv7QAeCdiZIQUAoeWN9q+QgbKmq99JNWLfT3yPhmySTtifMUwjG0wZGpZoB3knUt
xEgUBKE/L297f6fMNZLPOF5QN7Pus1Nemv9Bliy0hxDmlMNu7ik1wUXAZg/+iChC
wY/Uqm3q2WwH2ITh2CKiegw6NyvWm1huDR9FcCYhVxsLK8Bs6e/MCthHsVmPRV/a
8SZWal8DmEZGi5Dmlf6OqGTFlKVI3Y0fQQsSWQf/o+8E34X+Jw/skCTID6xaIWMo
JwHeOtQKGg0SO1nO+2tibiDwRIHmvxUtV0vBwF7Cq2CPbFwe1WbI2AZfJxS7GSvl
xluGfKNhLBWhyHP/bgjYmVRddKtpGJc6pFJIf2qYsD42+qN9vxuksrVykl2+22xX
H/wDrFbtnH3SQmbSvyKN8U/caP64ym6bypD7FSocRlpd7ymsggEV+q9M3EIDZ9gM
GHCf2PzOi2TzQYPVyxwrNcFbj9hHs0eMW3NiM/NTU4QylYjhcR+c9lMOU7fDJv3M
zSwbF4FYwMZQIJs52jJp3z6ZlfRElqwKXK6Y+NPRcxC+w+++gOZphZZPokBmZ3iQ
ubPx9GBvuGYXWLWl0HV4ItebvUeAyhwOtKKnUGL/68HCV45xDQIxsQ1KrNac9T0y
Qxx/Igj1CkclAhcpjIziRrxCeVjW4cD7SeTA1ebT1/NaUaw2a6L2/whgDMg7goYs
TaN6mdfK0v4wEkEG9WFbYlthPX3IkNMWtnZ4CLBPkta9bx9I0oEVNZYe9K7+cowv
ZWEfZpDYi1kXtm+4V4KFeHZiGNAZK1LKCTufJh3KBZexUwqh53XW0K3RJb7CnCcb
SxEoep+FVb3JNeycwT7JFz2HnfsHRo1uRcG2khLw8+yQz0ExyNR8OyEGqbXhQI0z
teLbnOF1uHD9S2Zf/fAe+eRXm2gKASPN3GeUuFHzGJpcuyGzZ7v9L/Sp+oJikHY3
7Q85S22rbRLJulEBC9h1z93gm/YvpAsJrX8vuZXWyOeg1Vs4y6B1wVz+KZ7T3z/i
n7C6Qs8bW45OGcb/xERWMUdgK8zjSFlIc2uY7iTsn8y564p2HahhQn4s9m4m+FV+
NjsI3SAkm7L9zeN7bT6+b7c2blf43Vz9CAoExTzMrHhIRGoehwrB5Ri6DegMHOAx
rLSg/sy7s2qe8w+uNuFbZ0wTqgH0nKVDsKs3SPY1PJc5otUtrxenPI3MpVjvXCRf
UKCTo6/Yzz/OqsJpFE8icxOyXVp8GNl/2IxS4BkvaT29C6PgA+mD/g5cW13Aa8TA
MBaNJ/GmvVJeMXybjvgp4s0z4K1n3Xo738v/DSbNv+GLRd3JWfkWVT3u6Ya0SxXb
xgSfbOoepRWpuP+9x5vZt05tEi3tPypViQ/CdVe51NgenP7EfCQVTUY6wYKubYfh
LfqxecoW/99wQLLcqu00POaNc6KG/v1gaXlqJyR9GYiSLOWaRF27hbRuvCeSjkFh
xI29kx/3huvCGc7XeTEyZrDnv/3aZ9YUV07SnFlKUpndFDYLK10HKJ4m3oRWZ8Sc
Dh6REtM1PxApUdxVsGi+R5lP/NAas7K0NEnqjwvQd89lfYAWdyuD9v+dd1QVS14+
EDoBQ868caxkLUMjbiIeGrapVXD5gK/Fn6SMocJJf1Po9ZQehdmpQIRiw+ZNNZfo
U4w+lvwIJODRO1X27FvWW0mF+RDIfoNmpSbgFAW/D735ToYSDDFdnQv4J9expaIb
JvH+TUE2W+R8ou02R1Nmi9hXhoxwNnJTnxr5iM+uqaF1gez8q9saMR5LuYQOC+ZQ
9/g75WWqE8taIG4uejolps7Hx+FT0ILJZpMFLz8doRfmjVAV4xeoZ732Ua2YzGlz
79fa2Ezfft/iOiSkRxoEmPWeBbLwXbXMVoxCCMqMp8himd3cEoDSBK1zWNKrQ0aV
v77oTVKqnRRfj109zjTYlFHtFGDk0by2Bgm6+6rGlI4NvtYTlddp3iFmLjCnA4bF
f7NvqsigwryZ1CigRtoX1IGHfLJ40KWYN6qMjN8++vX4L7cxkZAFOfxu5a22LIRI
OJhSLBBAZfVqz3qQmdW5w41gs6yINmXy5Y8lh6t/62gBdInA3UQdZCzz+3qP34ge
RbJusVzgvUwXR+BuccrLbeI5NJgAfo++l4ej9/2be5L6Dxw6oafR97HmQ/JIq9uQ
uezxyWMSj71Srft1UkHa4yUBN3CIEy/GXWKrJoKvibgWCZzrZji6m+FG59TzienP
ARDZsmDJ7wNuLOr1AmbhENJiyUC3+huCFCTLg0JbI2Exxguy7wey8FtZsqcVzAe0
UNXq+F0pVdizfATe4bN6CFzwu17iwD6j9lhq845EclRMVAnAlMsSq7l75B2fDovG
7fi1KgxaGBYO01cRnr7LfirsrKU/TGJhIs5Q7B4h9+l2SXfdbWeNyoH7vmsdNaR2
U134m0SBJPMP+fVKqCeGXblr10YDo0KD9xPPT5GN7AKYW6cUjhkUCBVV+c3efF63
7b1Rph4n5Dal/jv+2FqRtYWHVDl75RMsTzw5x4Axsw84nD2akCVpAe6rcZtf3diw
rlNifGCM2MAWAo2u33pSNFhYXfVZfG8yGmRSzW9vimpJRNXnZ4QTWO/XaHBAVAyS
SbEoV6qnhsoNLpQZtk210Nv0I9TGMBsONjePdFs1iXs1/1D1cVs4zfq0FKVbuhm1
rYhK7RFGwjeS4OIeYcJBhJMfRHy9eCUeVjStOK0hD/AgvVcLoNKUF0lfKs7B2vzV
kxIn0kfagfdHfatDjEQ/e+M3EKKxfyVgDfiyJGKC5kC8vA03OkNl9+1oTnZcVRIT
tdQkkt/U5sz7x5RC8AGVIkhqXIZhTKjbPz9t2KjyNoTulZ2Cg5c1lcVwhW9W0MDX
PUqwOwBrC+B0d4Ve57Zq1hMjMaPl52RSzbuEsdUllFXk6oLoG6slLSMbAoPMs56Y
LKNFywl6/sDZqqNmm6AAVTQHNG5oIyFGufVldQxcBDiEWCr0CWyZOByBzNmI6G45
3dzD+cjSmiL/9zSa8CafMeaXl9t18q3gxOD3wXyqPnEcaBq36PIcXYnRacNPthSR
ngQN50PnGWZeQ1HIrckPshTsF38/x5TM1cQJsr3MxewpbG2UtEQT7peR2inesBHQ
ufP3DJQ9oaB9SXm+6vpZL2N3c4KKVcred9f2B3Q5wAI+AQPcof1gF1PTErm+SDzO
2nwIoqDlIIX2hX3kXskjiobxbYaNOU054CDeHZs3sHYH1YSO4SaamzN5nq0DTX5c
NuEZ91/gYzqRdEK4Jbrw23bxGC7CekpMbI4jRkt4UpTHFNzrvAcqDTfSAnzkYOsv
uN2qL2DHK4A2sSaImk4S+JflTM6RBE2cG3sIXqESwWh2f31Wqt1rqwE1bhWd4W6q
KxA/5d6/wkZMKOqxrwm8pCfQ43FXvV7t3PEeZQEMCYcOSS5/EMVSwl/OavDCajLI
SPcvUErMcxaXP+gXMgW35kD8teDnMbJ3yMl/j1+Y1duv8wdk/+5mY+eMbCI+s9QC
Py0EIXWj4EzxKMGjwA2obwVVOcyfVn78kkTH4Wm3jJ3+utRNv9Mm6ZjMmxwKpIHT
rUan7bbDIBjjWF/Iw9gr+JtHhD1ouYA3AhoJksU6TnviB9e408tQ1LvkfsoxpbKr
Biq0Xdo6JqwsOdp0TFrOvgi0/3lGCgjQ6SHaC69ImwoqhpjxmT+pcLOGZbsTtVdK
VASNilF4BWynep31169fQM/qWHshpCEy3wzURw6DIZLN9pxMQSxtnQGXoOVbYP0W
kn/7wTB013K2+w9LaYO5OxongVEM2wqDpHPW+Tvyrc7MJE5/+jaqItX/GNQmE8Gc
QkwjcjKcOzB1sYwB10kLoRU5OtST2mqFJ+xLan0g/sXK5N0bHyug6kaoM3VFsrjd
6DF2GbpICajefo06BFCHL+DhRbzo18f3LjNmoRsWzHvMJ74mte2kRWVDKZe/d3tN
xejEdv1U/kPSPdjoTH5elSCexP92ODFqVVCDHc48xXIVBrbzdffNrkdHhmAdHES0
gm64r89Zag3rslZkyXm0OzWDym2+m+uiUgb5LNrI74CdqN/+yupOPqU0fmtR/gcv
lOEBFyn1e7RgBsuCPVpg7jndguC5XH+rDkIiog1aRTM7+uu09EMfZdtG4fla0Oq6
SuWRqii9hB7XXZhxi5JUahputzLSit9JOr6uA3ht0Y3TsJBUxFscMaNEhbULiPrp
KAJj/q7QRPw8TO+FPbcyw0dCPBqY3A9YCZhOUdvi6YlIF+9iB7PImIO8P9TCcAbp
uNr4H3QyxU80+lhMy/vEJpjTdZ8tzml/+n0OvBd7JVE6XNLRha8nFzN7YQY65/fU
niUTLle3jUNL+ZRYm5bjYfSoy7OlBI4S2mLt3oBV7JxgZhi9hyU80EqgOQ989BdH
Z0U/7VBb4ZrcZZraP/i58SQnS5ksiC+qpBOROx5IRuaNZ913X+lvbebG8Z9/QtK9
t469sBn9XAesXqFwPBU5Fn+kkYFfiwAG4EWOmh0gAYmcR2pXMY5xO3ybP1ayUmJE
DPf47YixnuCDhNqY+lvhwK8WmotbxBrxyaVLI6q5XO+foIWOJ5JsInZRE/8hR4V9
gqTMJBBH8WKErIuOJJuJyfW8FqHNxr7oNQc14MuoxslD/g2nK/KQroQdCIa6obCb
KagHCtCY8QSdsJDg6PkbxtcfWm0S/2ZZg0zj93pKJN6siinTen2aHt94llDRk2Vt
KnSTWRC5sHMYv01GnUk9XjLxOBE0lZbalaJxkeJtrBOTeuSHa0ajaa8LAaVinRoh
80BtG8g2Tgbv1MILreI5/dBHjNkMKSDcHuv+EgMPDSf/937gbQEQERExJZ2OOaK3
lSgdQ+qzSKCW+6pG7r0pmqM3CMD6o9XQqjS6N3OsHS4pLM0LIKtSfj8ZunaXJKIk
K4bsljayVyVdjUQ4aNAmhYLx8uNcORpAvdqQ+EmLtgQXF5oITgc5qfuVOU6mJbkS
74F752WxhmRPkxG/KrDE/OeRsST3ZQz5fI4fxW9O6ZgwVl9sC5E5zRMF30F6M/80
p6MHv9+URfHjYKltLvT0l/OE7Hi1spYNAIreKfZl7H2jg1Vd4/HYhqgnlfoUKgNp
vEXqvav/z2izRs/AoLf1Z3e/XoPoesVqzjH3TRiRsqpf/wam8acbt6CHhsWO0VCQ
MVq+bMgOtCoX8s3Jv4v60ZxCKF3+llcQSCZnMMh82CmQhaGVTySC4FqrQCkbESwM
y1kbgIMcFRADx6cT0L6GbAQet0HPcGJMdg5TDI3fsWG7SGHdNArbjfj8aPSS1PMR
jEwts1CyvxQStODMLqciQDI9sGRtG+s394FMDG4HomaoUpql1d2Ok4CLuwHn6DdV
XcFr/BKSGdEAAob1etkvtn73GmdKGnjpl+1o3mmaPgJjo89sdZbPm6M19XEQnZX7
bXKEnIoNY5PmiQaUv7cggcsKWj5Hix2KARsnc+89ArjGx4Lkmo1yvRiwR+hZiCT0
0kMqEHX0UR6U8Lf9qzcuL+OCKwJ9LBpu10EfZ5q4eLeadR7fBMCYSy84YJmwG4XI
EJj+N+37a7cYuf1lpoM+z3oO7kBOpxYLjE2ls6OzCCcxHflbpeCb5UpPZEk0M4G5
riUmMisx+unyxO9tf6ujzApslNcLpnEmFV4dMbxE1m06Yq9vvty2O3aoriHILLqL
9yePo+69SSaRCExanaVaKmPSlp5NN5dzfOSqNSGfwW0OhZejYacK5YikZC5yvT6O
3BjY1fcjyukK+u//nMhGZtAMJ2wFBvVUe/mR15M0sI86+Ou447r9/MGqWhs5ws+r
Gp3XgPzN5gAMe+Qu+wWOXUNXCt8btYAQlonRKXthsnhXRVS42B/Tcg1o5zH1l9pp
Vdsxes9f28tqQ9bECCj3UWu0k00Sx1LAHe+oTuRAMn3veHhvGTbzp3rKUlbCR6oP
rudjMXS2AvwoB5AbDf/Ut7/ckr4H+HfLXG/zNdeZ2kKSWqxRFVogLMIdQEAnf8T8
bCZf71oiv4c+7pQvQGY32/qk4CjL3cbBU9n5IPRPr3ANoClz9L3cGS/cakm4cAn0
Sqf1IrXJ1i2nZEOB754MZMO/XDS7oDuNyBs2gg3a/9QAfwxXy2l9OjxRPpcxdC+e
cLfITRKCsH3/GFYldIHXxAzh9VLGzUzFOo0rjNTT1ZW2tO+4NoYJKm+P4RtTLoyD
ED81HoJArQO5qObY3BweSpofsFSNbhymlnO4hDIGIo/xwH2LSOe52ExSe46P8Wr5
Jg3+33V14tlZyG6ugeBDgWdewb+8PY8uySrUvycXG/G3WU6plGh1Xck2Z2ZIJ0HZ
M/vfeRP493ThzWM7ry15lNPeQjL9iCJf/1D+ldd2DUo9zAEbsnaTCrqx5+c2wtV4
dnZ/r/GMVJ7oCjajlbtfIjjyDA4hokuBt+WCCC/bhKLpDUvxaj4Q7W1YVbUFeGPB
HUzAo/oP/ztquqmUhB31uTSsgl02wJIDZmoN0YaTWc7F0+6zIa8kzZgHiYv+lrWD
Dbsuj1rDlbR5mEZ5UMslbU8Dli/E1uhrkLBhNRqhFbD6tha/WweQz5SHQYuTNS+g
ZWaV6FKHtBh7SWperGUk4wT5hDmtzRagy9dyzi5eyQ5PuOL+c3wg1AGT3m2u41wU
twZbfuUkuKevBGmGbFZIRyXgpuGd7kGDjjk9YSvWn+eXUqXiGMo8IL97S6cElmOU
tfsqMPTuzfahrfOw8A0ac6zMVJz+hHt7mzqNFaK/3VeHTOVEH5AHk858ETmuXcYK
aDLy86aB5pi9mAQvy2m++2XZyk7dmjQ1OHL9L24I+VOiMuPwcNGxR0q3PS4FxVn1
FjSkXaW8LZdAyjCe9PSqzNzp5mtQeVTKyZ28GW6STHKwg54szpuDyuUtO9Jg2YuL
LHYxcLJq8p1FTQ5B17wsfFlv6ue0AbZGhx32VlZ2hGpPLbCFSlFa4Z5j+ucLz1Gg
+WyKV3mmBjhxXAtZlr1/9Zr9UvTcXhA/VlIYJzhls5s8MU1fcUnO1JFu/aER0iVn
no8VCtUKHoKNlZ0TEpKlkSqRJoBgqMXECrEo+yxssWD6gamOs6lJIQiiy2C8Hpzr
5Na3LERtVlNpxFNmgaHFJs1+tqyutJyiMONwTa/YU7uCJfKzwsxi51EVYsbVS84M
2TGW3hbb1m0c/a3e+V19LvNuUabXV8Zby2F3ZTu0YU/MxzQBdXZNdGB27zGp3dQy
us8rOzYp9XKJdq9N5NmMyvTVTUJ0LxQKK+VClRvcJLTy/fb4HUOHzUFAgqHvY1d/
jBza85WsBnQeIjqipAvNoktyj9iiU72Ey21NiqaI+3UUfj22N0O7j9/fFSZK3uAU
eA+kDluNL9bdKWBXin16Vpxxb961NNhuZwyINVGXTXr/CQNLd1fxlmIZnXJwl6lc
amJFiotyBC4M+pNueBbxRobYzCvygS07J92c16zYApx/1SZWaqE7SR4nA79MfRM1
igXdftbgf0lZCt/Jn+y4TWPxOwkf5HF4tsvutpojZbqDWoBrUkByYnOrlxWiO1S6
NPHEyNpHSEGYp4G4cA+0BnWBnOH3dBjkozYiqXuDCAAMEG5HJsH4vTVb/LN6NVbz
rHUNFUSBsDNvUAKqx/Yy37eRWCrt6J6I7rTtxb+UQMwxPFcQ7ormv5VqJddgnk9v
knsiQgTg4iew3nO6/72o9YCjd5/f9Jn8VTuw/PI7r+9IG1KVm2znA4AUCEJMySbt
A+2Ss+poAHCD0VhN/A8Gqt5x2+aY9pgOvWx8hbNhEUqJUXIrit+uO4lEpwo8qrdB
M347WOoVplPaxQTUSQfIi8UyNZ8k2RzamUdROSCfyXbw2Z9MBuu8JrvJloUVACMY
CRbKWijiV0vVEoaQXWOhIAuzmw9Q2AWoOk9q//rD0zlxSW930JNa9z1MhVP7T/sL
P6oFCVKp+L/8ZNJTI25f/aOPJ1txVV4NbisZ5igbIxtqRYEzaiKtilpT/WvOX3i8
vTj0gWQVe6kmmKP/WOrEltp02D5PjyeRfxfh1QaF/wu1aXPoUX4Lt2FKeNTSuWJx
A0EzSfMwEmJ3YxTp+jUgzQ0cMXGqw8Ii+U9Rl5FvJ6+Yvf1Syxaw3AjdvAhNkmOi
ELZru7rNLbxMcb2dMLT2p6+x6CFYhdf7/Qrht/5WIuEzt6UvAa7reytzq6j6Gdn2
6TNkdhxZksRlQDvfpTMnz7Sm6Cg9nYFiKT3T9AyHV7Gy9QWDnrqWzBRn9rbzugfO
gYoWVtDMSVqG4tpLaEJ4lFdDVaMr/OYJcgzVUFXkzgjcztTVgNbKMxKtdQm8xZCw
oi+Qf0yup1GaymmYKjaKzFdj8N+3GOAs70/SsZObYCRsBnHTU42VWuFffmbIrwUK
wAP7cIKZdkO0ECNrP9lLiOgwK+C2gvYaVbGHJ9Wg7gjzXlfrIy5v9kGGxhpgqZOx
4WTxXoJgTvvz12icJTEFoNy8so4i3NnopoxGHLaFyL2p1p4W2EbkP4BjfiSObb5V
aFlM58dDiz8cQJwVArhDSOb9VuDCrVP0vTnvuyLt2aFpZd65TH1vHRBeL9CzIMtA
rVd6IImoIHkeHlv+h2Y9acP8RbUi27UMhzfsKHOJ+8YoaXi9IqwBS6EsQ7bv0TpE
tYCeRb7XjdsGIzuMdSOZyxrZ4j079CgSgK5iIb+ZRSj0onHj0uxTXWIPaqnwEHcR
MweXyxysflroMKhJKqoIlM7rj94ogzYb0wXNUcvOyefgsrWrYbEhqXcRdszl61eU
TMmd1LKeZeGnJ10EW9DxVATtKwFa8XPbRUIcIFekrkOVRfXwlGSl3Cbq24Ytl7Pt
85kPmfbQJ8BBJlZ+u9pzeqwJezY+uPgh0IiAhBJZ0knekcF6QsceWV2pP71HEI7k
g8U9DkF6okltvb6qPGnAFVy6E6Fynv79HYa6ybjvjtrV25C0btBExB9LTp11xcyj
JVBkiDolmEvegGLliPGsuYOs0yYoqRxvBv1drv7luZjebquAWGync8uZX8q9Xhna
nFCXhrFC0MxnEtc4DEyls9P951vcymz+vBJJ06n8HTq6L3Bp08ftAvPA0mlhZ+kd
kxIzRWsFvxl+yi2wjGWYOrZySGVPbYJrLDHYKSj1V1mFe7K33dREFJ3c1tU9kI2m
ADiLqBfTXeFEUV7yiCR1i4QTL2oepo4dANZntinv4IXRMB7V+Kc21Xc1d6j6yyyv
DhwlurA5WhlCVxz/TdFcVNtMFacyIjZqBfuHNDBXYksCZ5w4bxY+eQQNT3jQ3CSi
DXB2o/IXM6CCxRaYHM9HWOA247yyAB8DuluVcDd1UptY0KtlKsvcGOMD8fJA5I7X
MQ8zATWqys62FyY+XSqAb2JEFi/7EvMFyR6DxXb9MkgvaVSWM1kzQEIusv4P7TcF
8uiDlA7iNHy6sdAzCZXtQ1yOX3RmVByyY27LXmmV34KcQtLPqEeLWxf67xyGVDDt
NeFyKX8t0jBvsUUndGq47MKCElF2BueQWwkEY2P36Vpht2oGjXxj+q5ect5SPh0p
ySENm5TqrAe8dF0d21m1Msn6iEtFZufcARPy1eXN67A4S2mKgy904u1BX4an4zHe
zy0yHyO6tnJuGWG+P5FP8gx0R8TLrSHe6n/nKbCo2jRHMEsx58BGXIoDo1zA0ebk
Q6OcJwQ6bXRx6wlbOkVEbRnGt8dsbkpOQO1RZaxY1ac4SVCKWT4pL7REmCs5qKOm
gK0rU7wJz5vjNt1YQ13kex71noX/8k1Ywq19YSF4qH4DZcy3nASDFwbdoSZSChPd
wZxL3SKqxz9nHDKdxjzRkLr9f9vsL3jGrZWNKv3OVntDVLiZrMCbKvlRQjR8BYIK
E2Aa+/e+GOMe6u/6mJ01+bD/iFiQf7LD2Ss0l8vxx8w+KfNJbefXg5htBXDGdEkZ
KTVSV0eUI3G5+VYEDoUJiUB8XHLxofQn3dvOOJTYpoKJRW1myIzhFWTx9+RbmtDu
PrTag2tK4oQn5supS8zuAO1AkQoUcT/ZdnNOwH/0pE8pMc2HbldnL1eJpqdkdacB
Q9szkYbRNibQoDglKBMAm5NMjzHuAJaePIr6H5SNuYyAKETMKPBVBQx4ONwx3qvf
+h8laC423lrPzE0uv6ICGQXNYr2+OflgYMgNJZsBR9GidMGuoVbYnqbuhXoFSRIY
BJC66ivuIZBUgt6G+ByYpB/6ldQeG9hXQq1FHDlO5ub+GyPJ2OtNmW2Yj1udSPAQ
J8P+kZCXdF14KO9tzRiGy3YpiltMxSDy/jqDbJFmyB+VoAn34/rkNqb0Xgv2z47J
0ULAYYQwIPcfApTeyOcqKIL6vYAaixBHRqYdp7ippPX2pJ1X1n9nb4+crFhy+6Vf
c/m4R32MZFn99G0a7QH6DP+umwjIDQKH5rbT1HWC3jVeDxhBd4i0dBYR4xkWUyet
hA+wBnYClTBl1s3GsjJcGgjumddO43hMQQEJvC1XJOFFmnJeBi+bengPRj1xTVIC
VdHk7zMWs+SdvIPY6NYLaOjKF1KfOu/6moq/ENHoKe0gcGA1c+fcEYENvVBAP6HJ
ijCqqrxmzdE7U17MxjKzvcmY35NDkzneQ+5N/aGnNDlctM+go0pFB2fixWl6rJ60
uVizSIgK6Nz5NmwAuUKDx8CcaK79i5A8dRex/NZy9bYFN+iDWSUtExRMexLaBoTk
kySLWK3JffbXiFYeE0axP7wFCY5gGoL8gVI+4QW1FRJpyni+S1O36+xyG/OyiuZW
9CyPyrUVM6y3hrP3cL1LMI4+FJ7mey3i9p5tU5PMT3SIFXUO4vip/TB8AOY23IH1
pCn+bEWRPqyy1aRZohA7ycUK+115c5G2vaIwLrkc5vZrGwIdwbiUojLZeCsjR7xy
v9Yur8MvXcAKCZEP0Y9eLucUrsiNZ7UrNvIR18Xg7br75dlPFFx1fTGzKUWmi8GR
hrWpJqJC+h0X0zrsDPYdTJlXJa83hbuQ/vvm9IlQ52cXMyDZS0IapX9Y0pkfU48S
746TwXOpC+xSmlUrzh0AO3l2GgHhjKnydaBVdHbj2dj+9tWxVemC1rVjprkQXgKX
fQXMTkZDG0GJ+fg6Wuty0kyVbiKSu1LFJHynKrKfvYSTmIcTgfF7QsJyAj9li6ez
0wfaVJ1pUS7o+MgFYGZYaGH5n9ayw4KJ0lIQe+ODT1rQ0/igYRUdbxy6TJQzgUVn
UkGto+7zRQlvO6KU7m6XvTHemvGorFsiaDo6zozXk2n7Mgpqo3BCa8Ofn9VVFWJZ
HxJtr73ch5enBlxBzViB0HCkTYwbLVfmCHFINUkMVq/qDg4Sq5m0dcM9i8bdR/pl
mjIRGvv4iPQt5O+OFeVgI1NzglFqycFm4L3xWK7J86Um2DSvaJ9ta1Ch2SKI4fZK
TJqqonHik4Lbsl8gtTF3XiouunYuNpm7O6a3algYXZRWR7RF2bVRVrio76hDqKT8
Hnx7Yk6Cz8+KcjvOzQxNLnjweWua3lvtm5P6R5gLCD9K1Tsl0RE+z3khT0+Z/k3v
o4phdSslgV6Oc/f2zjL/gWLndmXB/jXIuD5SoHB2+O8z2+ML8G2x+NC92dOibKY2
AbQuTFbryTlRsI+mJdAUOt0IeTBr44XNxcNX7ZQZgWdyDzAEE6rk1zXY38E6xPJY
/GPBH3hL6In3mAP2YGQJviJlVG65Gj+w9B7KGDNPEF9sh63JQTbuSaAflLX21sip
X2zycRzrZzPLsB8t7iRhKg5QODQ0JSL52zvMqijie8a1jKK8mkUEU4FI/cuaB9rQ
kPtMqsdxeUMj10uwFqvFut4XHKl5Ol2HEXYSqrLJGak1ngiyg5H3aiqACdNK8m+s
A2UIC4BHMvzke9GCusfXnKn3257HsimKSHufRjKuJhBJqfO/edJHbtAYaJCrqumg
wj6pB0TjmpN0cZE6tBvHb4L+pb9Hw0/m82uYO5DsQgsib0GJzBNng4jP0HQrb/Ba
rpfG1AOXmBbBo2nF14uOx3bUWLELTFS6AiLBNLL4agqLC4bXDfukqfvli8J/pJUr
dAVZhID4Wk/PPOorDaf4X2nK1bAvP/luV2hfBqI8SJ4HDH2cFrnggl1dDomwbODM
hCgYkgi4oQdihB0zZ7ZZhRo9OSZa89wEFsE4Tf6GWhImFNseGDQiLeg05ni5bvCr
qPzsH5koIwkKhDNJkQCbB50xUoWSTrEeEbZCUeTxUHS5kAD0RjEG9Sf5z6snXtNC
zE4A0TLHCN7xUOkxtNIVM4Xe8VOWAT09A8bRE5gxbioMq9U5p897iN7EtXG4rxVX
wBXWMJYPRmkYtXLewz5GGyb0ZB3Vej38EKv+qvrjzW7W2ciVUKDW7ucRldE+sefE
w2xhpF8NZd3EwvAKmPKzpgzjIzEFNHkhKWXBkD1X4jlY0jm2ceA41zNJUYgyN/l6
kCSS6gCQjAnpmVKitXI/yetUK96CROFgz0ETRX+myUUdcGseSTSCctmQKWl66XXm
BJ0b6k2SBFD3KlqsSkylQNjPGY2qMF9KG35j5sFIjXIJnD79usfwMmJdsUNRpVIG
fZi6bQRsh7zNw6slTqUAhUagIWowNbcQRCpFR2Inz+sM75CJjj6GVniomzwOSSR0
5bJJ7N5LifiB6UHL6lRZosLUyYGPshac4XTJHkk8ntqSwu0QntH+idfvLJyPfiP9
PMwkcP04mBtJF/Su8X5GA+mgldiHWFPIDSTcnqJT3BgAozgcM32nXxI8SiuV4qwa
ur8DDxaCjq1FOmToASOQUMtte334AA0pyizerm//DEdaQ9HBg5gfki4lh1M1CRfc
DTsqKQOmRGRQFOlHq1SCiQikqHbsNUw/YdXpZl/JgT+MrAXVlBhzG89cBW7gqt47
MhLA43hQ7I+UyErMS7SH8adHLyiu4W0NVhP2+emE38KjWtoE3N5KMqnk+Op232MW
YHHc6phVdJm3m0FsHshzWpFjUfl0w3vc5WbsSV6p9nVw3s2ylReY1BJQDvAg2Ajv
jYyKn912P+wWHJGGMo5Z058LPVwkPCvlU8y3iGm6/xfrO9UQmJbzWxEnjNTqx7up
J9aNYp0GB/JVE0oAHP96PH5Yvw1fhrBE1Ip1UOJ+l42SJCYtRGa7B+yu2Ex6OP8Y
dq4XBwYePMXB+GhLXHMA/YJ76i/Z+4jKAvK0qO4DoQh0O//4jPZ9rW98dmW/Vrlm
zRHeIJExVPCSfrNiLQxXpL1SAIFwfO6NfDWZkL2Xke6IfSUlOrNTzXw9wX8JDTTm
9JZHOc4b2J9rX+KdMSQ4uUwaDhFEjEEWpwKLZ86e7GaK+JbJn6o84+jnn9JKYLcv
bKFOPTSXzQHqGTGlqAn5O3v9to4HvnW3clYOMeWVFpn+kcArDg8S7U4XixcOb1Wj
3g74GDk1+e9CoSDxyaETxqbpwnxzx5PUaXs1cQDZ2jlej/lm43MLVO+nhuEznI+a
GshMZrzUsAOEufpOYednbE4TFa1v7iD8hbbH2FlRvN4LHldPE+xjCqLLkdHrMVwm
p/sCOMIOT+ItpWmUwiq+riJ5wdoB3sHUq4jTUrr+wTuws8kjzGgNreZngdc5ogHN
v7RuEydo4cr/0deaK7oySZXCUBS9Vurth/HGB6DGTmjmDMjcem+SgbHgp0XZNYhv
n7ulFnkU48fd/Jl9OyY9wYj2mSovSnf9Wv9RyxzW2+v8d58aZyQXhX2fz1KktQkF
k7FxFWh2+S4ru9FWpLeyBl2xA/hAczWx1Gn6OuZzvgBj0cbgg4LIUwqjWBbap2p7
FNSXHhEaNXvm0HvnK+cQjO6wZNdRf6LoPByLhqgxRisw/5EXBdfjdmmnSq3Asrs+
4wBrAibK6M7aR6SlGXWrDlDxIxV4ls4L8cqyGpF+6z8hFChaszWH+OATUqed3GZa
AqY2l2ZiL3q3dxPZV6bltMvlqwVJjx7Yi0RCQNrrldnOezVEwK3nuJryYv5CnCE7
W112imGHvJ6CGXOj21e5r2Rb2PRwOn62v8ITu3eJ6X1mhhr8YgruF3Iyp3Fltagu
ICoKkHuDybz8Ve/nRVG6DJeRnKGOYyTc33dms2iZ5SqXvzYif4NN6kSzAbIHnW1A
DmTS77XhJ6vRhgBgMjsXri/MD2eHvLs6ElFbOIE4TIP6WNx2G1H5hSVDxPgrJMpU
L+04g9+Lf6f9gVBrGLu2XR1aZXBS6ClloI+2GN88gxsSN4Kww6oKqWrWvwTi9Jrf
bs5T+AkBtjvmC13Dot5codTkfqi07PqKXpxO9BgT7y+/qhnke/dXTTN0WaqW09TY
1H7sAQNMgZcyPuR10fJcT2Qfr6EGVxSahUCfmBeSnUEJTz3cO1T6kPEF6I2fqFMa
S1fJmIV4pYiejt4KikHVonujhtDcwh6RJquoyE3gbNn9nJWuaL3fQqelMij/bKX/
7v/iWg9h9fpjBJ0DAMau074K6XuDwIOofe/9vk6tlNnjz2QtrsxSyGHXhUXactwi
GK/FZe8NpWNpgcT4Kpgmrtf9IK7jfVjZquDRcTVN+5zIsf9Kec2L3EjRVjXDDh/W
nPoUVJuFM+cL2+4KMy6KcNdcholYmubjPSOwiKa8L4kWgHTTdJrRtPYGULt6qEP5
1ib0OHpIrbSCICkGZXnWzdi3uaYlm11giRaWaBsUP5cST77tPu96CsPoy75ZpR+Y
BsKtwuX/hjxfj9SpygVf0FZgkfyE6bm0KPiuA0w+SyQ1fGJyBB6qGIOZ/ROfw4T1
1hUIJonhfqTpCtXx1FwXPDcfUNWI973hRTl8mOw2yvi/YnvisM50FWXKkguten3m
UWSXU9WHPNql8SrMOLY6AVh/9HAgBm2zrDnegRpS/jbxkb8DzW+HpIlKG9cN45/O
t/1sZYPlE9+TQLzbRWp3//TVBpEbkVfjc0mlA7FK4/4livUOnoTg1Ubfmhns2WiR
zF1q4P57FNaDeIJ7BYZDeltgjt19ArqFVh0CU70m2a1LCf4ls2xmaTy9d2VT6LOu
azzEeU3J1TRmOTuMOkTvSrKMPKD7O79uw6VJ42EOPo76B1tzs5SKLSlFZnN+pfAq
CvT2XGLSodYol+ACTGPexvuWCYk48X6dYiUIF4ny7GqmufcZVyCAjwJ0JWKREOml
/eq3/h8tyiZo6N+tw36zWnVGmDC0fEpK4+eCLKX8OpljaqXZQOKU+cZHuKis518L
s+NyawTyQDVcOfRUaxDS4M1kACFMckqrdfnBdnO0WAETmKf/5kcs9G7sduq+eROu
nDfkKtMHg0IyJ+UbitONtqZ91vhetSJGP3Pga1KasM6lx1F8j6RKohLvvw72g0dP
Q1o1bqPzjYA65XZ/NwMofx4XxNxVB04TdYo8P/RwbhFnGksdSvcjzqC5tFoeQnVN
F0GJlWfbi5tEUD94u+1TRJnPr+DdU8wB84oAzxeC+3UBB2ZVr6T6pvSm7qsWxWHm
Wx1RlMB1DjgZ0xLN1Hdsuxr6o4Mi55AZh0NWLj4NnpM0dvq+qETySswzBh52HSQv
BPCuYERLCcH2xkh5z0OqyrGrLUnQK9KTldh8Dp4VmutV7+sdm6QI1kzGCEbF3XJo
7Wlud4CBOVNwQCelgTtCURyAH0Nhtn/dJxCEKCPLm5MgFDCconAR8FHeGd7esabn
wRKOttuIN7MdO8bPHLRSRI3xR7GhVNpR4rF3fq51fC6QgQSAPThGnEI4zTc0lbiI
sedYqAuRhlfdVjKOQR9gLA+Istwoj2A5cpQYSK0lZ82h/sEUQxgicmFOv4QrKDKy
cSPrWjcGM3/nrsEzsQ+ryvzGYRdSmLj7KDPmnUSzyEXkrXaV/w3xOl0EYzoLebn/
tHjyyu/SdA68QCfkLBjge7JmhfLR9Ka7YJnGFV6FuviTyJgFCeAa5XJCMMmHw/2k
1xgW4pSCqtgYilMvxiwYsMCsY/Ym/70IUgSNOtD6HS4CzSUrnXpQ5OKPnqW9OG6u
5MuXSppWL4c8oZP78H/dRUzavVj3d1H3YQoWlFFLC12+l7zInbk15RyJaIeRv6+U
ZSfva5IpEEJIrHj8Fn/uK3+/MWVIDe8uqixlr22v6zFzfi6yLCEYkzSwPqgGdY29
dcxVqg93x7yZ5R3SVGEpOfyhh5BumiASC17D+5m4Qjo+MxrDvSHw0ybyCLTtluN3
YDcTzFxVx9NfTdqJImMYGo8ZNXylp+AOkLvUAIR9B4NKsSzRbJBBjT4Ecx5TxJN7
usHuY/amMpQyTpVGeWi0uRPyWbVdGGHudF+FKbzVJ4R++rJCkGL1NSLd7KsmbGqj
jHw6NjrOUfZZjrbfRvCAKW6aYQN9R75copl8Oaer3Sy25KPLPY19Q3JFh/GqY/CC
YVl8UyabUBnGLWrSr18DtPVBiKeapWcb8DJAJC0C5+XAB6Ip1vALS4KOIPhTOEIR
dWjxdM3mbDKZ9xcmnWQa3M2lubWkLxtTOpo/H+WG0S9PmlMqZHHYzZBrYFHWpck6
i8htDWbcEv+kzJPkvlQiPD65FeZJEYS8GYJHppQKf7vEDkOFceiqm8LgfnW5sVDH
wbUh3OwCopmGX2kcq2NoDS9Cbjh4F/VK2ZseGL4pArmwCPC9EfNRXHDdLqmu5COf
hpaPTc2GaaU4JbHaGSgWLuWp6TLt3rEnGr6mowjqH3/eGJU1CbY92RUYxvMy+GN9
CH0llXkVg5G7mVnl6tVeTOq4RaLanbZwHn3TIRXxsZpxZNgKkJyKeB0G9mITb/Dx
i6TilUX32ajh0KaPDLPh0oJCgSdIbyG8UWSqbRT4wLayjqM4IpxD+r3IH9C/rfbg
cDY1cmqQKoHXfhvxA+gZDeq6PIy9z/GIPA80q5YZocsiEpfUsZz+SQ/XE15Z/zxy
VJoLKjTjUmZ3vQ1TribvI5W9xKi17fIDNxsuzOHa0XMv19hNvNVdHg1u1C+QpmDl
YKWNX9gkpqo9gcACV23QhmhvtwXtLWcxrTn9Frnl1AYabFhe2Tmcum6oG1Ki+gUg
Gi4qTmXc7L5DS/SNHHFqbxKMnWViyuo+Ysa2XYFUVT8ZTJg9cxew3CJNBX/3LtRo
J6Y5sQ6hdESItH8sLzLSL6zs5M2ArOaJrlyIQg/L5ERqZ95+9sOBaW4jVmtGjDMn
n1vsnQzr7UyJQYE8wTxMNVDMyhbipFf+UEL5+HzuV49DCJ50b4XrkftrNEqBFcjE
uNCtPj+lAWh0thVqzrnwHLK/896TKHu5xmGLcHvMFDkThr9hNpJ2PLQh9VNVcqN3
BH4/UnUp0FmkCBsTEXbKy6+y6p5fhUs3u/3IDEQzPX0j7zt2ZQLnoMhN56Hbp48d
JFBE2FrA4BeFuSAHlmUlOi4pjonfDRJXQxdlhKBKsrIyIgxIGzu2ZvECRpbdwyQu
b1hPv8sRQ07XtCHU3gPTdYc1kmUIpN0T+cksNM4w4tqazl+O6JrunMe+hFL7gNA3
nMDLuSo/q1oo/62CV/433Z4HnsB9K272GpwcImACyJ779UuYD82CLCue25L7rYni
pWg9nbE8JclOI9Z/CCLIJ3/+3EOeWsCW0xFziPiZ6swwTJYByJo1PDeMJ19/qA0M
rAvZnXN9qH0Mpo1n9ItiO0Zy9mK6jbNLDYKdvs7R+V+mO3+Zggnaa3xb4YGhRcNI
+QaYjQch14+wlx34NUwEN6tFu4RsgHEu+dP4qG+UN+8OKdJRzXysovT6bJNmLGqO
3nlHd5RmDsPqW/Ccwd5qnrX24wqI5nWGhakO2r5yhBU/xHnUA/Wg16DdBqZedbkX
27a8bF86WurA+umFEFu0djWTKnKuHI/Kb40F5YeYXXtpY/URIQDvBfvpaoSGio5t
OLbOsL05Ty/FD56DCXChbyCWV4Jw5E9pmOUEm3r4mVUMZ9FY5J0dw7ti/aN5nfFw
+tCC+yJi++ameDqfpRVeGiftdmuBPDd2lHXQsG7TpZJXSDYJrzRKJsjSjNh5gYVs
JwUg+XSSHgD+4F7nr/ICs5g2NS6cErRpzLMt5YldTL57fmFStQBnKY1KH8ouLbMr
Fg9Yico8TM+vClrEaE8WijADEh0gTbGWswKK0gSyirXuk+voOfWdmx7Rrt75zZgH
yJe60c6Jxy+wfA2OfVFhjOxjvJ7poDqalY8I/Uo5WwesNrapHnSQ+Kgy7TcoY4iQ
pe7A3xGMwQT9DZPVKE1LXT2meLdT6fJckwmZtbFSxQottG/DwVYSab3Qha9yQ+Xk
9GHm4o057vbI81aOB9bynT0FOIeQ3HGQEk5pF0mc3VIkvsnaLUbWm8A2EpFaxzbM
C0McV32bYkGAFwTsTJXpQj0b6heoFJVf6HrNOxVCLtaag1n3qpRorS+FtwAMZFsA
lMyr6v57xsc6c2JhUH57kruY6/kO45ZqvZB93Yr4II9JdxlT0zZmvjYN5XjK3DgJ
i33s8robMYQgubxLkAmIVJNY8o9G47gQH9zA7eJ4xH7QN8ekAwIs/ns/p925MNgX
IOBHzUWW2hBn9AYj20Q3l9Wp9EjnjR1oj8MHwiHUbespYTQj+6V4eJOkjMPjj10j
SUW4INrdwroYbfB9BKi/QA/tZVypwfr5DZ8Ag7EMTYjRk+KPKFkHDk7Cx1/5v5xk
AGUgd9/WvuEx9UO5Xyr53mGNXakhyj4GOd+XjTXfSU2xyokVa19t+l++rz/+V4kN
m3iI7IN2+KyZ3Na3LdxPsitms3tsoUFeZXlpEmwdk716UOVABUwx/XL7+XT94lYY
m/jTCieQPy7YGAWqZZsXj6tkHXjM4acGMqIw4UB5q4cQNkhnt4rYJwGMLDhkZEqf
vBFTaFgtLHgZCZI8qrJPnl4Wh295+MzImFNvlXNbf+XPp5bK3YGAnNBhGmd0cLqa
QtrZ2Y8SSu85SwnNKW+zOtDO0pOfJTON1vHgKVGU77cNlIliTspq0kUtPGVyAHuR
/m+KCB41InhV23DxHuQH1clakJ7cc9Qv+7Jt7CkWxAk/J88K4r/8GMVQqYzaXCP6
xS2lzhq2jr1mtx7TTX4CHsI3zoh/Taz+Sl5mdH0d1GPNZKN9GT5RI/lFSFuDSX8j
MsGQeMGAWq64V74P8F4Kh+h/dVSDPcE+xQaxV9PPW2gAfi4LGNpSD4QNQVt4VpAD
gJSxu0NtDffUbuOWkQVrjplc0twFkJpTLQ18+XJoz8F/pxsQWBVs5QtSyaZdxwWL
Wgyxbjt7IdDE/wkfhkcXTX9l8CC6tzVBFDv4Uup0rCxlniSFH9sFWaYLijRwghRE
bsLGGsD+287wUeXIHl7mzl1vayBwRYItwMmd4YWjYKioL0gmyAWb4OvJACSKPdAp
mTf+ja/bFCQCnpoONTZ16j2ZuMkstsdNtLckZ1qxU9Gir7EX0Y/r+slFdM1AR858
iQOWPR+fqyD+hdxhEy3ZNUj6kxbKyuYUWxabVQaj/HqRQ9KJwphBcm0EsXvfJhGD
jWEVuWp4LuJlo9/LGVZ+DJdlvOnEPtOjGgRySTwpfSk41yvXSmSuZCXLUj6SC5E9
yPPwg2W1O1QeDh/1ZdPwzjYmkoyfQuSMLnadoQJaqaxVgJ8aFZ4Iit4YufDbSU7/
0uuX8tRTKRSX8HHH4+4hXoRjT+r7FSOqnKewh6uvoxpbASN/rGgxWK7zF+KTzkjW
0GPeAEMr5Zl7RlEdfSwxUoxts/W01KUxQdkaJub48SDfFz6kHRskwk3DVnKlM1Vt
gvNDwCo6PuRKQ5bRpQwE50bDjmmm0tUKR6OCo8DgkdMZ77BpLcI02xiCHk69YtN6
5cNaNtId+QTvLfRDrtNJJc8S5x+VdA1Hzp7ED7FzIuBc/35lFNxPhdMtA6nClSg8
ka3/7LK58QtgvZBMfi5gV9Ugv0hGP7Vi9JhDOGNQBfKiBk6RiF09p2YZKgQphKyD
D9h6whzjFdvmsJOOsUbAFq+7ucRixqi9IW7o1BGY+flPs8QvTedVO6/W2AR+LheL
4W8J2YmEH9KCUR5uCyWAqy4V8uuvKaOQHULFQ9SxBrF6ByMh1/P2MgHKQbHFSlt3
+dRkK7EBQ+VOHVE+/fDyJOHl/VO0wEhXwZlQ1BtDLcFwvhG1X+oPSRBux1ElKz1V
vVq8RPhmK5UDI3gSzjzZOKu1ZtQZA4yP1l5olzdTWZs7avMUTBs2vE49oF32DWFk
DTVWkwJaIwZh90QfJKuhJeyymJ+HsTqoD3vb+t61PUlrko4g9MBFBoArOFX+hzby
/I/4A0b3+jnvmhPuUHnEb8Cknjaxwi0i3fU9dXwoOuFA1Txep4h8+pkK+/EGGvY/
+UlGpMfTXUPc5UX7aoh21eRfruh9jcD7TkRjqWBiiS30utoqPt4VnCrO342aiT/P
hM8wIeAPlHMvnXi+wFwZKlyNo2ZFXr59TcCXKjQVW/I8MQLjP3dqK2IJmF/JB7+N
rfXqjOnbBmqylJri+yN9a5Slnr7BRrITdQosMaAG7rLj2jCffaI5ioRKiImm+ZFl
MHgferiaCMWbpLoaQ8TLfhjh8/Pf8BjYXKc3ex7xkwIiXY+Dqdub8u0ZJDfQjCCu
FcPr+At9ukkUEAb5p0RS6rXtZjA6uemdqAHRN1HpVSNdik5PD8KI3NyBQLszKx3G
bgMhAa1YrfRb6nO1yVYlOXqvH5E+mQLiNa7MMmIg1KAeadXs4r/mj3Zg1jJ8VJNP
8SOFURY0NLKHV8p0fwAlXrMtUoLdyCNI1Sm18CwUwrphBFvwErP4ex8H5rStdCnT
KVSbO1ol1J3oEqqmU9ujCnD0Bwfjufc7RMa0OFPCWIphdypBwApoiDf8+6G0EorI
+LGabuIdBhC/oqxS72mN+IxqprwZmCcXMKvcNFJ2zMbREBikgCH444XgxwDLS/vQ
R17MUK4E2w7E72JRkReZe3RvAOPOUo5CgzBWitOnh6jwx2i8p7QuK+JeEI6/5ble
AgvSt8iHNJ4YqtfHO1P42zyL35E+Ei3bECcDRX4v5pJwVYX5qGwj9AieFZTSLAuK
AKnrSe4GtoX6NRSRmYoaKHDDRK1yT4eDbvw7wCTtbLFGoghrS7qxkidhK6lqFr18
bAVp3o7o2n+yNzw6q88qbxEsiqzQz0VGeX92qhTEm1O2cWdDYvEH8QTUUOtHl0rX
Ce45xejvcNumBKmmjw1aAseWt0aQ6DFvoUpGuF5TjGnH8s82jl6OCjfdSnOWvyf5
Bw8zTzWQpXNuSc99WMxswg9GywcxLpE13xphJUNi0g2PWfjZDXYaQ7mshP6K0lVO
odVaySmuZfbodDZCT7dZWWLQE7nkGRAdOW9xK/9x5uzWg4fyrTZAyPOUKzEi/0z9
UUM99sSSK4t9V4Gxjjm1lWhMuEnw6fV3o4pzj+4WrOqaa2OIFEusVEq8p8FVJmtl
/wU+FSrq0qbD0OtCF/tbKVztsJILw3qlhnbCos1AwzJfxjlrwwcdkRUr64oR4bEk
cDRXZSo5gLnOILKq4yctfKJCmw844a9AanOSQYjQctvY3C7ouibqPYqsWu1+gdLz
7XjZiP8OUPZPOh1MKfREZEhtM0BRaQqI7qcRhFz1SyezBldCaFgqWrPoqTaVayy5
Joy388QqGazij4u8TV2lKvlaMvF0P87PbvrDJxR7mRQX37oqYrnJNlDMBOwgr8MZ
lCrEdB23qYxzopbOma7fs4LdWVI4/V/P2TDlW70zbfzwBp9+4bLecDJN7Tsd4u1N
VcsiSQg6JzDD91mgJD0hUkrlyMmUQzpjoFAsumyGn9RnKQk2iAI325ecrEyXGhUd
G63agUboW1CQYQNlLp+s3HDRZfaLJdCKK5o6kCKo2g92j1yDBey3jgNU1BaqTTUY
K5PsqycdujZn7CQouChLEtFOjNVssQKy5Aqzn4AJs8rmwl/6IjxcE1wPMRwDwpo3
7Q2dfpZVfLoscZOAmmtjX9wFWeO8F9Bdkcn+aYKL/fDrVGaOFy8MEgj1+M2B4w5F
VPIyNLY8fNCrWesVJBlo/JhS5p+xM8mH1zLlZRiAT9fg1ejI8NSwso4tJ3oKoqxN
9jaf0RH8JgnMSUX7JlDz9BqRxJgqglIutV3foG03t0awrOU0ONYJ5BbF+tr0fKhs
Hpo+SufBYPIiBCd4WBknlXGLytKPDzcj9n28OFgGfoLdDf5PUhpxZMC6B9jgfuwD
rYEaUAovqnV5AsG0Y4fTn6J5HvFTJLgNGwY71aGDf6LIeAVWOSxeuBCTUWpatLTI
bzqZBhQT7G2EBovggnMQxUIu8kYbZG6c7JuG23aF0HmIMqNseh76EVc1aPWXtd8C
AJUlLdfrXYtxIh6SXtlhnjM461ZZ1nVEPUKif8R9ZdnMa4wb7S3PQPfqe1HsLWRy
1ppbRolyMqJz8SOs4zSsgC/eQL0nzBEBG0mnhkhfhzKB/v5MxDpW6g1PPBu3jHs9
jgK7+0h9SqztIzHEalelDQVqgyEXWemu2DQfwNyY2SNHfWV8i1uHFRTdINzb/ZIv
tK4yua1z9DVSEqhl5jdnsURIfogYagTrS5cSLgpPjBzPaNi2rfWeqJ0iaVIYxeGT
ULYWfUzWadTvy8qu63fNNZELe/dhDvXSB02UX6XDBwQNA4xDaR2hCj2XaNBSU8K5
gOsECdnPbCgBAfmo4suWA8vGNBFHcYQvqQlsB+lJDrIQT9ZofYcFB84LdgYxBQcL
oYLslSfppFKpT2I2eXk+o5W0vp0KlcU+VUCZuaS461h7ANa4Wijpawg4vfHfNeJ/
YzN/rYX/7Bcb8tGgdo2HzCQ7zflL4cMoSa5dty665lPTpzsGvr53OeEG3XIIbab1
yAGkgGxpavNA8uLxoBa7Bnmmcij/FKMaLcXyv8lV4afLXQ212nkJZaTjpxTyoeUU
9AQ1cjLJOt5omPw9OJ9RhCcgSMzvxz+6rUEpZLYAqfSKNAymlDJHqKB7iYys1ANm
Ti6WKaeXL3S0tdGoo7NKcuD/V09Z5+hITqETTo2UQdE9Cnio+OR3bNY9GWZq4MXB
LlHlQ9vnUDPjAkWex1KRwDNVmfeZEOt6uFumVEIp02Lh1LtYOOer6QKMuAXaBIid
RY47llxqvAxyy48jHLKKA20Hjcw6HYGYVEj1z8rdunpDNel7LuI/1uJQOOImVpoc
EK80uV0zogu8tbez6UCzfiHLuftwpqBwl7reUrkHBNqVNtePZZIEU8KG5Z15HAUZ
nkLVcjHREwb2xiocpaOk7+R9PZFQ+exKkYfdWkUjmwHjGYZheCSBCt/Iqu3qaVSh
UydTrPUTFdF3zq+AXvtcfazxiBgU1b3lQwb90Igm8fP9xo+TSqNGEQ288e/stIC/
mTpz7ZKDglbp+qsiAasckxTQ/LztQlPdEdl78OEP7x9F4Ov/onvglqQ6sXcOtA4c
+F2oBXK8+C8wOraRH1t1SRFdJVhiJAxCclgmdf8osQUMeJ+M1JigwCJRRqhmQubi
afLWbaJyLjzeJVuUoayauK58jDIpYH3LppYnPW1uuXRkWrl3b6mMXhN5b49+LfeK
sCw7Uvxi8s9MLNKXuYGsGC8NTNKM624KSrPXT5uG2BQ3JRWFYVJMt9Px19mk+6RX
Xh0skCcrO/2OWGz2UY2g8acYB7gVQjjgUrSrrdkkpCwjOyOKhenrvz0778VsON8H
R5KZW0nTin1hSmawqXxgPqj5UFvQRGDgE59J6AODF7bfoW4EZxC8toFF6udQfZOE
9u4hWPwssM/6qs8dJ18iN8VD8Yk7u+glB8tjWGmv+lqFyYUv0OSOrfsEx7h5CEbB
+bPUV/bIb1Mg9H4cY+j+MwtKmh9SK6AOb7pMR7CDQ646lqPJSdDVSfgPV7nRgS2E
j5ulYf6JFSCNHXUEBiZ+xJF+b2EU6kcGncCN68zg5fInGvhKFpl2vzk/2KFcYvwu
lD+Fp+qF4O7X7kDQCUMibeGHPJgQxwZn20b0DjZ18pwmE7r8aTAjKl86+Q+NYnWN
UD6IMMyxcG1TYpUh1Et5UET7Vi9RegJaYhA5LGb/z4xJtYCIenDnV3DzJVeK4wAK
onzrgrZqE35GVSIPan+f67ILVhLglt/d3V2K0I/GJo70AxnFyU9SPc261dATE655
2KwhHQMruJFVwxlz3/HaO//4HOS2H/1SF57FdY4leSZ4/U7meoy2hVaelLsVoLX6
MY7T5TVmiLG0miBKkylwCPNcc74a4/T7qF/oddy7fywV7+gINwVpVKCM4klmOUu8
3Nx3bjTp4m6BVKyVZoWQhU918JeVqdWzRUzV4/Sf9OtBsrFG48S1W12ngfiCxl2w
UyFzl/rJr9302D91FarYVy4dF63ovdcK5KM+KK7WqV3+2QNbhoFm6iBrToiDVpK6
3dahL0v2e65hbAUcTs6b/DCoFv1PEOQAvVvIZzy0PHXw7Qpq/uerLh9sEClMdiRR
gXmiVo9BWp7umc7/dd7LHNd9OvggNjZYOXDxg+stesRq0NchOqAu8neS8bw3Vjoy
mwVXZsGLKQpC8JX8qj3eWyPC9YtrAYx5IM0We+0ZOiBVDo+8lbzxwdDCwG5BdOnd
hDHMTtzNH6oIjYNp7RGv59LnZl7Ug2AlbmVtVbAFHkeqyJMubcyDE89vjC8WSuY6
QtgWuqbgSzPYpvWK5FTfV33forEwhC9zVp5xoZsDInzcZd209gWR9263aF8LWOWd
yih5UeoE4ze8hHdh1DuL/MTI0GrjH6UPw0a5fqvNhsP2EizTtcY7gOaKlrXU56K1
SrTCKTTtiHb/gUkWvgm7a0sndyCvTOU5R4IYWe3aXUn3zfIyCMD6ovlQGTzee8yL
0fLkeZQG8hghKDS+jbXlI5RoIcXX5F5j5RRqH02M1lik4Km+3x5aIMYdbs59egxw
B1A0YvYzhTdDPno53OEl11mOTGEPgXGAif1xkTwxQYkXTYovKU4dX0gOA2C4XNnj
yM4b9dPJCz+TdAns+XqiZFHC+lCdWKSIOz73B3NjH5vN4qhG8yqnpWdgJ3Wncl7/
PhnhABigNhSpqXLAu9Vqa/371YGpDkOa/H1JeXFvyA43Ig3xx8gQc0rBMx8YB5Ak
IuVmnS56oLGqtJ0DuCzJsRlYtAW6Xc7AP/2UPsTaPedsFlwaTh9MGisqD+9JNikU
qmQ2W/hyOQo0G5qJRHNJbMEsVLmDzV1ukVcvISM6JzQUJV9grlmGsKK74xkWkwAp
37OKG7czFD9bddDzJ++UtoV+t+2SvotfKWAEukg9Ef6DuH1n9aBrZns1nQ72v7kG
KAslQZY7WHtA2InbWAVRvYPDv4fE6OKYUJZrSMSdvO80I3yTygZwGRhjfAj0bH6O
SiBjoxJA038blM9IOKiE5Ra8EZgvoBl+20ZFqM71Pdy/LaX/5sgzAWEZera5G0lC
khlRq+2HzsKak9XHYXhVamMih8GmX7XWda+Yf9g1gZPkMRt/85EdgUIwnubAwYHP
gMgsASqoDVcNVdvN9JQ4XW1991JoqnV1HHq+M2KSzG7B58WTtcUg/331pReiBS/G
7VKDqpIVYNSuxEfVWwDkOEdMJv0Cs9kHahMtdy4qd6g++c2p9jzEpX5Ip1j7//vm
4sgKSdq4CwXNxOGKNEdcXTF/NM4q4qKqyVatipRw4XhNrETAhjgeffI+BA/A1GtB
T/JWF9deaSdUwRuAOHh2NvrDl4NK4DUxRJhokJNuLHGM1Dg4MFf3Y18Zd7gQOr1y
9HgelbhYf4HXkXha8v9Xm36l2lfW99W5lTZ8IlOwu/vlV7eBCemyX0BvqA3omcwx
oPsQ/SFBwtlaWvARZW6GLzDXm/gWFhimXgdLwYZGciLtsvlSBQcHfYE48KRi5diz
I4VBORJ05rOla7uUubwAgHbGeqVtD3v9XwyrHG6p0gCZYcATn7Z69vL42efpJPX/
EiyrRhYjDG/GiPAh3zeGfaP6CQLwRHNswvjAeLbZ/GYMi2mc5XXf5nlSNIpkcHlO
RoGAyancRo2ganlqL7qv66G0iqb3JnrbVsGCxyL9WD6XpuD7mV5EIp4rXDoYXPvH
6bte+j2KklRubHuzXm6RBZVCKgLO3TSsGzra4qRnr0LC82nEj6iRDkNs7XzU2Nf1
AOJ7JpqT2iNFFCv3H5v0lTGKTWUqiOTFWA1FNSzNrkDtigEgHMrsm3s8+i6nEEus
E2cZrMOSVr87md8oFN/4dg6rwYxhXwPaL1ZK6PN3mRjF5MFUv51KhywKbBTPaHKl
TfNsk4SHA+f5kos0fSVeQRAgbPRVCMDYBm7HMza+CABwm8+w+cVhaZ6PWCK31PFv
E/5bB3B6Cowo5vtOuD+zN9IIIz79RHvux3+cfvTeWz/mwBIbdD8OpZmz5y9QxyNm
TGUrZ0qeBwT59qEmiKpL6OegElAz1NIqcZg1m81Z1p8kaL2xeRyBNmGBV5nBZs3x
/KGwRDBCF545gZedS9rEhh6w1O4OvxWRMgBbxHGs4Q03Vy2eMSTI7y7dmOu1DS0U
yKVbjKvsb6JaAnKu96fiuGn/wTHKwHMuGhcfvlX70BBZEnZpObQDMhrtPX0uDeym
x6W01n+ADWmeEGWGdxfT0uLY4nZ5aDecbz4R7848ldel3UUXOXfM9yUZi621xEgc
YEBDzPBiGH6trtCgHaWX9qfgrlUVjWoJ6WaW9rh76Fe0VrirIQ8jw6VqWZQS3gT6
4HLB3qTrBZmG6nFKUwkjvNMEn5T/Eq/f2DOht9OOSlgLvgzDFAFAOMQysDUfYAaW
icyC7UZ5hnGGs6lLKElI3w5yTpEsq34qTmjc2eWVJ0mse+yRzVyCDNXSraTxy0/g
F6pggXUIMfUAwEptwYY1skFd100LZofuyNE2MrQ9PK7Y0aKqtWfLmy++qZe5OflT
TdsvkUbdE/6Jh36eMEmaGvlvVX8gGlgr6zQkcxaM8fRi1oTNcuL+7WcZbXrjMwsA
S/pT7lR8zNlz7rKCKBhp5kDyR26+aD43hM3my2gU7LenHYRHjL9tls+YiVaG8gxL
D8smI/1pBpubjTCn4S4ErRWnx3fuYtiv1Ro2IOsdhn/B5/ioq5s0fARFtt4IUTkU
px7w1tUIELntZp7mrnwOrXOXJ5Dn0PDwpz0GXvybviZxnj1gWfpmZin6g/se768l
1X+Sq6ljin0vI8drjnjYvgaC0qOs9Rsg92LASVV2JsHk/7IuIaHsWFqaaFc+CGDS
xI6A9soqdUTQ6S3cdYJqCftA1SP38hSQqGqg1SrHvcFAXKanQV/7BW3oaCN0t/ND
kBglj1zlFt2Uyp2f73+c6H4/fKbgvLL2bijbP1GgPVfqsIAo+7On6JSbrIWJZ/I+
PYkeO1ZDnrSNd5BJfHhjogRlLvMQoAKUu5QiZIPx01jfDwZxOP7gKOX+eDAP/4RW
caTW/laAMIu3KhyMVtrr4VTKYixJX+5vtI6d5DZ8ruHHeymtj9H5nGiiXkcuHImo
HHg3klJA0+w+V9C1i8zfwuu44OPwc2cJPWFEtM8JevFGqMgtd0tVBj8wrCi8+T8x
+vj7N0LTCYnbQNFYNx8t9xMmcJVSyB9NEy9O/AxlB4NjqTGMeSjLSKsqzlqEiyXt
tYB5WfvxXwU6bXeFAkV+eqWweH0CdfcvMXRFZVg2pX4hS8Y7nc18QysBVHFrWemo
RxPkbWYiPikDQyfBfKORg2T2YiV+jJc2JKtcaLSxDu0A5qxHJob7F5WyVc7Noov0
9tHr+gJKpK9NwA9tjgvGrQ48WarnNd4djqS/VevwlPhrhCkyvJkbgYJXhLc7/f+1
oPJq6rJE4xXsbOVAtLkGCh80cFRH6dU0vFp+cM2PxtCcpM5qtuff6WJsi2o/EnuM
IAyvRvmvN7fTmQ6Vtya6tw2yEfE+3rK95I04bWhg3saICmXTlA5HNgl/UALzvCep
slQQ0SHJNYkk7ylyIem1UIsuZRKycv0+C/ZGeyUhNkpAdfYuR8suctNC5Hzk4z8w
aF9kGGQ3qoQnB45HyDzHyrgk2N4cchbcBHHeemNJrvkUatbpIB8Cld79IORJZi65
oLZUbF2Przd17AuduuYRr+TJkdUqa2VHSToPWhLz2864S+A0nRaWKsTs3dBDxIqu
8DA+pA7AALjgeCJaPHqPcnNtz5Hx3WWq0hRIMf/qfwusTTJm4FqBIOsKwJgYEIiG
9A29xsg3YWLVGkUE3UQK6LXdePBSmVINHXmbywo//WDKWc3JYpeKcY5vfdbqx0Wl
TscytcodyjdaW7Ug+c0TSscuFcXLzgCwU/tX2y7sjQgp691Fa2RuA66x+4AAM9Jv
Xn/DKgdyyve4QX26k6OIsN2IUloFVVOLitT3ovzVt2wzK6Edzfhq0jFbW/x4XAzZ
qiGzScnyFNZGksuMYOTMnIX17PQRqhQeuDzX+t61HYdyDsVeLioImfz8JFrXtxfS
Cf2r3PJjr2C1pW8szMLS24YRrTsevnKIgjilxbjqnyPCxxWAd2KcqbNT/UZDpUiX
pKzkKlvtFsx4OM7GnqZRsPUD/hLFACpgHYP9zIuSLv9fnLM0V7ngjS/JNJm/ajj+
Zr/4oU892D6l1ECd5oFNdl/KCfwhs77TlcPpIocCq4Syozg4wMeu5+ARAytmfi2b
HI/AaH7XIMHIGByd5WEg5KP5gEXw0K1JunkYGZ1IShW1An0LbGGLVspEPjIk0iq0
+8dFRYPDOkKIKlyExeQsVnM4GxJXpmdvWRzrF5KqjVo7D4rfRxhdrTg/oEpPTsbd
2LVodA90HdglKJoWOcRPwBkkntAlpskLr/Cdw9ZJvlmmaPf4PuCo/9NDIPpWN7DI
1L/+b2woQbmz/El0K1wTHAaS0ypnN7Tnx6jY5J83QtJFzrRv4LdyJBhUOpm0SsYp
vxb9Gq85q/PecPqVORDW7qaJXVhpBaeQAv3jYV3FGgr/es1lByWzQwRD+ZimHtiA
Oo3BpS8ObobbKeUTH/1g3BXv5K43qG5e47S/vViVD/gcuKI9KYlYT1OKjcqg/24U
h14+jFIpZpN6czBUyPAFhBlz+Ti+o+Hd/tbMixDrljwOnPVkCZZBT7yOhqEr14uu
9PvM1UmoRSdrBhvAz5uadGSz75nT7XxyL6oIWasi5ELttvvjfT9+lq6x+AvYQE3f
soc129ZqtOjWP6GbMV/SP6QMyRf/n/+4PKQRYR1qLj55ANTWEqNxsYLeQ2svoXrD
awi4kBU0A4Xqesw62CLgeu/rs6qs985BojaUMzLdmnO9EmPHJF0B8KFRLyVY+eD5
CRp9/+mhGWqhbfpsOYwlOodimR4cc0i6D1SP0yeY6CVXTDpBQejb5U2VaWI4CIYA
65QLFPVVkfKFa87elosGpyIXH14yIUNV104U08C+8D6lhje2MzndoLkifN1uU9fW
xPdN26H4/s8DlmwlZR0Pma8dUT++4CruBGhKCtd6AYkytkYLGeEtUfIkDnJ3sM35
3kr1IXT4H6qt86pAJOac/w/zi71a51my3mG/CbDUAOnUmuje6ioulx1E5kYjzbBb
dg5oBC3jgfJJfWggvVBynfqap3AoWAtSZGG37q626gt+RXexU3EHO0BEIwHW+Gpf
ExSavyMASp93GjhpjtwNLADjOP4kTpP7SvkM28kPBd8odILx+q4ssVzTxcB5LO/9
ZEA5fK4ypkFFfg4LrLf0HEbD+ugAAUFz7QPs/gjMzMePfn+3C/y1l9+RRyP4Ymn5
Fx7wwkwPfzTtXXrk9qTlXb53Vlt45vmm3a1s3uqsuVoIdru4AsjWcsL1gNpEYINN
DoGZKINd/CKnRuCZnscAvU6BlTCIHfU5u2j3iM4GwK1jxc9D1wrXn7J0H18tq7pV
41p5LxK+AM6SKsFWMxj8ePAujhTpJ7KG05EvKVRbKyjLWa6gOyfErKONE0FICr6V
Ly6yrvIghkR3my4AXmRz0bUuW9wmiX9MxyMYyTcO9z4DOygoC1acQap4Zv71g9n4
DioWMMjoELCqfizs0GBsE5HCk/QSWRaVTpQ8TdR8wcVRluQmwP7T0DI1twKQCay3
FjOO9vVLMiomHltZQp0yD51w07IVp1V57rMRstrcw+ehvdvEtQ0LOR/0KHmffIkh
C/9UcfB1I1vZ++p5fTBFqPsklRGdWs147PyNidCfkI4T0OHHbf4o5LsUt8AMDOHS
pEX053nFMm3S4NqF32lnE2vr90HHGHyuC0dUaIIwodjkq49XAzqubJgoax5P0UjK
6W+wa+C+dB85DxNv0OtTWKwrOv1vETeOc2kquvKyUjcojVaaDpAzQqaW3mSj9he6
Z17nMbVKi4zfpTM/+MWJEfvfWdeXUdpqrjas/keE1F8F0ql5ENpj9khgxOzmIapo
LWBa/baifW1RhsBLS+tm2bPMgOXj5d9lHHnyxF7xbUXgukXV33NI75WIW5O9fvZ7
y3ft2jOvRs5YQkTfLSO0CwhzL5eu+vToqMXG08AoJk1l6g6OiPM/nZZPVoytnS6C
ZrXjTKb8nDQYw5qE7e5ugWf14GNyHCOlR6+bCgM+11LSyBGL7WFB76LdliBrO5Qn
vOTcGwmsygiZOoIoIUhg3CLjY3fHpgd+ASG4+nS0hwTnlzh/xfYIfTIX0V5fmXpo
ykV3TMByS3AdgsHWAcA0BwbbMHseS/sE24FCJnHsk7ZJy9kj5fNAS68ckFz7yCov
025FtMcq6ARZUqHrmpgsuWcj8/O7JL5dNT2mQdTnITDMowBLDs44X4LCRonmaUlX
FxYtlorHYGWB6nTVVIAixo3x6+LAzjUkVRUkjY3ENShnXYphIA/BplzJqFk1iJsy
t/j3RDEWmJ7tzQc5zZ2eWEMJ156Hl2iyDieTE0b6THR8+6b8Ib7aN4j/nMwe1iqI
dvSwN7id+prjxg5FlJapQ6t4aPM0LMJswNEWfQ9D7y6iVLHSocbA0budUosn2cUL
OYAVqnaGtllQFs5hzkq1JHdTn1GYUSgx4ej73sYINhWnUr1qm+uTPTCJctOuuyQ9
xFLWu1kIPJZ5GowDWQvWH91qtmslUcoAoWsPJ2XNDxkljKNhJvO0tOS6mlcVruol
AtWnNg3coiWkDqlpJDm863f5Q4hEGzALS7R8wu17FG7j92dASu1cY/3aY78v6JDm
T8/I5U4yIq3PK1rkdD2SU1po9Onj/YehNpJnYT+1bJDrrucpz5NOGhEWXs6dlHMS
a+MJHz2vPNr7kGYdxtPAtHB4IfCAhKqZpwf3345jr6f06ws06NN5irdWYelmGYOq
XB7QpR5N6QZBxYaiK///l/P55Mox+Zw36eVXLkeSBf6DK8VCehPHmHhIM7JKy+x5
ipfzRhxlMXPsIaqgHo46C67Sd4aBgJEMjWUSBY7nEmP9H6ABpT7xRO7FxtPiMHmZ
79//rQMXflxuGDnBPBWJhZNzaEzHsTlwat9bN0BarHVAJ/cf4vw+RB5/8GIN/NeH
yIUhStP4+FtgvQIUJtKhHs/zgq/HsSa3S+tAXuC2oyG+zpstoQOprCY6go3+ShZD
vCFvbCnpuPjvDOZMlACvCFEtgfp7iV7lvVuq5QAGd4vEccHQeHHTTwtBC1ZSpw5c
BSGjhZIv7Vm0+mwIqp7460X6a9cxwyKBSwJDTxHznwObYdaI7TpamMMGHDqztBUA
2iPbDfC12Wfb3J1j++uxzJczNaIcwjfLbQYGCIsGPh0kvnWZ8cf3BeHvnIz5+gQm
K5NI2yKqXfZekMjrNYK5NuDZ2+8/ZI77CB7tz+PIQcmRvMOHjN2e/DSmw67jyHmB
o05ugjBfw42J8xF/g8rbr8vXCgCFxGd+ARUoU4B8JhWlCz7g8y91LNhqbvGkfiBB
zhWKA52wBziUYH/4OZrkKMTV5pljW352rtrL1RW/L7HKMTaf/jwY6BOwhGnRLwMk
ZR4q29ejblfxYGWa5lClfPmKNWrbPG0IVUMnQsC+4n1Am26B3T9UToCSh/zMnRtw
BSsEOJdSHHEiVJ3pt3sJCp3pyTvNVme6IuD9z6gPUCMYXw9qD4RJJW0X6imjyOw5
B3FISlAlChcdobrSV+g2qGf7ToMn9VdSfoZ+3JctGZ/bJJCLNWf9AiSpz7etRW8c
db0r61p9ANS9Vz0br/g0x4+njM08q4AWUL9ECEXqpW5hn96yb3CmRUn/9zyj5wl1
pBM+6hp92PTi28ay66rgraZcUEuL+IN2e+XeLrdgdm0zI7DAedKpcHbwWIHLZGiX
ucxyPHXojpUpTMAD3h16C0cVsHtBrJyXeQcuts9qskgwE4cj8bHB4pTQyjk2UelS
blvWv3KSeJq7qBs610t185gRIsy/sKnOjkAkOLbHE9EHnIMu8oYC8NsvOT3s3uWV
Sc/+dx5WqsnAPNTiyOBTzDJES3tbVSIFnhtiWWtK6X0DQZr3fg/y0AwGx7OZZqE2
ibQlMGExWPISTzlCae6N9OXS4XTSIuYd/HSqIl/CjuutT8p8G7Meq9G7K616Xvw6
4pczwE6C21Kmc7kbt979ZliN01QY4UVdDgF+yR56Xwq1pkVz3HzrqPvgBpUywg75
2YiXZYPwa9qZd0yY0nMqt4Is4D/izAh5lc02XjvlH+xi4Iui9K24yOZSltB3OxcP
VKcHF32tCH1aO74QetXTUxDu7YXVDrAc7ka6AYpHRTJpMw/63Qwsr7hzGierPVP7
xRsBXKXo4ifJ2CQ4n0GDo/1YS7WVLQlE88XhLvMHyYrs1FUvIZeN2KELYzIKnOHR
MnsDTKEybxjxLwo2w7CvLmhjAPqpVU+lHBwEA9ozuR43aTvIUKA6V7JEGypPj1fg
xxuyuINfgk2kKQ7prhB/TzkneDZdrl9D6t6EDfq1RtLnSC/1a38Jb96PL9/j45/T
7dbU5EyF8vXLnvp1X/bBx1OK2Ky6+ckQbh7Y9QyC8VQ3Pd57fHuaagnWy5Opw5VY
vqhiUxV3Hlnlh8PsXlPTNVqZf7A2vbO8PsEOfACvhdCAu6IMJfoJhQS/b4B8jg+3
fgjD/yRqRZJ84tO5rDzC09SCGXBVCoatbHsFloca+/+Dzzqje+WVVBRh+nnkc4Hg
9KEA8LOyV0PyeuL4C++kYk2POOleEoGZWYIg4rpkOXb4f3w7o+yDP83GVeN+bzkp
ITAK2+NM4ZghEo71xyVdFNT8KzxVs9/+35ypQy0+EdK7Hp36zCaPEQ3BVVa1epTm
eQYCmwfSZWQoaVOr5hW1L8yO+y63ZyX/7xaQYGky4G72GY9LrkeqsCuTJFLoZtF5
ho+t4Lm3oTZ2YQLrtF8MLR8mdiYjyWWYdQ719gkI96h9/AXXWgazShr8s9GE/cN7
gjjEMBdOU45asknX/2APGJUb4vnyjNYo9Irgc0hyz/PbJrWBNEHm7x0HODt4U3HD
S+mcJZJAEgSWy1rMgnnT5gsnCW4N8q76oFL864KNUftUJNjmFxvsKyo1KbC5traN
xF9mI10/bNuPvJ/xw+HSin7aWi3RqVeo30XqdRa9DpAQ8FNRwFX/wun2YrzAMtR6
WQaQ8gA6+qpn/XgCcpC1UDPdpcNRHglbtVdtYpIZFCuqZViDGZZ2hhHRTl2epFED
4r+PBFSqJ6ATGi3upJoyEzT4VyjHEFnkUZ7/auIQ94xPVFKLt+4dxi5/Ygdu/qO+
jwGozxBKMVryYrmkgS/5fVDpiiqMEtnhl6LPY90c1fL52GJN2HH1jidgC+x2FdbT
VrdewM60rFCOLjZy2ZEXy+CKuWPAPTG4wpF5qiuI+YDvdAxz8yjRm6P4+mxlR4WZ
Fux6tTEej00iizb7AmFrU4a+PLHmVJSUP9F/SqGI6EIJrnazS4lm+MULYzYUE++p
bv2x6bVJpYriumPxQUDikWjDUrfWlaVYw+GduD1fFZ0sP+cbP31fyNGY2zLAWj81
TvPGanDcMRqBCfR/40oEr3e1w9lSZRO5Blc5ZDeOGRyDEaRSzdXyXUnAYc63JFo5
NJSEmQgY6sJd+b6zVmsNlhbRGmpKj1mdzf2cy/LZRS77JjU7mANW3yEPnX8+nCxE
KYKyJivUjgUi245Vg8MCeOteLcLa4T0B9zHR+h1cs7KNZNecCK2ap00Zh4pK/tXa
nD7WOD7FMhintiMrK7PBSVq1yr5ujVd5SUTQl1l2AaWr1BY15XMwhbR4RejO4b7k
aKvTl0fSrPuWAZdRNNG4AkOxRMfB6RXofXzwzg1HRbHlfH4618ATWPg84fjU6fDn
KIvWwVRJjrVtGhWTjn9OOpNCpP7oHtDkFx0lrPmsh/CDdrjBUgAbPEfAubRngF7q
/joTUSSHHhPIJJSRiFAYfdqUF8/vjM6KrIIdNtIvV2m0FszwOS6DTUN0uJXlxaSa
5H4tyVSbnESptoWH+33ylhUuweDO6TESYEwZ7BEtGbK91uFQhLexcrZ5NXV2IXdy
fqMHL4m7gw8WhCGXlcA55b/qXxM/YYtxX9FIiXqpLkzTxtMIHYGdMtNhaTBMP/YQ
nMxPe912rUwkjHo4sKA5dym1oeQOI/yLao6J24rx03EPy1j1HsPRGzKA0Bue/IET
VwAZf8xXKJyVW685w8WfusKtzp23cSMGHaTwH2m7gM4EDpPdmdJ6Ttp09AaKBncg
2GlQS6i5JxZ9llMYuO7okjP+bvnNrVzY8uReXd6SuL6QhpN00LsYOXPvhwBXc/XP
EG5s2cS0sgtrajmlIfqSMf3ulznmaC5VS1o7KUtLW+8UP/NpRZ5QcdSnF9fFJ2Dq
F21N2GGnht1vv+dIjV2NnHTYQWsR57uNvmEAadwLCc09WbMQA5xAje8kTPQWTXfL
xK8F3JRYBTuZRsATeXB+gsE66wbOII+z3h48chDSWC1xpq6s2qVPzT8krgV+MJU1
/mh2eUvZEYeB1D09GhrhYt5XeC/dUSVkLrzMFfcutB1AsABMO2ECx4GcO3bJVwbL
iPxyWtjNmkUUhAjkAGxKBSYBLhJbGBhD9M/qzFVPBC2fOJDAeWxP1dZ2oecR9Jf6
xDc6YUOG8/vUW476t6AIJI1f8zF1LXuYysE2f9ewzG8qhKITHHQFWf5+3h3sfSlJ
a/haGIq6ZmHC3lcnzsoRi8Vs/amIiG527CjlH3uOhFpSxmS5sLH2lS58Dwb9muFA
vxKIkwjKMFrEj+ozCaUyQUbtD5MXH5ALwR37YIojKUpSZZnWdpjFpy6hmBCoX4H5
1eNyF5DjOBrKlymn5laDWx9prrr6qVvlpTKHmB5FlrDlz1EQ1pWHIqiYT9HA70Aw
EvzYlTaF5UG7xgtRGuOYaQevR/uiBhcGawtfI1+NFcDiXE3ts/Iw28yS27zQuJf0
RfRzNcqm9dtPAo5vhQ2BoDQKXn1coJ6UiJTUXTCQhk0EGMD/hEPhYHoNa3oryjo3
eVmqia3OX8tBvZoiTxO+tJNKTInVQY472MIB6eu8JxSLC1CnOYXb0fqzi4gAZfk6
HEBs2Ceofv3HIJJfYA5C/njV0gkG2Lz/Jw741BZyL//7uZsKuu9JCLRtSFA4YAwD
Sl7JgpfvHMiZ8blYpj/n7zmAYsBVF6ezHfe521fQi9OuqFsWFtNPSXtbTnrbsXjT
eftXqEx1cGbbCzatU4QpaMOtlVuQp84GBoDSftrFYCd6lZBEOk1aD+D4DRn2Mp2I
G6pla3RjSzxzvrCWevEnMmIkWxiv60j6k2RKqRcLEvY2pIWF55X+dpFLbCfW+E/B
SfbTObCYH63SgB+fpN0+EfxtkrVFgxCfbT312TjdyPdhS7xs1UcUpWKHvwBOA32r
YupzzY0Sx31kvUWSzqkHukSksf1Xlo/Rze4ADWH7tR8KggTv4dPdWWfkynyjnA8j
AQ0gAGDAkpJRJTnWCGENKjcAMw/Nvd0KKHopRCFrbnseeTdI3qkWR4x0MZe0HTAN
8kv8deA+ADC+w5aJOuto9kUc6HFdscipC7zbhvf2zVSxYOpnx4VWkHervs2lKXuJ
bMS7+jhXnJZ3ZyE7SBtfTKrAtv/a1lP8p7uKtwJoreyxJUpovbWfVCRdoSBCDRz8
vca1V8cRyD0iO/AiNXymCxFPSSCSvhSlGhO8mMvk254/o26imPcM/oWv0ovLCeGB
Q7Mv5IhJiuXYMRnAI+6FlyegbyzRhzYnDNTua4N6dy9B4p5QIfFZYCMChj9J5aTd
qIyW7Wp6y5rw0cvCPUzi4UfoLOWvaXGOyhIS/dSnLX+NPPP/fDkC5PVlHicpTfXM
flAS3tB34QVxajEyMyfZm15xEWNsAGYhD3QEcyVum3gSZBz28dA+FNW+PPS+TP/V
JoCJsxZq4zjd+pIvOnq+2etrtpWk+hGSegBOb/PgGTgrTj1peeWZQY9LGeL00+4S
1dg/Qn0oPIY3++485Iw7Gc6wFhZ8CO9954QafqtDbugeAgf6xpZlBoleq31fACCW
9xEdOX1eTNE9FMo6p+J1SP0F9t7J75PegHP5/K5nozZ3OKz7jNhB9ZtuOSOPvLOZ
W0M9iTsrdXLEImIr7q4jojQi0XdeX/Z1X/OeXhQ/BjfztOJZ+NjjwtwgZF+tuFQa
rce5WqR08zjes86HLYqd/+TfzyrBzjYs+aQ4x54VvRd2PF+9cG+fJhqXDttAoq/G
GIE5U9q58KNl9sy3AHFSVj+yaXU77DaTvj+QwBwmWciq2I2IDAacBfo0YOphexzF
xtB+rITDIWaYPHngFKqnCn1Vfvt0duFlwye5nyzG/h345IuVMs1L0qykFYyEEUj0
UC0r599J23kifgsHIHpEk6LgIF6j/G7urynWV3pv7h39F803V6x8vX5bYZfp7W7d
1ViC6gZHH+sO+MkQ405usVuBFIZsJczJIE8mQDbXdZTnIfboM+JXQNAlhbpZofbn
JWdrhK9W03VuWK3ljXsI6LoKs3vgRckWa0KaDSYAoC459isWGwugZ3kE8OKJNvWP
Mzz+lMinsOfB/s1KqWgYTjzmKf3kn1nY3aqyd8LaD2wxOFIdDSuokb4oYt2i3fFQ
2wfdd/mdQrV1raTMFL2d+n3C202V8g1g9EeMXf9E7Na1HHXTVLCfTZPCdPkDqUu8
H0jgjfcr2jOayX7rgYzESMbwzLuXKpBjUuo/xjClZm58b0ggajP/2jMKucAMRVKB
R5XKt4Y/4+yowZ5k2K/cwQjQ116+1QsNcXEJaCuE1zs77NiDRxQJvJetq8xVcgvT
aqnxPAHZwfxVRGiEOdlqtJXMVLDztpKKAtuJ4u9z9Rd4U9u0tUEd17D9wS1HQfg8
XN1EsxE1LhhNkvUe5rnIUeyfFXoL7tJJm9spwwchppPQVgm4KFzM0LIdU0XfHO9q
C89oUHVaZ1aqUwXirLsOkaV5mi0NG/ObHsE8pCvrP3aA4MMP1FTo9vO5D3e4p8/w
FpACkoAz173VcsFUulkmpxcKGi4lMWVdTifj+2Y0xpE3sfNRIMxrU8e8SWzyyEkY
NA7TsMQgK7tFwmZMNW4xr7MhzELIfN0FsvwWt9ONObQMRYztkeHeEEkQObeA3riy
R5DLSp9TM2i21lD42NVstytZJtEpGlVPEJUt8mnvZUwbuobAXmRwC76xZjiNhqJD
muLf9Y0j0RzINhy0Y/NjsnX+NIGaG5LnTEjnZWnnfRrojXWUWRGDLp/LPFa4ZgS/
0muuap/v3+O7sGNHgCSjca7TCoGvLPPptFAxVJ9jvLUAx8vjn5Xoqc7b3hWyWaTc
x489EVkBKDMXG0w7o/Y7FYb7Tv8nNiKO4udQpXnJt+tEiY45Bk1jTDowr+Z/FZA0
tSTAilpA1KhMW/vq5qiK7qJJFwgV35PhlmO6qqfj+KOnounANSHLC0s1B2lzPdlv
6ngRQA9o8tFrEnyr9Dcx3/3EyKDeCXc085IVL47gnznOWNqdO5wQQIW/NMOiFeYR
7pr2PKoPLVtcJjRshLuEvcYXAlM+3TZOqISjWhPGLHt/zmKn3tS/r7sqPe0mcEqH
khzX0hA49PKmIqgF+0v489UZByaCE1B5fpYxFRrIBiro/ZzUPZ2FCwDyP+i6PSee
19m3rAVzs/2Vi0nMiWLfhoXDRDNNqPiMsl1LsMVsHxPupuQOCU+kKmSRY4JL84cq
zDFVWV0QndVvjEWizJzdRJPfIxa46wQbAVyWicAdK8RW4xvj0wVLrT6GS5FayTy4
nwsoi4TvhadS/tl4XVUUe2JK/OzJ9z1M7ItPsVCTSUNkKHttHsASeAgLMSFAzk2j
HuTDcJzc2CGW1OoAOqdLEx571gVNTeJ8vP0zI1AprCveAmQAbVSvbfDup5Ftum08
qHQ0MrjhZJyd1ypKQHgoCsUFLOsLn6bATciaC2MRuZVeP4+uCa1EH4QGLit0Cwqm
FdlFM8DspdjVQJ/cQDrSmK0loaWmSiyHmylFD3C4lxpuxMKALgRSta5PSKyvtfPr
/GEc0lHYkgSvhyiOiiw+A1Q3qN6jlwTjtvsYMODgGQzcXseTbVApIrihBGuKJhs2
kntW4wOspTPYVpyzwyjBvSIxx5c8tBWBgrcIA6K21rhK307k4C1xISYwUfFmb7B2
uPV7x+R52BsKcVqwfWUxW1WJLSCq0vW6fHHCa4D0Ea73xzB9ubutwDGgLjtQC3EZ
+/WqBVsq8fvfKVzwYai1mWdFSOIh9aeDsqWwQekl1WhBUwIJktDtw3i6TxgTyTTO
8iFtv5u7+pMsqcnzTkuMZ+fSjJRueCQDjFbUcGxeJi+d3DoeyR78nBEXrP5m71X4
4/kh1AzMLhqPKMH0DOoCh+QdA0/NvFyVKoqP4wlYo97mjCfIw6P5ml0X7lBPPcN7
ebZODR0rgcZ/XV8lyE06AZYd8XnqPEwnKgyK+SLV8hok/dVdHqdf0WASJrVXi1K3
Ew0SqXBBR/4vW8VYfZKDbMCwsYKwAia3nk6fodhad+gC3rethlCYoN8eYYQ96Ppc
3V7tmRdwCCgTgs1WRN9AP1R9bChOErc/s0aXK8gKysLCmIOEEX0QLxtbDNxFz03R
6WV+C772bdmYLlIWl5RYmYnxw+o5Yxl/euWaWUf/SJyKZzmvJ/ab6Tvlwpn8UHtV
RvDO2vA0BWLknSLIZOT9o4NEippSvKIiNghRcurXfYOJBU8v7D5b8QxW0R5YuSRL
pMhdrA89lz/90+2jgI+HXlaTdqiRnJ9p7WJAyJY4DjTKF2jApPz6bKQkijf7xiAT
v9jplG0THeyi2t8BrdOTwe/IRmYrFHv/2yQaIAxAOEl7uy3g40Vp2I2maQA9xBSQ
rb53o8s6uXDpHiiVyz85hzBo/1/BQWUPDFzJJM/9CceXOeyCcyynrtYtoaThzcMJ
pfJ/BJ84VJjcm6X98jbXKOuNW8Km+P5/dxYOeYrNKWnIfV0VPDrHdfWlefXPXtcZ
fPDjTVtUYmrn/y1S2iu82e66Cyqe8HACoHOgRTc6RVKIFc+BiudrnqxQlYTUgnHk
Fx7pCqY7IR9M7GnglqTALSrwe8eHRA+ocike0/7J+Q7C2qLjpzJHHDCpE5xO9U5p
sYutL04S2ZGCFDA5lH9njy0Ezah9UDT54XclaahqHr6NLK/oSBQ4VQfvU5GsmmMY
ExjZXbHnnycVp5lb+ZGErwP26RSvYCsfbGMZ+dlk3Q9skRTPv8chKbrQwPjBMFBX
bwAnQERYCYToRo6D9zo8ItFWgUq6EUS4ri1K7NGFhdfWSlqzMzZKlsx/W2kFuSNq
vCsi9sB7yu8EPaWEmQqrCd32JXrK2rOifTknpqnSHetIscG0DvLfsZVEpnqvrziM
UPAqiJDtXH6w0WK3oAaJIRGbG5R6IIH+/LPZlMZofR14Q5lKG7VovbsMuAQz1WXQ
Jvn/H/C5VEFNGxwsTxAqVMnUu/0LJUECc8yRKnpk8+2cPLD5gvad5oPxC+9tV822
RusXrvCi5nfKJtG538zhqfq/oDIHoW9OukNTRl6XkiTrX+Vp9YoDGJMZui1TELCi
p9hCUP4TLiMyjjcJBZm6LWdF/ynFyY391zpm3VZVz6FILna66dgbe/9O/IimQGYI
WTifeUafhV5OljuXo5pwNrH3LNxlP2uXd5+F2C6Dioy+On+budttIVLlU5X+HXNV
TSiic+l+0DYKkl1bgGjnxus2wg8z0NAOCxi+XHNP6j8Jc8EgA7BYFWYifQ5srkQF
ZSc9eXX1XHoedR3u4lEXtETyA4e2wdkEilCBebv1FGCCr/imLB/pkliqyFXhQEuX
PceGMR283SYwro+NdTEznAdox8DFTGlo8BTLWjDIWAxsRQXRJ7KUmgzRZMAKg96q
jfIGms7Ljwv0Nm9pvpNNVeSycIEX++UaVBj+DcqH5129hnpw6dh5m5WEU7/5J4pK
7Mm9ITfFnilw95Ecjhk3RY42Po+DI8qupkZyR4BkWaw0zdsoAhvxYbH9BEfUJmoz
foR44uv67vx0ejFhEvzt53IlEhjCSEa8j8YgIgIylb1/5zS5m+phfbXXGDgeHbso
N0F5mtAIJiTzrOymMpfZczZbXrqqqv9qLUsCqaUPatEZnQtYwkWDIYM1t4w312Vl
KEkp29mMe67V1zIJ2eaP9uX+EsOFw4duOjEFrbu/n5BXZ0Xum1EJnP1Vl7DrK1dI
mF9kREXAUoViyMT+Fs2Wvp/2V4COhEb61PvDdCxlAQtBXCXH6pZCwuB3KmJQn0BQ
O6dpGYNvqhr4UZT3CzyxoHcj2ESX3qCYMcxh57xAFPdfLJUtiawZIwii+AadiQae
fEKBFP0LPZG5DwIaOTIXGF45b6QlqBSBYOkivUw2oZJAYIXiesH0WnG6gyL43J0x
YKkLsJnKBu58v9OdsiInOEK1IkCWI9lHmu9XNfB8709Ra8ndqASUaw4q+ogyO61Z
V5VaiJBkYqL90JaUBA/tRVYZow/Gn91jNXAYys0HC2x0v+6fAdz9P8DvRQSS93tj
g1P2S2NsfBY0pcWl+JVcLK8NGxliiX/FTjbV4Hqt4zTisNxoJBm3kue7xZm92I1Q
mwEZ3hq8H/gHyzSFH/7dPcv1QUAGcwQ3KBf2OgRpqFmofMBrFslLLwQB/FwbmDUw
UqfPjVJ1Sh5TM/eCrVZtEA0vvAYi5TmmtVpdc1boNumaudP1+PhJq36K48nL2fab
ASSsIK98Lwu704FQgEDIQCx16D+P98Z0tJXDfFOGuH4XNdz/zyQTCHkNYE7gRPqK
l69JpAVNCQ2eGx3jADh6GmwSfYKkwy5ZwVEXjRDUPFcJNoXN+BPnL4Exc3RyIu1t
w/hybYqbHERuvzeIuM0qsRrOShSIjGBDML49s3zTS55xQq6b+sw+Gxd7pWFwgzAr
3mF5Ch5MVhgopOoebz1oKQYoOshvM+1OLu63tgQeHNSBkeALTPMDqncQf9MUCTQn
k81JOvVpPiN3nSzS4KlNGh7VQ43JDRytPp4MjH+mlKHVE0EaoTxriIvcA9Y9Tk/R
TLj41RO3BtztHIUg6icO5bycH+xBvjpRttw/LP/JiHkKmHH2k3aZGXZqApwrIpDV
cxUyG0SU6jbI88RnD/7ot4CAvHdslBjI8Cjt8CvQAVB5R8hrn1DvDkXLmp8Akfc/
+z94BEsgjOR9EKzSrJ9O6Tv4RnYzgBMR8TFW69V/uMgiEW+wfAycYcLcZmYYj392
Ihqcy6eb9x9gIrez8HcGdG41f8zCjo//ya2W4HC3mA2szZtB6nKcPhCES10vmnxi
v0XyVqsKNatuzLw7FCzmcaLX4yuVqDSh3MbqHQjUYqkv9JdzONiecVT1EUOp2uH4
40HpIR6SCJ/vjcOAfUu1N0+gRdGFplQXq4nkN0wrnXsQ5U+vyhNXwB6SUVle9cFI
Co13DV+qLMhkUPlkH/YYyxs9lN3XDW0Y5V1x/shhiR56NY70hSo5prl0vd1hQbun
DEwRV0k5z4IPWSyKhs/DreGgLj2Q60P3TqyQyTAf3LBEL8uUILb7GV1q3tIVWWuT
TBe8lGqPS5z/VexOx9FtsGcNBO3qveQrBi/3AI2NDdlFoNAXGBu9p1OnYsMNHt2d
av57nUvAfYLl4OePonX5ZwuL2nmza4+Pq4j2A13XE0Th7mHjuKBuNui1/mPeVSeR
3k/l77paSlWpoyWfLp36PGetT5WIEnYXDfPKpRF9pr/fMstOh5uisv8njX0/1D88
UTmjkdmswiG3+JwIgHXKFgSsSp8JFOD1hpF95+gldlm1g3TPhtiSSI/S2Ujxjv6y
C2Hxd3ckWMTEkXLMX2+66U5NLcyyvlUWkNWPMzMjxCnidJ1aBU0/tNZGZG5ES9Za
qOz7AP+g2IxJkvHCvyPcpt9zzjq9/qww1KmKvEExaA+7Z6mkhU+i8SgLzQazWe/9
m5mX/aL+OUmJAqQpSN2bh/XM0PUYPsjGyNKAbDnETCSlE5rINtNxqmQtTi82t2Eu
Kae9M5Mi8ydvtRPnbYYW8QWY+tsw3ReckERw6UOKnyOJuvsc5bnJG4aj+UtyiR0a
+omZA+xkQYh/lG3KCR2ZOVcmqk67eFpaJvxC7fTROXpE6JQ6m6T8VIdLsUYWajs/
tCkzbPqTegkak+Gy+7K5wq1RGGyr5nN65UIPYQ7RTc2z9uyaZo5gdM4BQrs6MmpJ
CJZvLZ7w4d1kl7MOvx9/pB0vQiOEavmcx+S4QR4agkQ6tSiDF4b12qLqzsXugZLs
sHhvPuk4lBA5dtWzD/D2kff9XYRg6e/ERBfEEpXxqED/HMVJ5kNN9y96SRzo6y9i
+TjX+L4PtuSWgTdOuapr9yTy7JhsqUQhFWxwCZW1fNKUwN0lFokTv9I6qAHAVIMH
bqpT+y4Z45mFwrFnr2n7APPPooHJAXaz7E26RE7UoPRF2VSm5HVrKzCKBlPOM6gI
Al8CmLNcJdADakritNueNl65MqdPwH1uXxSIpnaliOqXqEFSI5+hPR2Yga3yj5tb
tWPANbQuddN8ooYUR/SCc1IJrO2ery3SHMG4FLu3LGbUblnncO9sLyfpC3+rGiTk
oWOnBWUX12jFDQtt6dBgnyADNuiAyU/gGnpPWtDvVYeTEySrU0cM7iWbCDZSALaA
YDjsGcytWJJhf2t++5s7Opr4ixlgsdmVvYqnos26gHkdXKlpN5Aq6/O5RhYIOPLZ
2dK1UevmC82m8pBaWIG3So4u6WTnTFctfMRhuR7Lw8QwxtnHnp87gtNzxtGPCc/w
x2WjRsm6DOruKjSrlN3/7YSoXERdWbnKoYIsYPcUP/LhZfFO8soJcO5n9xAQRrmW
j4hcsHlvqbybm9dWH3NfUhD5gynOGdCgtzKQWL4bqBTrG24HRsVW/uc31sUCMigp
H7QxZqPChrY2UNFSSuBsonT/9rEzzflvcasmLXKQxeFPtAoD+76VY189QKjSWxR2
TOyxby4NZsTYvgw4byH5JRQgF552elQOjjuO2MVr3ZIJ5Mzwn/xXHU/eDduGW8IU
qnRzOVXwkMP2OOotKBPt+6TnVzvm9MltG558IOy0M6FnfQ8V4i59dAiFIns0pIBI
CklSQPPXvbqpxCGG9kLKkH1HaAzFO2mIpfidKOdK7wYAUZn5bY9+EWKJpDBhqh5s
j7Qid9XJ7bpxWZPDm48P9zqVS/B/VN7NQENFhO2kBDj54GhSf8pb9Db/h/QFD+b9
oaC0J7Djhjkjwel3yi6OoXZKAYWHRzJ/XtRFNfaHJpNoiKbINMcST1p/Xi8QpYl3
7SCAphSDPbvT+GIvoMfPd4hv8fRJqEIzX7dJEuBQxynTkH0Mru1iowFLc+TWzFzq
`protect end_protected
