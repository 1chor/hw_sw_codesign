-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2Hc8Q1vu45zso0Xvo3qsCaemdFuNK0lFg+ZMbCN5JBl2D99BlS477Zlhr5u2sZmv
JgMzUVfPMFy5Wmun4cIP2ATZPw1Cyb2xRKQc6BIJfmYCs1VFomKMmpYJqZ8oNLyo
etIsXcXwzsUnWwBQJF/8u6OWz86MgHzyblmRnWzkzX0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8688)
`protect data_block
koMs5mQfvnGkE9Y5Qmf5nnS5TEc2OPKvM2jkdJ4Y1zjsy45Q8ykt7ma3uZ6CzHA8
rZg3p5eHxsL+pYylyb/0lG5t0HLyYK7iYp59y0PkmoR+Ery48xvetO7TRokd5agi
utS8vJvRd9exZXUxrNtTIssX1PMxhbKm+8PY8B2IwwiEb+698VN7OsujStwjGJn4
/05f5uIySS3ZIHeKVVxMtIqaJOQw194HDASJJchSJ++ZNyGv2W3Vy/4WmM35yAA1
eVoANDfmMjIro7injH+NSrG0gM4CP8IOxDuilvbg6uKK7yEq9bSObslhc082klV6
RLeTiEkqCpghdhO/7Xp6Px4xjd9A3NW/zvVIvmkZFJ1R50OOSYQz+2bnVE53wbbp
rvbhNYMXKNMm5GqS0Zm6CRynMAEQLdTHfDaCGNEj8P1/gWr3jeQjZCH4KCde9TRb
S9skLksdmkcDO9JlNrE3cCbWw5+vrueRMbm94ZXVgEgJqJN72fza7B4H6msFF1z8
zet9MrbJbereDybezp2p1r9CNrv0ME/F7ONxG+Zcym8gzT2e6scnYqCnA6+YxJTw
YWBrRmrAUx1BqsfpDexMzc7ryjk7Ny/YvBFErjuhR1moIaP53KqJWvN5ohHnQt/M
+snt7LYyjfGSO2dVdSyRUe4KXzPMAHk6CIUu1bTJxrpEZpXpycE2IQeDLFNGHnOP
9QhHa6c8SZe/1L1kUXIntDnIyxniP2+UaO2CHhwlokKA5S5zdC+pv3csPfWlSF9w
g8ZqAHL/w5ZW8fTbCb3cMdCLfUqz0YGh2Js3qL+5ygc3g+Uv5W1VpqMkMxnJkKXP
P+fmPvKv3LgK3RUZYfoLd2eKu3HwheiGQ4FlQF3MzlSokfIu2M/+4loFh7o5ZtAl
XP8GOe2wHl/q9fUPcg450UPRe4mw1GAiTDSI98l9ZACjvYDIvjcYI+t7DBgRW7pi
zJ4Ut+mNENLuF2F5v6vwUVZcUHLqNiohM+arqlp7DDaGc1FBEcnH5BcVzp0KjGUS
f/rMCk/oNIibpo/+ri1Z3FSLVagpVwzpTnmLqJcLXGo/ulXqqcLh8EXEbRD0qoBo
em7/F4zfiC5KjY1hxMkPoRNL3RRUumNdUYxRGhFGm5wLmkIWyMQi0uJ1LMUCCT1j
g4UbVb4Lh4Vsyhqkw+otj2Ab2EEYBJutafyxq1Vcv+QxJMoRxFMqId59TzuSvcCq
SCbRUjOQikOjD5CtbrkckB2A084JZjczs6Y67OC2egR2+95IEl1gVN6ReuV0eV8l
pZodfIgz/dKmdxwd7cMuftVFllu9Oj1Fa6vgKewxl1s/7mnjU0RJhGsB/nIZ9Q/p
J8DqEIlqRV4wsZOWIGb18V2Et3anFaFSoJaE/PgxlyTOb+v1CRjLLL5ltJ+yOGaA
S7yx/t98VLjtQ28qVcOhp7Hoac6MnUX+AHPcHPbt601gh2N9E9mgSIvhuOzkWboi
pj5Zll9qMF1TV+0cEwRJDScncfbITZhUwNmIvn01A6vosGUXaqmajnxTshoxiu9A
JJydM5GLacpdsjgFUl/vqv2p/kw/76jRn+b0NKmmznJPAf7IuZlAgU1yKbiUI4uY
LjA2CLtY4cmPpCzcLPyWBMGqWP8v8FVMoADGekRKIF7B99RTC9nTdPkcd9o7Dp/i
Fq9qcVF9bz33MzlBoMe7EZ8aE3Ft4ZccyquF2kaE4C1k9uf3VNSHGhOP2FBzLXFx
64TjN5T7SAmd622FDUHcQoXjlXm37uE+QVEkFMS1RPEfsyrcpe+Hf+K4AnAYS/Ko
6Nw/hEqUx59E1MflDI9/5N8VxO0be5pmsgSJTUph2vp2oq1Z5RxZN035UZO3Y4kE
NEG4xlB3ifCWq+N0GazW6G34vQ8tsYi5QBgHXifzkd01QuKqk02FcXoXeMBhCiom
CgBX/QgW1Wtmx/jo1kn6p0uhYlcLG6yZ1iy3cT4htdVspxeKcKAzvQnOrMkGaCky
iVWoxbT48A+L8cuvkjPsgztbhG0fdBzBIPoTOBMOxMDfxGDmZqIDKyXYjjLRo7oR
dlqidDYJOd7tSJiZvBXdevMwuN6WPDfuDOVqAz19b1Y5K+1lWfTS1H9iBLF4y0/T
8lqnSWF8K/22pxw+sPb1OMuKCotZEbJSnZnPKZGpkIaXdiB/+VXUMYwsywRDzln9
ikP54aBvF2M1Fc4AItS4nniuBpShgclxjn6KT4x3pDiB1wcwtL79ITiRVTN+XrGe
ThZfJ9rxMi6cwMePBQpZH7IuRjy0HOw6rj8L9qfDLCJTG6Madc3iduEEMndTtzul
D5BY0ocdIqpEtHi9QD+QOahHRnKcWlH7k0f/FuHFrOdyOJFUwaBL9p9xkuTu5cWn
ke0uLI7kCjmr0rzLVLQqv51Q07oKwjQ/F1PUf7glRRDbzx1wLe8Hc4M/XXDikyVq
Wj4100C9K/TGd0wRi0w4V+nL8s9ISkfSNLF62leaLud1841J4gqf12RohY6LUjUe
/dnBtIJDnw2V5CtM5+rPBUQYRdGpL+JWUsGGMwCNqcZ5iPUfP2ZFL1ofIqFwp/qS
hJ/sKsXBwnH7V5nqYoWPfGsrwPBpdfPClnIX6KlDcUvyVD4mQkt9viVbGreLcvO+
Tnhzu09cAovZCm2XEU93nKIaNHPPOaCZpKQHHo5v9THTah9dwxonJ3JbtzwMdwgi
NFbQvuIFV/70ipEjKEY3hO3Gft6UlJwdBpQmdqSubonJNRUMMcrXImK/J2w2D3rW
Ah5lbb6Qnuux9g+BFHpL9l4WaxJA6si/gND4TyqVacuyalYaSS2+fFUIK4pTsTs4
Nfhb0TuIjddoYHJc/ZlD6HyFc9JURnEfCzufydVm98D1LiMoAyH8ta1Su8YXxlrJ
z0qvRhJHfUFj1t4zqGoKy+1SiSO5bvZ9VcBD1S7GW07soF8224J3RJvHrSwrkFP3
IQvQuw3YyKv1knnzsHIobKYldhIc+AvoxkIK/NXmdbY4bxB3H3OD+KdF0NG6vRnM
K+jqUtylrVZAMGpSVOta5/ZBeb6TWadkKcCXKiSV3OtzUrzpcSk+IEXMlVlMV0Y9
E0Fad/YuQ6A8wUh1uQknaJ3lVu6Uk4XUvBsvXOjxkgicBrze0SUYVJ430nY+A79p
ys8ArqHa9Vgz1LVRvQgqyDXKkOqKHm3MfoAtqrtwa1xmAZgvYcRQqB4LvCqVNghv
H5jrMKossk/5uqxD/JWQs3jzhFCEFPIn3kaMjZnO6tsx8cy4WoZXxyNUfHRm4dgS
hcEClByz6RpCDqHdUPDRisgizIZkGkOz6Ohj7FryQGZ0SNUE2Vy+9LUEcb3Tcbyz
N6bZyNUZPgNURcBg7amPxnbrfbM0Gz4HsOHw8cx2296udGbS4LK4v2Bh+yX04tk9
i45x6WkxyQCmOZULtFN2DG2neZPHrVkN7l2CtkAuVMJg5xOkHw5DfKmMCf+JfOG1
f+5OMTCxxsGeWhWawErtnScVI7S5F9pR/GhyN3NGC5rbTbsEpCmg9YqSogPWl19v
gMojG1GqLBZX1yAzR4uYnR25pkJ+6fE+LCkeNN291mx2A1jarSHfvIafYQ6PgUy5
fJ08cwoozJgHvQrysWiXoN0wPq8XFgR04SpJuOSGdjKoLtdu3Ftrcu9qC661r+Z7
oHgxPeo/KcZAypeIJuf3c1/GRHdDBhqHsJlltP/ImZ3Z0mbXCFDFWcuG7gjrbtYb
htjZRjZLu0MnhBfRXxRBWYN6Ca2fTzuO9WQESJrQi//d4fju9KEgN05+V8auyu1N
HvsW7/wZgYHJpJXmxPADBTra7Q1GnhPnWgHLDdUzunDCWUKncxhQ7OHbDVgvZSPw
hDKyrkt8SfGy/C0iKw/hyjIf5DXTILZN9Nu+8Y9UhdiBXpgSKAWxwXbV2gIm7YSo
9DXy3hOeYO87u5XOARD2J79OpRn0Oe/kt7UnwvJghgvBfvP+SD3zM+TNodI4Rqkz
sk4xxifsif632oRgZqzaKss1FtRsANodQizRbdy8LAb4127uyASvQuh4fOfe5VS/
IwzHnUlpu6wXzk3iR8+F11FqkOj3QAH90jqKutDSKPPppD8icaFjqgW3YXPH89vq
ElwSq4UtkUhh06+gECmwHR5VLsvCZQtirsUMN67+igBN0Z4w5CmoT1Sg01uCgRHL
cGIyRCQa2QqS3YVgGNgM+Rhuacp3b1/gMGZfWy0BnbtgEW/+Mxog+++kO7wOvVyC
m6PVTw35sQr8Jrj160M/JTSEIagd3NtRT1Wjy6iqI9BWVJfjUpuKaVZdkUp4625n
ypVjfpR/bcKTVzPM/4CABMUNt6AsgaiaEsvHZOEXGXfr2SliZGU37de274WEnvGM
v3yM1ydT+hxZ7lbIDN1FjOQN52YFaCb/dqDuXU2xeY5iScNgRqYB3zPMF21RFgDU
Q575mSngLdWuzzbJjIt7k76pzV6sZMDA2iqY5sfxD3IH7rJJTeql/EzLkRzXqEGG
6k1V79M/HEIeXbRY+b0fWdvqT9K+G0KIuEJc9vZvXLYUz/bnJtqTkA89ixsVi5wL
djCtPpeHgvR9sHscyFPWUBfBNWj+eSdgQMCP4+5d7RHf3BUc9w4ISBJV9GDxWxj9
CZWaz/mnxpidqddm2+3gEsBZOw08k4QGplFFPMSZlzfHmXv7GHAjo2tAq3SkcKGI
Gh7PvLjMG/jIEsOibxVLeK8JGm0sGaVEEYQ0uvd0NU6X8UYVgwShlWSk1LbFpr8z
2k6EucRdEeiokNyT77r+fj1Js543jnEvj62b0zZU4oEfDpievaALrW7rUk1HtW2D
9NrwJ6Q/JQVyliM+mUHpYp1UCSSu9YlMJOOlB6LDMeU5Ippn5gCe3gRwVQdbFPSv
6YiPrW0oGu0CJ9rQP54FtbqKOzM6b+ju4/c5Drjxh9Uk4Hq+qF6Au1TsyZHKrybg
cl1QimfOyLOVpjeEsXgUxPYTFByTxAEs2VnvjgG4qYYpzq2+0xVmnLL0NhpKUYGx
ryh/BkHgd3P3eRpzKvqdigxJMdoDqcXB5UyySdC90WNjuLnFPn0EKZfUoQDHV+ZP
793yyqegAd1CKtl3KB295SaU6RyXAtiYrwlgvnHb2CiWJwZe2XMw66Ono5yKZru3
PKUDL4thz+Vix0jT0a/dDYP9OKMmCPyXRvwIUzzspNISpkhA9Lo4KVtJYsiYV16/
S+ZmT/QHcyntnEZp8qfJ+QmSwgFfVr5FldJeMI3RjewBIytMiYowg/WMzp9taR6H
wPOtZHI1WF+lPWxMQR7zwq2cLWJW8VJY9jBol7YZ1pNLHtM52oB2stiibfwmjktK
YU76XW8y66Lue3+KWTzwJr6PMTqwekmkoypQvoHcqbehfG44GKZevrr8vd6agWNu
xPhRyJq6jzx0ODsM0nPsPgSYw8aRTkfRI6cX/7S5dzvTpB10HcVU4p/G1bihwh/Y
BNZQOgCg/EpmmIaEbiqnFR8r9w2DrCVBJthGCBL082zIcJ8oPAmDpq8XiRi2xwhP
1QDJaUWt92wGgVU9pW63exXF8foU7EDt+Riw9+/pXBt5stjbCGExPlFXGlXp4tyb
jqt+Lq6JKR7FfB6m0oJhLL90MtjefhBqiJFKosEJeYX14y4wld+TKjdczPzeHXph
Oo4iNqUSsSk1/wqgFhq6Izl+xCmSBy5Qx56xVQ4WAv7QTpabgXbdA2cNXWhQdKQK
DptPGP/rqp9HJj7YbgeTPC0hU0poMXnbmXDcBNKIyNqTYpDBVTsb3DJMYF4thUSV
S0WP79HPGatFWyArBCpK+nVjYYwd20H6kxfRumdBQHEG2kXPE9O78Lx8ereZjp72
wU/bNey//xYC4/hCo46pTK2lG4v7ycdgNj0dUQC5GqIVLkkHbKvmTGtFkglTG1Il
jOp1zLm69Cb9HNGfmscl2jDR1ZTUhVgiwgYOjglLRoai3mavPcs8UiAnnkwllKyL
9Icyde0c++/qg8HBOlJgVQSss+NHu3cUgsPYxcOpnUzgD+TnewOm7a98YUR6mxPO
fIp7rEArgFT5cv9dNAXGyg1DQqkHpakdRhV2+jF/BnNqmF2OLQ0B9Sf7vF+svKQc
huVUvXykh/5IgXqspk3Zp66jAOMamYsaWlsN/wOii/hXRGFwjBlL9rPPY+mkg8pR
VEZsBbNq6Q/+0t6kgUWvZIF3wNvyqPhLiBUp53xewECPMcVwqVPTJdGEid7MZJO9
k7hCFYzE4IiC89nyuYRjoxVVLq0qeNNZYfs4793GqaaFB9Iwf8lTNthAwZj22Jqo
HF2uA1DW7fljGE5pphpjB0BvCAGNIRm3OXurYnrMpw1OY/jMzkbEKvL6+uLIDgSD
nFrWcY2zZk8hnqnYiwh9jMg9GTmz7ugEpo73oMRC9piVo5YWUVk7E/c1Io24Zr6D
QMRiLZRM1kI/SBV2phyviPs5Z3/GXEcaBEczjmmA3KHUZpGrO6sjcOgbTzjJez6K
ey1bbmBxD76PAv5jYDXxrEWDmJ9SR53nQilVN0HhHodHDU79zrrCckHY3BxQBbn5
V0saJYzfAmDiTGaZtiSsBmLfY1rAf/18UZ5nzAy8+kykh9w2ZaawJdVN5OIFb1OM
+8z3Ts10lvlTKNwt6EQJnYYMdUbLL2uKg+NYo0bCCTltR7Uyqnf7Oex8qFR5MgfY
+yab/4G1a74VH99sLcYztrsqxGFgRxVofqSQp8ubTJf79Y64FZQZlVKsryX4wkyb
gvnhyD6doPcwnm66QG6E+p/4Lu47+zCW8D/plz+icPVLa6wPBDILhSpFYv95EGw5
0Pue/8+mco9cG6XAGcseQZCvWJN49R2DolZASdoa29AuIwQUIJbVL1aCFmjdO9ss
9zDInsLZ99TMmuu2FHNlBXvvYnGMQchoxVb+j6FtZTn7kuZOAyh99f3uBC1iVum+
xO+NHOGloCmVkT9Xrz4sbOlT1hF6cWjkUnz3WOe/GeHDvgaZAj5oTLxqiqBrn4MB
9j2lfQT+NTd8x4LKDHLhRrtKXjuVVdMAwkfORcMjF7bHBVjeZZk5S2R1eMg0F/nt
GT/hBiLJE/h9ilf0i3z+avFc3fG7tXmU0HXT1VigefwiEDVXiLhRLXseA4jhDbkk
lkM/p7hoENmbwgzlo3aJKwmuN+ieMisnBeL4rR7eedO3R2vYUT+RKla4NfBjbYHv
pWtMn4ifZuvOcPj3x9ZeGYx432ZFaLHYmoykU7BIGNFIp9DSI0E2NgQFurWIrdgz
SRkMUEk3akgTtkiaYfb1ldkqNN4ks79xfkeJn9y1FRf8dfclRAMrXYtfSvaK626j
VnuTt/aYlnh0Cr5EFvVQXir4cTGCb7aFZQNv+h3q1+wlARx1H3MPMrPPe3S5z1p+
rSpFIAxLqooQ66rFCcKYdizXQ1PmnikPzlQPlwROW2TCh4Z/Wmdz9SgXhKdW6vQk
miw6EQuDufIs55V/UJJyR0h8q658HXXbI2LzXnUwZbLSc/s9n4c2X+KGkMF224ta
Wxy6Y6wvi1K8DjmqG7x6eTKsURhyM3bmE1l0nvf4oGzrFZw+DNJPfyJTVxujwB3h
k/xa249+/1o7yoCUmlHrw4jiMrwlghyJw59r/YDo+qfmlgKgoQuNS/aToIo1k6nt
h2mhHusUq7wPszhxzJwqVmdg2xuDz/u2tz2hFu6qqBI0gjmV7USuRumHM4uDNyIu
jWouXRqQ3EbmtBII5TOvSeE8ClTb1+E3zATRaYV69D7f7IAOwX7bH7FueH2dVC1v
wGoTcsFd1z7gb684LcXcA3dpCI9KUmi5kWpBQtBuJ7ANJJKQwRPxOVB1lVAjXM0L
wIkpKHRJjmHlV8TSQoWjqmgFw5oEpMitzqYeGdG9VKUnH4eCYPKbJ2HLR07XupJ+
wh7I/XyCT111rveDAWgZtVUpRiYkLJCvScEF0vKUgSE5hMJyOzRADCo+LFCbDglg
ddKYKzmYX5u7rZdyyL8JIPLsjBDfKuUmm//4bfIYlXsI600pCF7RCZr3EO5rfWue
v66ycwi+pjlP+js8FXonr9TA02MRMgk94MeuQyCZDPvTWMr3f0bDtk4cljTII4IK
FSghWCSA0f9NvqJsIWcIyFGtZHQ6HLo8WiA/GpsoIFJ/7aRIVATIh6gIaeYWECZh
QM82SqBBBhKRfOr2n7/KD4459efYAZpeuAsiRK+8lCl6rCyZ8O3juLUYYGqXBj9w
pXQ3/S2HcuHzyEVSt8DWqNePGftoJx0Z4ZdWCApQuBA3VgjJoABYAhbwRoAHoW6j
MdTy1DdZVPUo2/0BMXFaa16t4h7KR3h/sj1f0oH++Pzn8jqlnxTX8EUdB0mWi9HK
mOU9yBC+wwRpcPu59hLE0cJozD/hv5xhUk+6Cae7YqUbfcIxk8GCQzAM6ZLnqar8
Yw/nEiquBKrMnHhhKFwrqgY8mu0jpbvhsHML9zPxCmeipBk1Xe+/NUD7OlHfPxSc
7s9L5iT7xn6mVKjCCUokZfhpzM4rVukMsrUQy7yBTEnPzpZNqwbX9Rvc6K0qFc6V
2NgtN3kEOJ5WZ1E791EM8UBDAyLZUG5Xa9ZWJ3PvE0PqIhNZ0AIzcx1QqxQ8L/pU
fStBKYRz16JZLSDi8rqRiPXuc0tbU+qp5vWP+Zx3FlmJSYtt/DFN+S1kBLwjEx1m
y9zjbRegrwwjtqpmv9EUGA94ycXIY6nnDomXVjpR3oNopeSw1VoEh6da1My68mGD
BB17XcVVGK9QTYSn4tS8ZCckjHH7xuxQr4Ghdp0P5N5JLHy25zJW+onTsuniCUVW
mRTG3LVGMMZhw7lPP1wfwQmuxnfrXD07F9cYLIyczTflDGhrYPFobqYQ4RtCS17g
MFCmL0zR/sMHX2V38Y5VNMMtLpn3b99gxUU0M2DksWFTA9CK4L12EXLIWqdqAE5b
miLyuqMN1+ji/oMYkKvWB2iS9titCXtO0oPjtCb36G9gAfPJ9hFL8+XcrAHvs2CU
vRuK4XVfCRC5gqU8KYrvYdiVSozAZ32+w1/A8JlnGfGb9kLF0PVOedAAA06fCv07
+PF8AiR0RkuFAaTfpblj6FSWdNzntAvIodPQMrJKL8s0Iv1R7whY90O1NXwD7rBL
QhNc/j6YUkzEMGCqliu/Nwf2QIvu2ZlsQM18jIpyVhndv14jEiPILC2+rzVFi4ue
Gwb89oVP15c3T8oDjJ8XEwEtgyT2j4BPPP1SpBgSxlX+WNQvudoj6aOlctnbq6y1
tE+ENqQUGYqk4vxjI9pA9IvNpEQkpqCY2PywhW9fTKRY8AFUI3c+rmoR9hIs+BXM
4c71JU7082MyEYA+64F+Vy+wvCsU1uDem1fJI5anpPlF97fmX5ChRjKRPVt9PXhm
EPnr89el67QWTLG2uIJbFs1TlzmfY0rv+D7+tKmZP1Qed2sChfK5qtvTl8g64H5V
k3OXdtQOsWA+UTLYwmcAGWS1gZv9Z4eNqgzb8gbfNmjQSJPAHIJ5YNCiJU+XmBR/
Vf+oRD/De5XBRFWf54mkH1UcJP63gWQ2boZ+bT+Gk9K0LNr+1hqmUERjaCc5oubz
ikprD9S2dESXpicWUEnG6b5EuWfqcgA6B/XQuR0OuJBghmAENaXeg8r2s9EPeBhu
AahfVJ+ol6tX6hnUBRlwDanLUN80ePc7ZkCvP7kROIwNyLv7kO8BAXFy0vspMLKh
/bs6FSqhJGKq5y2MTF6QUxX5WJQ1KqYBC6mJn4bqNt8DZsCYxtTuDJUsgZOoqQfr
7FtWZxvfxJQ1AW/pfYUj0MWIFwLUoOhImqHV8tZ6Y6N5Euu7NfgH+5TDA3xKq2lQ
IQBcBdVBUMx5As+4pxgnCY27sVhZnA9eN+FqXpZMMQO2Ckr9AOd2zVeeNSmtzMlP
6X29xjpeER587+vs0WyWD3KdbCIdksYD78UFrmzPf7ecBb7kZzDqjOkJTKBHRDFU
aIze2KQ3HckJBaeByw7UnB4+8VEvyPqFEH3EqyabBIHRmRCnnR4U1j4YZsIV4l/g
po0XnD4TswUZlVa4MpyWlUA5DvwsX5EuQ6PkkVrrqv1+Ps5ayP6Dxz7At1wuAWym
34q1uYpqEJdZHR3jT45WDpSj3lvzPECB520pjwIdESCW+gfjmZlBDurz5DNFA9uh
LohB6puyhs9PIRBJT8iB0Xg+fpwq/0HqQIVkqDYGSLwahRPgcc6gsI8mYHskmPZR
++lSJizDNsbwA9gQMJOrSpnTPvhAJvHVvHyIlhAZAVg2hg9zUtZ+YG+bAiHm2gnQ
nelWMC+L2lS4RGqzp3XzPx7x2nhF+eip4DqKGQfegPdgkNk6Ds1XA25CkW5RzMX0
fSQbLuIkDyuriLdMxRa1HhFA/9c9E42GHRu2WPI7jec154GdND3yDOx/Nkmt2RZ/
YrGAOyrZs9eQC4OuvIwLDTLcAQxOHU+Cw+an5yHi8HoPX10DO/5eoUYghRSf8k7G
RI2shr0RBDPAtK8xNVRAJ0bcdxzTH8/aJXq1jQAHyLs95pD9l/Sct4uWcyGZJz+j
LGbOLo43ca3qke4SB3B55mzYuyvkjcc84YmaBDAizr+p2GQEdvE+en78PuwzJm3B
1WGXXIC4ff/QJhHp/O7bbF9UiOAA6odj5leNwQoq5NsJ9hG5iWiaGcO79ve2CnJ2
xBe0dYr8V/6n6YCTG8j0yuVVvvxt5YfNN2rWokdRedF2bk/j3vEAvPsdnh5toT5c
SvgbQzzeDTiYtU2Z0rx/epDvTgzP3nqZK+tHgSvCIwD/NHvIOLzurzlhUNASgxso
wz6pun5UqqlfAd4tVA/0GQvDrhT/MZ/d8iftDYPupo6sXuPx59XdzFRBDXVqS+DL
PhGDQJYB9H81D4MIwdmCvnEtaue3Tq5pNnNadrRbxn7ZDpsG1GT+xssm6OyYxIIn
VcOmKzfDxhA2tYqduQvCVrLDbITI0WL9yKUjsMDtL9nBzKwdNBx1qIFjxP9IocNV
fT/USuHMwSDct/3QLT/ZLNthVBU2tCv9oddv8AAxP/LX6ClpxEGgb78IiH34wPZu
fKAqz5iO/QBvGTrexPVQfJM1pG9Vcv4LuuTCkCMf6hkb53iA99BEdDBvedHfrMK1
IxXnbumPgCJQo29fuDZIDfQd7lRTqLZtxRWE66/MJ4F7WBUlC644IuVx1J2oBkfz
B8Z1IfZtHR7+393iycOJo2/HeLqshYnr6TvYUtf9MvnWvwsJrqIKaZNzJ/hN/BQ4
Hpr7H8kwunP+95JU0iOcFNcDE2H149/2D/iBRUSRYpp8q15xqA6TfupXAltUr8sA
jjetcQDkoa0M208bAR0jDc6CAMTj1qR32FyG/OrLUhNFYWV7XrcRt8iucgBQQKxU
oBIymVQNgJa09nrOcSmxtX+L3JBZo4V/6uUQ4s3WWjk2XPLoWPal4G0vw8mzWO5f
o+f6rrcxQSTSfaNEXI1koVlFiRtw4DfD36DEN0KLYLgzxH5WMN6WaM4gXmjLbxkh
B1SglXqdjouQEQ9oAe8wjApggkcut3WvvkWisjphWeHmWH1gSyuukXetijd3RS0L
UuUdIYPmBtRGGsZQK7UdvYvS9ZTjqU5ZMj60gpClewtvB8j5NNTgt1+szxahn43s
`protect end_protected
