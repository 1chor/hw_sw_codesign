-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LzIE1sJb151FitQG7RZrXVLlILZ70lVZzLMcMFy/l+EvrwxqBc7tevwUwPndBDmomixKX+tctdsD
IeK7oaBruDRj3m4PUGUrCkK48JNh15hNbrH3KnDqrPTKYpW0S2AnZ1MGOpSo4gHQy4gCZHQEqjTw
bGrgctUp4aQVlVeRAWodBukjRLUvCl64E+zMSv9tZ6sys9hgs1cfbkvZtHFZ+6Y9CLRpDm85DwA+
OUqZNUOS8LoR0szhhmYPU++Tn6rpkW8z+Rzq+o4sI/QZVT49qx8FTAib9dqS4tKQ5UxMNiuDgOkT
eEIDa1iOVqtwQFb2JD1VI8mWAXPBEhS+btGMFw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 19904)
`protect data_block
6W07PH//vHfr/FlSqCXq7K2w6pXqfvGA+BLJV115HrkJlgMeWggDR3RF0SAs9/icupqQp6LY6Gxy
ciiVInZzXJOBBykKjrGRgExucY8hUpLKtbHXsee40cBwCQEj4V+Oz9ULK418KqvHaPOGwoXUo/T6
n11eNsUGdsHpo5KcITkZaCfeGShgrA0p2wvPF5F3MnXcucyav0tRfufR3qZMuKN1PlnDXJ+YIKpZ
3cBohxNU5HqXD91+vWDdZuFOYPgMyqlmIplMgTGp0cIFiF4aMWtE2+cUFDoWPC92vrf+0CH8/Jte
fph72PIa5x+PV5QRZA5uW/5pbLz5vINAeKrsWG7F/z1rkykPCottIXGc8jmxW1RqwdTuvMI7iAhP
0NT1kRKoJH2YO1WP9LNSdwbSY2uwmCYuc41wexrLFbmnrWpo1gaDKCZN1PT1pP18dvh1v86gk+w1
UJqFRHMkimF/2mJKPyGwFNC6TEVcLkQ5z/MieOKmRATpVUKbWl8U5HfHJwGY/D4FyRFPUEIMALqx
J7KQJu6fyST2CeDfhVrKuUfyuhxpsfziz9fzXwhjlP2LxMoJbMjEUMYC/t28sN7VplXyIXL9h1uj
y+q+7+iYqNuw3EkKBPSLGBCH95DMcjD9T0pMC+3aiyMmt4p2fK65kXLTdT4Ddms9zOLhpDWX4LXw
i9L/iRpuJGW5TvBGfoDAQRYO+no2pGfvARBdycIHU6Bn7/VINyVqBvJyqWjVGNr0Y3i7msQ3aVNv
DFbSIZwnM3sMNOIz+qzdi1buyRTX5xE7Dpv5xyq5hffufW81le3LHDpedRKmcheH41liF3w/sZge
pjPMKSZsf5dHcYCRwmQ7zXGwF04cKCa0r6MG7JNYtQO13DOdnlJOBT6ibU0nYwwoot5nyiONN8/S
M4tqdh90gXevFURD6Zw20TA5DKtFb5NusXFcQiHZzkFfHwI+KEFZP0oATeiadE7QXmWDK2OZ4gkB
+aH6C+kJDxslwP/IZe6KI5NoIX6m89hioXFVIFB2M+llB8gqSSqt1GFHWfhcDHv+xdREwQnY9QLl
PjM7Bibw0bv+wC3V4ZfvCnzYljF7vL5QsgWIze2nBV5UcFEcEr2M0DZyXeDpG1vPfeP8fj7O/C2z
E9ZmF0XBSOEVm/WdnuCciCXWvOpfwTmmCpZAalAPf3s6VKiSZaOiAvTBrcGHRr2YGpZb7K9IIEuK
McncHcBynOFPsHKiUT9jJ1Ep91DL3RBUj7JWxwQ2d0wpX+JKZ/KxxKz10zgimpyHrzH29yrglgmT
JQsEKsXgQlRBZATwcvgAUFqzHM5YtujBQa6wQVKy+sCUKD6oOOrB+e+qmmYYGiu1XRHBo5nASUUQ
Pw4gGSsyelhWj88t6hpkNcYgYvCqwm+6bHjK55aB2olc85StbCPMJRsxFq3piNDEgsM1CnFBNmdb
kjk1q3XFdvpEpLiS/2ksfAJG/f4z6E7s+YWoiTFN7xpRLtDQPEvXDaCwBKskJ0k2CJkUF2IStFFd
J9cyM/aE6iLNyx+0Af2i6AiFTXVvJEHHJ18XLx6QJYmt+Y3dN1PYMErd5uwXW1TwL/deCLIF+xeM
eSs9g73pY3Bi68S2WUJjPGvFUtzCPZ81KtexVo7z0C5PfL/V132+vpyoBp9FdgoXs0MGM/WKAFlO
e6bqeB892SLZwg6XNPequKQ9bSU80giDnyvquc3wroyCmhxlNCdSCXITZaQvytygvKJ7UZvHLvFS
MSzs9fFeFw+zNzgO7XdclGbxRsVDFzO+JW+0Wmw6QKy69ay+Nv/g/Z5dq1LI9V4udliLv35n+RYn
cZaOkRhzyq7VRx1nDt6J6n3IiuI/g+jHTtUKILlYxdoIZUPflybTcCBfMRX6AA9J7TRyDUxdiAXt
IBwdNW+Sh4EYXnhi04ZthpNNKV71XemttUsDeZCGKGL8cPpQHGIRFmvWspMNvx72fH0Ofis5M/AZ
Vl3KVZFI7yJtSooEBMbuOryUPW2k2/ppBVvpv3LRhNQ/JS2bHCpOgjIoAa7aD61V2oawE6UwzeOU
NuQ1fgr3Mcv/1GP7REBB3aZNg5FHGUt21EiQQbZ65jQu7eMTlzfjdksWYm9mXFs1HbWKfM8HdT4K
0bu4xWBw5zWWD/mfOKUdSsXX8XKf0KCN0Blmk1n9/ZDV5RWmWJyChV5vHAy2x4kC72PJtUtTMuC8
IopDDWVnl0k/zVcldlwyiKk9Y5+ZRRWqTYg8IkoUsS01y9NP8l7IsB+Sh7BAISUddQqyXgdGAJH/
hXYfzfRueFlQGaTcJV0tDFdGOabcAzTBGgQ1Q9izfN+NJb1AdxWMQLFOR8oi+aIQUOQpFvLtNRlq
8llBJgCwkrvh39n5lYR8AKtkdx+QG0oU7NnqWndLO4S0dz+2LW+VNPvHKAWrgarp9KuprpU8/f9I
0BHtCqcHejWK1C3fGsR7pOJG+7ROg1bGpqNUrvVr5YuF80Lb16Z+O+GASP9tAPGn4FonsLH1edFy
fr5q5TCzgtY/F4TosGB/sa85RafYm7vYbkD3odZLPG9lbJ0s0YPvlQ/DktLmiyj0ZicoqqoZ2QiP
UNEM2GBEE17QnX2llxn2SPZ1zC/uXksdITlPCn3nkMuG1N4RS3of6bC/CtNMtY1emDSOTBcumDIV
mE+CsiDT19+tVN2B9So9n1NK7DACg7DiKwBooAPdMpaI0iiPvEAvWg9/VEVyXYpjVO7ZlAirnjLc
3MtWv7n9FjY/Nghd9hOkQpeSRs874cjgpqGCZ9qFDBnEBE4JVNHoxFaMl+a7Lbq7L8XdX4CJlIwh
7PCzvB8O/Pyj0lDiOotw0trcLLJvn+czW7pijRLek3VqayLqzcVn9YqClcyY8pIn+qtxeatjFnUe
BoOLtepnb0Bxr2QaNXuKbEyQApCPJSDWFbGVkX1HIxFjik+q1j9+d3/sGsqtOfQDHViIFLQ+YH4+
4iu1fULdJ1Dk++zGq43bQA7efLJdjpffZGWsu+fHOnGV2y49sn3R08jgrgfCbeCogciu1uP5EbS+
uzNLMMRqvngfi4a73RFrLaWJKUsokO8/xGpiHmv1vOBes2eo27B9+eL94zS8iuJQKNgNAkDMHCQX
LfSX6K01EG7q6CnysM+4N12Ii8CkXa54nfFiTgKrMfJoI0lu71jOSfmeYTNw4SxsMUG+IEmPw4oZ
xNcozBSCbHwNd5xcJCM4fuXfOm2oKLBVYRMu2rXjz/9Lz7w0lISsZWoZRcz+jKA7FxjBXPpLxeyS
b3NYQsR2//95t6AWnVn+xVxUh4/Es/8Q59wnN8uSARH2mtyaTVMpk9cOR37O6T32j70KjAlDepnV
KY5TlBBaITAynkx5j0r2VUm/pWI54FDF99Xvg/To4gjLk2MdgQQ0yzH0wI5DHu94Hg3HwIt0s3Fn
7eeO4QO750IfDZY+55jq3zNJrix4Lu1xrsWWlfykcLYZpP3yxxn3y5gcg+YLTqREE3J5IR/aHA5l
B3/lf4IX+dqaPZdrMZNhguUaXTMTIMYfnfN8AkJJDL2mxkrq7XGJr1r34A2cfFL2r4RhkOuIEfKh
+k10QACOY0dJQ+ioEsbkEkvYeif55NJzsfw4XhlGESff5p7gUzt0f1wbAmC4MJvOro/JFDR5peCh
xbYqZAu/HyDdZsfzLbp4XhVDJs+0RqG2Dwotv9wPPIQ1z9WbNp/I62MZnVNfREtSoyK/b8ErrSpQ
FpsuzBIeHosdiW8p7Q59JZYzPfA7SGDUo4X0tAyPsA7aOOr2cJvl+XwRSdyJOqgfb6FWyvSfRydq
CSK0k2jCCeBuQ6I59VjHQSw4kWWa6DYwWzACZ7mYRePfqEbqPw8tq7GZRLOezQU0rowYKso05QlK
fCQF2rIvmotY9FXEeCSdsfmFd4XafZL4+YIWbwLv9VMjrSzmhoWiWkn+AvEiF2/bIJTCVPl2y13H
5Fu2Bcw+ymR9BykVs8QX/76gbZiQXtMDkDjhFJVh0sICNfc3E7sHL4XzDtk8ymbJ67KfeFLaNjQu
7elU1WwUqps0ZMMuddIcSd1G148BliJ6bFEGv3Hx/O7ftRxPqrkgP/ANy09yJDjW+GpAX2kL1nT1
SWbxO4qDUqEMyuQrvqj+okLnwPDNe0VIng9HDbhQQ4pIUPKCMhmt3eQbSsNJTinwKRI9NJ8IDZXY
C42vj2FdwSqGhG9sI41RPDSSkWJ7xvirP2AVXAXvKFP16XAYBNS7+4Zh877Bfi+s8B3ELHXMrrjk
FYGkzj4/eDD5Cz9xTM/dMMDZz4h12agnSmHFSRuA7A75+FlZ5+KGJzd7Q3pkEqiwNNaiGZXqoZEz
GiXFuKMD2RhRZC7QD6S+VcXEav0Qv54fp9KHLL9h7kH9FZX1hhqSx4B4Ir0Ycc3mKVZRYxgXOs2/
CtE6+3tPJI/hZwxxnNZTJRmJPDvBWVAW9ZpQZ3MtVtkozLKvlWtfiW1t8dYbLdolnWhonoUT3GsN
6Tjb5upIYuC7cJzEzw3Fhs+Em6Zb6FOrhjrh5iEdj0AZMV/nVP9duQCYRG6EekxLO7KmPg5YCTDO
WtpnKcv3uqk/M9duYyMlPWM3EknmzOkiZscOPIRiVdyyDO19JiPZSDdn17Pnv4Z6VJ8SslpJbM6P
XwXltWCiWPWNzyhQfYDm7LX75DaYJOk9HPpWDMZK7zvOC7iD7kw6QWoCKJcFPyDC4slwx3v7uuFW
kNpCWsuBaX/lJyTkkIWHPqADBk+cqwkXt1r+WIrTMjccrJYrkK2cjeeNBDqnJYuOrJjSKi+by/cz
Jucxl1AtOpA59p8zcrYucawPrwQwGBvRIQGjyJI6zZB8zcnan8wi9pJcDUb/8uV2P9PRcG9OL1iC
6+vlh7pXnHIq+cquaI9eXfC5nWXDgPDwTUmNmiyUQuexM0qNUsQe2yop/yNEdYkQG8Dmm/RhBLqf
QLN7Us9Ac5HnFnghLBp4f7y39aJuk7MjYgvdyU5ARawvQwyTvy6fuTy4zQleFV5PDHwV3hdwGOUZ
UMpqaTuQeWygEdPXXVngFyJPdF1OPvvTmuEEpGM6J1FbxUkuj45Xf+FugmyhwRhobyhfQxId+Cl/
NwbQZC6OydDnXDE0gLCQ9zWRws0uLAnaV1eQqCbv8nGiZpT+jM9urzBacDlSOc08jZOOVKnNBQZG
wgkxOigInBmFfpJbN9tItNqC5PwNJgGeP/bvy8nMihFHWMt+YWABwejjQCsW9rUZQZRlf2gJanQr
e/I7VYq/OFkV2FJXMPbmvWh263rkbHCM4RyI0kP+2qKUkbSOh9ILCsdgF7XlxvoDCfDbBFfRRJwz
fxe4s55sRA4MwwCHatmHRKnFhm1fYIXdNCaknn2WhgPH0K5pe+ivUEg/SO9GsJAE9apZTCkW/NTh
tqwYVdyZ2dFE3zhdvb8UMQQz3lX8EeFAWKd/JBlsp19EMio6OGdx/ALTkjvsxohZXQspO4RbE20q
MlaZxLgAvihCkO81w6cuGtcC6zVfaRjxs0vp2GFdTRiQHXLhvbFlmSMsz1/2DEiPm+RgYVR36B7I
j/buElQl2tdlCEpUQO6OPHD7ItIac7PZ/NjFBO5mqTmQWJl7L3QW+ALoMLQIi+AcSZV5BKWCxI8r
yABwW2FGhfOGVlxIa0t/MNcxVii+xq+ZjFg6mZ3eyCSZwauQT0fod79mRNVOHdseL09R2PZDl+fk
GjT5RrKDq9WZfbt6DtiVSnLzt+Q85G1HarSH+7R98Fnf33ckXooKD2Ule1DITh23hSGwHlDhWIZP
dbvJAKL1TT4MWZGvG3TG8hVu/MPrFegh3WB9t+9UQjnTgp2mXVtRKwLMDT93nBNSCPKrWBoadh5u
4YasTYK+srZ5lJvkahj5rD5YiPZJh0mnng6dMiyRBrSF/KjbRNuyalkr5kgjcKkiEgJf7XLCi6Ue
PhiKNi3HYRo+9hCUMKfwxcYgDQ3Skwt6cCa4omBvfhMwg2rnM2yncOldPnaIFsj9aydLnj7Hsim4
lF6ST76hnHqQBvlr9CuOPZC+ubq/h7n57m8B5gBLblkD73ppFSz2NeieR1MYUc5TfBKymMYLMr7g
Ect6owhasBeQ6DiuJ5R8FVQ/U9MTF+X/QO2lLc2/tNKXlRmP+dlROb+tehT2CAosySRXVq6Twy7B
H0UDdEOOrR/qC/ld18S20kedfSnuUpBu7EZpJy4mudsvpFHyd/2o/cdNloY5QK4RYNKvuX1fKXEJ
KxMylLrWVn4o6HzxO83Luh8MyV8O9ap7MKVUN06Q5GysIPdUT6Iqnw71aIBBfe6/3aiw+pkiOL1o
ItZEPRrNH4gVIpH+LR1IwLZ/rhMsipaH5DvR+o8pp0MjPTYHVUKgiKSJOfqyvELlyTrX/bq4MHTK
u2vOVusUJkGmhJKM9tBNK1vQX2Wln7vibv5CUXjjCJQ7r5Ix/J0rCCsZqZ0Aa+AsZPWk/5Op5FE4
Y7qI+mHXM9VKdQy+VQCLauhK/9pgw827f8K2g+GQfN/N9zlMZ8YI3A+b1Y6xTX0WrhASvb7pcXu3
bspkBjLZa4B3VNd2R4ZfGjlO2Lr+3Bus2aVinXbhU1uFRQQ4fOMAb2rnwCgQOSZJstyocDO0NfRM
ZBdCbaBUw7nqLNeVo6D7AeUzK7ZbOhCyJankhxOu9DdTDFQNmPJEjJ+8yGNSfzO5Z+iHGcrZKnZH
6EW/cOCGXi7EsaEZeKS4n5hPxRWBukKfG7yX1WTn5xals9Hmt+2f+GbInNjhQyyXAXI3gFJ2tmbb
i3rv3BytFinzDIPlGrvxMv1tHRoN7utv20KqoqmD52d0u9hY2gQBLj2c5iXoH7StRsjJ9UfW89YY
y2qoPmkQyZAC0OrlIiBT/DWRuYxafNc72+q//Ao6Ph8oGllJpXS3/TlEOGNS0HLD2PUhJxs7qJTl
ohXsbqbm0yHQwpr9nsNxS8aW35s63j/uRlXLjrumxXrusTVULhQnIkcq/SsiTPKeIdkvwPmTv8rB
KwpsZZYuTo/rOnK/5hWZgWYLNrWx1Btdz2nuzkfaqqCPb3NSGH++W0APURn4eU3WGn6bAiZi5dn0
00uABnhve4ZT6++k3RjslCY1+P1R2UZmnkoyMpjHqQoIjMJt+fVAaYbJMDoRvMnZi0L2lE7LkNC0
oXonidD+eR+1mBsXSBSqPoFZi6USgEBxZaZuzHsSBAdo2vXWqVIljqHvrhFEzaKGW8FTUxSbHReu
ikMMkYo/nZL5lv01q6u4j4TQt+UK0ILoiwd+FQK8+zjQS4SHaA8iOICrp1/yDxzdXwJHuuQgPNur
YKBVq/hTmt1d84AprvqI1RWAB6C9VIw/GhOK0mqEFQpDBxajTaw6m49vDzbQp+drndHLFQyGL8f8
i6JeKW715Y6XqWJRI+QtxBkLbZY01LpybmiiAMBmMR0MIvFalQLoBjrXOu1w5Q8RvYDJj5EzDiQ0
UBw7JeRukfXu5OZ8+7JS08Z02e/fEXfkdofaN1w+qdb0Kv06On2Q2zHeRqQwIlHCVS/MUu3wVekA
pNdLtXCrgPOXor9CM6uG0NaUa092Lv/SKTRgvNqNJHU4V09tnKbERzfFBzbg7zj9iBQF2e/QECTA
/rgJAfItIldwPkvsXpvNUmcKp4XwVdsGQdUfJCGXAyk9STjeKa6INTCZp3j/P26Z63SROYGYxjX4
uyzUhTTn+TZuH9103e3CKAsaP1+DiKmemx4KaKnCdCxL4XE44olMgo3ivif382TITLvSIJ6K2C1r
ZChvHqP6WR+oMiv3MgWqiBMz2sKkhEmNSmIIEwNR6HgSeN2azgJtqSXp13nfG11IHBc2zDJC48BK
ZKXuU2hw36fySudsMJKSi7Kz30HxaBcdu+4JoJP/zZY8Op066xLktJP+FUjGrCrdBugJXFRb4vhx
OuR6CBVEFaHY/w7DM6BHwSgUhtOmZmuXMIu6kIaRo9LFFHn5edOzNeweuc4hICPwaMlvmAr2nZKs
MZDCykwIvRNMajJT/bogc+ftQ8uMHyMazjkeCzWFOijoX+lYRlpMDf0bWjpruobLRsWrcnhPGSNc
tuBHKfTTrfm/LRqHI27CCQ3KrH1TfIfyx2ZqMr9xrHGjs8jesB7AM/rbEOhr/n80l5Jm0LQ1is8F
IJgwlWjaiTozRGLi4oyec9oxCKJznWS4FShmupz2CK4wS6LreBkdhLUkrTLk7xi8fCxjlLOaYExb
im+I4HCP8UZ/0x+8BwSCcWyScWokJ7zRIY7YzMuxbwQzgBVhJeNLvgLUUS2dQD5vntp2xUDTvDZZ
gja4mgi3vlMkZKWpKhL4MevisMOz9jH9mx9Pujr1hMCdmKYs8vYARFhukbSLgMv6549TQ1DejWXT
86kR8ikD0iN64hFMvIwHD1zWvrTwH7blPKXYSLBXcNklpHzn84jgKiYkygcHYLfS+qxvXUnJM100
uw0RtPcTH3PLSXhiG/Q9+Izn1qLNVIuGWB2wS7nF42A8HUod+gljrLlpAWj4lMgdTkVcXZ6Gfwva
d6ePKj2dgwfl5GM57gywHTMMK//XbkSLSaCJZr+bgDM105Qn25j9dVw6qFPcZS8aKtaG2L5Pc4oB
sqyFJGbytpg9e5E8QqaluyUlLE9QcYnffTPzWZRwybWuB9ZtJd23KCsO/WJei20o5myUJ0kheSKk
tcfnS8L3gptv66Dl3j9QYv0SpJAajCF+RJWrH9nvpx9lRCv2RPR509bH1Law34h6MPyzuad8UoPG
W1ZfzKRiOXQgfBQx4c18HZ20C6M80P8HlHUkhjqTYXDv8YfYpfBUD7SCvVZiLTXiQ9KyAWdpirRO
QwiacBLXmXd6GDdpObQlwNftnN8EUfobVlbiuM5aJWWzdkYFQ/GCaUTgx/wV+WOgLkdNVUy9395N
NLAtL5O3s76DJyY+pOFuP8E6aCOGVoeKI3MKI9vh5wzCBkth/nto5kaU+NUAVtrccUpVr+GhQgpT
B6cOqCM9V52ltME+UqCWYi5/JsUA02PN/U8DZz/+P2MW/+q4tcdy9SAPBlob8NRmsOOawrVVRo66
1fI4Qrf/dLq/qia+ZLOM67+3jk+JR1l4YlXgWhDtekFrrKWUGatSVMs7Z5yLDqU6DS1/swkcTAky
54CTj+02Whc/gQT2wk4Ic28eIz7a6jn1pPa6yohMpO+eYd7CJ16LnoAf8ypXTw4K3yTKXbRVv5tA
FgGoWvDd3qO+s1FrQb6AuPHXlJ7n/BZudD2MRJ5gVmo8PkWh78qubISlpABtApX/y5fEVI+luxTq
FO7lytvyJFgjLl3Ws83PD29vWLPKyxmmxrHU+9nJ61rfj29VAdqI8aiuYI1FZtICS4ZupcNnzvH8
7kJITzcpD1D0ePB7L4h45b9ggWHyKbpbk8hQ+Q1r3MbJ6R4EeEiiInchVTOiBb//Tz31Dr3Cc313
weXhDPibps+DFgry4FXJ8HKSLbGySw6iP6OPL9U3F4et+fVp3EYftb7joiHF3YF0HLpaGhrVcjYj
aecAWT38cUpEZB2a4AUDlhtqsCYrb3vt9YZyKGEZX2MmWexwSNSEsB9IGB3Cy5eneb1MjXYiWoZL
4TO8HpDVT4YTUb4oD6eekjm8cXu2P3v1AKiqL5g1pmRAQ+ravllpX5zfQbLEtCZ0z0tmdC3LNaVc
elTYmNbf0o6GPtzGd+8p9BWzAg62dGBHJ3Mu3nSxkn/i6gevyPlu7hg5ODm0Kum8Zbc2+gFmcPkJ
qIxQ+aDP3weJ8I/W9TNDyivqYMBooRqZ2k/NQ5WNQKz2kdsN4ofbVtMWV7bAZ7klVIgVwHtcc5UA
wGmjLe5zzg84EFhpLf6WIIYtMbxjuP8mV4nLckNr1fcm6IuqeuA3HikibrZuudtKSbcX2o/OQU9G
g1abHJLwTkW+4Drq82MHDFWD9h6+URswm+vSRrjBpADFXb7iRK3jxZ6xFG+/1gUJIk6XXTte8Ls9
+yWvOaRbo+q3gQ/4Qlel0gUZYCN4q2yX77rFjAnBsKVxQfOO84R9W+5xOY5qSf/ML3PJNVBtOwcs
ikoLVXXuPtQwMgPVb5cYLWVV4zLRYbadEbvecJKOfQlsjau0AOLg3PyFRuQGM04bE2xf5M8Wnowd
AP2KM89rEMGXbe8tgypGrwur/9PgfO20aaxt4ZxJ48mTNlrkPUrRLefqqGAwUWv1BQdWnGedVbre
ntwFEbls11Tpr7HZa3v1IdRaTjiSM0IUcEG3ULrT4OSoW8IKdkZ1QAaT8vtI7IuqVCCP4KxKm2T9
qYe8pYHu1UaTnmAJFpTucjMkim41BAwtVuo1+wgslWCtrskQ/EW1uHXQzJRkGQl46TXJdqpJEM4D
5iC+FTGHUzVt+zq4SvVzO+imllk6sEph6En7MaZxMBruqnt5IdNwFTX6uOMtYZ1h6CEo0grIhJdW
GVu62RWQB8qvZBPKUMGQOsgwYn9rH3nZD67y7055y/o+ej5tAjZIi64X+MxbxiCMjTnWW5nMs7Sq
mN1Ie4kesrL4r+ShuoWDRfGwWbzXVa7yzqGdZYnZoX1h4siINygbWFvv+r2YqR/b1H1eZ43zGWyH
XW6NgeXyWIaZL3A8h0SLF8UkyJfvDMlNodsyeCuQMi9zjQY/ikhMtvQpgkvz5IjbBvgddey/zr2V
uPbyaFEO+jH/1FnTEQrATn4fDZGmtJbJiwK4bznX29Hl6Ot+EVHPA+7IznhB4vPR7BlfhD0Umt3K
B9qQp+vk1If5+Nge0iuhF8eWDUvaridaISLC57wSC0UlQcpAEYauTnRYqWC9SyNuffr2ORHka+qp
bA5cX4/ItR9vo9dtiIUBeuDArIhPfT9jhOr1q/Hn945nzQ4KsxrlA8oLheXDU7uBjY5NACHQ7mKw
edYpRW2xAuxm7v+tt5xLE+lcy15XIgiQaUlRLJnDCB8SOxxqN6uJ3IHExfbH3oz5sMBDSxXj+ud/
Fg6j2dzILu6tV9eLmK/8vZ9xs7YyyWuGc2v6NUaBJknZ9t3p43KSLzJVkLrPTD8fWDOYdiaIlNJg
Mr0RefBeMTdrbsxvKtNbE0/Qzimwg9t+xEFEsX1phtYD1IKywxYMMkJTEShnPnD1APu0m5+gR7cv
w1tP8Y0SqeCYRcRQk6b82OFWBp1dXgznPrW7wq0wEEbksJnryQ8XbKR3S7d2JQBi2bT9bWF1E3p3
cs4PlFfd6WXEbN9JOml4VGnPHIXkwrSmqZ19C6VJbqKA1O7BpQDpRQKGZ8LFaZ9wUxv6agatJ2M8
cF8ZRtPYESAAewTVcJQCzWmocuwZ4DPoJ5HdaQBBVajPG9uIzReWbJt4YyyOjz/2apTdUy5mLSOU
CiKvlDI3TlhwIk8bkFgiDP8e9NLDHtibOumLqz+0DhoHnP6xLYNNbc0u1H7vG6ONM6dSVjdXvX3Z
UQHHgGkgJmtXHX06mjqdlJBVJDqG8g+F3YMeS03+beF8ofNMG01TQzfpZXbf1jrKXOfjnNYp1SD6
EUnSKUfC35wMLj5S3OluV0dKHMN6c8mlvZ/WStANIXT4pnNpVt0DEPcRrB7cXi96V9nU5bU0UXm6
0xAxX3VzHAf/7DSfIgaMx+cl//e2nTu74luhJBkip8Q6B2/ZjWpy4WIEpvI/QerKpsbkOs4EHPcw
flbWOE8powv5CPGDWJt0dWcNka2ATTFvPB+WIBVk5jV0VgURRP1NUMVh8Og9lOeW/FvzmfzuSIbK
nu9i+mNGdyXMD0T6PdUgw88RGFXASj3orpA/6erPwgT8wz8t3W9bydqeV4FQJ41Et/Jle0g6OHG9
JivM2rnmWKRX7Ujh3L8Zyd1T4ygaEQHKfVmvRC1XRkZ8mpSmMxT/uF/DruuT8pl33Dituw9Sf4oH
tHICHFcc/sSymEIYcfEqveCJ3gyg9w93oosD28WN+1fS8w0EDlAuwQKLUZ9T40Hmp7LEc33Cdnhy
wooVlB2dQ9JFsKiC2fZrH+fuksmhK9nj/UNozBhyJr4KCFR+1nA+OnwzsbM+5TSDZPVYIeSG6Y3L
wC8AB+iD1endQVM9+9Na3eSTjPeCnAwOU1bUTrSmRAtEnrE9vx5IfKQovcp8qxycO9aOcTadlRAQ
OTksIi8uEvdEuZqMT/VgR/hmtdCXrBw+hmV5Q2wHcRuss91amELEP4WUPcdAI5WYu6I4R0nf72vC
1QoXnVE1eFi3nDTomyfCICl4QkFDV8TeEJxE8rN9xgbP+V12s9ozVbi4BlGyBukUUui1FUjVXXn8
tai2z7qqbMKcgU+IDlyWGQcLGrfsNFkElgoXLJe734e8V2Zlqh95dyQmRhrmlx6KC7e2XNchKZoL
l4J3cviQjpYJa2Mxiijy56toW8zYniXv4z7+bhaLryH92mMHvGR1OVfquB6jbGKw3omDBKoukDBv
IMjSx5Hevf5922pfLIK9OgNGtvX+jfYDjBTrQZMNQ3eM1yYt8kuZyi2O/ZEeMncqF8Wchu8RkAHR
Zzy6RIHWAOusDYWIUdatf+rpLYKdz5XF/m11bdPPueFlVJt5qQNlAwyLK5RQsexl0pPpSbq7oIMV
TVjO2qjrwjwDXy2PoaTjDXettmlGO4ZLoo9MG74PamgJ3Efb/1rbtYLbXjhf0kzYUbFkpqsbAfHD
0ej2sqqM2fw0ToUE8eDEijteJPrRCqA04z0UNUF2pdNR2016QP3JJpUjSF58TvS1SZyhTYpU9DwH
NzDnJ4/w3BheO/L5OnLJ8xAspZWNmiFq4S5LdQKwg88rR41PDNkjaGXGwycd02Ml+Rr4QYpjFtdN
x3PNNXUIKT3Q5qioHmH/jw/67p8FuCSKkz695AcuW5ypIrQpZ6EewuQlZLaCAs3wo7iPGnk9pTqN
JkQyUO5H418IVaDoldOaeG2NNlJR0OxxU+gDV6PFou3JjUxZcyddSyaIvGSgvtOO2PLwSRvvimE+
ut/OJMkOt4DtrkL5IpUW72CjHkr6rj6n0Wk9/3AZpbFLVSOGC/9Sc6dqmxd/TtfZpi/3fb9Q+Fwt
gYwNDBca0HIxilMyoZ5BePXjmGZnIuq/oLQP5Nc6mgmG/SzgsEupCH37crS6mOQ4NzTc4xrVIsBE
TY/gkCin/uCMpZKiaBI+dQlgtBe4OxPOcBv+M9JLZ4zocA9+FXzZVAHrD39qJXqhBdgEFLMQDEqt
hkXl4nmuLELk0kWQhAqKJqO/Gqo8zYReCy1o/vyWJP9ETxk5VRYxm4eSv87oDtR6wARI26uy0sOm
WOiuiDo0BkdEm1887mwoDHTNRMg5jqZz5p4b2Jl7CIdQdV0Vm59RaFppyzkxmA/p03jvnp6AG3e2
y863JMA4mr0xMqmimMavHMPvlCJu7wSUPJIDjnbjuV7Vx3CnfF1wvsYCespTpk7TnaBgSMkpjq7D
e0Nz2bvUNR/cKym4U/Ek22rqe1uh195xapM44IGRlZPUZZ7r8yMr+DmFIpUiulrfqsTEugLN4SzY
wV7XSmuA3sGQdgRxdKgSkaQzeTJZtZqSENjCgrIg1PUNuj6tU1NQeMRjOZUC4eZ7ys0KllwHQOme
e6c7lPfT7M/pcpb/nkJmPBBks0RcVTA7MULVU62DtUhHjJ9V0jN1hjJgQRO5dHxvS2VK6694As7Z
DLuCZHBtKyBR6h3n8WYnq+6GCok30cf6aA5nRIvFuiea8c4GOLfEktVnSuG0zdDgbB1t3SQbc2mp
PM/GghbemtlXA+v0sJq2AWFvN2+ol3kUw1YbpmXJlBgi6yv3zlUFDpkyfVq/yDu4M41GKyZH4VT+
/II3sv0r+oCOFns89XnOn16EDR0HGUSyYKVxvjrXOADZKHAgbsySTEdT7tdhC9ZmgINNO+cYATTw
EirhJexYoYpgupuNVNepcd7fvfcYNL6JtngOqqqdwzYsDXPbpTaEDgEcAPtRMisGeWgdUMwOdvYK
QI/VrTI8NRo9/VEGpyFzTXlL6Nkaw+ipPgxS7MrEjOJNrm4nh1sBUTJ9mFRLbG0RwOgJmxLBfQFK
RN0YxxzXzuW8RFggA9iE42UrsLjGNiq4BeK+4OFgioJd3F+yMhDXWNgukRAbTT3TlrlBs8iNa9ff
n7DzoBBjbeMS5c8OfbGfiHQyUXKHjdpu0W1ApEiJg34QgSPmCXU0gzsKn3qvpIFsb6TAJLtw7Via
FbprfSry2b+bQTNxsOIsx7oxUuyqoWr1lD8lfqHG/Ganm1J7uORb7CrvzY1iEcuS2BtdfpjAQBNM
D7sOVlmNSZK9WS6+yJ01XmhSN7BHsmF7q6z8Wk+n37m7PoJXPB7GyQ5VE8sqBSm4LJYnpcrKYaDo
V2747HhFg14zdRrWbVadHz+evAskQp8Qj6ELQhDzEBgMTOFW+cT9Dzmz+/GAl+r2BFYvjBoOMyC6
7jX3/ZlppSvem6iYvW20FVXzdqrQaLPyP97kPxa2EVDma37vcArsv+8tkvmQkYktG+5+asEcHTPX
y5X+0v6/HZZqDD7BoZfXshIF+ai7Q3cf+ae/zJN+arLsQrXRhZ5VB7o/kP80SH212OkmtSZoojXQ
dLjapMZZ/V6I98VryFukA7UfeS0gcXOdDSlyUpyIYZRseo5aH4cBquAaJKf88wVM8ifhSYL0e08e
1c0l8jbgV8QzbiJuE13wkWqrq2+fkOGGUcBt3h9BviFaqh0ZqHJtFeUN1m3QByEeoaUtHqcqkXhh
fZxZ7UaWyy7sVP0c2KNSpclae1hLwTXgSjqJs/rc4pC06U+VbY/4+P5MNnQd6y25uFSv62cwL/2e
eUslIgLtuVZQbTOt8eq1IzUb9EdJC5c4R5L4PmK9mebe9fSueHUiQ+APk75Vy3P8l/n7u0na/0DC
gZWnFPs/FKIYCtGMsA41d4CrVWHVz5FnWxafn4UOKevEtsoa6noUJKBH+Am7KRT5KkoZbzRD2dAN
GegbsNZZQ2KXxJ7m2i44fNJDE8INMRHflBDUnBHFlfypf6wjmEEc7d8Pfz3nsoa2HxUEh690JEH3
b1TDcJm2aF/njhAgAJwvy0VI3I2mA++ThrfQidGbahRaYoE5qf4QBE2ziVfiLaztEL82iFzQ4P7X
sWeqHJeSwfSaCdorHminpkDjqXp35R7ADUr3B5GJqu8/3lcR0r4ZqUGk/aUwleZXxVT80KAaz9ck
QzEfK2urxPk8oGkBV9XYiiBIjEwOdqL+KfB4oVaBw8V3XdWiMjSJt8AN1qJksaR8usoT88gcRLCb
QWwwYhDhJ9wE7CGQ6sNleX/inVObPg+VAmuT/TbwhEjCCgb0ZBQyWgmS/wjjR6KLPMM30/xI1yJD
mUBX0d6HYnXNy6vJ/2hlPTi3pFQJE6eRp5JbENfwE63boLo+rYbVFcsv2hLfM6JHVD9RkmMYIYKf
uZntAJbeD45+QUlMdIbg7+rOV1J/VTZ1VN3rfMplBwethpz69cbXGSdzXhQDoW88qhBxSO0ty0px
WqbzQEaxkUrnbxp+VJ5QbK13y+paSmDvf8Rp9idCQ/cxJ2Vpr1bVh+PWhzfT9BAOxcwShmgQ+5/c
PYziyYQgT8mkeVMCoy9pFCczHxXVeH/bcRtcArMQHkfA2GezEi9GiAFUhvvLHJMFtenuz/eSQV6B
2z5d91EHunQ5U3o0h68o74+zFG7XynjTs2+r4RtsWJgRYx7GlipCapgTHTTQqa90tV+fauTqwa9+
c6Y51Nm5/Nq9qIQqJulWyVXTC6NoYqstRSkNblQ+q9tEfhqTor012xI3kUEsiTt5IvxQNiE+F+eK
LXliU4eZIUaOkP/yKRlt1YCS2Urf5oaiKwxypBJnOp1cMl8xKxXobOwm5Ji4yXz+Q+M9IGkXIbKL
BGLEv4eQB1aWW51WtvpRWTBF+5XhFslBUUDFxmF2BYowRfGThe6MbdAB3oo/MSwvwJswQRa7ElCD
aoiiVpomtFhDf55W2l3ajpufpwJXwB6fdSjKydRMxDXUSbSu1/OXEsYMSiDsaeBJdMwLm9qYnj0V
cl6d34J/I5opiuuJUPeY2te1kLdqqAwHMHlbMqJnkjUkWnGBWnfKFz9x87+F64oCHqPWQgiFtvcI
jurEKeQYxa0z1RlJc2tHlPKl56oNp7yoIulgYZm/bpmtux7edO9cD/+5A1aDlw9ADdB+4UWRKsKs
5xtmHhoH+4Krs0u+5NBzKjoio9C5V0S98cjQ/rwte1TjiIvko8jKukIuzCsjeIVKxxXUzXc0y0b8
lmlno0Vs6TGJ4yBq9DhCp/oRvmqbEk8pexypABINl2gCVC0vcQRriSWmEe3PGNV3DgAGowufcbQp
hTwlF8d4fqqdyXutNyyvGkPI1cQxlMv3wdGSiV+9s7ZdZuUQnC+KKSkAmnqcqtdTEpoKyyLK8sdR
R119BAfXd7Ya7/ttZx8tDjZx2PuMWIzPEjK9gOPx5cXBbkyB4EJdiR8ZhNslMi9+k/mecVV82XdA
wyW5TDsBkeUVIlftYUal+GODqKLG971z4ExF/pE6XyYtsYadkZ3lnMcRzPlUgHyjGeDodoNleUSu
EoqcV7HtXBFIRkX5oDhMxVAySirqnju53nxXi8VxBzu4AbYR+C2yiAKeW5L8rxIm9x5a+aFeYO2j
CJ0UTEZwQVPZg6gSB2c+Ui0f50TKJEHr9YymA1k2sRLaYKMVT4OmukKhVYSDsG29pIpd3qHEsbbp
E+jYjaHWpJbervc+UdmniV62TsLU8M6b5wfkkaBJA93XkDKFU9ZSPAzZOzEFoEc3/y7t1ctPsM6y
e6DMDcrNT0CxxzMuZUQT+A8oLoiON4TubhVKFk2fymYiKXyBsjKZxpugOC4JJsuTDw97tXHHsYSS
GgBZRbht0mcgM9rHQzOMspk6thh7lSi5UmKcFumy5SsEONmv/PdI6c/4rhsoiYzbKo1mok88Px/w
dBHQvHzjoWPinFuQNDCCGx6Ap8rWoS3QwwGwDWWVLo3343iPJKeIvYIEfEj3CVpwWsTyd2ZLHNv3
O1qrmPLd4ozS9grxtcQsVSB7Xgkn+WKXJJArHCsP6LT6wGLgGQpXGKZQTNEOoTgEQRHZt+6rSs0J
s8MXL/BlQBJZmNGQGGaHsH/R75oZkLGM5F+8oNmhiEbl8HjLlJQZix3dreYRg1Qdi5AVQfWs+ZLW
vfz3Yy5ynERNWf3TwZ/oSwl4sN2BCZ/PJevkpWM/ivOYZaXgsdU9rKYdWlWjLRD4hV+1nr5nwWqA
zppRScjiGz7yFIxdhO1Tm+uUcIyL914He+aYGIS5pXsN6DuP07GXnBLjNDKj49bNt8uNr7SCcIgf
CRHrS9VH0z8wgzcRZPNKeh4eT9icqNksE+qTCPIeJVKK4/g2mvHN7ReakK5AGins84pcMA6v+Vzq
pGQzrtqsKEUT3Yd/bRwWe3P+MrCJZfXj1buO3rKpxvmLmkQZ/lDDYen8URRPBKwgsn3TNRvE86wY
PDYiKlQCCSrm344jrvGJzg6IsXrU7wljh21HgAAC+EhK8qF9YF9YWQHEFUJT2npBpb8SHZnvV6wd
X84yjbZ+gosWJY2KnmnPNwTGn2Iz9oqqHivzTIotCPN6SrK3RcV2XWZyqER/CPjVdLhLIU4OAyFd
Fa6tQT7zICOzwSN4rNiaFvZ4rYW4E+kceX5GwcP+zZ59pyGpYLIHhbjVlYjpoM7KNJEsnkYG6ABv
3sD+ziX+KBAjWJuMQWT04FhYRorFYjLe5tBXh8dTV0VDJ/DMvYVIOkZ4QzBsYD3mg8y8zJmHyKXr
EIpKkQMGZmBbaZ9ydXuxVam1tnBpwIaC22d4nnPMkkP9JxqtoACNybFFIJG/BH05pOkqJz7Vv9B1
DiDJGUt6Pmiza7CqJ2srccMT6qsbj3xAdyvJkdOuHEF2+6erMn3UobTS4cmFfK8F8F4rPzeA2hJy
cS/07WMZHDLGfEubuHc7+VSEk7MgA46Ns2Lvhc54DpLjdnahjye9BEY1MGKlAVXUDBdEQCLYwjL0
Hja4chxSKFdzV6RDmlvgQ2L7bDomF4mprjdBBaXXb9QRq6SuzeybukjPj3KH2yeJ+QZ9A/7iE6sd
gDSoqyBEeb//GOK12Qwu04zcgWcxFW1Ol9QWoPgfrwpYt2VTuQ7Rm2yI6Jyko2qjj2gSU0578YkS
0Ux/K7tKrpmgthpSjNsIlbbkyFM7foPXXjrbj592SB7AUatOTNr+6UMqtUKMKlOlVQ6Z96JntRvR
AZlF/ehQJ84FbqMpEwzZc3ANHgU63lS2eESYR3APK74TgtR89WQZyB+8p2DJMjSkkVrE+gYp1BjA
0OvNHVmzmMBGFjQ7yCglNIJnZzxhZCabdL3Has0l/lNT+I5KLng7X+NNI7gg+6sxlGcuYVi/qdZy
2fDuk7kBcddCDaiaPYkNLx2ecalJRHBRt1C5IH4kcooDEYysW49MBCZl0jJNy9jwnxbTxxBH897L
d1gWWGnjXU7isr8HhKtAgyFb8kAPjm8VT0cOFyroTmpk4UXTpJCIGZUVxiX4hEvCT5B3eT16IVo9
3gieUoy8hefhnTfreCk1amQQuYkHfD82yUd354M2wrNE5ibSpYLrAz1vmfUO/i9jnhzaOBYhwkDo
Z1Nd+qKm8ptfmk9WuVWZBcxDtjdvmJQZszATYac/WLQli+rpLUuwckNQ80T0WAvBTV8o1+Ipa0Ze
ffv3dEx/p1VeHk431mRmfNJxrjhb64NgQmiWzFovN4s/iGaYIgbYN5jOnzVWjlBd6535TiRAIytD
L87VRFdcIhzFlqb/mXPCIhqnq5TwT/QTxESDONfpq9dw6yUhpXdszfgQgBfWP/sCu0zP3fYK5l9/
TBCr93Pc19LqwQTeKIIyxirMa+D0jARTuxk/e3g/eOyJc93NKeVVDQ7wF8qaFUDFdWY3SVxeN564
WMkOFJc2g1kWCQW/ebLAf0b09Am5Iz8Y0Ccgb4xD8TcqJZzFmyryjG8OpSGaBoe1VCDNeT/+DtOi
fjM+7rAuZ4LnqvSgMJlPk6OC0/ZnQVHs3PEF3+QWRw+UglZwM0Hj3RtUizSmuAGpIqLmRqBW/Pxn
rpwFaACF/2SKABCpBv63n7XxF5fFW5kmYh8Al2j0aySrYyrp67O8nuTVQEw5ReIphYSjWmRJ+w0F
SDe4zneorbswXtZrJMUojqQrwKSBwpvJS9JVWZTw6DU5+EJH9Ng3DRIgieKb0KKEcWjE6A65GVXV
R8BdE4hEC8C6QG+2If3mps1+QgGIfyHFzriAj4LYOJi+KY8+TdDBOk7TPrudiSn770Jxi3PbJF3+
8XpHU7dR47UEMba+RWJToCXQi6z081uiqqqFODvCoiQWoRp6BE0cG/4oRhDWd2q3Qf3yhkID+Bgv
zW6E/Q+KxIXj3f+Hl0jwiA0gYgL69ca4BpVmO0Fz7eWzNvsByLujBtTZ+vfotBj7ERDMSAc9HvfU
Ngbr7uJ4aFZ2sxgHdISTjA1ezMtVpqJC80HXwt8u+H85tg+co45zp70rVM2OwPyPqdRUVmAdG6gN
lu0i5/cld80dldHP4+wpz4ExY/opSGVHbnqcGG7s0xaI6l2lFvOQthRmWdM3Orsbs4uYyLR3TrR7
dNYmnbbDUFwfMFecTabcOh/XaG5ASSW7PbndiHwJOsblIbLHLrV4zJB/z7kQyyadXTXdIcrNdl5u
c03X+rHIOXzdKsP4+5glZP9TWo/UEOJvjC86mIqQda4VbPHMWCODCVVOPH99SCfQaqvtMZ7Sgr2G
+y9S+vCMSTezL3rvuUFZeYG/p5YWiTstUEzgVhpmT1wsLtvxB37/6Www3gZGKffbmdQqEd+Cakzr
XQxBoZpFBw67emCk0W5BveTUbVWoas3KzuHXM4G0LTYtkUemEtbXiWicHkjrFW09i5GEgclP0ZCK
kGhjGkzVcAWIvRAgQBlWoelLX2YU706IESu7uZ3yfX+yYnmY6tyuWR5ZKnisxx72jGQg/DVzreNR
gg1xf6jYI+w3lLK6uimkgRQ9hsoOSUGvoF8VqpzgBP+5r2lG+n4Pl6MnFmQoeu+QakmBQZ1+4LmQ
UU++5UvVeLNfwX2VZDLlBLKftLd+xni81Hg3Twv8q3D9WdAdLBn9er4OAxdg9C6q8GI/iHUAaauM
yp/0MCTtE2KRuuBT7nOJxpQZHa7JD5NGw0ppsRU0yfFVN6vz5jB+LSrcDu5wwdLobfMxIxLvV1dv
DfVuorgKo0r/JKm4+KITs1DEii2rM5Ipe8uCHvLxYRi2VYU7m/4UGE5it5rT52AtKtOUTUvIzoGq
jOTnbxLwMKZtJ/v8MuHdGcgmeWZsDNqrkdnZYehj2b948XZMG0+DuBrOs+mkWx4vEqBVR+2hzjnt
/GF7R2a52LvtxxDHfc3E6Sp+1z8GNIUEuCFhCqxV/1aVXl39bgPJuHD7LLH6/HgH7d2zVbjWNpcA
P3/VRl8tOF3m6IOtC9EJmHi2GcYD+Ekg9qtKL66ntBWQT2AwfP5gAda8okFPNkz9FfUxc8/gXlyu
TKyeYUR/jYEo+3+JK4MO7ydJP1EZgbzR9JjeVY8xbcHHJ7kNPiYjdaxxht0M0k9d0mpiZTrQWw14
cSnwj4WanDuqLitaedRuR0yLC0FTOfa/lDHdpmhlO7bn+ZOWal7dj/5wZeF5zw1prRIMP6UC5tWQ
QwCTMA/ZNA6NZqvc7DvMc8I3nOITiPDFLxg9nLSNJufDqKJhyHft+kdOqc1fVh8mPODjGYqWi71r
sU/ozMVP8LN1sM2/ZJeasssjNEI4d3SaGjVPmzqADGe1QRPHiVTRNj3XRii/8lvaL7L89fDbxTcA
F7o1HhNTUy6pc4XE4dBgXsllI7XIf7T8DHm+s11CsJAFfuxYPavJ8N4uZWM6KS1bRt9jrFqO1uWY
o4K6B/B2m9epfqBvlhwUT6FpbtYdskcyDw+6ibTmP5VVdQ4R1AMKBJJMj+3PBVv2CZYsxRzPDWaw
yaWLwHG2PhV6QBRy+3a2viZ7WuFlr0pnuC5kRMOWxvj3F+HkgFuG+lGhz19m/wgGznTDOklR9hym
8x8wK8lRAtEvlxmnzp4N/mUZcCR/lSEbv9MASNTHIWqNj8AQ1hlyBn/JOa2baPyA8msi42Z5dTll
ZL5ktTUccJvAGYm/VkHckc0Yy41ysz9vo8kR1jfWG/XzIAt6G6mgs+iHTa3MR9C85nkj959z/Z3W
Wp7Jp+JoqXCQBndKaXF43M2F9LK9XYVivRizAapUD15SV5rfFiC30rS6HrLRU0lct5O2baDQipD3
tceV4JhsEndu8xXFvY5mjSIAp4vOFp9h03TBVXuPi0uG4et700szGBeG82l6z1tsi2WlG//q/zZD
Zmc1M63k0yaDeVi5ygpkmCgDMYdxG1uhFt90jKiT1c/8iUDFqd3eJThV7lnFskLCg+LdA9350NQK
DGs30yI9R7YqxFsM/G9EvSqHxvYmy6H5FhEug2jk+93ufjXtanUteordWDWh/vuH7amjcukgYrzV
cnY2teuW0dDFBvu25SmMcflZ1RgSztzqV029+b7NjJwPoJOehM/D9XzoyH5op61TKDMtZ3xcscDU
EV5fw0sEuRGR98uVGhOOWYf8iEQogc0+hDkItxExzgSEPUcqVGh6Ck9gaBEJj5b6OGTdxIHjEj7C
OqzV7KFHg8c91NJnu7vFlyuVd8xDUN30p8A8XXUyL+FweuaJrs5BigzF36ZkQ6nU4cJlpwl6bonP
cSDZVC2vMKcysEDRFWlpSF2v6vrhdgb8KGcYqTujbnFLcAMHO8avJASTet+TBGHHBdpeDSqKHm5l
SLNh6R+4fzG4xRYsU7I4eVXJmk9KMM/4R/k9zzVKPDF1mVZXU1xqi2ghBohsvwu9YCce8sI2IAAp
Rr5PAI6oPlVDaq3jTBB+5r7Tx6hh0B604x8GhyAYQdG8hMCWMEauxdkpggWfMZ/kXfbi9eY4DNfv
hjI/ouyGszOGenmPWbwvXMuuEK9udCBULDi7BhJhawnrSHatnBc5UKQ5darEOgb3nHO6eC1RLF9b
/pqzc1Rs8R7RQ5aPRULHGLwBrEZUpcQtcZ/WhRF+JK5iDOLWf3O7C8VOujXZ9IFwEyyYzKYoWlc2
KvvxREFoYBPxktu6jJorLXpY/pAxWmDIn3p+TcSItDslf51iBvVf+JZdoAfBm5bXKVFtYxwwahyx
MogykxjRTHA7MVMUMZEg76QfSst55FRyjMlqR6jxIqV0kqX+mLX4rp4xabzKNlFBrE/fRXu7w63m
XVkQ4GBmRYGRyGCOMuG3p4lh7qu33gw4h5KT2Ce0Ep63SI8VZJdl3fi38m8+ZhE7eF6PAUrO2o9N
jf8YO6xWBgtzOxlLsMGxyORjBpXLuhj+ljHZ0CYRaCCaAKnEvdlMvqHToDX2j1aSIxrsDKKim1xk
9lWNB4JwaEYnkI8JJFHCiyCV4NfUkmmP9VcO1HGyBNXsQwa1o4NpG0RevrmKA2KgjE/BKhdjcljt
Au9zVdaDA2GKoobrwznwCXokgg7yPao8Y7NkF40XDxtbPr76/faUXlIprRWZpXuwOr/HLqXB+QvP
xlXj8LJMX+hVu6RXcKFZJuT9EMgjyx4QodROAbtsISwCotZaEsGx7ev4ZChVddJNnpjzmR8NJPfx
o+ecEFCQSa59ZDcGuiOlfPsxQF3jWvaCSy4Ao/Q4D8zJ+dh+1uG2VtGwxjNLsfzyCRC+oOGxuFFz
GcAJCByR8IyJPw+oWmcol1YkpGXGvm9zLf3FhifSDrWGLFKRpmqBDU6NpTxM8TsBdW0bAZVDrHRt
lMGc3P7tnblmfxFfziM6UnHwzZDTmZ8tbIjPMZ7wvt/ncEtufzwu+GZRWMMAAo/VHs2TGNugCyxT
aVD6KlZSKlc8cEgUKa20+AFYn17YeRYqxf8coagtFf9EUrifgEBiliC6wAXIUwSmwuex4dZaIeEA
sfzSHV/+g3BWW/v1wNddB5MmzTsaFjeTppJd3ZXrpMjWJq9M3mKfKhL6DwkSMeHpq1/tFj50aOMf
9J5ofpgjPMdaUtQFHJekc69nAIKlXtZEM6T+ifs8ecjLGtkggiQaSNfWO6oj+phD3fk6vqd5kEQ4
j8sL+o+TW3gVL7SULBSN51uWhidSCDw6jhT94wPeKBO0GBKvDOw6EH9TyaI9t6ZH458DFo0WgwdU
92x0Pte4jkhKbMtaY+6o7rL7FX2Xv15cYrX/DCQappE+MMlx8XvtT0dU2pMEhwAT7Ck4LZR3KsEu
veH0re0ZB4MI6TATLpMAvKeOK3xFlysryh5BqRgBB3e6twOxyAZHcCjFFky3tGdmjau0IwE96F5B
gmorbu2XXPIRQrRVWtoDOqtyQiQNByeSmWHFGtqjPH8bZEpFUUUtQWfRFjVtPnLVkg3sNjv/kh53
iuoi3Gt9x4PcA6lKJ9AruIpGNZaEFUQkH/M068mS9WlY1/5k+PfHMT5V6h34svR1ShrKxOdhC4yW
lwycu6bqS3R/TnKw57cE7Eqyiljg9MauiNJ8UI+13s9i3KJkaIWhD4g0wLeqidVGsIrvOWuTo+rx
6Wr2N2TTKloXQHD5uwc5+X4zDG+GK8KomlYCll4gY+KIe6BtI6leIQq5U1Jsxhs4+hzNOudq5d7b
KACTTjx3rRIYc2HzqNG0qA3ALjMgW3pdNpkBa2Hq98I6ifUNcWuvqZxfotu65Aus+DZbbvnOLovf
x8FpvAlbh2X1VFwHD2mKtsFNLXtPRJ+XCfXRT9cbVtg/V63aWMqK28F5b//lPhw9CD1sxVtpW4SN
aJceXIL12e4xCa1MG3Q+/7gJBhnCXURdb8iXwQQm2KHkgOw6Wtq9MyJ6kYvlLNuOQoY8De0I+InM
weiwRhIzM42RZx/x0SFw5QCexlHhCUXAf/ne3abfnmzvw0jVRXFJUGQijFCu10s/MqGIAuv8ciuC
IvvzrB+vgNQkXWPAptBxRX06Wx3VIXA7imYzQ+g2bY91Oxtc3ilN3zpIjPPvN8V0D/kfUIlR9b4M
ZwOf/2GypdTrG1+Ta8h5iB2dddDpwpT/KaIXG3lRprvwXVF0XJrl/XdRXUzQbYnKbFG2c+8hA3UK
7B+v1Odg+VrkpcDe9CpIrDXE5oIDGi3poy3OU7BAycjYrXcOTCnEyVxziglS/cCPz+Qiz3/Uu0qI
YmRtXvNK+Qmtvd3TdUiE1Bc68D/jz9HFJB74MpC61EEG+VQmzP8bF2P8sXYh8cHNR55ZJjYzz2wn
bb7utKjzPYDDwI8u5M7MciZ41LS0tUrzCTDnnCUCUiVtVCynIQ22mYys3mydfzTWFKZKvhworEJw
nPPxwzGpm/F6FVdBFnv/N2yxbAU9v/pcw+PNPksK14ftkoxA1YhvxyC5GONaXDKGunuKWu9I/M7m
cHzUbomDPeWgWG8TkpYFcICa7jvEbN9HUuacB9xpx4RZ8yagAWqorK7j+CZqKcfgx8tAUKFWvX1a
ogPEHL5RzFWNyl16nwth2zD2ezZexdzGqTjhD0sFDe7v42pd5Z+wXBSgfc7KES2DD5WenO4qEoT5
mTIwtAdk6I5NaXRFvw+dqiDfBrLpNLaY7HLre0G27dWNuBLFPJjDbqdZUBLjdkekNDffge7/9N2p
6ElPxjjtMWFP5CZxVp6gcE4d7YAflrrpYymhw6sbyNPePgI2YrhXBm+1I3s/E/J+PjZTGZGb74Du
TOuEi8/voRwHXP6Sl7YG8E9FBt2t4wxthLDHR1CbrofqmpGviIpp3eQByGulh5r2KtbrODpFEMbp
pnUMg80weJr/R0yEaL1GX2VNzhoeyab86ohVQbq7yCffO5TFimRBxDvZXPOY/LAXRBIgPu6sfEQy
yk/2eSCxCi1Ngn1CRlhhRBipFMtsC3ZloH5Jqm5EuBSzkSnw71xJgewtwnMz2ocVSUTh2NKD1q3D
AKHCXh/Zlla3zUAQ5DrDuDZIRRl0/3GQ8OosNo7/tUB6vQcUm4E/qR62Tc0l9LPJXKqdGTRqDuYM
ExTFFApYVKv8Ve1hTpx8ZMYHaymH/IX6TVKY5mu2Vw8GRgdWLtUOZYtkfdcqwo/bkiarP/WMyzKc
qMv2b3Ii0iX7Xrgwt36tmhvgEn3R4GAUv4t6c5p76GMAYCATWcG06ULY0cgoeaxqw4lQXbMgkb9W
UnlUBHCEG5ncu6nydLFTWsWfTPFHpDyXx7QrlpSGCgrXSD753mjurDBKUzDj6+pfTtNMBR9zklou
/ctF5PcpxCtolK75u9UbMM6piadDyc5zWQ6pDv96He8I7EG178cKNwSQ2vP8TZo/X0LYXY3+HaiF
I4SRm/+xH+RhzFKEDSETCiZuaa2x67fABhgg1cPlbNFa+TizO57E3hsjRat+CvvIm2qIoW7lOoBA
wPbceEvMOy4DEDJRpNfZkA9cCxAcza8aSEqnxI96Lk+17DIVkqUfKzn6OIbjYYP7vrEe5XfoSziu
xSP7I+iPzuMfLcaxK4AfsCbUdO8lOJ8+f8k85QvhaXb1vAzUOY4/7LHC3XliBlbjK5SQ7QDEgTm2
DlF1wfXDf84arzAZdB3FpJnmRqQJa2LO39qYwJsPGt7SFP8kLmqxX9yyaJx2MhDC/Dl+/zECKT0f
dKJzHAxJFdeEY9YUVv2DHkQQcTV5eBI8fpXWiSA5Wm9nrdtDsaHBim8KZ0WHy+BKK4Dz2MdfFbYr
XFxUe3EdUQpwYR3obZogaRQck3NAw2z2aYFrW51dlvHzJmmAb0+poMP6U415ycV2EWzNs3m5Y31k
8VUSDy1BSJJeej90cmMrjVZk+uz+C8699KZ7RpSRj8PaYyosbSUVb8QM6VDfR6R3DxioOuOlIW56
vPkYKXyGkck066akgQCTxfWAtHSl8bQP6cy3sT/wWb9HXq0tTSDUxMLBZzkrK+NusJqZ28BtCTXX
lY1mtc7nkI4WERBT4gpTjbPbGmq0TaPWKBXul2IgZOlfCyhkQSVr13bhOVRPue0ZanmQv/N9g24D
lpmbd4KhELImvzz4FQ1SPI/FGS6xOrFo7V67HI1e2LvMs/J6V+3BEs0UpIWWp/45HXktpqr5XkL9
H076ujZsJHWgSrF7QLAbm6OHY7A5W9FSTw2r19fAetAEMTZZVIDpaPrfAFJXF6q6LmFT6fnm+TQ3
MIvav1puICQicdORJBE6fPPXmHiYjxi7e4u+kkBX+7AtfDsHzYNPpMlfBfJz+74qC2oVtFI4c6ar
Gx6k9f8HoO2Lp6W2LrUMt4WqcK+awykYKHA9Ls6HDkRHvAzyajCN/b5+NT6Q3nNj8mfgAo76P4ma
Gt1n8EEkMBLf/B8soJnbL/ig9RrRrzugpMOCSJjC2B03BN1x+M9SVqk0DjFl8mXFtK2dh2jy6Gjx
GiEYq4gNz5tQjyNIoG1DUuKix5Bgoz3XkwXvD3KB2xnfzo2mOFCCkHMm5A3UuwIN/HlAkI883Fpd
PXQRuQz8Ev4FO0QhABuVbAae7s1+gpgCJKyNgebhxz7mQHVD/LOHjS/OqC/I6A9Z96rGwIaG08fD
z/1C3YegAlGpzWdWRi9N1lAr0Q8WxbfTni8jPAi5nhiyH7ft6M37/NaHcYgudzUriDdVxmgzgUBc
73InPfr1HfBuLtw=
`protect end_protected
