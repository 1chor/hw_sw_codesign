-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
oRQh65u/H9xyCHnrRNMGEkGm0qMlQtkIxVUKTjhvPqTWyWoUV23n5p+N3QTmymvR
eIPVDBXrdy/C2cb5W3LFsEXA8j37QYG8TyKc1+JBrdzXxHXxzYcgr5rEPFh7v9M1
+pdbX67tnAjnzBcQFzL/WuZ4OaB8U3+z7wIuLbPdmOo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 116336)
`protect data_block
90BVbFU06hB7aihp0HJxSXpGtfXcWgSx5dGoahn63jlH2eI4HzrSmYt5jca1QI9P
lOJtZOYvWXxgjyRkGdJcjLTj5zL/4A71FI8MGpY6hSYwyvQdwiBD43H5HLl1a/0Z
v+RD20QCrrbccWmr+7eYXtoKblbg98ocjaApSml4I4Zzdgj3uBTJJG0UNSS5Qbhj
YAbmO9wdAjmZs7rUWJKQwJVT9HvaK1PMhMsv7BGJMameB1YYlkcHl+fj9QYC6/g1
qKrp3eWe5+0LIW8cS5da7c89keVZWuDFIkLw/5JDytZik/T69o+0P6dSdSwK/+aF
8/wlfqbmoKet1LEcpMKbiRbafByt80vYIO4EG4cMhmLgGR6qToScWhH/stMRxQZF
MXpVRxjagRbcPrSzgI0kY+YtfWQPoqabQpeT2EqqgaUOYPVI44r5UwbSAIeveOgn
eeLaRZRPLT8/iaG98LGysLoaNsbJJsPpVKaAGjRswSL8JvZAeGY7l//V3Os0O+Qj
PBp4+xTioe59h0qIeOGlnnLtWZZ9JrLWOjZvWEC63eLwZyiocfgMXQBnIS8d0qPJ
4QlurSihiudyb7Es9UEQoR/veBWp1lNKEXbZ7wcumwqzY6e+rrH00cXsVr6jM7IA
Qf7Jh1iAZcoe5jnNTeRdCBNXyi0AlMrQSfnccUDX0JJTLLZm8gEQt4iDQ5brFWdM
Fj5LIxK19UY+2Oh9scQ046upUiqEqvoXpdJTRf06kJ4qVxe26VGembrFPFudnQHd
AKrOi9oEUTq6oBSA+dvHYXg0Jm/VdXounqBbxmLy23NsjuOkRtAeNLJ59G74Auvj
jduh8Euk5cpNFkvi0tkSjo1lN45RMIDQduFSUmyoIZXo35TdpAiysEYgFGARZ0G3
7m3JZJPM6m+vqZShyBAw9V9BaKjLFgkyU9GPV1kNlEYUQuKWsK/8nlvIX6MNPs0/
bhd/D52uoE4udDqL/ZAn9Sr5v+BC/eKFheeAOnz7xt7X7YOLJ2YKmiXh2nujSqvj
XIzKU9P96UwvenDLwWKtB9//9iAsStkO8xddtg5OJMgApsN7UkzdR/TkYra/pCiG
4I1HALCxdZv8s0LpJqYHEAC0TD97t8RD0Cv7qBi0DgyhOJrYPuMpDp7xNLmBwztg
FLBvMNsG+XEuHjsvmAens7vrPeh9/Kpp+3zyu3qAk3iW2m6E+GE59nz/G4PNSSRZ
mmykG/3kBOztnTSUW23YuTQu3xK06DBDTAqESfNx/IkrYX5TmIVGaLxXtb9cJE0s
AdQqKmCH1RnweoN+/yRp11diMoeDAtOAQIB2RnagT07nqAkQBYTqPGCVehga4V5e
8angI7edC1FuvsE81FwRrnFEoHbV7yIBdzGrXH5Zt+cm1XjL1QqPKckLS2EfMH/F
TBt+nKYdG0cf4rZGsbDZdykP3kdcTxOvKotNEzjQ2+PR8xCATCrLeDgW7QB5OVQI
H2bAmQYnDo2bcIIS89ZM1vHZqx0otXpgmfvJ26lcsWuLswmWlhEp2cG8llz5QmwR
OyFyrgH2EhiunIJMReqU6qKQyShKCB74b+7UOgM8cusc0Ms9MMxW+o1MH/B22d9I
5AixIAHWCIMi3qWseN2TO3VrabYECIXqFTIC9szAaW3ehvRSmMqzANjpa9fDbqGi
DvrW5qSY7IMHlW+t6zDu1bWDs63KzMo+BJNcxaLkGcd1PjN2NZrwN5ZfyOY2D3bK
Qxru15h7UwYUoLfeR4DMbkKjb5ARQqtaFQ0zOcSUclT2za9uO+ZoOz28q6Fu8IKx
ahy9OfqhzXPkYrxCz3pCh4LqgDPF7H+BjGXbs65yk+xAmXD/MswCyWERrDCRB1hp
PVfOyTMvLPVQXoMV7YnMh0nZ6W2ldmsi+/d+TzGcGUvRuoJ4HHfqjPzjGiG6OuEm
mMnz7aIRK8vrlIqmLwgYXljN9WH2XmsrPuJqed6qCTOKx1CxONKxu2MHg1RLzYkI
HBollQ66PpLVZycvfHJ9I0K/y9ncNrc1hADkBZ/HV28HgLu4d/qN7YRTzkegxWCf
WUr1J4eW8XJTeeqW36yyQ25cjUS049xJyvvh7oiZGHI3vjapPGk4zxXBBTeR46NM
q+FU5xicldvsgB/Axa4Ggfd4DMPEDG2irtAI9sVrgo5eezFSnPpmOHTPmm5w6Lcb
Kfu34S3dK9nJPhq38U1vwEpi0v0QMRYKYFisO4defS5CDY99kwtZKvyIKc1QqDEL
XYUedNebQDR1FoEEJoQ16fWhGhNEiXxc9AcyaAM5M6F/tMTF0qWADagr2u6TdiFZ
k/D7BUHV5LDALfoIwSKuYEO4wtuljltKyN9lj1krQFQQns+cL9QjN8YU7eC/YnQR
NDKCoWdu6fIPIrZmFl3C0dSfv45S8nLFbJlI1mA2Vr2OGpU0DIfcCQOtxcWiRxsh
WLuO013Hrr42hLarpIoTkrzfnLzR3GDFrULBJxsuifkDW8X4RkIZi5Y5jqq3uxYW
d8HVdIfnRoQEuDJbJN6XT0+vnPHDT2Qji0iwWfEJh1YLCFvTJvkGVl03WMbcUqbS
Np+VzVXDqWRVn4jTAaXEKt0Zzfab43tkYBBVSvMTBJfzxoN8Qqkaybop1Z1iDEXW
LWhf+N/sTpa/R9jpbb3lqG4A58ITeYekcPva2IA4JH4NRdgkFaF5rjuZA6q0065a
h35572od6iia81GQHsnOjnjI+OQYw36ZxG4+6JIezrBizCbaXEdGlpmvFHyVUAeV
oohrjEy88YWhaaAa0FGN44905svaR/9Wv/80KtXdzRFKBzPVADReSFQywuSAgVU1
8PiK6RgBftuYELjw0OdMmcxsET/p+Uamffa1tF7xgBktOTLvevejR5D893mZZyzU
bMDFyjTnCkTXeHC550w9gqr7KSAW8W+HRlBw6k/BgImmWk0zkEKB76M7tNUOf4yO
Km7NIHI6H/e9FTFo1A6E8fYdzO5ccUl72I82rpnY08V+MIvZ9sQbYGDUorv4lhOV
V4BDBzeVszswSdO5TCNz886xHw4XipRJlst+yfIWYdbl72vZ8TptKB5ZK3ya++ex
eQ3esFNNZZe+Mi3aw0nvIAAPwwr/Hz4XyQWjDm0J03dDRU6gD/QcvPIpYmoSJ9nH
+sJKD8kfVZQkd3j7N8HGV1ACjWdVMR7YtPRLt+Jtm3NVxE6dWQFaQw83E/k4XLdU
LGFpUcwVIJQy4MfgBkf36/pJYPopnXx7POydXgN1RooDSOVfacEefPyX6qcmwvll
hOIK+kPxZ8S6ktNme//kr2BouCm0ol3ewOxkxIuZGu0J0n079BbaTMDCGsTZZEKd
Pu821lCCNX5qcq7OEOHDYGhPLdLF+uAzU7G5xVp182CRm+NejWVXIcZ4kWwW8uYK
UjoXSsJZjOf9A8s+0SPm3LsaG2KEUec1ocBJLbeTBDYaEUXzPXVMVHr33vR62/Er
feOWcq8cc3rwZpCL9/fb8iJxz/UF2fJ9cZX/oTBMFYMKYkUxbqcvMzzezVWBeecs
PDkhJjKkRdYf1azCG4ZDWDiq3atfjJvhh6ZjgJHrRXDfRyBvWky9GiW4h1XoCyTq
fto/B5YsLsGe+WFWj0S4fLTqRNSHRsv3DjqEuIvS0mNSGxgMXpGgbfNU4TqAufgw
lyYrbfTcPZvpyJz/irwGRSxQhzflSlhumEmEuLq489U9GBL1uzFWg+ObVm6NYrN5
BGdsy8VFksb6PuQbmGrWpYPc24WdylZUH8YgslgPgFgYezUx83i3k0zXjYCVOBVR
umD+hENvrG8jBhxIPr4FfbAHGXycGsAeRzuMI+5qE/GeY2Xjd67rFXIG3B93m2c6
fKArJkmSt6hNzAWCDsoybbykqLn2lgxd90PSmYh5aX8X/DmVRwMyjgl2crstmojT
/FE7Ik/VLgDpLluAHbrEP3l5edwtGZKDP2XgjQAIk62QKy0kHgFdRxrCimYixynf
3Ni4Ku/QZLHklgtif+om5DP4w8/BxSPuW+5UD7JX0iHEZAFzGQDNUV7cRoCQqPkP
RkWmEdfAJ08SNlMkQVuucRDi/xCaK6Lyj9gKnkIrMrrDFImqqDntbKDjSj/pd81b
v1Y02sj4J+RB9zgJMJJWAJgNbhiCF1u2jIeTnvbf0GdduohB9oH+m3CEb5sPYXXL
C7TlaO5rY/0IpO6J0cI+EWvIv3isQTwClAXUubAMo8iO4ES+vul9oRYw7AJSTNHu
ZlwCkRS8zV40b6pwVtVAwfxnC0E5FwDqrXv2fXXUHJmB6kOrO0UFShW9fhYi7KQZ
DTGqHSAtow6MC/Dgv069Cwn+WOYKplUfe9fOTzygYT7FYUfw1CccJVisQiJCBnfC
091/XLElfxifh+kDZvZ9DWeMy14XMZudd01rKQzjt5nE+36wg5qUhU5BzBBZrdw3
gE+EXLoqU4ebfTwOmvxsabV5vS2ksT4r9Kf/ax5M3cpg1MucsDz96By9yGSb/P2x
sw4bH5BIB+C8l1yKI0o9+GQmb5gLG3M8Z6fgCR+QB9IvdSM6d5EwKBaeOWbb0Mmu
Ioyf1NgFiO/5zti0L+zKeqQWdxQVccqEttKlQ/WZ8ZhmwPSqmCyGLzCZSDruAPo+
IjdK+H5iOUxj1/6O1eajWwqHGH+dc/svDrC6oFyCfhGIkAVklHCfuMTzwPRywzp+
hQl6hM9HzOZecPLg2gD+VcFZmG1JIufV8G7EFwE9/8QmSasUFrqB+b5sauW5uTcn
SwSOwXuF8lTfeKWVQNpZkKCO301EGhcpHhUy3aPINcHI7DnUh/Q4gdxgRxP0hY3R
G0kZUvq9NVRR2DlfU8lUp3Mc25+mRHz1VIXGJ+R1I/AZVGEXRb5WfPcTQBcLOLRU
NKV8V9ZmXF8JF+qxugIYEET4GL31R1qxzsuWztMUVkU+MtytyljDl8hzz57VmL5P
G31ET4wAJK4aPOaqYROyRcgfWgTUOnH8LEfq3arpwfj7bzgbsPNzGOAHnPQV4Ec3
HuVT2xMm25WpJo9BV3lJXEqM2FOXj/opJlN0otKafcECz0nyAWejFZ/Vio/C2nXO
JXNbRHWI+rsk6NpX9nv7YfLUVk0zSTzTdidnJDjcMJOPAivmtEgqoOmym8kEnGtc
uvXtzdrtSwrTwhqHlkjuK1O35TEg8XsrKKT22o1AL4qB9QGijYD9rkmWED6mvKQP
yoSp1l0kDp4l9Ha20Cp/CsfDOssvXsCkvb0f0d+cKa4aafvb6X1HBdvpWwexKUsA
iEZKVVGnkAM5olaUQTlfEdfVFF2M61Fv6caZF2bVjdNu36VRKVUwAeevKbOXYWkg
6EjEZTS7HV/CcWhYE4lhEYt9kk/V/LNUvjgxMjobRODsDIYs9kkzwAhTfFS9CqyP
f3QkDElSr1oQzcerCeF3mwqVQolniKG5F182s19En2tvSWPnZjxDUXC96i90RBRQ
9rC0BX238JA7nc7STKJ02nZhZfsUuNdQyOMcFzY7oIGDs1acYoQEZEEOBfuL8XbT
ZvDqVYQX8sqApWk5ksSEm7Qn9/S6QK8kT0EH+FyjllEVk9b3LLRJBbBKLjMAz6uS
Mvy6sDGwWR6/mQ4JYyaYFF68d6Kup1J5KQjYBg1Yvuo/bfGA3Ogi37uxzou0Su5C
JIwHRtmHk9OqlLCGz8sLrmpJ4X61Ts2+bZEI8F1vIditqYnkRNoi3QytgsBgsuOm
oLZL0Ce8MFUl9QUl23UE4HoQVVtFrltyi4cIJsBWuDGRdEaqEudQIy4tAERnEnu4
5DVsrXvw0BPmtFmDp4fP84R+vUfXid2l7MvKgGGkjcsVugahx5pFKFKuvERKtcz0
MH6k6kWgIwbKo3vhTEOP579xuHLeH2838PzADuCIRAr/kB5TdRAfmk215TeUR/IY
3ykEaD3rXunhy9F1SO8hcy163TLt/APV/FE1DfE/vM+eUGaPurfmyPR07m02tAzn
RP7KtPbTN4uc2w67s989+09YqfNDUE6BCA/JvLiFFSSrCtieQtGsc41TXjzgNoCl
dIaZpBpZhueWxRL/xBuDuyCggNZ75xoTC5BB5MCYC6fW6VgCTNK5MiIT7Mck2g5w
eOOOK0Ai8SjAc5AiCNZ73K325n/2CsAc3Slhj3X+yIZ9lcTh5PDG4NW8j3SijSn8
o17qQFNhfKltuw9f6CQm0Vt77QLoy3ZOkt91wlsLgc8woy7VR7bvpjK/eYLks51y
ya0EYAD+TY9GKfZANF8aPPznnaWjMNvAIeBSgM+S8rt6UJwnDSBCpYyBS4mudWUh
eNfzXdPbHrvra0lSNQRa4gqrm70dGmTiDC4SdQQEnYkXHUJh07+2CZWHEEuf7j1M
oS3eWSoaACDb7NB1mhEPGD1M4OEIuM9hc4ZMwCxKz93q787M+R6LD90c6obxYHTC
B1m34aNPM7OBpwGggyt9SLyNGnC4lpF484snMhGzVVAfyV2njhe92DfV02cAKSdZ
tS4ilTtifPeXaUUGqAsW32ioVz2oYzCtKCVN+Y5J3tad7Sz5+vXAdQGO9WmVgHPL
OWoS+Z3UzfTLLy1taanWRfhsavswih6eK2tMYzhfXMApE8rbjq5t3zwjRR9lThka
TuQ1KNckyQIs9BXFdAaABMwTkObbYkKjEIZkWuiNUNIhWWPXsbmWtFXl7CPzxhAD
zyfx9Bwpi5KV8gUW/2xVccBS9T90Ndhy9jPdAd4xtrCqnoPL0yeQVMzS7Ulxzkuj
l1XQUWekKNUNh8HfPECKNgh8hp1XHmSBqSL4vn+fGW8NDx1Cb3pq1cADCOtp3HRE
mQLe4QC9F4j3ZxKZVd4q8hvC+nmavl9TTM0bMFIZYKXvMdyRt2u6ymnRRzt2y7XU
SRgF5XPMIfvLm0halohxcUn5Ar/S0KVzd28EwcmjvE/tfX1USFTY6GUSHhG9NrIh
9q7o7Bv/e9Av3NhzacqwbmpSLaAlL1YhxGGe/huR0049uGhWtaBKH3RLLasCjkiU
yKpIcQLml6PZ2iPoDM2XPK7vaeUymyXI56hfRTW0L6WjJ8+acpWsTSqTFDSzVniA
bCysUWJNHMB7oQ07MSzS412JgX1LB/8/qK84AX7X+rBpiU7QJy2ES+3mcJVetflN
QxVVfIUnHRyWxDpGhbw3tFUbnwh+thfD4qXI0WySeCOwOu7LLp/yhqBfjw90GoK4
xGqoekzpJdL5iQZ+++WI/vae3IGT4B4rhThvpgaBDTSpqBSPnIuj5XXNQ7DaGlW8
dhfljddt40yVk8O2uhCvm56PfJGudC+ERn7ByUs+jpVQViddQGR6oTe42yfx7GTR
U90j+1WJlfhT71qhOMK7VlR5MWz+bNb3LZxMPUK4jeCdRLJ/29FLdJ1VDM3b0jG1
p8+zfYCzBmN0kPkAjBgkRxEzAU+cNbqY7drCPOTsne+/eCsMl9J6INUFsnTAeaPZ
UVTAwREMMjJIgJwDChFWm8IainJMON/9/VkcIYr1cxR3p7ug8mQOcuUcop8nI8OP
yaKmWS4SSD0/zL55usVjZvrHp8IimjNggAOohX6Vyg70I0RAK52CSSR8hF1uPrhx
ImLRTKQ6fxyYohiL59eJ98w7gb32tifDAA53EAmPkLgrYdbYgYjhFVL/MyHN8aVF
yx7Fb2bRVH0PNFDjqD+yvIvCn9r9b1XoDp6iYk2WOeOf41e1QbVbk4dXbgXA9UBg
YIalmDZ8TQG2zMVPjLqTJJYXlPrwcUb3z+oVUvQzu4LDkrY6pe1TE5QxHcygly6k
/tRUGZamsrH9RwyA6UGn1/owstfW6s0wTRFmmlygXc2WABQPvTdgbdr3p7ZsDuJS
LA0Il61u6wmPTxp8SShvkmz49bXiS3DFKUGjS+Zd3mN0lg4cTOy84IwN49mGKNaa
C1KvYqmpoH2lYlbOK3VEimdxP14MSzeEPmayi39+YkFI14iluwtyeV8dBDLhhFEW
cxG3oUcUjjLG5hT1mq3mpOLulj7lXc5AOdic5OwKuMpqJH8ocsVJn6uceJD0moBE
+v6H2ZgQ0oWpTIIopdJVRPJkraA4uaJfk8DRAB03k6uj7jUXlRvcTytVCZoMccXD
tH97XqfojlnXvf//FjZNWikUJoyaFfqV2mW3mz9WG6BAV5u0Qd8U+McqMdbbZAyT
PrvZ4Z00/SxRRNIHM5JXlKAiHXMFbV34CZFAbN2ooCSlHMk0X+gQ5N3cdw+M1sNm
orygRcO9xXBEBri2h1hwg2LTVUlich2fH+a5AVeHaojuBycm324FpXs6J3Eg1Am5
0/+rsWNkFzAf/soPUq2PYo1/ULWC90+9XD+jvXIIVtJZOsfAIPLV/VAqEGwAkpVl
HtSQFYFdjKdvg9H78jKfKQdsbzswXiS+UIXp2/OT7XsKjsJSeOea3c5W2++Aml3z
Yinr+iAirUemIdpT8NFyXr09Cs3Opq4T2fa54wPQbAzTMa8kE2vwCT5DzWZvfVJ/
mVniTSxin8Snk9TwIiKVcAKQ7340nkzK4eN2MH4m7WNh/Votnbs7uuGaUGZspw7l
muIugag4xLJECenJ5lCULN0W8NZUckOGPz6p0tTngGu8mpSaiQ2roL1IhsqyD0uh
MOzJhLYe+B1eWo/cGxA+Kq996ce61rWRv9Iy3QXo0/RqB4/amiWNF0cWLkdl22+N
T0ICIKL6u7idN1Un6mjC9U6lK7qsntr8LgYs3geFC45p2OVM2DuKAo6VKufde+nK
c2x0VvEvk4f0qT9vzDUZJrirb7j1b99kwo/JK4uv9WHzgrwOfvqUxJWNSqfr6tUQ
8BC05BtxHDoPTGaByz9tzTCGbeaHTCQEe2QZOekYYUg5XCOKpOtBhde4br/OZwAz
1H085OngdmqfKEt3unhzdwq5ag9DMiyG60Elr077hllHnQypwkOWboe1H/0ubD3A
+/ZHT4q6qESG/qEq2PznJ7tYWi2aotAJ0nHULvuuZ/QYz4yeYpKKUdWspSw4TDF2
SoRzueGs/dQ29ujpdspEoB81Ixs8aa42m7H00zaXNJGb37yBTEWLNxeVnJsKH/8M
UYFIoLYT0+Ai7Boe8XozRHsqMoZhANMDdsC3SaR6iSYhSYV9P8V0xl0c+h7qSRTS
hBTuaC6j6Mmd2msVf4EsXn6OjanRl8oLUqftjxEgelvCOjHneHzpPeTtWCfiGiJv
71M1iFDtI2T7rRhjMNBDSPGov655Bunx4cZJUSeqtyNK7/BmdgD8chBNz0cXrAnO
WPPS9+9C02Ltl1RF4Y/MaGfmXSN0YL/ErB0q/v8usPUtb+W+SdWsCaXwJWnw7sOF
Q3Vgbfc2rRqOtzGITcsFnyEr7rZvjBpa8R+IaG8wmqGnIbjj1TP7QFS69vBDHKNJ
ldv14JHsZYvSoHFJWGLL3uz3qRuRmocrr7mPfAAZZwtxzSqruztbDq5cmh+leCgn
tWZ+bFTBTxla7ibRgTWDExJDtTaPBS45NmXqDWTfblkUOQskIavqiJe1Bb+FOqOA
ribXpPjp3imiaVXzkBpC+10gxAD2MYKbQT0gYaMlyVCltN1dipu6/zoi/tBjWrSe
Fn/vKSPNFViucuXk5EnnGOP1mT2UsLT4nRXVl8fxdyr6VT0vEZD/1UHRWpxm2M4e
xnMaK9x/qJfMVfbsqY7h2bzy7EqnUUz5/l/jwy9KdKw+BCUAd7uYTERHYlLMp7fN
5M39wbVPUEI2Uor9GTE4ryXcCbFXY6ZfOkmERwkY5ijc6qjzer1hPgV7TR/2S7AM
ZN53gLvAttgQQeaUjmQw9WqIRfX9/kYSyPmYaevYHvA1IHT+Xiz6+Ow0w2oeM7aY
lni+fwvTUWp3OkEKri9QCDMLJ+tyx7n1upbnGXbiBmuGITzQLYjl7vyinT8A8UpF
IKYUJ1tK9QtTlgx9FuTHbed+g3yD1cky0OGqY4iHUzPYMQitaCC109+ruJN6il1n
XwZN+SK9ggoP6DnNTunDX6h8ULoMsaTDSeIjlIhHZbmGxxfm4YiESInt/XrslBmw
XWk1WAWAxlWfJpTy0+7TX6JNy1Psl6g1g58OCVWkyGTzxEZWbd/EvcMj8QAk32Gk
jwSDeWTsjnks4ptnGrwSdnG8k+MD73+KQednsv8Nj/JG6dLO+BUzTiR7FDoW6bd2
w+2bhcmkefySOHpDYu8x+A3ANQsNHzUc6iG++9jiWJ4Qmoask+/zr6tTU1Vqkb6b
po88Z2cY4oTDVVfEcDz9L4pwTX7GlN/FcEraorsLaKNwkxwlsnEhfSUBK+jMAuFx
GWBS4E6WfPNdQxAjPR4/ijRI9kxVd3h71+0cl8kZl5BjWHphRQgf9kZ0xvVCXspP
ZTgJdZWhnsdNjGC1G39E/37exZyxuJhgie6nQubislUC+bj2skY2RKhfZIpLKJhX
SZAZuD2irImcLj+ox9i87vDJ5E2kvhSQK7qxmWj4qyG/wuzhzfFWDBH9438zwmaN
RpNZwQE3bI8MrWKD088kIKsCoXHOQrpvILXnhec546c0KmzsiWztDv1VnK0DXtBm
m1kEbop/nqy5uMa6TKKkIbnmH9UG02DQrqWWkMic1p/sf3KSvWFu2FUBk+FCvaNF
bcrRofWuapI5X/ZgIQPk76YZYmNQkdJSX6eqGdz+bFCW7l6Bg/RO3H0TeF75vco/
wBAgR39V3lv69TsosYNHcNWDz2Vc5ULOkV+v3P3xthRoErdfP/TVcTZhPuP3EyHw
4byZuIXQ+yX3oxi3buRg9SlJb1ly4b6ioozsjKI75VT2P+xI+lz2C4Pf8rwUZose
DZ0TD2QchYqZwDHsF4VpoZXjKmKDPIxMP8G4oOtc0trWIiQLBlTpRcfWpAiVyM5A
w66NHCMMG4Rvxd3Us1K/mYxlHEuuJdeWAr7Zyok1DxcC2ydD4Ngf8QrvxspgsfCB
ZBL6ejwBTx2HVn9FFAwck3l0dVh6WaihHv7QL0DqbxgFehAebIkambgGOBZGF34i
3rDPKq0n5A8SRWE/fWv5WUtYm/0NpFVyhSP8glewfxNp+NAX93N+nd/31oB3C6xN
Tf2mh23jYmQAW96nuK17xGxhAzmdzSz3IRIjbQGA9VzjV95hJ3rEsg67osjljshz
d7JR6VxZF6Sd6CCjGBN41fRLde6XH2v1O0fL8wyOxeh7lOtWTmhIOnuYO5hO4Krg
VSfNjMv1lBvGInsG6U3LV4bCmY8GhcYEDMGMzfdHQO7HD58Iko3i5jsM6p8n5lAl
tqJ7y23ihL5ifpr81tbfw081kJ66fZ6RPfcrLs678iXkjjBl7BJ0iCra0R90lC0L
YYGyxKHk7uk77ejok/qLIdDxDiSMbRkB6qO2iU7FRFhkfCgNtJBg7wf2J4sK8XTK
x26zgp2RPH9JhoVfnYQVFvHmHcN4E++dsitDrxdro2oM0WkjqWNu1lN3RXCActfv
JQmMv1HKxW4sSVzHI89P9f71Nk+BpKiVJysn8aFv0oHeTWmRrli1l8ToVpDPwqsu
fL5jOm4zOJGNREVjy/64QJoMhlVYJYdBUVL0E+GKDx6p5MDoNIMFiYJLDCmgs+BV
ESs8MfyxKb7YRpae4Zl/XecNnF4gyVG8uMro+KxBniXXrBxHcpJ1pzK3V1xFgOlj
siW6aq43O+9pinsTyZW/nJqB8HH+7mGY5DdNiNi+u1DTGwcQNzvG6Te/2ZTCw5GQ
0QKdlYQinFKaKfE8eZbL1nuMzPIVbZbnRKx8oCeCDWL5EiGfmb1tT9AGKTlJl4s8
68JHZe8WLPgzBDGgWFQWRYqCzxKDQT/3LyDnjnw40LKQunTmYQiJTVBTC4urcL/L
lLENIv5xFcYzjhmv0N0upBVgQ6nZi7nd8lMJk4YOBXJIL3Q9QmAHpEb3kaHw/335
HEzFglH18UlSRvOpezXj5hpj7wk03B/McvJLRvrYFPEnVvKznSqYVAwcbgUeERCr
JwO3yN+G/hrGZCtwUKYwsw/TgEiJnrUZ4+dIni+vTZe4ysA1QkRH/lYtjcCWFmy+
mVnZE5FiYFuRBmiu0D34bvEv0XNx5eFH0DM+y9DiPri5Kor/x6tfYNoEehQIHGMV
mdDvATk5gbbJuWLcg1yMhtVWn11DHaHSn9Eh+7K31wbFAh7oMJFsasuyxU/yZFEy
Uo+bZ7iAAv418yZCn4kNV2CtlaMczhW0gaq0+FGadQF1KrA12l1E6w2w4hzPswgk
9h4jeVFZ1z1A2nZ9aa8okPkSSLlrfaCYkfcjpY0fNZh/YaJ4w4YewXLiLoIzOyhc
ffjkVGCIciGYfHdGIsbpR6uovuKuni3zfV2clZ/CAHf7mgB3KcbyGP+5Z/RF7cMe
D5gPNVAgGEaB0Wfu4QgYsSJnBsYeXhCvMQevFkhwqkgiOD1mjurNIyKTU7Ur7EXv
H0WUoAgYkks1GdBX9eSyB/C+TwvO20V/e2XoHEaJ8Mf3OBkSqK8BWobJ55EuOy9H
SpzxYPL3BohlaLGkrP4jKxhR44uiKH6vVdj0TivQPatpTCo3QTQ0NAXHbAAxBx+v
LkaOFJW19mTygh3feNVJ9hEhmEJYIdbEI7GToFz2LxQOPbnP7gm6z4tcCqNmguBH
mtoDH1eGrACZbgPK9qWy2/PzLwMQEiBRa3xnw+HKiQvLhRwZg/4cQaDb5fZiJ/zC
MtUEPCowKAkfjNfofaIP3HEtKXfePE4dbtjgDfVQGheld/3C7TCftA5rz5a8QIJG
MLBRgWxlSNOfNw68vtKFSL7tHBk+a4Lw/gAgH3ErlvZkikc9y4FPDqin7A078/fC
Vp9LN4km4j4R72Q6XAWEjKxZwLpHUlT43g24mhcv6chP4v5sTJFYCA/pn+X19Wei
9SHjdFoh0lre4OXqV8KuG3FI2TdGGwHf2bM0kg6ss7q6QmF+r1N/LE+a160bhkBs
RA3FCaNiEQocAjJhdUSj3OX2VzWYyBI7BQGMV8oEZOA+EroLemVwopAmK+yNMYkK
p84zi6XzfilylMNOs0L3uLmYamZtVOFKFDhNe7k8j0/utvMDdX+X1MflVXypj5pj
4MEBoljfL37HvuFRr8UA6CwEnc9EcLEgqSWy+Xt2nUzlR6dh874K1hcM0BIkmING
lH7zTkainHaOL5sdQ8kt+uMaiF9DpT+kD/wugl03+WL8Tz7sAoHTEd1mdpya5sNz
8PlcZqGgGb11PAjdLFam75SXQJMtfm+AiO2cpMuPS5wIDmd78Iyj5uzj6bwtyuhK
FDt1b6yC9PFMEQz8gzxmZgcvHLWUvvXdDClUIhL93pZsS6H/WdG/6btlR/GLDwBC
ISJhd6F5YWFDIBgyY4r2e7Aq3k4Ox5BYGti9SgtHPm8Xuzf1u1hU+M99fM/GSvXl
/n4OLrJKyyZ5Mj0zit/oQbiinf9TjYC41zidduwpQ2etuTK6dsg2E63MRNGGrXYn
u+tNZUfj9HwvZCCjUbPN+jPHtY8bIU+SSSmKnNY5l5ENtb5FhUvmFgC8GGbP8Rgq
UrLu6SQ/foSbT+5k7RWVA8C3ihZzEJMhEJ4bhKh3iykEj0ZXic/qnB9dBS1Xpkn5
xEv9s3sfa8Mcd4rRgcd9n2QL30G6JsCQg26munb7jiurxWPalzJtQfmAC/BKypUZ
yTPbAYYm5AiHEYz6HAgf/c+aqJ8y3vvrxBbebKSiX2HY8maiB7bo5YjMhS8N9lzr
WcMj1Ip8qj4zrACq5lmc7EyG2oMrRLeHGtVb9gdCcoY8+ufk6eRGi+nDhxu4aCPx
+f6hnunnsGxDzmdcRfJHRLIB8pCYIyFbN+iN4AtfylG0XWjTY7PcUocZU08OKMCt
GqPGQrj4ZdCoqPRlvt4dzwZH28odz1pcrV1oTwboTx2XQbKbfTuPjrO6xZ1vsTt/
A/M84aP+TnGcBHUhj1WRXUos4tC2hje0KGUv9jgSdOAn0vYqEad6+1+q4+/M4kKJ
TI2Xxsbu+z021+SH/enDKC6e74jkof7JiQw/Cs+aWdmZJ4rxdZTci2NY3icAQYOA
nwUKHx5CDlUTvbizuwt4lX0A0s15UtIJWBM42Z5dTn/fIWQIfQjIA1vuGswt1vH4
fUlk17HRu9bXyTNt9we2KvCYvYxvPQSa2ffo0l5kBv6jCXvs8QIkIvb5OrfC/Cry
GRBoFsUUFKEIc8cKdyZ38IAbMklqESHkcpRaHy5vZ4flsJZ7aAHwM032dpluxN3L
ypx3T+DXHiLtAs9Pgb99SdKnayb62kZ5ALKYqAwcvyxXVgyD/fo64oYSJ6uHR7UC
ad6czELjXX/D0DOxsd2thC1ykarUVVq3jJebPHIeE1Mmg6et34jucl40WQjX1URG
0+2hJBmkdYhFE8Gv7OWAnWclfM88QkPjatoaZJ4jjR9JyaAUsJopzRlYoJT2UYON
YQ6T2jxqnKkj8USRjxvgOhWro0NNFGu1u3ITiG6uuEfTRFEnjbfuMrf7w9wbfi++
91fkMtRbR8kByLemlLjcN083rQEUGgNkxa+X58C1NLsbr2FNqRl4eTdKvZIy2hH/
JD2RutknCchZLEd2XGIAwCZd2gfJDOkRyHA8FcfpyycSq1ZcRPSwNxorXpDqscjO
IqyCNUiUnMq50dNJvnhiLnc0NlFSDM4RE5KMZ1efmYJU6QKc0+TGXPp4CBgyIy/v
cTwjNrLPOLA07RU24i0XymcqC7n58YOYCYscciuMd7ytOYlkXvBoa8cZPHWfjxbC
XEn82ZFqSXe8+gEG5zOzfG4ke2YP4ILrDIvMWqpZ+mdHyRu1SekK/LfYKdE1lp8y
ERaWrQEw1COZg1lv2Do6omjMNszbfzMHs/bU+LFgpUkG5/BzG0NeRWEQE9Cpaek2
bL5nWxt0MvC7YhP960AlMtvVy+pNhI/7QyBTotbhy03m6rnLDsI/C5aXoO3CmMSn
AIVQ2RfcG2yxXUlAJ5O1aJRr5+z70JTjdHiiKb+8bPwZm1hGtvQmFfxwlN4b+Aq3
Yvr9p7KrNrUsTinNJBrNibFHnnG3RlzbtJVIOymCdKozQFqbS8iy8ehcRD7zpKo5
nIsGy5rIe5BttQbsmRlZDvhwoae7nGe1TwU3M+X2J4aot9QqfflKVpfgNW3+9Ugv
qdudi1JuedC1qPuGHOKZ8t9Sb9IO7pk6jBJRc9SrD26titUsja/3WL9gRR2cu23T
jYvqHhgceYm97HZ4AEPdQjkinBpTXzND0VdNQKm5VmWF0glLmIphdH9AjX0Snsts
ifeaXmv7Rjr+xrASkn//UTGErC1nxkBTpH1CkxcPvVOL5GUk06D7PXDfHdiDaHMr
YPqXsH/fbxalO6NhoCNHiD8xyBeatbSbWEdtWbqIXLmiSvQ6bGv7TlFGnWuhOb6P
23k1Q04D0WZaEM3YzemxEOjLjQBbyZE1rIu72NxyzhI5+D/1R6Zrm9ZOgDGtVvrL
abbzaiM2Z39jCdSP3Y3Jd/SU57Tvtyz2HMyOyZ8ay1JSfEyWTjXAizC++OZB+WZq
kpRuyKC3k0Hl/CLbjtO0uhkYfhSFwH1Hu7SJx9cJQKmZo1YlT2ZGzy12IL/UOlLp
zR+ynfOuroKpiZ1Ln0JYxb+c39EVFs6nDxoqfnpaRhBIi1OaU0FC3S3E8/63Iyar
GEB4HEN2Vq0nzHh95ZBRH89/5eoEE4Y3oBiGN9VkhnWS3IaDRv9GtHvHXicDvOcp
ICzbNfL06ZzKF1g+K5INZMvaqVCoT21Ls5WTubeTjpl8Yz5lZ7p9XFF/2UsSlZew
emSl9+suhzjCyyvpa932Wlxs01DDcuvGkiL0haBZ+xOxgUPdDTimDIQptuc1CeZZ
JTrudBdP5pJG+nDSM+of9hVmNciIAfskwlagCHOI/m8LXzzuomU1PEZ0rJ1eVd7V
WnPHmgGjJKj3tFiQxu4cZG87I0uu2A3SgCARdPPMJGUUGPYOBS9XP248Ci/Llvb/
TfzYaSvzTNJc4SS2NbTJWv/0rU2pXd2YIvH4bpYqpurCaF1+1xTqN9AHvFxfCfkH
yjZlLl7JmAAQrH0vhssuUcqqoVssOcn0a2X+d1iYaExdIU8VJHgxWW3x4VfZZZb4
hsxezIV3xAORztOXQwfiaTd/9bmEbsVXe4d5sWGzT9PQWNUUdQUYMKeSG9wY0OOt
HvxtaWp9tQvKKrWWgIBzgB71o0aJhLDsSlyAd/WLiAi1O/s/g6y/Dzlt0FDupxIP
Re1v0M2+Pdnd85bUoJ0uodyNzvMQrDAV42xRgkkIYfJxqhKOO9yBuxfUYyoCKU/T
zDh9zGauvp/83TxMNduZ8y7dVN2YjME/L0gzKML3IqOFCPLNNWkiQeRmAPBq9ybD
o2V8Kifdvy1DI5dk03UYstc8ibI0nmqc80d4neJp7qmucu6XhsYad1Tk0zQ/w3tE
/h6TFcS7FSKiPx+YrjQWyRZ9t3MSivs4apSIMOBje8AJpjgG5QjRK+0rVdPNsbso
GTPK0Xz1NtcEi5JdpQpiebKxPqO+J6cgJSl8MdIZDjVKtmFFN51xNLrkZWzgjJIB
y81P9twlyV+QKdg1ncM7fUuhrB+jH5uTOaxpQHzB3V4WdBPY2LPNmusyoaX2g5Ko
zPxTXv6Mc8QKnw0dUyPl5W0ymelbKwSzpPyNgGL0hsISSdOgXvIN8n3Ce7q26Km0
HZdFHgKZ64ARuQ25wtM6HKLJ0/pmcFGmWZwa3VP4X4L4xogLtMlE6teUKs7S1L1p
jqH9Spf2suTrObidDxZmhfh8GNlXBXkC9M+VqYVuUS4TRrAzd4zdTW5ajjZFjqvo
NSiwlP7oASHnnDT+GlZH5g7AC8DHHgacVj9RDw3+Ng09RpU6Unjfd1c3ypiWl/4O
HVO1q/qGdVGWCs40p3hRBCaTU/H8R2LRFNdYlrmTrzmRBYRVgfM7EU9KUDNgfs9/
dwYw+dSOgMiiT5hdBqhtyoZL8TzDRbI7YjE5wmpdIl4KrgneIRAOxxXN37fltzlk
Mh/ZNQyWFzBTKvZ+gHcM+ZaIW0kCd2wGkkDWdgkx3rJ6I7qer4ug/aW4zMYQOkLG
32Bdvd5K9KRn/9+rtI1SKC3AZjfEpvEdrsjN0lgpT/9qQovFJyDzwXtIgKZJNiAd
++EMIjmVLnzLIlXbLbrWwu5GgGsq13zDOUN76AsxXvsC8/jC5QeclRiX+Xs5LQJ5
FsxfDxbDzKserq7/K2N/YH+hL/uk4TEpuf5Fo6wpDML1Zg3vuUMXIddFALHZ/6n0
v8BHAl/fYwIoAIa0uA4yezAlVKCFQsxiwzuOZLguitivYA/w07vY7SoxSgR69KtP
6bzbMeatNKEsni+pCUIO1auTnexK9RKsjOMgKrVZBGAMqr+dkTc17PN6Ffm26FGc
m0NVVaJxaO2RLSdkgLfte2necgYkTVPZqwin6HITUzNr1S7KcLEUTUysdOljO5AT
5IXEHPwMGxTYo1/QdhyVhdJxoX3Fsdahle756jPSXfd3UR7OaybBV+KGqaHaajDS
3NjevQ0YJlORuWDmTDl7oV97goVWP017bIPdQuqIHg8Ek7t0oTVPsmvZYlYCHrM2
iAHTFgygfEFJv1W7hKVJaYaTZ0/HUYxKEmqe2AP6xH0iK2eOT4ocEscLbZFzuSTv
6yV86WkmCDyioYsUMHWt9tg2bMFsCQBPnFxcod49okUGa1vyizxONA3NjJYVG5Dp
X1wn7XrHIFYRbUH2IFCmzF6FcoZE4sodmcTzEzjrIqltahg+sX4z0hbs0z4byWhL
XgYFuLUgtZ26pP2H45iqdRCAu3l5vO9wQyfqerBo4EDC1KcKa3OgVap3u66Ak0tY
I7SKMtp35u7jd0T+xahXGzJFbTmHeSFJFYw3uDfmqXB7U1Ds9XWOWnD+K752rTeV
XmtdhXTTDBBIzbxjqI49zc6HNlQhzKGeo9ue2GkCrmUWl5iSzWJ579xVT40c9zQU
dMJ4XA6ysbReaoXdbaMarKBmFnBsdmL2eJkPKdZk5k9Q05xoJh9Yli6HyCNVJLL8
4/Iw1cRB7JKhIYOiR2MT1jiDWpHzbqQy+bAKNFaL7YdV2ZD6BgIH5tIhRZjiHsP5
PuzjVVlC8pdliAKpiA3javrSPniGyNggikWXWzsbwlq3VBhYW8vGXonjCs+4WyyX
o6GUIzIBAw8J5hoKs7VKRWCgSs5XG+LBjWiOU+YcGP7+GO0FM3cfnx2DVjlzBpBH
G3OIYycUX827oZ0AokNF1KH+tyuxDEpB51Vt24+25djLOQhakBkwM/iOZedV1lnq
1aywYYfcNULVySW/roLD4VA86qf7bmtHUDRv9FbLGh3m/vZXemjj72HfKLFZZ2qn
oGV1gXNChnxJ9Qmc34l/5IyDg6niWqWjtJ6zH9n1fiHzjFQNc3iZNkkqKVgO+fF0
YqXSG/wDTnFSzHY/xOtJDqQ2VD03DbkW8QaP1AvARklicK3rx1EfBBjmcaq4cg5J
ei2B2y5Dsu09qGb3JexAyQoR6J9P97gsFdbnIwf3LlQjuXFnp3LS/eT0MeAFeox8
MBJ/Y667SHq2jh5y44PLtbmPgG7Y39M6YF4t8e2Go2lFxzMkQSWv33AqaYwa+wLX
dekevJrVePhTqXOOSNb2OZeFzSZmHxbVHeCNo0hRgG1tc4WCiC6zM8qPEGxl63aV
y2n9Z12oh5VH2AlTBn0qfohhn21DT5YPNPAi4+fumDCGRG3FpIjwqynM0vWedGVT
wrbCvd56VP+v8JHmd77Ro6depDJPVkoWSQH7Tvc3WY5NdwhLZ3RGVt0aEyLUCZ/k
fsGLeYE3bHoFjob4O0rglA1KVSncFQ42nAIdg56lLtnaBkD0YmoVNxhD7bSQQ0lg
Z13IH2ZU0dOylDJiA4x6Beay2Ep2Vubsw1uCNEedEROizzj2pBOxcz+GKd+smj/N
ZdetOpa42V7mIeDxvl2cmNQd5I1DQnaoa4/zbOUamLh8U8/gMkaflfcI1+loxkSM
dIExR9YdD2lvGdNZQwcJ1Sm0VZABJ90NBxUXUYVlujCot2yj4zFM6+jZ7RYnfQ9X
OYUUUitPbD95KHptQmb7XmmLyFzKbdxDqxeqmvf1684y83v3wGtqnk1z8VLJb2E1
W4xRtGbeMqCIdBv0WJX06paIhuNtvFdD6fdev8ZYy1oREogITlJYyLp8nghddGSO
YVRNn3aXF9lfyXW8oQN/AhSqGxnNdHmGyI19uJkvx3LvmsWNuYKra8vxlZk3EbfV
DQASd0J2mXOTuOTuqA0c35/qFpYfVMkz4diZQbJFIVDcTjn7+0q6UbLkta3dCZTQ
UraLymdZ6h1lYdCaqmTRfL1SQcha86HY/4+tvnfAM7Q7Tp6xSyLNwXfvWV1cwtJJ
xikvOG1UNZ3e6vK3Si12ioLd6Grr42AC1I+VSwih+QnvVrxad7GSY2Q4Qj+xErsj
hCjEsQoeaa3yz1AabRB0PjForZ8pvhxHWh5XuCsqot6z54aZAVgIeiRuVrR0xtbu
rMLVV7S3xclQNKlz6Ap/rbMiBX/bzWigBKibJiwyBm1XwedYws+u9J8w4CtHjc2s
DuAqkVtrlguhV1cuL6QTmSc4R0OvLM2zovZ8BvI09i6UwNe/Yn01C7j5tAYz6S9R
ZmLOFDyuiT2NbQgUS8pFV26Yq4YxVM2/tM6KuJlTLj03Zd2qttYJSEmsHTU68t+p
mFf+Dm/dJmgXPaj6znxfqqWnkta149QpfPZI9XIHqoeCBE/5ILTnXb0UJlR47dOz
o8Sx/Bue5YTZNEcbP8IEyiBOZgmM3TxSf+qoZz0fVq9o1hrm73AVnbK91CAMQfAe
6lsgOGjmmgZbWen1DehPbPartYyA3DP1lwkVmZl9CTrPRBH1tsd3gz3G0tXIk7g2
mZ0SzLUOwwFVvLIF0efShoyxyiqAK5sWXzQYrFf/r9deyiE+ghZDMcLscd0WGNLN
y2KYKyVOxzFk1Kw+9b/s4cRHZxdqd/6dqs0x8BbG8up43SPY8Q6MAkThgD+Knv20
Q9ToJ8unahJjvTGtOdmAViuvbALkgNwgtWMlMjAchNTX/JuuEXG/eLoRstxX6nlZ
w/gS/x9fnoo+E3GfOhkUpocKNJ6d9I2Qbns1kTjpn5OkEgRQl8nm4QE8xS1jBYub
Tco11bA6drt7pVNXnFsC8wVc0tQMK9H/9iO5DUUt1UdeIDhmkuDBkkcjpK+RJpAW
U4KMi2eZp1xO+0mFpKb0n03zduYmr+sO44neKPQOMp19nGz8h8/NiPtk55nppqMa
rdm9X/EgTzILLPB2gFk3bCvfGRVhR4rjepICABYO+VBGxMpHhzcIDnoRjIZvuqyn
zfBHYMyUEMDbcGJsOrucT8GbjO1pUpEcIEdGduIH+Mr482OS6Tz7TJZWwEqjCvR7
T5GUxdWxKYsIuRUUf/CLTODBWjZi2iyF+FuiVnad67deSz5ydvUdntK6QWfSNlxk
b25BksQGNRCJvA/XqKd2wUortfwiUhy5mxWodDVqV+CcLowi8JYJp3VSgpiNBHKA
3thPHQdmK5jI+Y+o2lmIcHGPOM6DBUWiAkuINzBW5q3AKKbsVpI0FBovTOjl031Z
NgiVxoTtBe1AYj+x0WfX6Tp484O/DA1yND5zFXjZ1MFxH6HmQyodKB89JQUlwFpW
sjszZ82XL5V44jneTLTNqOKkA65UKqqHhIVNxdSf21ReSVe8lXW8Dy9uzakPrZkj
vscCrLV7fgMWd9/WxoBbLp2jfYlWXeCfG2UmneWJvkEK+sMda+nIG6ejA1SxP4ls
tVvfWkSi3CEK2mcnapUNwIEZ1U+hU+8ef6KvzDS4Cia0taeUvP1zIILeTZ92j0YR
dCRQDIXFTNnv8ylJaSMWOXNHLs6mXicHu1QT2bG80cucNBQavOqoOg/FbSA0Deri
1L3OS0VltIJ2hC6z0NiEzUrxKa7uoqYzLFs7iVPQkv8vaXLBu95q+h0nK8PnL5IJ
z9pNJhH6MsqpEi19WD/QEFkGngHy1JE+EF8vxEfTMZM5sq9yc8fSv8l3uoEXRCu8
1pEnHmPYBA6IiqNvFqdJFmb25WjgE6HPVc6AqvxsCdv8x8Y7QU2mq+F/kX332cFt
BJpRAMttg+jqUUgRBpI/SD5usPP973B5/vWxF6xuyELBJpc1lMj8pqhOawiAKERJ
9mlWu8yJLW+qFChQqdCxDtZJeNx9P0n7CL7EGv3aKgpVdF85PBT+aonF6H7AoIPK
T0toMji8N9mXaEFvtbESfrxbiLFRC+OTxZYxg68RceJOgByTYr8E2iXCKmKttaG6
dKVNGkh799Y50Eoo8ZWnIuoaXpcLmsl+DupPtk1XLlVH121kevIYYWTZVag2nSub
fORLUQjoJMukTb0gAMMubfMqBvU52Y76UkeVmWG4V+h1AX7KXFemEAR7xzURU9nD
2SaILwYC54dMpG/OGhtL+8d+juxoo5McFBDpeaCuWs+pnyyzSLP2W2bcDAyFaIwM
3El+r+KLkIQvN0TyHtyBIHOImdI0uGQEL7A/0uRKGCbdB1+Rl7k70mbntQv5ccAa
edisqn+l6W1XGgZtuYlMRppT8/26VFuCQdLRyIqYzgrtjjQANGlTsrHlfbC8baRO
dHBQbd6C7azWhRCPpobsNmYUhThgzcb2Uygm0l+SbMFEf+XZRvpKbv4kkswNEsob
DIzmz/ll+Aq1/9ISikhHmTgdvs/lzbOT+pi7OeerJDpUz1yhL75uwsCSLZVuqeTi
1Rij23kguth5CZPIfIdXrKT8hj7lCP1WAK4zxtrZxMv0w+eHEPiJo075ZvZJVGh8
RHFOFD8AEQwmFZAut92Aji0ZwPzwq97W21Wvfs5lqF/znwejOvmDWVrlruRW6X44
chgAjea1ALZRXRUfiLEACo9Sx3m43LKIhYp32RG356io5A7RBaGXdt66aOHx4+8x
xXD9ljXfLassjqdYbK64Ifl3iplTLDBLiNHzHl8NDUF3XoaiL06Sv/G9pRCaeFwA
qhtE4gXmh/jpycm2tgS42WtG/cA7cE58az/Z5c1dZB0sbIMbY60L/4MjqF5PirKY
rdKcDE2M7QM3auGwJZVezelT4++bEAhMizN0M04H7QZZDl9oGqWRwgaGzMvv0Hr6
I4B1QVsoda9eJlNP0KfPcigtVG61be3TUjdoTif/CPu7q2Ag4xzCNrZDN0lkTZ/H
tUvsxICb3YIpxsFh7RLGOPOg8m6Ysb2Iq2uKIOXkN7rr1aXJ7no6zs8sei4NQpFV
Dxj7bSlurZQcqjkXjHAohlpngbQMI2JlPOOLIoxaIrFs7wIP84wWrz8CWRSv7xqc
lxRxup9hn2fEW2k50k4DqXjDZcb+ezj2p2jgP+lmzONKWcEkBXJzSSz5821Qqcer
9oJPCFrH9TkwbcQ8MOmKzD2URR9sbHBum5eUyqGJDJaLHp9/hiPoY/Jkoro3nK7k
dglQl/4Ij0HfkwzRfBiv7YRzDeXNET/Zj9L9o/j9iYbI8+9x+rmV1WXF4th4E9sX
SyniEURtpFrBsdvH5KRHMoRmWsesUvsVOWacWuoIvf9d6O5LV9OwnQ9ZcM8iyVHm
9fZnUVIZXwbK+EnhMKyLUDsCSumcM+GeUlup+on23TPCNG72RUYMMtnHTDnkK/8h
8r4Yd+Moo7j8I7qe9cjK7HQs/AFI+sQIwVY1TJuePoaQM8H+C/5l3q7qiBdyTuox
lpvPGLJuT9j/R7dxIeskAnDwmD2p0SalVSA4Eq2tM+B+jDdnkQbRA7SIOeRiTCYa
M8dbue/1U9kOeMXBC5wxDcvMqb4VNHvY3JhrbnIegyMTJLTclzZBsBm6TePIsG3a
iLi7LWpDWhsMYITUDWi5qfR3Z4db/52riattnyPWpo/f7DAa+eiCn8cc02lRorJA
/OVwEX1/RMAUX8wsKjvoKPWRs1Uzsk5yBvamFaa+gxb2gf4NAolKEqcaJABqYJQD
knGXk1MqHY9Cvv8eb7k7PduRJmuI/D3awplmnQEhGa7AIGG7GbYGFAlVpYRyKY9r
/Rq8Omso657E+QMvEf0/IAxfyqksryKMvKR39YsThKOLrejP0r6+UD74c3AssIse
Ruz8sIk6eqeiR5hcuXtcD4V/OHsL32ybH9greK7IE9WZUQLoYZV0VGlL7BI5m3hw
5c1/rIaluH8PXOEKQ6KRcIjwC6GQ+Z+MGoHWlAuYzWCPBlntwFO23elzBtTjM69G
hiQSuzFfW2a6QdWYjKVhYJkYV9+eJPrljuD7/jDDVVGo4E2BupcFEbFA6glgr+lO
rKhOgXmuvbxz0FntD112Afm9GX4LvpJpNc3MnoWmKjzR36aGbjHTvi7TJNTttyEV
rVklvZSn4VqYQhM6zOCGUTHko04VxJd5UzkaoXumajL4XL0hJqgTBHOQZtuzsoqC
esIv3XX5gLyf6dB/DNFxjTZfctoWnJNSt/SCs1vl15oIYdDOI1Vp89Mt5QA7NtyX
HJekcNnY0CWEhH6skurz8dBCd0FGfvJvxZnH6fbsUEbnUBlMAegXGvv5AQOWBe5B
akbYNW72VxCaBgl0MfW61Q4jpigPGU9KIJiNDCDuuw6Qq76/hKSeUYLO7hesPrpc
SNIpg8BLDgqgXBj3LqK/j+1+hjBCtoSCS3amPBUJkPIKaHd2+JECXlnLX86UCgTG
oEpDxjOx3ruTbpy733f38WAS2rcDgQ9YfLlB8YwJsjTShkT8frZyS4/ceKuX5cn5
KOgG98qlaZO3RYZ953i+e1ld1FdgFDfGOQTf3htHDHrqc2G1SLQg/gEov1jwKzXN
nU/0OKyOM/HlLG7K0Q5dYz2o2H1GNl71nOLxkyYoHBXu/iUz1w3PmHLwPrPH1K4Z
Pl6SoFOqK+P0rcWhMGbWTHq3dn71AdabVlZ8BrF/qKtokHHqslO62vNsPPnNdDfS
etvAa/4ctI4P5/QROopJSTlnUEuraKtaLWDvTzLpuyZ3uL50s8oLveHZnJzo/vvC
Qi3nS5mYOVzi8ZKMqZrFU8Fb1LbbsqKobyuuiSRy3ifv6/80MOtk93u+PPl5HRV2
+lVZPM7AwoqnlA7nphYKMlIr9Z3nZQL/fwSr4C4pesXBRN3+GdUKEbESZB1z0EiE
FXs426jf35LnebAXGBaihaSxUc3bZV0YyOtT6+iM5Kw8UDAbvWNSHUmK6OhozbxA
PyHFlguiAHIWABRsnjJ5MVr7wW7KSIj90U+NFU2dLFH12MO8K8+leqIUCZM3j88m
WrbzYUGm0fvsBiyPpZvI0hEV0984GA9VQjQi7BIoQ4MTpV1VXlT4ehWXv1X8WiO6
rpXKYZoyYlCx7d4qdkAK1rgDKCQonA0Pu1l637YwaO1d0b7XmSjA9SJAOrKynJFL
ccvMpoNSbMsWp4bmbPurobo0SQHgUhv0TnoN8yUBE/CMNcX2fn6IZW6XOn9R79L5
8BCEQjWMs/vhyjOfeXFaZ1cmgxcnK3I+jcaDyfqjN9IEK3Vs76L8WOKLJbg2olk+
Bg1N3WIm8oFR2SR09ATymyZH6Frl2rOhHqvf9dz1v7TdRtLHw7Ws31YHIvWoOVxw
Yw54DeKF+1yx7+l7cpc8ENZqskop2O5OegzY+9E+ZENcY+6dMJAf/dm+5Ki/fucx
mVk53oPo7iE03aiXFsBADXB5sNVU0E/pUG7iVR6cKG70wWId/b5VcGpQ983qh/NI
/IMpkXmBhBgvZGYHH7cIfUvpz3X2GMpwcmYoEGuOcyXVwll7IsQGDDE1yHuthjrD
86L86ByGp9BI3IKvQI7aYhBGGrRp3dbcfYQDNn5FKhqwxgWk/JKqJDc1/gGoh4ds
5C8giN17NHOUxg/UPgSINsXA3Bzuk51KDxCSi2CPC/xPV3Xf5ql+LbW4m+puFv98
j2H9Na3VZZMFZNUsuTrqKIVSwK3Twr/ooXVBOZDTTbMyjEMjLa+DrMn4y1tYUdlW
bv+6sj+zQ3ErR2DF4iniTy1FN84N7tG7jii/emDX6OiE1LNHh7A4BDkzCRYmhong
wHe02qQGFWyFiPAzISmF4MSF6hRgbuN/NmhyMSHfEMXNvI3ukkS3+FVpUwVVWAdf
lg22afibDfHjF38/56tSvHvrecYQzF74mh5/xZF508fKfUI3ecwUpprktaVbhEdg
icOewNoZtrIetRAMEPdvrjQVgSbfPdcptKUWPoRpFufOA6Aq8z+wl6qvQ7qurJlH
By4LH1jW9kJuaKEreDm2W6tfo9g0EjPjHT+L3fatRpBKnuWlFsrKA0rIKaekudg6
oHQVrqLGzQJNfR7rJxzvJ4hHHd91q9lGh6k1oqrGxILEdHwhET6ajiSSbGAzhPGB
vQ9cr93EEIOAqw65g8A+A3ZwR0MsvLIgno/O5EcSwoJsujY9gnwsKrVX6EuX4LBf
+gWATKcGrkFWpXwX/aQw3NSK4p0AafJOJsOGaHz/rz6LFZVuol8ecPpdw0QzdEKv
b45UW5WAv62nBeCwJSNd43ZyXP/OI7nIpRftvhvuH9Bhv+s8letZ8lnl2gsmtelM
bmFnXH7VXA1jQIuyck8SfAApg8NAycNcN7z/xrjw/OwWsNNRavag9YkafPEskYt4
mAAemsPISQ4dfMMBQ2JFTMocrSRUyFWgR2TZhv968TK8HaCfLHC0TWxsiFxfUSuQ
R7VpGjqNS01px0pW+5H5/qeHbqHGqUIZR8dwcrUUPH1hfsKu9SVTB2t0QTBzknf2
vEyFSz++PDu3B4WKL1xkZRKTX1sWwJGdQY52NPORiQsLjBw3AUCb6FZLx88WWZjf
ccGmgzLZi5z3zChFdliWHXckMOVhhYGcdfl98HaXTBxbGq6fpDoQJo0R6zFv6jhq
zjvk4kl6Fc3xhOmmemX/Rjtb9s5SgKMQnC9nPxjJ1rh42It60D9zVshV67gJ8lXS
TYZfjg0r3P/c7VbiGASygUgigOwuzpQExcIoRpqODaWyz+P3Bgg7u+zztoWrhNPj
rAPfu7muXT1wf9MXIAeI2a4G8DvNUWFMsMN+MxXiWmWRDXPllbFs/NIx9BHBHhNb
nzlIOQ4OaIxB/M7tIfHflpqr/yFBBamSgwc0Lc0ply+yuMgvJTsTHVY5gfNHOL6I
mut1/8mLMbnBjpU1e5ccomxtBXa1Y+Z7ay/QPHj0syvy4MJK0BAtULen1EsTcwEB
YriS7MhEsdqcgsA4oWObJTqRS5rpPf1JAA0XEG/fqxjs1lnjSsoY770ojWp6ojr1
0c3/k4NNQ0+1y4S7PWcu+oBdAXotT5vwiI0ShPCUal106THXMH5rBSeeo/dlYjN/
as4sh+F9QJQDZ6y24ObNBd1Hc97iNAce5oysIZrf7i27WOTmnOF3hDwLH2KmscJM
zSml8LeZtvnAmpDkX7ayR3atm1Ydz8lRFQJmYUxlwB0JqY9gKZT5+H9QJLPfWwd1
H8s1lIE3i3vXmUEOCX1J8Ce8yWytjImqfPslhIAQQrl0VDN418+c1/M3+P6lISMm
vdqEIm6K9cVcuxbjTCvmD3V2PliN4AOukgaoJIPKWmxDjT7rRLeIdALfjXAqgyh+
oM8FdwYF5cauwoTnHHwTvmnR9llFblMrxthJYRg4uRWtX0gs6vJPay5p2jR7Lz46
OGIV1w4ATqigXzEvyyF958k4asrwTsxaMFbyrLITkRikq1MR77zseYxq4NazjgHj
GBFQsTvWzCgZXYLhyD/elnjDvDB9TiqLtbMQJsMhYAoZjvhI5qHsXkTP/2WjgIKJ
NxcSmfNnKqA8k6//RFod8s8S/j4LlIQBA4kxOuptJNaDboD8nCazWXxssmyyDVhD
J/kBOHtJE0KyKku1J4kBo4FdmB/iW/sWt/vKwb7esBS1TrAwxeSZPGLAbw1pw+Ix
4wqaw1xkQi1I4ZekFeG2P2t+GXN77ZDKqxwk+3i96ypBw7TrRcDIki6a5IbVR8/V
fXzt3QVHSRKN0AJbJGYDHNJycShJUdsNxXGHQ08hatqn6HkaTTdgdb/RH7GBlpPa
b0kHYhxYPKbee4LGxGfgOYjvqANKZcvSkqxbMZ85U7fwR0SIm2tVCpJp6ScRXm2M
/rdbYCbtQocWTAqpC/cx9qOazptAubh2e3ZjHcR3X91st8rc95ZfCTNSueXyNsYS
9+aOSn4JaFX/MEiyc6U/qyvpsYDGFd3r3VdgknwFLfaqiHoyqzas7dwJ7n9RSazm
BM95unhrcUIPrCW4TZKYAA4lwRIoxRLDeez07SU3ACwAKjsDtAs/4NqSg/vzzdRo
pgUQLPOeO4tigQ6Evil1XHAsYqSw52HV6QN1eC87d8cj8s8vZ1re+YzIuysQJeCx
s5NZJETaahYAqsIOHA8HeRedYSnf52bNK1AgOGHhtaYP6x8wiiV0YmjVDlASSZ5a
rOgJ+4MzM7UN7RLyLA1KRlbIIUk0KsLzKlrYJgq5KrAteY9jQtjZXZY0pcf6wrpU
t7EZTo7UaLXN4PrmX3F0zoBgNeEORV32KY0aXcFvRrp7KFtSkUuUhbCzHmi+alhP
CQk5IjLcBtLBUhn5nOTxWYq/0jvBRfoP/HVfiO2BtddckuKARrnkK0v2h1RrQPsd
ZLOvK/2XNt5u5CT/Ot3DveH5SLEjzpxGryO5sXxkuZCTAkynpvl1hbaiz58N2xJF
8LXaaL5ea8OeCmp4IYkokQDGgeo6JsMwEm7JjFGgJQDSp8A9QC9jGcQuRWXHsjd0
QWCrRoljI65uvLA3/JkZhB6WzWSVX4NA+hTyn+5i3DbNDiuCUAqCJ6WRz23bTDpT
kQBgfl7Kz8l4CicBCLyJ6a+G/iBvlFpg1rC8QNtf3JxrOu1DdoDfZYDxE5NMvD/8
gXe+LXd+X65MYKtQtxGGT9NGWJYVTZe2HXdk8LQAb9+LiQZfBs8HG3bBmfdmQlUg
5jTvbYyBSuhnwbvgKcoZ1aSbZyn8ZTrAoL4jkN0sVe66dje7xXwsPHgfz6d5ZZST
lLnU0Gh8DDugQ++ZDQQsfQsxK97bIHxCrm5B6ZXqLQEgdDueqtxhViZHGgWtwu1h
Poqf5+yTA59jWaHbcvCYJPCAUrwN9ZFGlOinf2RlU7XdZekRap2ZAwtQoWaMiIJN
aWDB5sCUmL929LrgF4TySiRywRJFQTKTjrWhGwXe6cz0HutJz0Kgzhekq0fkn1iJ
oIQUAt74Uw2FdbEyip5xbR3E0WjmE6bz9vLRAjjJvFhPzlhnn7HaBLIYEgubRFoF
XC0AxX11Mzw/ycTGQOoYP25KsIB7fHh0SM/R85NMWUxpYtL3nGSheii1Qz6dofw0
YqkrUEPiNg8bg2TiXZIqAFvrw3qWk+vOBEQkt7WX5YqO8hC6U5RAeuZs6sgAB21v
i/xweKj53TLjr8PFgHrAQcs4twb2vv9I5yPz6kUwkWA6w9BtE0M2EMs5vImo+myB
pRtJJ1+4d53U7nMFTmfrRBjB/Q+QDhSD/FHbZbUvw89Z44wsL+lOy38ksptQAt6a
c8kdHC6rhBvCFGLHjC8rUZe8b3au3xKB34mxwZBc536xmXHZi7ZyKlBSGApvtgS8
JH6GdFiW/d7s+9Mrt8z3jKanSH0egFsyoce6W6O8ukhF6y04DK2X2bpO7KsjxGdW
9Ie04Gpfoo2fo2L6ZXtC6t4E/HERlN+mhbK3joYJlSGkQVBrZ6wb/+CDcLA2zY/6
HDYe/gBszAiNaosajWg7uhFV/2xUuly2+i3OA6hkLfSuTf/kIMCkkw+23w+IhX88
r0h04R+/bdfg3+AmAQOwHxo+zJZMd+JfwRlGVN82jls7ug7YR/W8o5+g6Sgdg47m
3B40WDgGgQhpiS8OHGjU0x/Re3ylK0KbeNF8lA1j18mdqsS2hFlzGOf8N1MFmlvs
M0CIXperBtTyQ+/9rU0PiO1D+3ALmEcgoH/n07EBSoYGB2CwOWDVCbJzbW78G32l
7Yz6hgqZxetXYQNQpV6RkPRWNJEgIOyD3WxM7ctx2KYOmEkMppuFUqoHNWP73SHd
/qM7fonYaAWbmn38E5JPmF3Hw+2cmuthBY1FFOGA6mRkn3l8GJfdUmgaBkJbEF1D
Dd2KYg94FQmjTJkdL2Xhhb4mkpTzxxxhaAfsp9bsR4FFSbv7NP3tonrhiN3ZusId
FPnMR2opOll1nYS8+RfHI/NkDHMFAQBU/HskjzRm9hfvwI1qEmDzYweG91X7QeZR
YBXSN0MO0H3dcowKtw7CXDXxwUvzzWtkoyNgOn3wsXNixriDJ/M045cfS6iaOrid
ovYNIGMWVcaR4uxhnuQlKZuBYVUEf3S+jK813BrMgiQi68vRXWBvP4CODySk9mkE
Mk4o5yHQ+fzvsEmqn4/eyG5CwwWb4cQfO8BdKLCyD7vxQX/L6YPcX596LdT5ISzs
hkQ80zaYjAnaMZBWAvSgla6q2atz4dR885PXTKw+dDWBZyJPLyIzr8C5LjkQUWHM
jU0nxIETPKeQzpMh6k+DcxwlUAJXOmpzJhHsPYVQswPR7IyI2V9m2U4MOF/Lgnto
09gxqWTQq5idVUb/v/pdqy3p77Ltgj4KvoER7bZDLn2crf10P18eIesj1p1oXqlX
cW/1maZ5nCIyrDph4RFcPkq/Y7FINAg7q92MLrFNzRfVA46vS8Z1ePLGErO6xCh1
YKIGGriABVUGHLu3XnjXql3qb78FaX3slpkznrIe3xe8TYt0lQksuL5qk7DJ9kdI
7IKjueanbRoVLnsyKqEGyTUYCt3a87N9hbqpi12m5MzgQkzwycaDr8d8r6KcuJVZ
v1R8CG92RUQkJ1VjjJIsBBnprNZkCBtj9rhaHJQLgWQOxV7YQalr9NiRvuOYxUYZ
WHBf9mkhdtczPJwGSK8ty9VqcfoWsGNzXPafdOXaBigw8M5bZDR40/9KkdhhRWbN
39XiNkMoyh9q5bDL0ktKhNacjbBnJ5gqkOMdkle4S4WNDM2zG1e7eTxzZmIEQ7WL
Bd88UMM3VLHxMqyV1G+E2AHUqLOb+bxH/eltHvXcl83jJJ1tgUkVwgM0a0jesnwL
37UmIvdZspYaKwXjD2i/dILldI8ERO15IQNPzGI6wWPVWxZNifZrCSpBHj+qj71Z
TERz6tPO2A7tnkxqXQpJXnpcRZEqJfus8YwqiKUltHFHrJvQ6/rX/dSfXt5QQTY1
ipkJBz00sFkcvw21Ay6BY6F1KQY1AHm226ELQlfPcFrSnS84mzmuTSQTgZMGE2Fc
mIdQrq79erayNQbDf1mjuso9WX3LTXq8kIJ5SBU6PNDvvvHWimjLhMBzuORhBsNX
LROpXmOuuSsRi6GuinMiTeYBHTXokImFt7QL6Fc28pf/zImJrtvb1brWZqX3op/3
ktJH2ViC686LvMtwJCqh/9wfkJzHcHuNLMX0oIt+GDHVm3ym3O5SUNho8p1PACdm
ZPBkNm6z+NPeE4k47GM+tb3GdGSBGGCIJ7iaHywqepx9qyWPRJBKJgFsXk25QtQF
PqidlSE491GJE95nSuA+X9GiU0WuNffUWJie1lSxs2TuQp8HzR4ujEdbIfTgvXgi
smaj8Un7LziSawSAI9ThAkQbLD0vUatyCY35lhh7X40jnqbpNFKmjmGWxvJrU27G
oEHQ5G+ESRG/JIRtWjyqYL9ti4LJB31BNa7Wrlh4LeDvI78f3ZKDX+heDtxXq8te
qihaybkxEQhafUNv0eptXm/nDnaGRu/OtMWtG8jhsEOl3gXu9HQq/oFBE97xH5Ev
ceDpTill/PKEmbqoRwGaXYF+wQT0lt/X9JQtsGvgcnWp+xinmZ6zJ2PurNDjhkB7
oWQlQrY6vBydNw4LUOQslFugWFLc/zotIbaZz2CM/wsp0NBYBm+Xfq5Z/+8PhsD6
t/IWi7LldT4WKDMHaQKPqWK73/kvEPZgs7xLOhVc9axyImqCUEm1cAq2dcisHyBS
kcz078ege76T2NQolUFyjMWu8hRKJhDiEoqlFSGpc7CZmvAMrsCFrdrzt4F22BLk
f7rKUmGOZi+HrfG4AFliMI9yXypoBx+9WZfoBXllWptAfs8wjj1arytQB2eEK8F3
tJLpmYMSzmRYZO/8nzCu1tF7M3+gNg//H6SZqzEdgHidYv9oZiNiLxUKEhXYsVZn
cjOdQ7HMcXmwEaUzWrf4DG5SxqJPG/wcbKVR4rvtrWuHcIwkvzHqWxbZQOABOqXn
Ow8eaAxuRUBO5qvDzRN1ausBx1XvXgwVeNKqudLHTMhWIUUYGbMBbjbhYFDimb1e
Ja+yetIErOmzwR2E7bqGcBWXi6amPMyvG15RCYyF11dRTBT5kJq6cw/JfeblXE15
/AATmxyl6PyWvkJwzSCELZFjPoSpVUM+n51folPe5pWV9QHgiO/QVooFNHBEuZfj
NNsAf8rAzwG7TIi/DEYA1bFROPZQ0ugJHS4aGu2XRm22/RQBtIi1p4omjNVvG1zQ
MFn8sRLiHMJUpiXG6ydKIB6UikuWtrPUMPULnoJCFYBvoW6wQsBNJY9sH4AWXbu5
WDs3s4uOxJ2Qv0rE2GCysgXlNjAaCB0dnDf+e/SBJ3UwmNIe+tzWMQv11LsDNMup
bkqF5cy7P8GhZtlCMvyfDiKpO4j95mCLiNz5ZhvAl54S7hM1XWMuJNrKT6h+3KY4
zw9t/h/25FrhYsoXjD+M6Q/vXoOqR8/8/XpYEkAyxNxJbHOGsX/D251L9fSB34d0
w4ezKAHYkdiuaR0iGBNRup7BDZ56H1/sfJK0MkzZxqh7wv0oX8POdQZDdi0M0TZw
y+EaqSaFym8RrhEPX6gedSPVjWJAi5QEHL3sCbTpgVuXnGBS1OStPGiVagRZVAbV
oGsxv16YTXsLjQTLGNVEOsiowmdo35CkrPd3CXa4g2tYhAkWR46OMmg6QlWnYAZQ
d0P+WQVBib/vOGTvVuk4LFPILw2bdNwRpIm0GGshCU+9cxoDcWv6JHc9bFqapUmo
leEwz4XaiUEPiPKI29Ag1h8ro/sLVFVI1PblTa1nqRLBhooxgMqnulTbDXVk5oSx
ahS11SrsVe2pHjl+ybxQum+0yp/DDY6BJnVxtF52pkdNBELfUHSxLsJoC8UhSbJz
yctCLRsGBdxkDUY0CtHRAd5nZzYa30iP1E8VpOTSrhfZyIVLVO7QIhlDTTZw+k0A
t24alnciFLp7CvWe6zXBBZDImTVT3x5PknEhsP7gS0Yv5lgTuPCP8PUaJdU6HVS+
RdTbJPRgZWapD0z44JnlrR7ZoOq9WJJuhNHDWcEDJB9BAG8k8UPtbwDF5jwzWfMA
krbtI8P0x0XCM24l4WAWsYRN5JZWvPAQ6e9IuOFZAwdWU5khVOElldtTRqmYKwCH
Dlw8hSyRplOmFHKrdhy4W2BjcfGwRRxZCbW5Ojhwm0T4Y2ycrLERXuI7eynDTf2M
Nrv1YvWS/9UtKW2BmX4mmjTLL6bKrr57LXJYdL3xRm/0/HIDQw7SRw0ZORRouZcl
avDaN0/9R8ghd0m95WYYyL6+epvlChns9eS8/DxfkKz7kIfVwbayW5uhRajtlhJm
M7aqv/BU00FlNAbyH2HVrNq0D2QRY65Sw4OJuf2QkQBt2vJnPZqE+CGpMe1RGCT2
rHGoAVCv4BKHAyVNqZU5PE355W84iptOnuFyVwEum551Rpw21U8C/rZq6EfGX/Zl
ascNHS+2PxkLSxTSHD0hM7EAxRQTYlKgWyOluz+1eXD9WUC6OY673wtWdNtk6sjx
4NZxYn3RmHZWnAcEpa28CNp5jb3FUdkk5EeLIibzih4DMEQ9qBf8C16V8GKmzCn6
TwbGAFTvL6qeU+sA2oSAnpmda/oDiBvo7174gwJ76iVFU93yhXkFGnwYQzzwRaJo
cmJuBYyLlQyc6xu3xR6pZCLAbU1o7MT5L9OwhIi8toXD8YPVpU2jZa8Xof085xbC
0zz4bVs0qEtzfwQ7WaFpLFKJ1q2SHze4mQnC8h7XelU8fG5UuD5jaPqasQXaV4qQ
fe6HjGqrgRE3OP1mci8/9CeM0o9c3loMWvBU5E6ySCKlHve2zNjcm29XX5tvGAiW
dVyHMqhb75GXnjulnqxUKJ7B8fVvqZsU1rNW0e41lGNj5Zyjc61qFmR5SOUQ4qzj
A/pDB5MugZUiWfYAKCaPxrlCUXJa8RSQmI1LQ1hLQfTHXCmpFwjd76lO2p8oXWCN
VpM9u1PxHSLyDqKZJcFPoa1U1UnBsmzlC9zmS7AtRvrXF8JbaTjc5y1fK/Yt0tuv
QLHL4nVOyKPuYy098Zm0GuITWg2zPngRiRUtXMXig/FvvbNoMSzPoIiYX4qsmdvO
fIJQc2SeTwxWliiVsKLOtRf87+YIc0fJ9m84ws3ughltiVfzFTkEhY7EbT6DHBmR
CVc3u10yjGP5YXu7Bdo2Qfb2cmaxfiwG4uFV2hWIz4geSIUoyfshxfbiBdBLlAg2
8jGYh+5qv1dbZ5tIRXXCLrnx8Po/PnwN11m2J0pPJErYV/meUpmBdPtv6Z2fI3CP
Tmf7AK5RxfHE8MMU2078N4jAAB8dBXgXf/kKvZjscy60vOrdIOVTiIz+kujR8f/4
tfISbFbTDEAaRll5PeadRA+7KuEbffVr4Y6Q6AqvW3CBF2kgAS7Lpp4tj2J4fdwK
va/lKL+hBGugATe7CajZNTUvahlok6CDjm8DHA3qhIIMoQqUWGLvR0G3JU6rb6Gn
4fATPAB02VI5F1wthx0mCVGv9r46GDzvmGqQwQGT1lrEB8/Wt052YNXjDL3VoJ1v
+qUIFdbpJd6EsB7OCh6M7rnBjs+fu6I7H0T16Tb4EDlauO4ZUe1VjJ+WROUpcqQy
ral+nxrwIa0yehfkZiF+K9RcXGR1f8LsKv1A8U/xxRhXGsPeO1ZQS8F8+tq28EHp
QnozZVX/FZMUNfhBj/GQuSSajKpnn1jE1P1TB2ytKS57R3JmbfiJUDUwUbM/PCRc
Lmx+0vNk7xdoXjmOowh5T1FyZSPlK+is0HUo0/hwwhmA+v05c9cjnP0vIdlqyAHb
pniqVrb8jbjCS2KAbYm7W0lR9QR/6KIpWCxXMdotZAvPKmqpJEHDL1dA37ZZMBvO
1oeYBax/iW3T8dyxdFpDEaELx1T4xHjDF4sXsTOaP/LAOMXb+p9TC23+N9Snc17v
m7Gk9sEX3WdfteMobazuZ+JpB5ojdTQL5CliVOD3KHpTgLbufWmtGDgalZn49c0/
/vBJCMl4nwUnIQ3iumC5IDp6kmzckduyzKZQVjiDh2Ndvbng9ufLAgMTj9+aPVse
UBO9zNsGG4avka98XUg0bQk/jy9ZjlLiP9jdZF3cUaaEQgbXYbCz/+ECQpzMb2ST
X8fXVI/UFc2We3mkweKTAtiAUOlgZn0eNW64GomY1dKqOmP5u7CSLOxZscS+FwVo
4EhpNBjKhSum13KQCN2kK4Swu9D64tEvqNrfhVZcU50Qjq7NKbRViopvN3lj7xMh
3BaixSWyWK2dccFOOQyp31GdoP6goiemNjOPPDooIOb0s62WOgXR0LBQld2DXF2m
mg2I/N9F1v5aal7/DzkMtmDE/9y4AJQZ1SmZnAcwcgdjhvblo3T0fobVBa5bmXRQ
MKWDXzg3d9obBJznYWnc4R1xqd4r4lOdAUokhDXOxt3QMIopYjlqS+4ST4klOKhs
ezBOxCU2v051B8ZFUani2honbkfTaM2be2CejcpSwsysBSYIofuQKQlyGPBQ9ZFw
xGtb9cEduyDapk+ciuRwfbPjHXyc6HYh9Ul4ZaxTyEwaYxWMm04hGWBqe9JoW/r8
Y7YjImGZNkutJoyt9GE5i6vaep4Pz2w0B6usrccl22UKEcoa5t9VWSn24Yu7HTT5
X5HfthacwUgeW/e8t8njXlJL4rg5FW79/ZEVSAbT4OU5PWODqVA+mlI5KHarrm6G
/4JfCYI4aJ7vAAJwSClQ1xu1IHTgAaVZSyY3X8pUY3F+XLjmNRpTol8qzmxCzYJZ
/YgDBDv4GFmD0Z2UuxBYMgpVpieosiigzHZ/7qiMqZdqaupc57xVEcIi/bO0BK3z
8YyfqFZU3wIE68sq3LsVvpSS9koxmIhTmxLqXn4TZqNnHRVa+QBP+tGkG7hFEyff
n+jG5sakjYIrvfphZZdmTdcHgDdB3EdCsgR6DZ8W2ctuasKykuQCVcjSGAhW2JTE
N7FdUyF9yAj4As9ZQlGY1PxtC7hUtwZFdE88m+MbBsXcQw7zC+JymVsRPbzmfKAV
9M7j0t6kFJ+W3UinQy9MDKsu9UMD497upmHcMWYqvsOLk90qWPqIpj+4KIznFJp8
dZMccFHj6llTzf3EVcjt8qCRoMJh9PCxmXtrbjIBlY85gVTd6RzDWd//yRsIzn47
1gehI4FE5v3XKWXS/Lhs0Iu9eMqd3V6dl5WxbnAKId2AlCHRjzal5714gH3GW5cl
0YfUdPb9+7mkW5FFEUUljCjkIulSzTpb8PNDgwIkPf945PaxeN/y14SeBrP5LYZw
Rj4HOBIRx3RVhxdNL6oQ4nCuKaDvKJPGF3+rgyScAQ7FGbW/0zwZqHeD3oHggD+E
HD0yvxfIsv30kRq9IcCcRr8RwaHe5xsJ9S/5g4HtRIRJoPiqChaqtCJ1EZ2uAlOS
fMADwR0SKyLBqTeFfUIK8L736sIL2Zh5TKHkF9IDXgnib7tW3k5Euedw0JhN5aWW
V9AUp9DYtHUH3my1a1hah2JQjFrqdzUwP1QpaHQpTl/FLGRWYTzpAXDDg4uwVxA/
e2CKv66Xc3Cqr/7k1R7q2xhFpLTC/BD/JFCLH+QqS/LX7JZmB6aHY8wm1us+LVmb
q1mxxRXVo4Up9Goik1mwz3nUonYQna1uhJ9t4/nfd4WrnYr0sN+h82YgdkGmY9rF
n2wy9b+X7wMHZnWyPLb0YLupSPPKHOR9mPdB5xDv1Qk68gkWXifuVKo9/Y18N/kW
YwySQJbkiaKO5rcmn1skxSHzfeNgaUrw7t9a8RJlNINIupZiXasilOfsRMaGbt9W
AgQ0zikk1oloWXhqYVTVS0WweLi3xlHMrMbAZJ84euk2XYMYFWJVTQCaxSPwF/WO
7dwA+Tgsf1yqitcJazQrNy+Qry9VDmKDkQxV7EF2SKOUOXgeZoCNxshDKOlrU6tc
raRPvpsy4hUjIB4V1QttMcsXGm6josbkWCKRf0c2GipN17x1qZDHfmqX1zFHQLYa
cfB5qiLzGoakezZMVp47DtAVmO5n4usxd46TQs3XDmlhbhU4W9niC6QPCpYzshUv
aDZg9K2AEi74stAIc/n03fQCzGXKC4zQ7y16kVHXtkg6KICYSqL/9X48YFb8vxQn
YvByiYe/yXT6hEa/t5j3b7dCYabijdyND+Ug2d59lmUHsmkD6A/VeWxntivWZ0Wb
BPglQnMNQ9jYqx7arzTgSiwaeLj32jSYL0dtTElIc5wfohM5bhr7SwLhZWWcGkV4
7eRRhW9LwDYpKZrScOi48XDab5Ht2bGGP+kaPgQwgyryLrprLrIK6mjcby2mfPkX
SvxlR0yolrxl0R6zcDw5yEFpSnHoYW8k8ONep47I7aD+KbyGSD7mSMAxbb49vpIT
IKsDa+Hr4AkTYpKJKprGI7pdLvWzDoT9sEpWrKrgpj5prjzABqm51gxR3Wxg2r/3
fizkhLeSFJ9+HbFy5g8tbxH+SHqfc9YQKDqkL8B1KZfA70DW/X/iAzAuOADpfi7K
tDocP7ZBFAth6HXBiDWP61Hcm2/uGTTiaGFdhvzOPnKyXqEDad5V83GKoSW4DYK0
uONgqxp6nwQavonWVuScvACv/IjTqAJZa0nq7JbcS1i452lnlYKi+L1VCD7EHT5u
U5zqTDNPU42GDJXs3Yj2asjLKA7f4rKX5cHoiK+DGxF/daJ7ftuWieY8QLbRjDys
fGAqyFjn1aEXW3dUuFcELs8y8749L6vZeXOG0kbrbaZH4RtH3loNhDXNMqU3Hkpe
Dp8wVDGViT+88thD6g/Ueph98ivb4HoKkQi0ts6E/cznin0Sw6SjYffm+eqsileN
xzr7X0W3JO949U3Z0TAQLaDySL5wdDXGaCMBgZ0AkGoi80Xod88k74mHr0mrhyVT
sPGU8Ipc+5lAGI6Hipup3nEN8LTxCQiLpa8fQVW69j3bsPn1r5KtPoSPYXCdEqGA
D5EBspvhJ21HhdI5GPcGolLOuvbtl+Iwx3M1xIMzaqvY+Ic91mTkXwl5OXupWmAz
zldR5LqHyA9EAeDyIuMbWX/MEOaeHpqo8o1W+wDgPPdSW7G5IehV/70Y7A/chILQ
yAnJ9YvR8SS42ltyYBLZ7mMNq7BiIrjR+G0jbtoMbJwA/W7wdOyDxnTCcSBn05Zs
E0Om01bKa+jecokSZKhWZYX4GLR+8UJw3f8AfmQceH0j2CQ/PpHwKx/WtbNBYevF
RYshsMt/VWYtG3Bsp7Q8r11MpREi52Bxu6o2qGadosZItK/59BvJNsKnP3KKX/n2
MljDYAbffwHTcBiDp93TSgegNyNXmx1nL1gVeZGGbgZcT5pjm9KFtZcPllJ3o5pJ
qAOLVnyQE64ywngEEzKoQWnGYfcbhS+6y5tTF/IYejb2b9PKJNyUumAECBesFkua
dYUFlUizu9mjqJXq7uUt/0DzgX0PhNO/kxLnXWSgjcymm7n/o1bMrSORxkvn5OzG
vXSk5f9SkYoA4afFxbPgpDTKnhB0U9BnHHeiyk5WP6SGFXZTzpRXx8AT3A2/zQo9
YuNlj8yKrvTPTUE3KEI0iKT/9bTUcgf62tutIDvCRewidOGGLdBWnstqBOud+dzz
PsnHenbo1Md5JkRFzKG98taGaFppN7Serqycut01vfLHeox97sOqsY5YRNFrtp9h
hVsR8RNUw1z+skz5HkDWpGGE4RFCDyRBjyZBxv11+DgQPGEFZF4AcHOiRsJ7IDez
ZXdnaMOSm8gnfWejT5ugzzCTrvTgd7W5TP8O86TAkGIvPznfljYAx5QofGYyYo3m
FJnhIlrioY4hAZAZbBqXG/p+SH8ru0Idbyz5NwRxtOrnIydmHr1ad2GBiI7oT4YR
zJso5xf/TJm1G670Ona+T1f10ac16OR7srIovau6Tph5BXaWiQOysY0F8E3G9ZYj
v79WA6pRJNgNVNnHVOokstqVfvIPgkuzaZ4rBPmZEXMWI7y7WA1powCO/sVQaOtp
OXhXikHDxeRXzwzcmSLo3BpTDvhpQcobmNCu1wieNTGxM3qoZmkEP2xkQOYnMSPV
k9aA96NFWl7yc1IMqXkY/XW1ogU2aujRi/3mFo1qR5BW4geqO1MIrfpMTXt6PVoi
4Kgy6St70MVn18klPCocIYJ+115SlX9ki8hRPagBR40OM9G7jgf7zAwX2thmvOe8
a57MdzyvElWRrKTCuuBVELhu1O0f70b5TlwAaim3dwX2vaoqAUn8B7ONWQSNC9Sc
w9tRAPFWQjMFeJxLsx42i3K/5Menij/2YL2tb9M2DINzy52wRVv9T3E5UUfpIAfd
Biagr8vnk9KuBs7xUzcXY/J7jkL8u5R/1ZO96G/kjSkzaMdoIR2rd5z264SyIg1e
HaZMGLCzW5m8TMDMcwypWSakEYrRYlQv//oaB3j9/JPG6VwHbjAFitBsmoSieYod
JLeRvvXuZvixPMClkBVdrJuSMFIi44ucOkfMIRlgWZjVzkXlRw8TeLyL1O+HBc6R
Scw1ruUb2TRBtL70VB7VvQRPzLKAwJGVNvwGBqzwGE1Um3UjeoBW2htRgHppVCWU
/EMngHHEvDwHEf2NqJfKOkZyMmdAClQ1hsEmfOhpAjam2/pL7NoOpgaI57ilO1kK
GDiEnmmQLc2Ranj4GPL9F1ftlThD+L7fXOw+WCbc/FS96oED1+MLpRH57b+N6wov
N+7yn6Q2y3B53ENltkOcrdyePu9M4y3IIDNoXs0do0iWxBLI1Epnw0o2Ujdkb15Z
cLgmIenS9GAOeslwMVUoALnGRE3D6j+zAng4cBXWgT1+3qzFFoBlG3kbW/QVF/qa
QhzhSwERHeDt8Gmrj/SY1zsYmD5+PMNDPeoyCGjE+F1ObPcuyaRCMNBX/2I1U+M+
uuAsh3FOKpaav0WwidDCznVuTj7JfD4luOZvnjr9sMRs/FEDN6TCSMXYXWBh/9W9
O5JBwVdZ5uPx10uQ2VXpoaR2uwdnNAonxPk7e84vjjMQJZ8ynbhfYe96UyrZos0k
i7Ls5p+MAKsdeIootP+8jvj4GJotT8d53QB0x9kjfxzSums5q2inTwnkrSjZj9Y/
M6GPf9Cv8mdDQ1V2gWJEanl1Rym7BxhiEb9V7sBjVrRAkOPNCbsvkJAANrfMThIV
U+DEJ5kJViSGwwnZYqNsRWS49+LfKrRiJ1Q+IwULoNodLcl08nu6faHm/puc1S0I
tmbF4dOPCVbqochni1rXgpVnBYhOjfqFbIRqz48LqMdI22usNMdYxIYzMNsqrEEu
Z78eEEqgTqJatJrsEO+Sx5crp48Nnr9JwIjwOjf2hfjkPdR1xn1N6YPgzNj4kz81
JH3lAQKimn8jx9QjukxIU0xpLrQCXaWeCbp1vayKz5DGLsbi8OwDNC6qcf2owiTY
HFLbwtBwFF1bHQ6EGu7YoYvDL1kLxNGG/G8Heq5qfk3MJInsSrKGhElUXy8zpZb1
wFa8DkmUNNm422EjphWY/xm3AiqStrZgZYOA4/m9dp58sXztjhzj3pWSlYLO6IjM
G7Z7YWvRmbtGq7QFn6U9BZHgrbODDpkZtjv60/kEPsH5ZckwdhmmiAyXG1HJBqBP
Y2z3dOvwz6t3tjTnfrLUEMU1x9+TlsqwCsyj/iX/SbEcPU/jbGOmvn334vhhG0Fe
OmU2tH0QiBb+VOPBYN2rCGfvfi/Jfqh8JlzHdO/Wgx9vugHeBdofvrGObnvRhbmt
gHypV9JwVQW5mklGEByflpqHkjAv9EOURXGQEqEqd5WQSBSxTivjrm9SlNRGuLmg
34Gj/Kzsb+drAdwZhQVxtpivWSj8WLAnTaa6/Bii5w6gJvqMEYS4gHJUhfVA72Dt
dI6a9/Ywm0F8J3IfNnDpdjmKCyVPobb+mswJe6GSlqPrMpAhTK9Mt8vdJLe1DYrE
4atpnjuNtv+Kqo0d4fyjmQM4UYRHO4l9xaTjTwjQPpuDgtZvVyPiasYrmDpJSuXJ
+UF6RHTSvjKQ402UFVxef3yNZzcfHbZDF7XmchL8nAlkB6UEaWL0MZgc+EVMQ2rZ
uMSzjENJYMzVAIPx8DAoOOf2pRoQdwOonMO/4ayZBwNY9lnektEOss1RZFqtbdLv
gxHPccd8agYY+OS1XO/8IjbbRH9YxHe5FlYCGaGomVJhp4nU1BHUfFa9ac7uJeW1
HVKlfuZ0BS6fKl1ekPzYa3a9LKtcR9k3GZMVMvvx6OpvmREUTrP4kDKgfngo109D
QUbVzkz+7+iUM/9G1x6zxRVA6ugjLMRGl4k5dEsCIW14aAZtVbKxy3txE0GFPigs
FCVPpO70hy/M2YtYTMPyoctS2PRy5WCZSUgcqa+nzPL5ItBNe30Yf1+4K4jGycef
ciVJlkbvAykYEtBUbCZwIpa+qvsAPjk5xd4k7SrT3MtJredZ9kGUjIbijsefoJ9S
UTXmbUvqdZSusm2OA3rwEsk+g7aszTh2/WuHKSh6Osuxp/0wahK0Shvw8rW1jlu8
9w8agOur3+BkMZb5f6peV1juezZyNFrXhWLrvmTZ9Fg/L38CSYS08VXlpaikQgZS
MGZYH0tgZmP/ZtY1Om3krD+3MIr3KLIBF3spE1veaQjug+6EX6mqDg6JWpmHnVXW
K1sLCr6dNxRI0vhdiFBVdcUR0w3nMtpcdyb/iiyAShwXp+zQ5iobXZ41XAA2EXgB
7Cqoz7BwxMVaaEnj5qd6Sam8FGUJ2diYKePrMe4HssBaIeCgMJqvDJNpJXP+Df2+
iAuAyqiD9W9Wbp7lvZloc35+z67tqOaL4pJxe1gfU+qy2J2bfA35KQh2stOQ3Ozh
hoPhhoXHLJqp5QUAMp+eK+YV+bYxmtTqd4MIom9ikgBxCrNcvAcIXU6cP+mxOMjw
y3CTaJIJF93+5CHYQW16w+ibumLZPTtmJVEZmadeqpAH0+d55UKtgafUujTjoZxI
Yho5hioDN+kGPQ0A4c6/cyz2deFTfz5X3eNEbhQ+9hhvKgB8Pwy3Ze4JEhxST5XQ
ZefKz5GtRffli5jD64b0jldNvKTStw3tU5LH7jVg2VEPyV3KRb+QCTIUKI6rKfvy
DQmEJOlzKa4AsUbTJMPi6LPrnLGxkIvQCQl4sVMT+mWY9QDHbNvbQIzqkmLiBhl6
JGE1cl9czuQd8J+N4SM9Qvocft4dTtDZsQmzBuLCTHnouho/TKk3yXtFwPIugac2
N5q1lsuZg3MCDLCbR7vSPf0EdTXO6FdRhy/S860ckN5SzFKjB4uje8TyCPMO0RYG
61xxzk//fcl8+3P/tfFOzsAcKXn0vH2DnVUz3IxVmuqwl+EqGgNj4UJMJWhrGWSa
e0fvgwGfc74CbOvCg3PtXjAMQo7TaIi/kfeJAOCPGo4B6zn82QtPt3ZzSAw+0oQQ
0ZPy3mc1ORw8UKZNfFL9P9bvAzcld5zgqxgn5FFH9yIDnCxrftqomwEc2zBlt+GO
B130WA7eitBRwN2H83GqFhgnD/wgE9xPxkcMVusVC8oLTNz7U6NCq9D0qsRDWe3W
a6O5g7jOWMlNEzdXLikF21vjDmj1PWTj9JKx+riFO7kXiEGTjavGQbKmYoAcsOBq
vrx7gYKfa/Z9Y82Mq9W7pdbd9SjZ5ziaTdjXvSGakheDL5w7kxcxSuDVTEpAbtTC
pdzUapYP8lm3NaSx7y5sAVQng9QfsnbevWfoyw24pjOrUiMaCHEWlRAOCPjMUGSf
aQET+2mCv9gCYbQpViYD1N/NpwzWGdrv/lmvJ+S8qN9wa3MshigsdlXJIJvhyPrX
osmKTftI3Ev04n3yUclFUdwuhuOM0m2ZPbHHICs/g6Y0q5s/eHO1W44dWdFQXDDg
xm78HQk2v7mV8NfhmfaVh3mf8vAQtN4de0Q1egcz3WXfwSul+vlWgJ2Vqu54FZWh
aXxWKLn2N8GzWoGBaBSYxcbAla0B+zJFxqiHrM80cpNJ2SOrnsrE7a5oRK1Bml0o
2E0fUaCcmxata/2t5efP9+i5iFLXkdD2T414cNgfhF1G5ha9OJa33iYQLw5f4p6A
f4o/giwRc+/wwLQ9PHfPbxFRJQrgHLICBoxwL3dnT5uywJEi917kE32h4FclrYFc
JHpif42XJIXpML6HqtJcMOHbNvQO/wgAuea9LmhZH1f/GiQWdI9JXFcrlms87DUo
4rvp+IwaoVrPKMGOdWL9TlnHDgdg9sLWuLE5YQVnuUkHO56mGKiL5QUf/F6v/BwT
WGMsrdKuTUCohHPdsgWIX7PssbMU3eRVhE4aooBedypO5K/ZYezvvCsF071iwSfu
Ex9LMV/y7T0FJPPUQv0b/eMK9w1wVFVuN5MIhj9W/tybriEPqpqzhySoldIs5NeJ
UyMK2yv44dcMux1fKqR44qipLigLun3eAHh6AwUnV5YppfZY4C4YbHFLgPo69bGC
N1xjjtKAArE55V7oWEzyVYD3MXWVttmjjM7GegKUvq0smOZUHWuelWOOOfD5wQCo
mVMUE4ObwLl2u+baAqqHgwKqC50+k9mXjGfAtwfA5aLXQY1wSFiM1x6qfZmZTQCY
uRi54ZykzId+pYkS+b0LELPDLenJYBZ+JXJ0MenM+X5frv+HYs6Twf8PfUYlme5u
gxoFBTSWZDloOG+rbbRXyPx6P8xjspOSQ9tnCMatEGOUYyeIau9ThKmdMPiJdj1K
cmiA1Rbuec8gKUVOHP1oqUEtUP6b/vv/k2GHZkvhzpMcnHCk9oFJFUebKml/tNK3
DuDgtvBnowuoNkRMNLVDsmdclHSFd+bGWHLsvsxzjCXrcwjExUFH2LLlBxbMMuHI
fLUve0BbT9Hbv9FbQ1IdZbamzeTOyLrOh3mfqUJrnFWk8ZdWLSeL+CMIH52tDsuH
ksKx9rqlqJc2PKCsZcf/JbbaPY0+7B6XB6D5jaQqFyMR2+q/osatF1k9IIlCwZjY
bZ5Vfmvc51UnTZdhoCYV53xby/6fdLWwYGYn5diMBvIR4K611+yciZ7Gaelbp8P5
Ufd0+Fta6Y269q2XtzjkP2urV2luaONH39ijJ9VwaqURHY0Q2WM01lqG2/FcliWy
fcs0XPaaYlI3x08KjOqGLbSmNrh8M65kK5xrfFeWLQZoQv7HKG0PG7DyR+MfM7St
rp1EhkMPV6OIrpioUSxnV5CYqxbnQndAu4gcUK2gRxqO0hRckko1SSvUy3DX5You
ju6uNbDGdpDwS8xVb7RUepUTW8uCS6Yf4iQdx2ogCGv8lCFSlv/SX2LtWSwRORZD
3gQ85Cq3HUVWMig6SSu3FVmDSqJu/NPbx5pn4S5Lzsq8xmxCYUFuk/PGBWSAHKPJ
mufMxbbanlvfDlZif7OeGM5FkiYYjsJJ+jnTbU9Fl6KLMT4dW7f+Zw4dImDYQ5DI
MtwwpGgNX/AOuwbKHepoEjVOtG178FaIOgvarqHPxWYP40kIOp7i8Zvi3wlG4xiH
QOvWglHhJjZIAhRvfhQac3C67TjGjezBzK8RyhuJshj/DEkIIufCDhrbCahnTGbE
MsAe41BcWFMLcInL+1Wq5yy4pVyrcSg4ysAq5F0HilI9eTScKxxIgXvQDN1FTdUy
yFsQm9Vaklse1Nn0XrjMpJNCdx4jQDki277qbWj87yNxJxUty0MormD/67URRlIG
e5Yo4lOQ3bS04P4DPyK81aEYfXuvOQAk/IAEDhCE0vkT+cpoUrGBMcFPH7XTwYtn
6j+D3bMXXEqyFN+AZBNMofZLs4tnL16wzl9GjrPWEE3oNIOjqeDHLqoiieHWZKeK
CGFKYsEZZ3wxY5rzcnxuKAZUphPvhnoUsV1KJUOJLYoXOpQ7kv3ePO2IFOtY1/wx
5nPMNrW35tkV2PSNr+q7+hJSq6t21g/WbVEJ6DMcxtC3QHnXoWLMEIjf7MXPdxa1
h39NU+HbQwKn8FngMwWOvpDp7kolOG/ctbuoG1nnTnPJcD3ZGXqJrorZOZpP7LMo
sBWiu1yYXXEvEFph1NsQfbJg5P75nELY9LzeNAAnkyOymNoxW7DLxgrgl6hUI1md
uJiVPAp51Im12xHrhzN4JRg2+XScdcV/DhG9cpjFTDbtwvgYO4al9RNYj+Gk3wVp
SrWzWeLirjEjNJNUCsyWQXFtRdLtu9fBroF/FqXQvVGUZAedEfx6CbKsIww57gbC
fVpyHkomfnxH5FVS3J1wWTBsmmrgDZWfR+zo78OXn1ofgCQSWaPmGRE9QMkCUGDr
++AhQewRsJ3irgwx7Unr3UBJ5kVaz5T9lUZ0BAYhWJ3gONAgiR7N8CfAGgMc4YBC
3bB1xDVWNGdcV0xOBPpSnlZ0NHMDOCES5n4M4ojdGDCYmC6AVMCwFkcEi02eJrT4
SJsZsNu9/5a6rUkrGjm1+gtC5Kem57e29N2PduHYkNfPxx9u3UTVduIAA9JrzmSJ
iZcsxVMhcxYD9fiV1pwyAnBMke4WqEtkEBX4u+aY6pox4Wo8yOuIAcjIqChel7E8
1IFpXp/C96XZDCocJUMg0pMDbcZSY91ubvgfsS2cZjOKa+J+jzmQmkXkkrvMKjIb
lY37FKO0Gaog9dPZ6Bv5cxoAGGL0vFYTw3USUoVzF2CPElc/XDfkPQHiK5CGci6b
zdEi959RgwI29x20eGhljpOkNGHaIEjY70rctOeif5sbx47olYZQuQfSu7LS8xJ8
XcrzBdB62tVM8+5N/mug0UZ0hDHDP7NxVBwiZR8WYeWm3YFCSfIaZi58ZQunPo/E
3H7n0n8BZfyvUSYe/vEZh0wR7HW0PrMIs7QknkoNLz7YoO3A2n+fACkMaiY+rIpn
1GcpI8+VSizZrnPoLvikzBAXmvf41jZNrLAFxtTeC/YZFYbgimchzuphhse6Jdp8
u0r1pcFjFqJuITxyzrgHyPn+j7pONlj/ZflIRvGDQ0Aj/R+uCeryeER/R4ID52jr
wiMIoBS0Wq0pkXJYS4yZltaA4gk6y/sVn0msCQfosm6Ap8veJ9A0vXbjSpo/tvQ7
IBf++k3EkIV0b89rLz0sqr0SsIqLcP+cA7Y1uCuLwW78pLVoMZYpM0n+Ej8ULLqS
fOWiSHY263GDLYQBsgUVXjf/5UmMfblDAfzOwwxqHH230udaM7WreaczQF2pXT0j
2puKISaIKY3hbpBBbze3MdOkqAkGGDAGNx49gYDcxRcRQxIcplJGYK/rjfhy42ao
X2VRI3dtzNfEHF9xoN7pHoCOvfw3A9xq64nhaQDr4oD92ZSs0Z0qOPX0bcCDlyAj
xmLAr7Cupa5Go08JU630GRNeDM0O1nebGTC/WxxmQ4iX8G6/DgdOmZ3I8jXr6f/V
gx3NNVp+oiKDY04/nH8+PPlI161t3lBmRjbC1tq8yJMip0gbig0pZd4VwWlMfifL
FwIGDgC4etPOcU9MJ6Z8SMBAsLevMGTcCXQ0c3bxz6NlgM9lqqAXg7vDIFqMcQPI
uuB2JslWMohNyOv5qbbAIWaiV+xAWtQBatXrle23ulZKcAgPYRWTKBPejsH8EP7m
+pkFX/gTecGYvYtMe7xXPfFr6OvKdxZoAJ6g3lMgQB8S4jNDvE4IQpZd+WaxIY/q
bAHgaha5Hm7av/bC+9LIBrqhuZKT1XKrlXfYUv+86Y3c9URLCaOY3gXQWV/mEsn1
yteG2MnP1QbK+V5BhIJeMbfjPSsWX6j5MlCQR5HqLMpHTrNGeQ6iLnP8HrlzD5Oi
dbkyLCjAegAa4M7sGGwDpOcwFgA6a3hl3mRXedjc5p0YaVoRCGjG7m7MtlW9tp3R
iGmuqVVx1nC2GvjkbaHMJIam+BKgKHvWLyY5utEmW2EKXXLB75uISCEHJDYUGw63
RyjmZP5eJgHTSYd9Aiw4Ec8Fff5WDPsOKgfwcIFk5A4JqvODq6AUuZJ8Ud7Uq7VG
49HLZ6C9OvtLTf+Pa5VoLB6UIu4TgICTujSsRj/3UaNFtuhZj356Kogjl2S808G+
bBMHYFXNtvOZ2xJ9idxN0oHFsh27E1usLM7jXYMtFa6zmMxkEf0J6+wL9+HFsoXQ
RvOvSj4J4a615LntEBjTRPdBNxPYvtWf3X7DzgGJU6uQ+YxjO2glIHQk2Dfs+rhF
awUJ5MpEopiaP3PxATLgT2QZ+fDHETje1Rgs2kHB/S5vPa48sBM8g/4ETkJI4ckE
4f4uyUtTG8lYtoVhSsKPA/GoHIGrZodehVRRXB/eseR1/yWKlkNvG3GaBg9abcN2
RuSYj3JvVHV8QrHi4ove2oW2aFrvdTJZTia+0j4AGWn+Yxk838QdKmH+pGJVgzKv
1vDBA2PbpmK25xEFqKoySPaoEgA7RDcV5wo7Sj3YjDhdz0MZFh9tHLrU4SoL/oSY
QReRsgZEA6hx5VvbXKGf6+qbUVmG+e62zCUYTpwE5wS6XArgBFvGwBZGI4P0GGYx
NAxHCptdr0UpoBGGK0kHnB8mwP3wX0ioXhti+E8Szmq+7dN7ixkmyBuAkjR1ZmOY
yywsMeyTW4X6WHVHtjyX3DlYXtE/9HKQyT9fz8g2luj9A/XT+VM27w4uAOrk+rho
3VCqPsFf+V/94/ZihqJiHLW59vmPYmLySncQTHBu9dp5IxQl4aWwX+bC84L31ZvF
iyQD3D4T1wThb+JSP2+T2QF+9qpnuZU1r+N3w4pBGd+NEsSKVvo9U8XUnh3N0phW
ypOc81jHwEBQcm73rCySu2yVsrncx9svGezYx/rH4wINm4Kw1zppXAZ6bTSLDyUY
BU/J5Pg06eSSv7h+oDesoYewNb7v1dnKnL/I0QdylnXmjaJLT+SvZSsENekF2c2W
DOqOh/ORJ77RrndAzZwgsYlobB8KCX0UE80hedncVg8V+8bh/kVCeOAfYZD/v5CJ
zoIBzoGSxy3yQKNRb0DrOPbFqVpl2hdQ4vLnmzg/O60T9cU3Pdj5cRBaRenx3K6M
b2hKbabzkKqpPwbpWga2s+fLLacyNzSgiLWXx3TXVZLZqEWIUpEqERq0RDoDKzmF
juXK16uLfq8T9uZXdbiEsx0YbG+qho/+0LlrNdmtGiNAiQh3uI6Vw8kxQ6GO9jGK
QvL7jZbeY3tGnrn10yxZ/7LTAtVc38GoLnG7/tAY8K90uBd3YRcd6Fg1h1BqP8ul
SgP9MrAlV4jNP3OMUEQ7RgS9QP6b4aiepj+/ViMWSOXOYisZJ5kGFwLfE/vnNVqX
bjlxF0fEEfcMt15gNjk/O1nQa5y/LT2w3r2v6SyTV4q3pP1jA7b8ddPNIXw5EXca
Z2S87hvRyeha+ZFEvJxN1zGMzRRwF3x1uYaMEHVshJDdYtoU3+84sG2e+iDuttuZ
UbWqKGYmjH8F3BkMvCahpuSSkotC5XQc2DHZq8SPxIzBoBIDMBtC8dlZ1bl09zh/
QnIA8ebGabI1JjIIu5ceYzvSFpS/eZarhrYFJqMCnUT09IDqHvpPYlKUv0rnLfHV
bDF9R0+PsjwmfSh4WQel5J9ojW+2xEa6T/4mAIh4ttQNI+W8QNIXJI+qJDXSSnJa
y+qESrMDVVr+Jbzb4k7PBGKrLfG3P8tZAPiMcSh9QmBC0PswlKlaVulJm6fDhI+T
rhDq1eBZSpC6pJ2uw+g1l3hy228WMZPuKRhjH4aA6onLIFZJB1mu7hikK+ox3Bpo
uyWStMwvSHfeV/JACeUcYzvx+LS4yTmTjWvuH6Dy3aLXeYkTlyMxlzuaLpp/tHfi
AdmbH5tY/PkxnGYKULqbLSJLCGU0Mo3v1Rz/nmYY0oC4P6Lr6vj4djpBNd1iuQrg
+J9uvZxWyv4Cztyj5YOhmiu4NU5odX55RjPqPTzKBSeYH5i39Pg/PfjqE3UZgmCP
93inWP/ZcSttFCgrgx+EerwXJFbVGG58hyRDD9Y6hjUEVs130hK7PFGHEpgbuiGD
ImM77aazU9XOFkd+o+uaOFAGT0NgEdiXGqqhDLX1/cPELQpKBofKs0RryJ8cpE+g
d9hg83mrLB9Jq4UpWAn7EnA6IR1xFaWwWGaCrRcaVT72XbucSv/WgzhAp0utJXo6
IPlu4lEc1iqgEH2L8AySpJW2gciPks7B3RhsDBwOPH4bD+CMk1CnAj+3AEDc6EWJ
/WBCcgOyBXicrHyRxuU6/oX2etQVbzwGcO7YjLTJGj3njYTki84nsEEYvKD5Z0qJ
UpJ+Ui/yEIG9OZ4Eqm6ZFQz0WjllfX6rvBNZP+dc2+RlbE1GClgAVyxJkkcnOl76
6lC51Hb41nR+774abqB3M56dTU8SP7Ru8O7GJ8mJMO9l/sNHnoT5TgLAeGx/934X
ZJI+eLTcfgzWKGLMBwPoAu3akDjQXCy4qCU0RSPR/sgFfbAi8Mq035BZU9h0z/Eo
DsxN1otTzjX/9Sl/je+pwrXVLvp6jf76X+CypHD0W1pZAUh4Jr+J7UKXz2XawhnX
92KB50ZS5FTPQDfCihEhx4ZRnB4vVPZG07aDXyvQG62lf0MoRjEdTDQuwA8Z6+uQ
Aq7BkxBwY6NsM69CDY2Y8v48+RSE/DXR8UPGEVE+5B2A1kaGK2hPhOFnQ1q2YNOK
VXu+WqDMt4mGcijUWp+2/GZETqf67JUbANHnbuGhkK7h+RQ/YcLGQNJshDxEtqUZ
6fCivc1A4CASoRrdMg5wKcBI8k7cVLN0O0AD/FyqvDf0CuMcKskbrJgb2SrS7OX/
xGMNNnm2hUb4sZ8d4P2bwbpbRKazXr3joBSgghf9Q7yqWePZgnScwiSItY1wWY7O
zpdR8g6f52dYNrFUwS7JOA8N9xoOSxiC2MuFldHdfZZuop6lJZbt9BPDCzxdNIWE
jGIs89BGNRK85uajIBjLE7AakSc/PCQbUu4EUT3i8u2+8jHIM0q0YBaRx+FOauLD
tcSNbV9yenekFn5irUosf3ua0bbXIX+rX+MZUek/Frm1iihX0mysX2buczK9vln5
1nVqA73TD0+VF0StOPvVRU7n283YqB0MT8oxIVoQhbZU3sdqM/SS6qZ+3AF9oP8/
gF+v0/HjsCdc33qT3SUlhDKdtxLCB2X5Xcc3LPfS1M8p4GsciD1ubBYE53HeW0hy
ShtiFcYf/lgNfSeQNV4YmPZMfnXRm44dZGh9pNhDAqjJ0qSuKNdbMmOALAs8xizl
tTyzDoLalaw2xSvgYeBJeF/GpfIMG7iLG4aqale8ehli6jbt7jquyxAkMXsMovRk
q5B7RlUh+LZOGeL53qrf+3JUrW5XkTDxw1qBfvis8xeFmThG0GQmoqPR31UoPlzW
MxzZijd5X61rZjSXyhUw7l76D/rYc4hYxj3nWAgPsqm/TMZ5oZppXLWXleaKJuP0
+l2puc74Z7Sy/a0b1lsw8IDb9/McRAAhTVi9PeOzEXw7L9S0MoaqHcr9gcN50poF
pw3qwpsUt7aVxrJyl8VNk3V9h9V7arL0eGieJ66uUvoSOhLmxNdTYRsaj45H5aac
GmehYkw79c19snjymuT+mvd0a/alvWJ2awMeUAX2YxNfJv/fKK1iUhwvrQqHrZ7d
JuQvVMZmiY6gHkAhq6fbvXw9z+zC6kTfWPovnITk8Wyb5ZOa6tuxHaw/Hg5rEaUC
2lrQiOGp92Rf775nOWEVkaleb7fbqgHV8U5qe4lesLIxJQUQn/xg3KtSlDNz3Dqg
WTJ1G4FhwQbwrr7vPdp877vi9GURIVBoakj1ql+4VtP+xys7AYGROLl7L+1IZhl2
DeOsf9hMxYe/zTc79sSf2vVJK2Vze6TV6xEk0oeXy6gLcmw93g1LyZsvPkPXdmay
jCgX1EYGAJ4Z1VxQrHEPQ1PhLKKrWGiR2b8/RLaGz9ZengSsonQFz/fOSbL66PSU
ylGYAxvKURMb5FZTY6NSV9jKRG8CwlYCkSnfiOR0jZrYS+qzmHSYehxRvKI0Q298
mRfisuw8pcgMFHFwGheC2yFcEJuEHaMC3PzeeA4f+zVokYaEVIvlLYWOpuxLko2D
sNOI944KnAB2hkDEm1ECcF4n82C+qTTuzs/aYXVgiRogYo2qDIPf55cxAlt57X/7
kKToziOc5cC5PZ6XVdjqvyCxIlxnRcgf7PtcpritNgBc/kvTH07U1L4q43bsz2zX
EpkpObcg7jVEX3CfBTElMIVOZFTGSHnf1OBZoeZ2y3VCB3Tm5RMwmfaiwgXopuxe
8azmXLh/JaoV339nzjIn5PEDSP9lSfNQWFVNDS98PjtqltXkLvKMPvlRxSZIEIXE
saszAVIvj7KIhI5WANT9LkPqXjL0u9M2wGSasF/cdX3Y3WPKLsA03aXnDpSGQMAW
vSY/Hn3tTjohQd/oCyRQv9lpe/a/hMRlK1T0XNQQ/FPblP1iCioTvb7Vh2n6Whuk
KQ3fC96jKxoxDFq7E9ItqXd8uPI+nTW/74f051QOwUw5h6TgQLeX15R22zWXJWbV
qFD/0rWDmKQGal2jHd51oaCbcubagycsgGm4CpC1/HdURLXRBU3dakWIDrsZOPqd
UArjSxcy10lwhImg1VpxVUhQkS3rZ+mPiMeYypk+aM5qJMoX49QtONDc0GVmQHEp
dEx1ZgTb78r2iXAoYK7Sk57PHYuS+uF3v10+9Qh+O4/JaRroDmjaP8ZkF5fzCEsU
gzBfiWA/cJZEzliu6vQd9H7ghboKgumZRUQiW3UCIGrkG8pESrjHFcfD/v9K5hnz
4p/ugo17V9nZZLC3oQf//5yGcxGAI2l7TWPC8pl9T+xRmfnF/aJaEnTrTTFmQksr
UhNrnGkiD6N78C+hzjjc6LfYiOjvCrqmzHCfISqDkctQbk3FtLh3wqNe+UvoDGfi
9UfgKvffjAdqWq7FulE6biyjokbv9oKSzVt9G56nU9YaqXJxcU0HhIERLWTtsDlx
cgdq1YQJ2lxkexNE4vEyT8f/2a8Gvk9MjI25S8dOH0YglzeS6kI37TZdvwrhcItz
jqUbArgQUTx1jkhceaYsp30NhwyUuwus70ngS6TIVP8YsUuXtwMz/FTTV7LFJ23g
9edJNRslh6WbMYVUcPVnfx+nK6zA06gwjP+YXhVkvBnWMpQvgOuF1rmhWLsbSz7x
eFMADVbUDoOyJc1/vikmU7302TZqCW8EyaoS7Yg7NkkqgfChTw5ifKEigiYEtFAi
xrJcCYR/GcV5fHUhcLDGSBsaIdokmbQGxjcfuEMCPafFL3rpeAJZ5t0Vj0EU/cB7
Gd+WbAc8a5UiDfwgu3LoZzCPOsq025kVRY66/sYkpjDPYLqZHwsLecGbR4pwsvW+
ZJxPRjJ9b6h0mh9XJhEg5R+ODVVGKWSZpD/4twSvm2KyZKc9t0y2arGwFFAcDvm0
SfT/5RYw5afTM/AamnA9jcpgjPdzWCqg8WJ5W1za5fP4xRDSoH6fwX9utHjd1SM7
LIkDXI35w9dTZUTbQNQlP6N7XJWkaUM7ekPwqFK/wVpyPdBxKFj6MBuXIa3j2W16
C7Mc+M2vJjGSr7QYbAKiFCxEiLlQTGtHU51IPDhYSVChFp08c7bGk1okxZ3LV84t
qbrgB5HezSndTbLxIWNQYG647iiRBq0Sk0F+OkN8UQnVQOzOcGHE/oMkyZ4hXsrv
LjqE+mB7+ATlT53jwoo2Xb9gqXEg2bK+2GvEqYo7tuQB0k29v3RokR2Jz8QcgJ3Z
xZ1vjRzC8NLXNB6MxuWKTzgeCrEa4fPPa70NLktJgI1sIiMGq3BliaREkwm3yO2z
isgrSqPYi+zC865OB/COOcfYzFLY479azODRKcn0QXudIkOJh3UsEalS4Kqb2P4+
fdyqR4LDmDSwJRkUUV/DFoctUWBizOXa1+9p67Z7548vxr4/3EAzrmoGmEu/bQLp
8T3iyxWim1SBL+zMgKlTZtaVY8N7fxKA5UrBA0SNBu8V8JHvfqYGFtYSu6jDyekK
U81f4gOteutnsNylX2gdZezc3/nbDy0R+q9wGu95xDOhvOhSApuyhDN9WyKTQ4+5
oxBDpISHl8droU3Q+Yr+/nEiryGuRsyc2xjIF32sR9hiPDJuUT7r1L2ewqqYvEnF
YQb+q/+lWUtE3cjuNNrziEr2xEQl381OAwQUD0a+Z21yoP4pzPt5jaj5X6wm4BXY
rbva5IdNoykX67Z1gsHQCh+R8Topz0WGpj0JyMVc77wDqBdHXMY1ZbTc3HRhb1xg
jZTcM0mxU7gi7HTg/xVhthCG0yuYF/qG7TGaCL+5V8rHsXFLux5VFQFT8hqhIqqK
gChOip6DXa50rQlxQBpaaEybk6+fNNB2IOLDzkaM+BG+Ls54+huDgZQz//6QopYo
NYHkup26XPJtpLB4QFOfvn12zl2jAYmCrt8wZYF7v0C/pepkAbJHLMUzCHUy1T3e
Xu31f+aB0GAJNOUhY3Q36LtEiNqCrxzi+/S4EYgwkqQc3bfxAbPY5z3izdz/RYK8
WfZBnusPB9yL0MKcUa1rFphwAMAb8jyxYsHjU5EyHDe0ZDmjWMPRUmVUqtE69NbZ
pgz+dt79e4ZsuT6HR2O24C1x101ZM0Ris4948UaUEZNqoOYdQVkwfMAGHw2JMXR3
KERFosyvw1a7HKS4YKWYscHqYEQ4iGjCpLsxH8j9gjBaznqUjULgBgDrm/qA5Mw1
+IKJ+sNn/+7z0UAl+ks6OT4hQ8WL9gV47/WbRnKNk1uZPMALEk8eFNe/isCqFRDo
CWtbkEL7EDY+/2sLHyGC6QN/kOsCkxFqafPVfGhOjgkCZH1uiTnHcOJVk6qqdWK5
MIELjofg0Emwc1gcMRbkKOREZV9bSInRTIbRyONR2IXq7/Fis6FexzIz6hhCjN/P
pG5dt7G9pTolXXVZoglzB03NCCRwI+lG93Io/WbRSSG7d5HmmKZUv/CkFmKPiQeb
b1IjqVlYOU2zIg8lH42ks7NVr0Xg4Za9UyoHhzeOitJeAxRrOG2vLwjjXc631zA4
IQPdR0IRwPRy1Gb0lnvy6ArBE7MVmPEBsZ40spa19d6KjKpb8MxyoeYQGHM8P6zY
SQR4g1d/4tN+tzQQ67dMZqvooGfBYDQu2nSw3g7E7AYzwoyDFACG3SkLEvlrJQCH
pBFgJOt/+C+lb9qdj0TLebtnTVrfjMJZMA3sNzBPsXH0qSqnMz61WeHG2x29AgZa
V2sQrfHC5/utkOqm6AzJHGvrGI5H7lboGaSPA6+YEQV6jsvgbTiqlefD/r1/YzuH
9k6EqUownmSO0rlIRPYQzaymRgeqHwKSe8668NzUa3ukWiM8+nLMHoaGqG3uqqf8
fbReWXUEpTLkdvoyKI8lEJTsW8KR5sdND3lVhyJxtVXv2RPQjRHg/Ff1dSoBxTGA
UoyHdzVIzgzbaoEAYB0wzXHiQ6hvUx4KF+YqW6pdINTcW0MMGpgw1fi384aj4FCp
GBCWeRKMq7OGDNrKtJ+6WU8I9VGkM48D94xySUmIwgERMDo6HqclELtDa832JN2+
4wGwsWWrAHfFLVYmQwDVxCi85ZGWeuW/F2msfH2EJ3j3OyTtIap92oKjL+IDERid
AU1wbO0WNQN6hiG2mpE74KSv1ZYAUbhR03yTAkNdGtZBBEgd/JF3/rqLtdkA4TGj
0YIDjBg4Hvy6eRbtlpiaC3+8gMmJxKCKOsNixVhja+nutC5JXL+o8dgHLvlC+82P
5zujmuq8PoVDkqG37uRh0dRKn5rphOKKgY/uUYKLwp8Af40GOk/ffGLvhx1V4kyi
575yAkX6cSblLMgn609Sp8jJ56RM6RgaECHf1BGJZCYpmZWOGndbPDt1aPuq2zTM
n4q1NnXgTmSmesajqcOUL7WXSnjzV7TwBVlJGj6dfeM+w6algwFaZ1FDmD7IlllA
Igz9VOBbURAW/QZQ7c9vEObQ2F9Dk9nyBUGeJD+WjHWP5Sz+kwxQMy9jtEQf/evt
KfgNSDTIvJdFqvjgoqbsWCH7lTD5RHdSM1tShg4/tB1xuG90lpvFcjnO6UnON7ZV
9n6zhbcZ7FJhtFEhq908N5tbZJaWbWEIgTJpyL/XwbOXPsvokgVORdYJc27Pyghw
xfc357JxK6lAOrvU11MHuokSoQBRj5zxiYiVxRISiYH/RQ2Q77fXiSe/WkGC/WCJ
y46tLZs0n7NduGEicA8o2sOJ1JKHqVtkhz070HDUp6yCPk4tAKYBiVh1k1jozMql
J+rbTdf/KsShC6zprZ13ReXhDIuI7GnYD2kdPRZV4at6kex47eeAaMX8Wbm41Ns2
tBalSEkntAwrGj8UMGWVy/F2SVxeMx75ry1TBuYAq/h7Cw5cyZBV0laC2q5uVnoG
ArNwPsL9qdDGzxrBRlU6T8J9wVomPcUO0DH3EIe6KXVqZ3cYURfG4PeyTcOO/A7j
VXi3SjqcTiTj9cjUA1WWf+vyZD1SknuDhVJjs9dGPuMw1Zj0poZjZzycQRGW0N32
RSLDDWNXHlKKtzOPTlKxp1VAli6qHpRhGD4Ykx9KwfZpIe1b5j21sDarA+xLerqI
uODRqW/+FrK+AWlPiN9O5soNffQfbN4AbpZxSv6SacU8mrZmlZVI2qmBOSspR7rN
Pt4LpwRZ+OeHGx+aZapLPB5X5RedJYTm8u5G463x/ouhV3/PPXmzExZYXCBFBQgw
ZsmkHVqqu/QEAWRElVcDpYscBvMCPM8jfNbLm/YehdNSjWGTLLzq9YaQablFAwbr
bjpXNI8DnDVmMBLg9rJN+NsK+QHCrb7H3mwLM+HfrDz7dD8Kat8EFtjJq5B1CAnr
aO0O49DtbBYxtsYpJocqQJgmME7Olz3A1wYFX9DdBRV0qdFWL3jagT5LdNPOFrBc
6wmq3jBwI8qXicteqU4ZOqOI1+4Q7WwttX9QNSv8ow+R5L25amEd1LKk7PnPaye7
nd3y8JdmPL0xoVlZqkoeXwNaVHZV/4kNLA7D1wB9L9Hedyx9XfwQEZ9A4Z8+5aUR
ilw0bZUiX4C2sBSSkpZPeb4YriLjibRdb+aG8H1D76tlWC66cs7fvI+trWXszays
gvPhawGZedjre+uCXbOSAPfkqfoThwbJVnxKucH7NiMB2jktmXs1EzYvFZT3I94/
JxPmdzhJxydDcir/QitX/DcsNgJ2GyQD9Io+YzWJy71zAU/Dul4R+hCS3EZOpXIX
gNAZIIShlg+1uIa9k2BPrRtLWD08Cd4RCOUJRd1DO0XCTvVHnCrhrgGt6YJKjSWD
mOnU8t1+LHhM57H9q6MMZrazHjsc6VI0K/+cDH40FK6YXUGeR+rw7yslAXoppO+H
r4lsdOwl81AzLNvh03fugwY6IjkT1tmpvP/Ca7l+8n76LuO03hoggCcAvvxku/tG
ksotu4YPKSSEQvVheAyLEGoun8owid6JDSJ4+IW9Ome8HZ+fnDpNdePPrmvbIzEC
xOC8kuHK2HjEJ/r8lz4LwiT0PoLwII7gTooqYFkLhfazFlm3Eh1cE3SsJah+VwnD
jch1K3K2TjYKa6noK5SjVpxKnL871aDUfiAP45yTzBOI+gGOYgDtQIboMUExMHgN
ELpK9Czro0IjNaMVq37dbajBIe628C+WkdLIkOO0TW+K8sahePsPRFGISN9/gN7M
mdmyXnRoMapfBH9z1kZtFP0eXvxCm/zkNM9wQ9hjNUZk7X+0HkUc//sKYOy7hAtC
RrM/U8trtH7s4+ZAlpoCzwGNLESoKZg8RgfO1h1r28fjw5oGguQj5zVr1RqikU+k
w+Ed6RMorXDoXOXky/hSci6sIO9Nt5JXTUxu6kPSITVd5x/w8ZleiVLAzvythfFo
QCs6uW0vg1TM9G/juPxBsdLHtJy5D6pwxEWKpvHeKk6dtbWrmyQbUm53q88vpXqV
BkPAiQsxiYz/rBCZwAFJ4o/A2vq969qrPDJw9cnitqEKT9LMaGs5wpoZVE1Y+5Pf
xJLCM6JjczpCAT/wxoqODTSJp6XhqvTxutq6eB/11HFwy3Ixjw0m9hdWKcGATK3q
lBKIrs0U4u+8uUlp25FNOVrGcXBqVhTMPlegmJnZWa0CKuaM44y6VyZRoM16KVkH
96y7v4RPqsuv+wXmH18MWIc+7QgR9vDHLTHOnSUNcEHATvViSgxob6M1PyD4xd4F
TGoB+iQd8piq2s5eDAHekxaH9ISHCIkv2BGTHn68TS7fuwWcVqlxGrSZT33E49xw
jdDgDu3vKMo/no1aRWwSxktsYiqsmkEwbb7dT0JaRjuRB/CNHT/WqdkyAMoj7+5T
UGQZYspopy32UBu380BOpDTcHuzzlUkT4K6QANyoqEltpyDlnpSnLv0Xo6sL5EQc
yzRm2M29TB40kScDSMQ5kr7kuKXNq//Bn8d6dls04xnVZ7rmf7n8Di1n/30HML3u
TlqHRpy7B65/tsEh1ykymjHv1BUcRjxzbPC8QEv971foR05w1QHsX9edg3OHT1MA
bjEU0+cuWzsBamd2FEO8o2WcQcN9lwEzg3eJrIecwfHFZI1gI8ZsQyr97+TUpOgj
TQ03dPLBovep0spiHlZUqCHwrlZzmHridmveSUFiZHfXIxDH+IMXlbYETUN6Wwgv
8NVRx2O2RIqwUOsQHicuwj/wWWOBjYCAIdCIg9nXeG7gMfnTXBw8Z5Kl8ox+uSyi
En2oc+F9HymMxwXec2AfC2ggmAT0CfXUy7+udPgmpwClM5THoznlhEIzzNa9sWlw
+w04L9XaZg0ELR1gc1XerjanxM4Us8mkw5cMuHKJk3ocw3f5Xg8k++UPvG8WaXv/
AvuZLmimdWNLigejCL7iM5D5EjT1J3nZlY2oEa/VjvXlUkU5zcr0bKDDA/SBD+4z
ULxqadQSUyLxbl/MeYNbSkZuAEODnM2gmhEphG359NHfWdKq5dfPSahewyRUFFUn
Co8oarQgVSjjpcawCVnDb0e6B4Lc/p94S94G5EfJAMir1vrDQ0VgzutKYqygQCeZ
rXxkKMGIY5Y4mZFIiphqeHyrjvrw+nZE1PMklHffp/dEh5EEXxwHXhljvB8TvEr9
c9ZeNKcHcj//0CgH0ryr2XxbYnwRlpVpHCBWm45uGVZoDR2c/ViEvRVrHHJYY/y2
ApDo1a0DQvfaE2xSu8+6S3Z3cczGrjNYpb7arnDmEVY0D2Cibu0basKA/kOO7VOP
a8oNZkp4dyA12DPSpdE/WH377lqD5PPNPCRNKC969xd/UDk0z1z84t7D3m4liRUU
27/2LCmPkXbX/LxG7hEbdcfBatQsRASWfkjWplmqVVuVpU/uWzHXVb7lDokUAA7J
1tR/b7NvC+iX70gJ2JuLm87I0XEYccl1CsW67u1UYloVym3OImwKbPBAVJPtbH/T
cGdYSXIcMW4EO1W+tvUh9P3xC42CRFuGIKk2z5HyeiV69JMgQy0U9Zkau+sVg6Ny
FdjGxwJ3DgnEu5aXNLIqV5xXxTbZRZkF+r3R4xNLovfi8W4uFsA1B1sBGvQIa6UN
CAjbIJsJ/a3PtPHwrN63JkXqiWwLLfQsVyPXkr3iR0ZKvhepf74WR9pT9zA9TorE
j6LhiGQ3fcIMn9Zwhr7i9DlVHL/n+29bthC8Pa0zNYXAQ/RLXCEd+LRSmeujJ0TX
uoXQhJ4oI1dawO1QMurNRmzIcFn+cH0AiKrH3OHcOgTvkkqPrJZDzjTZC5FrjS75
gu81e/nJHNzG5RVXKaIqjiQ6n0SgiOn9EGnUChOItmqj1vfnOIwQH+r8SZZoq25x
6+FNml5KaKmoeJXfxOBFEOfH5XTQkpNzZOLe0/Q9352fFM1hcUJMUpWZzLo3n93U
Yo52YsWOAlsUtjcs5Vv655mb5ZL3cdFHW0LVANGlnOMtcu6/1Cpmoozr8WcNS/kR
IzocrQ5/51xJ3nQHfyy+/sw723/ipmFpyNcefTXiSuZnbkwqHEixgqwnngkih3Vl
ndNBpt6oiE8kgCzo+IMXy5XUrMjY2GATvt/b57RFdQfcnLneAKJd5ketdzM5cpbd
7fD45zA/0psNK40A/GV8F0di+bCtYCpk1RTamldpjx3osll5XydwaTs/GRqavPIU
lmf+NeQYZKvlTtTQt/0CEYbh0HHM0/Rp0kGBozo1r66ojprmqRGUWfkVICkby2OE
05/uno99rA4J9XB6TMm94oR7F69S5ocmN3KBVs20iT8kuvB7EEL7Ty0hyIyjNBls
77A8mRZTInGUTXvzKazHTp6NiJLNGylF5bG4FX9VVzYN80l1UGRqwOEF4nc7hmrS
O6zJrxScudm46lmsxVoPOAMTa81igy7GqblHQWHq1jnD/li9wfCX2v4+4QUt64+T
OqwPphaDeLt1RyruzBe0UIL3NH++07VIxQDBti48adkTuaLEOwqQnQ3PxUNoSg6h
zdjOG3a/GT45iPub/1QxCRxY4HEsrtFTxj/qRGhpmhPN+5lz45ACd6Cjx0LBND4G
kUdHsaYzlZnrCNdQo7vW/mwi1J+QqqwlWD/11ZY5EPdmTHlinJ2Ee77jkp2ortYZ
FZ3mNaxKAAzDZ/RCb+RkgaTKR+T6uB8kxrPcd4Fmnm+FOlmV0lhcwLL44vafuUsp
cD1/6J6aG9eDJUhJ/y+Z89Yr3WOY/hfB8SEmEhSgGAJi5en+JQ1/zg6BQ9XwfcGv
SqrmXdICUIG5KHXAFNNII9t4/9T9gf2TzDItQDpbD9sXhCg3gP22JQNp9E884Lmt
4Y4LwLXNLyV23rLLYcqJf9EwrgjxPGqQgyVax9SMv3gGmvMO2nmnWMPYz/rbp5YG
aIWt709wlMsJbDZJ6UV9HSTWjHDMBw/NWwaVbbmCs3NwJkzpVOYxVZYdxVNIVKOf
uyKsc7mM4HCMsoB2xpLn06g2L3uKR86ySsYvMqsrfJyfqqsIpPf5PAyL+CVj7rDB
SSlJGzcF5ZV2myZ8IN477myY5PctItLRNxAvQaLRs/xMXzxGzhv8ttkyhsebjHVw
7z5/R2/csIKAP/Gsfm1eY4rHJ9+1KG3VTWA1xu9mw7NoZZsw2F+djhiqD4qOtQRD
MH0m+rJo9SCapIHtbHlWm7uu2PV8mN3MbSFDOVgjGy1XFfspVqVJAWKtm8su3hPk
hxH5sPOfIiZTvVLKcHOtSEF8b4TGIQEVIJK7Jdc1bFCO9LyXMiOE+78uh2BTSrm9
wSm9nCHY5/MQkdi39Ros/gweIQ7Afvp6gu6E/Gkp0RymnfhNMvFwn4fT+RfKhkLb
PIGM/uw4+CjOhd8Ku92e+/UODqPBJv6a1lGbaZnK4/NNwWhwtGDY13C0egeoJWEI
cxCaKe04tvmg2LWwiQWsicYKIaXfFJrT9lKFLoh9qwaG6K7vly1BuBz0NBiSyJHW
JyiHgTwSrSfnWJaF/IVDd/kEuPTVg3h7tAyK1quahr8o1vn5OrjPrXsbEnau+4UU
9l/oK3FO2SMmlxxDdifBp0awTQ41jBtWjA/OuebQ44KUXVQc/qTR/UOJ2gu3H7TZ
FgKAVE7DXZZkj0S2j9F8I8abfXwiJD0axWcaJnFgySeIYhmzDmkT4kMePk89jjiu
QXQJ8UNsZwNN5AuOc743LE9sNSrp820c/f9uXNSQkga+1/KGAloqXW9kyKYQxcQd
7k6IfqnN7kbbfY0hx7H/UfgpPRZQXLTj4jLDYrBQxLpbydP/WusvbRjm2lfp08Pu
ykC/aYXDZ4ebpMegmfXGzVAEXA67pisxWQIezWztX58+VT5/9PAMt5pebQhiGasp
6lrCBkahR4l7VL3m379CKr9rhM7MJkXTSJA4UvSZZrhCaWM+t0f3+6OPLnnWO/CX
6A9sf5I2fn7lWNjZqhrxXco03CV+wbh8uA4tuNhD5sQuhHFnuf78Mf6+eJb7yX58
tXxGypOWyaMEDraVRrUUeNhlPw1VkzDFv8rALUpFqx7/RgKPTOOhDwBTj4S+KDIv
2ALiO4isRmckrfdzDGmXCcKhXCwEI8xJaMpeetRMi7DT9Xg8sezzzdJrO9cQYD2Z
6x+fjKIC3kdGrTLe1yYvgO2vjsGes6ueRgCoNeewfg644US7SmVQzqmjG9QcRfpR
VVT+ZESQhOJx4nT4ZUlN1cLV2TMBV8pJvNE3kD1H2gxMFVghJjs7oM9YsGhH/p7M
LUudZujtX40Bva09vmYcj34Ry+cpLHJt2UVWvv5SHnnm2Knf6+VPO3rKLYATABig
lZoIQoExNs6vjX7Rn5/bmB9Bnh4l58uOpIm2N/vwSIpnzOv5QWelhZsPUQjb+pPo
m/swKV+8O+BywVDq2+E87R69I1TwPmf3gmk+PqMCyfir9BVXZYc3zyOQoo3szpVs
M3c81h7QE/GEvFdeJOCchJCxGz9G+zLngYvzMjFf74JKpA/oJ2XIaEK+plV9b0cg
qK3cmIrFbCVvjnjd1+QFQgTKsPYHnMy48SM/b10FWaxRnVKUwCoYk5RoP890sbIq
Dctmbx1zHgp6/yqurfp7M1mihRrNVc8O1RMtejitBDvxiD4ISM1qNTafDeauw8K1
qnCH66VI4KqYxeUrGsl67nmmSnoeBJJxXjBI4D56B9RnlRo5Ra4dS6/QzdO08azI
vm9llUmBVtkp644sS4ZajIlFevlp+8bWMXoLx/6NNlNep69bdY0VEydOb5bU2ei7
L34l54NS/nZ3or7WgkRQsG6PbviLSqhl3FqVvPstkM1Xou52KXlnEJhxLf2h3h+0
5b4fnYk+Du6PPetaJt1EHDgmVxWOtQUICAPJoYWJO0l/dFL6ueiMQT7PkiwAeO6e
zDifRHOc9YZSN9XSjUR1rxh/wfG0ozgTo8GNc9DLBCRANb3TN1o7clYcy6A8xcAS
9odTuxx9iONrh6hpFXi2ojgW3Cgys5U3ZpP9uiqXETOZ+l9KY0H6lMqTGRFtRA6u
kEXdgdUyaadWxYKcdGLtJBmAoosdGWYIMkXuRd6mMCZAJgsKnYQvBPkUJ3d0dONs
hLt8hqH8ukpXIt5V/ZRoZBRKcwbNOGtS/awLQChjRipPERLl+iKFbpmY4nT0zx02
KvuHV8pmQEm0l3EH9hhCTA993+G3qeFu3OXaiJVM72wcZnv9u+fIB9gZ7kb15IIX
+DG0SE6KhpFoLKG6dQkbXDxqs5ZPTU/y+DJmSadtSxPPhoMuVHs+xHP+fbmD/OOb
nuwt1sFhTwB4cdsQPzPVlZDmhsV+LESTd/F/rtTx62GhrhwKIc6hOisQebnLIHV7
8fhCSjigPwBr2W9hL82zwU3JCdeywt/VakJoP3vyGE6wwqjkq1h9ckA94IkodOY8
DC3s167NM6WNP1WtK/FYj94KeNdC1ECoMAWNrilKXyJ/5ecHvHcdbT1Wy6UjJBvi
8eDWG9gy+AxG1IemhIuwrfn9KCByyEVvF8C6l8Y2mF4mb5VOMRjR26B+FFxSqimG
qIeYn69AviMzNW4s0UUpd3aY2Ota4ZwLMFPMlDaymqeSLWTrJoOvNj0qVdt2XpGb
Zm+1GZXsLJPLvqvguM6NldrWOh1YItXzAsNussJ+IQWz+sQr4/X73xrH0eBGckJ+
LDbW6Wec2woVOlFCxUDwgwRv/I01GqLuW2YdW/OYDZcNiIENNDYqjRKXCsp07J3v
hY28aek1r8/vfT5s1hnTKM+7cEUCHpgFguON9dgb0NKDw84kjx8bT8IKtwBgFoJv
1CkslIH+oCulZ5XlEcgsT5MwD6miEO7VNZLcquE3tOWgF99iO9IiLd3abdJdoNJx
tT7FYKfj/gzVmQhMBH3V7CcQwUCG+HYlZ6Y6aBSMswWLarNSRiE3evqnU5yVmqCM
KGULrZyPBr3bpqfqs2DI5Kh02EmBpDGMAwjW8qGzAx6eAkVModMPiSnxd+SqXuMo
xti80P2Ruaelb/y6NKzupH8psj3Ck7X6glztJgVC5DaAa2sddJbW2L/ed4w9t4CS
pZ6ZHQSLnOJkpblwN7+wR8psz7wSgI0+SJRS1sRMYLrBveDmpxl8s6zfGiSGZK+L
auMDE5q1RLA5wAGKDJgIMFuiw44EailsyyRHZNlR1ve7ohs5VrJEobr/IKPYQgst
/2gYVjzZY32ubb+5tNGHKsN9XH8BMz1H11JyiSypD1VbApI9UZGMGa1RW/+qhMFs
2shUAU5ZM3ysNwfmQJwBoJ8OYLFdlTO5SuWOzL9Q78nLTMTQ3dzm8YrWJXTP2w2U
g9eL+sHtEB77kwBh2Gd957ZlXWx4QFe+YK2It1f3EY+qriNgbVEzXL6Mt+Rh532Q
mtaqXHZGp4jEjV9t8hj+Z11SBN32pIQ62iVwQzLQH6kMFc/dOeQ34wKzNBpORjjI
6prtl2et6AKOtGMmCXwvIGBjyvQboBt15lsA8w6twm9Vkd2ZgZTiI5RSFYpQrkEQ
Q/eDewGcgllkmWuEuHXnwEh7xvqQq/r1XGZxRY5u/4ikvJRazgD8LcUpr6dhc6UD
gNUQiIS5cZsHnJYMDAYoIPx3/e/e4bagVGqXnVBje4V4LHZqgr4DYLvxfbq5VFYv
Y2vcQl0CQzO9kwdAE21YVCg30jFkZS4PfZ1ZFhHmAgiBkGcqsvQlg+Ssv/RrODAd
DJtGqT/2vTc8ktmElfx6XUp7PErkrRsyKmeLZWyU/2bCmg3D0iyB8Go1R4a/xlK0
Lppd6qeVmpZxrnXuEpzYRzZ3pMmL1ASPwWCUD4Av9OtaNbMCihccDkeca3/wMx/W
S/CJ5F5oBLR1xojBpqarzsDzf2WCt2VZMrC+GxqHu12t9/+G0solm8TS7fTmkVtu
OnyZ7v+3S8143TZuTOg75NfTv5sGxnEsr7OuB03ypzblwl4Mh7mhTkN1N0TjKQe4
8DLJ5xo5NJMC0bKZNoaqfxgkgD9DqBDNWhWsLNA8KNAJtfq00oWLO3R7rqCL5QCT
MFCTUfuR6IU+neRAFYory8iBfnPH4cv6WbZ7prFt4T/F8xabh89Y3cuSg4Qyvx2j
BsWbKA02368zNA9EpfGlErb7aOQ1D51EVBeWL5YbqrbDpSfcut7339OuBatsBmFs
0tlBAAVBRscw4Wise0DzPMGf7QHFc7gPyYp7blNhUJPNgUlPNOKf4nurL6BIDwvA
Yi5hhLbFtz9IO6sMKcKlhcttVR1JNksqmsvoIr7xFx6e0Wbhp+3+J50/khx4qGNM
ujQ/wc9yDz28nD0oRwScDUYAIfbiwalmBMqluptvbS6TU3u8MuEM0Uv15kXkgKgd
uhd1F2Ec+NBp60iJize75MYjcg8vJIJyDYYzXqRPd44RvrCuICXutTJT9am3dfZO
lRwRNF3Z8EbznuDz4FU42fURj7DBfOLXTfe7FX2DYqEk46iIPpPngbXVuEF/PQvp
9VuMhHs02zzYXPMOpySyLuu3qnYNUpR7NV0x2sEQGbJuat8YZxeAMS2Tthh9rbBa
27xxaehrzeQhtiw/UyGpMbhiJTISc6hEBzasbmNQp5CQems0AW3vmwMyr40Tj5Yb
2DQGjs/VMDptkb3OoliuO4xcDsTFOcmaE4BNVzVGHviAWa87QbtPahcnsQ0eBCNR
rm8Xnp8VuFU/AQcGKitCG+JzKqtjrtUqh/KgduVElz4O86tC9bFR8aPD0+nOv5hC
6dWbK+wN0gRTDj088kl9n0gmn1fWMvhcxlbroHx/rABs6q1MQ68gglIZ7WnX2Yva
iee3CucX9eDDn3h2dQyHQ5u138GbKgOvLlfWs0+goLCenohhrmSWoRRLgxNbtKB4
1IG+JrctdI63la4PHcU9caT2YwPOzeEedbb/B9cCVv2YHZPAsI02LKp+L/NTjC7q
AndCcRubpSjiOVh01lw5BeNWe/c6OwwzjX2DBXouxNYH5p5kMM+TGqrn7TBkPrgN
gZyc6el/dQnHRWV3y7TyHNktcEDBMXtWqcewTxEoN7fqFaRp+Nn2/RryTv2/Z23M
i5oagYsOj7c/vUCJyoJ/ely3iRKPLUeQyx2aXI73EvaqotEtWubQIebWrLqVyW5l
zzg9kE1xD5rSpO+yUd+PqIKfizswO0mc2+VJOUXJF9gjvkPbRFaQa9OhZ51VbT8/
NPc5tj4d7tTue5ni6p58DZ1dBZDmZRaPyQ1ZOL2x/pCIalU3aY3F+A6zP3hXUYlG
kkqQxTZcSZc8FTQ+zKF48dilXbfr58777kfyhz6eGTPYgWslCLrxb0hkE0RYHL9P
Hy0MWDThaFMzmLNTstVRITyULgQOH7TgHQcL2GKNvgwpO26j4b0IWWWN7+Hxfbgw
8hQtgmYpw+y41ONiDehH9gAwW9Nus/BEE79mX66ybrqhABi5q7wTwqlbmLHdq3ik
xY+NLKTVg8aj7O28OSJEDjJxUZg9OYkjvwOnKhht0xCKRr07bWNTyANZswmy0pGn
vzNYAur3U2lLC5Ij97HvOHvjOTSfvL1ulf2xqQAhlOuk6oR7j7rTha+3GZPttjxb
KZ0AefrDxwt8sfXh+c5vhBtc+WfEyKCnFkX2rPicvAqSZCn1U2+D+Mq3jMYW27Pn
KrO9X2AJFTG8g1whvAgB0KPg16fwCY8TS54yTAw6vWdfi+jEhpwsGt7KRLS8pyGu
CNm/jGTjmMvKAwWrxOXf6riwU23DT4c+OkZSYdWeM/GobKzwd9sTyl/lc75bO1Cw
B511Caflg6W/6E5Fy3bSJSjVwz6gUwLJasU2YziNgd8A+JGIffAuhfZITp81gHjM
PrcVocnwkp2WnmptWpDQAu2R1K7Nr4O/cnL0SD+rY8aWT61d3uSmaqoEJd/4KYkK
46T3wiW/6xrJdvbn8nUoXoWZu9HYsuS47QQ/S1nna6JOr+smMHfdwKgsDktTPTjQ
CKmEKYUCmB9oooCUFyOHXIjWNzQd3QhRoBkOPCOT5Ek5NTcguzYcjNFZOJko7Cfd
H0Xq0G/OBA8zA5EPaM2wyMDTZ0gY07M1BWtmb16d1IRNKLRZ/6nZfJ/klbyRckjw
d5fcaZOtEqQs3Z+ERV4/Hx2+vnj2BP4zgkHlbxKfsPbOLItghqDqjOon+8B0YTHt
2+3JJQSlpePF2IliPlw9M4FBoVG/u2ILz92+c5P7u+4xrLe/V7H9Li4K9yk/6Tqx
OmJIGx32jHMfX88T0KWbzZ4ZcGNXH81xocV0Ch2NH3sU5SxKoppioU2mCo7yMcEL
LY12aFaLz4bTKsAC3pxlphKkdZE4/gZ2lDUD838ZkxwV3hbybObnFoCD2F5tqd1G
l9ZR0R2IlkK2K/uLfbUxYS5WLqwIApIKM4W+GC/8UWyC33aqDLQxstDSAWO2SOPT
7UHlEfEaxxyyZ3M1tnHHOa0FZ6FYf8l1tY+JPCZThMb8NnF5x+5MqkAUTU+4IDnC
X3+uVal+IYBmVjMtaOIAF3iV7E4CuikS5fWYfnRWMzJAvrdHaNVzeHNfDPs5o0tp
CJbWheBbXZsi3hmK4JlKm62xKvOakCDbtQtWs/Ix6sNMErsV4LPAA1GB5sIMQMLa
oopFNayCSQsuc3BN0PbOWL3puDZWms2wU60Gnue4k6imrm3HGNtqyuQ5hAh7p0r4
FJvbuOkNd6yAT8PqCuChRfwEOrBXeAftngP6ApXAvMpfaAWSIQSKZ8WDaD47Gakn
0ke3Njo/aJzlRoo6a27tGfetwseU++nm0Bsr+RgLrgm4S3U4rBNNBET3ZhgLuU/Z
zXdkxOVICDw+jmqxPL4w/U+JY7WQlan52H1ImCM5VQGlJNiwcf9YvR3T0n6kXdQr
/wKn9aEsWGyZ55u95Y3ofZmEWB2Lip2rQLg/wef7AdoXCsRhxokXi3xmQqg8NVM+
2Ds0/X3ufCFunoYG9wRCGJmbnrlvVQO68mcQiUhWpLuICjma8kHAcNWvQamnIfbZ
jyxGphDSAX7GX7a6OMMHn6FDckKMpfSIGgFuGMnHewHK4TeL9dQSqcOyrgMREf63
JDb0ObuPVy+7Q+is3aSbRp1CsS7lIBItNYqNKrCN3HI9qOzL2jLMMOf03tWyBDhL
doW1ip8DeQFyPWn3ZUjl529IQXv0osikmUMaglfYJhayAVE/rwQD4D8T7tYiYOBY
3klOH4wcIBijY2hjQvR6wVnk/YxSuz7xEcIbGiQcdVLIpW4UYMaljfKYIuHXZpH6
Cw0ht3bSW4JoY6lJV/pZtHu9oFsima9xWYh2fJ/iyl2gW3KaJK8w5l2fWKmTipAq
rQ1hJt6r994lkv3828UjExvCRW2zglO1cyCH+tUS5VLqdHs3lHd2Rr+/sFijSDLB
xslZFG0Yh6xTGfV5RNBPKRi4LSfi+sbXEHksEBu68pDw0Y3Es8te3KZB8JvDR06D
n5et/P9w6ekVC2XcKmf4tAhQ2H6ExRPm2LfnoT1WYmVq+GNpr1h9Z78Mel7hNOTv
k4nyTl7oG9glecUpBpGbfxBsTxNneUhhfjaMFF8tub2KNRElkJ9aaxzNdu2Qfp2a
APLAgQoJBr36XnVkulFYX+18pzwQPq1RsiXfzRXoXNn+/vX+W9dhXDZSxNFnVxN4
L7lr3EWK3ZWCw33NY7RQgXq5pTX4BQdCVbiUKPVAwdGZTSd8pA1dSx/bWsgmdKls
HIol6iq8qySsP/r0OhE7fi72yMoVG9TDwqx/+L20P7j8RLMU8ttSDaSwLwuJ84h3
nC5Qy6hNXN6s0b14H82hMYhPB5P5x1vW+QLNOChb8hZAEUUHUWtetrqyHdAlEI7v
gcWEtjeeQD0D843G0siVqA8dpv/IFb8GN7UmAAebZlzy0OSXuEx17IXD+ddwxtYl
KO7U6xGZwLEWD2TUkrRxWbAlSy8PnT33tJ/wpXOmdG424fobuV6lMHND37+tK01x
KD+s4kOvas0b6s27nOvinUqAD06kYoi/oOf+DxkMsigK8RqPbCPT29a+S0+bVPgw
htnAWKkiqq0y5DcCj+PgtbaK6+J79UN+ku14QEnlfVTnyGtKBqfjY8zTKTvwgDZM
PADEMlPx9rxUE+AiCA5pY9AXPPQw2XaTNCOgy1nn4OS0SH928K2E8KwsuWSpMGuy
cbufAUhIJ+syyDaXBSq0qkZE8YQAsucFdp7lkZH6lNebJGLSgj0C0XbPo5pl0QGE
3z/uoBZQnjnJNOztzWNrHpkrZMhGshNjL7YUvBtf1tv7u/EYIadSP6CnJ2bRVnQt
kdPrTMyoBRbiMD04PjgyfZ1BBObFbIZRs7pmGpFeH2MOaJJ87Q3R6C+WUwngZH3Q
hETFUMNDfC9nrlv6FE24baf4wFUTxxGfeu9t+9RGjSOvLqO4TxiBnlJZWBWB8ME7
gGDEopICahTwUTqRMSXjnoKdOvt9kg6Iz90ox+QdfVw60yNmOadA+ppO2vIvhkCd
vEgqIj0ktuczZjcDZi3k0EZCJVQ80DK6ljyobRPmhvUS3Owj5coPKqPb/G2q94zl
+546+xrC1ZDNdL4Beawv6H7Gs+4q0oIdBFGN/Y+UsG5mWaa464DfDtKyGAinkZQR
+mBpnVFVGl1MEhYxHrthNokFr1hFqzxhYHyfJDzkpv9CVObIIqYORlfJxsvt/BKa
8pmdakcR/Txa7AGYmkYqFEyrAskzvBJ+6+xLfSVB4bs419jZU3e3p7UmoBIrNzwf
2aU6BsDdkdanj8IwbK9WiCt6bxNGtNR2yGnkzGC6JxwSGlVl1uZ3DOeiQzcMmvZR
b+/w14ByPaxVJGU4OFLbjK94WMzlNXAGqQs0sk9RHJPAraAXQQBqL//rQVba0Pk7
Kw1Z8vf7S3TwI0gIA3jlfQkgFCrDjxUeEUGMnyebuA+3xDRhCNCDoHcykdvVs8RJ
cRkBzTq1/GmnK+BqcdaJ/Lb7Id7se3R8hHjebVmZsM0Aoc4eFU0Qx/RDTsTt4fT1
NQCSmra5/5sEeM2mGqJ3Xua8pQWB/OqLfAQALScVsBCFdk3Ny3tkybJsuwD7Lpim
Gp/a27jDbyf9JjueJqW3nx4W3WSHcF5OK7RGXKheCiDFkQJ44KJV2qT2E036Qxli
qH3Gl/JkXPwJzxnUTtOTXTH6DArRtMuPN3JWcf98rLM8EQo6aNrxNx1m5CNGT8az
x1L5bHh0HjwHogfhNqnwqv9UisSn05YQm/LilMd9KLvvf1jgB1cwlpqusHjScAai
PcYNhoF31has9THKmoOiKKo0m0FdZ03oGW9egGE4jz9nQAVVxr93U/8W9kzku7jE
GYpzhjsEvI0oT7q83CYBtMXDob0zs2Ldem4AwETlEumVUtn4lgYQL+xRd+ZUy3Hj
e9FR/g7mW/WM80fcyVvVqSH/dhtGxmGltFoBUO7f8WvR+91kI/m8DBMMd3Kcpe5c
JzXTrJxvMtdlfO6tXLI+8vDQulTBM4S7xL9DBh2SSOEDA3t/RfMRx9iwCqIfUkzT
SyQ6lYqtmrLuZlvjICwksoFDuy0BiDhJyedAdjwQHLahQgOfayNwZVJmfW78hvQZ
okTSlfDuS3p1r64t5BheYDrdWv4qzlS5UMbnTu98gAyOZyrN++KROQJj9ZkaUQ0J
02VTAVfRjmQGTBoLv40qZHoRs9w3P0ukd4UlLmxoQPPFWvug6JpUhQ7reQMZ2wbi
0nChvhjBh4UJI6DUAaHPJ7BRAeA2hD1eKRV98vnQzZrML5djrYFXMgMLU+Riw8UZ
BrI3VD5myTTEg09ex6j0J/L6bo9KS/dnkhv91JgySdSEXz4E2+B7m3B0nW3qmaWu
DEDPWDJW4JNQNlNKgctsmPk4uFAOrB3oW/aV6cM7PgQRkPXj37prYN5czBI8iRJW
5QNohQeUO+MAAXX20uBrm8vd3ia7DXmDX0FamR0ZzYRawbv1wF9BT+svG0g/+EsZ
lY66HMFZcddCwSseoqdrqx3IoOCJPpTdFRMI/UMAnUTyLADeCqSUgGfYjT5QGXc/
wVHNDQIW7h1JJnBzdopNREm/xYpXLLzVraOErhUdTCahLVAaQmUhM+ZabWwaiui7
J3JM4xwaOwnE+q0KrZneRMA5Me/dzxs6IBmS2DFZ8RPlUOGZBKlBa5AHh+ma45JF
IuWnc6YaEpo5nytPfO6IJyGGuXxaNQPgNVpmAkCcbvG/ZqYuA3pYX6P9w0LZF20W
hYZo76QfIgul0WcR0tNXXWrzP6yvEAilXl00TDTdxj0wCAEwwWLw4rhwnZAnx4FJ
ZQLbj24YroJF2btmTTrkeGVE1TzRN90eG5FY9gMoGbQaI6ZIvk6PB0KbQ8Cm3V0T
VLAn4SPLL/dMcI253dpx4jsNliDLIfhj5skeWTP0AsnxDyB8kk/LdZQjp/9WdNXr
+3C1ZqSAAfPoWQKzpwDuFBLDklpUcpg6W9S2QzfhmyB+pyfM3KcMps41ijr7qrUW
i4dHWzhYxVy3fGUibumfEVOO5UOzTh0bZSK3/y0bX+ExwEXhDVfve2urPPDFkq49
XUIQ6f6rLlnLX57DoyMQOkPN8SGk3Ijg/GKtP6h8/Sf7d/qyrqJcfjWwdTwVv3vL
OR94ZqPP4NeQBMAj4tg9WmeMCChVf/LRpg+VluntaP0TSosKangRAdn7wbnfRVoz
/gyrCe1U8ztaSM6MBJ+uUrEhXUwyPIVDSaTK5JYBUfYBk3FrQv1cxLwHpF3imeit
nFq4FWbWZTy6dNs6PUHzJOrkuiDrJnhEl3m+IpOSeYpODpO2SF9lMqFQWSLnGUYf
pUFsy3RPh0+0PpbukrMnz5ZmmjpidW/OVvtNfjdwJe9ocbfyQBpLCuJLsFkCtPOo
Q+RNMYrv+K9yXPqlJEGjHSx7cekhbaP+PyFXMzKlUO8DJHU+cny28QzO+AOi82ky
So4K31WEw0Zy6EJ+88zZthBh47D1IYHQc7yN+Pc7FqgQ/Pj1k+e5g6z4Y4yjQj9b
C1UC4wAvMKaEhZ9urh5xD2uPpN6RBGU6W3LN/m0sRAmD1EC/Mu08MbN2eDx95NZU
AU9GSKEtJR0sewtKsYm3xEVFYVXuv15db1lmlEpwlNfUh43dhxlcGK2vywk+f62P
Qs37aJIvdiKV+iEyKYYwtmaLhz1MFYzd3yG8vC+A7M4WiFtkaZZ13sJj2T8rO/Hg
ochEb42Da2cvEyANLitzUohDwEgpBBG1iH3u2Lia5MfqeyvoexvR5fKu1sFVzwpc
8SQcixA/MWs9AZ6n33Ul0nYL7f1oZiPQ3SXR3QSPBWIoHBREGL0ZBgDlZkGrDcN+
6PuFLDOh+UHMbRMkAGoVjDk2V+xi56dZD/tHNSMhKGledmNonr5hrNaJ97t68n39
kt4byLbmOm+8r7EQPVdxoex3kwwk9eSoX7t2lJMnwAASEe0NSKrQrZPy8BGieZ/U
UxgG/pzG+SAsXsa+boiml2NOHSm5uAAAGwgiqAzFypqwYHm4r7819OS58fP1TdkP
pbPC3ryKVMgz7O6KGo8OLmgwshQ2xvkoY307dHP284QG6lhdIOQGTZp6xjS/0waU
jtdT6ZbhDb4kKpcrsa9JCrMJuglQzIbg8wTCdj5m6rtbBsc8Y+snLDR+IKuF81mm
uPVJu/c6o8BkrjHuXQsUsWAuOdJT6fCBvXsHANciPYrHZ/Pg0aX5Bvtu0eo4Pgsz
B7LdQs33HjpEGKwgH2j76fQkTucZphb5lphJ+l1Ecuof0UDbDrcTS7w9mMAQpeVi
CjHdQezxM8MNl3w1nRyGA1nbaeEqe5wf5c5/OAOPSJjASOw82slr/dmpL2gkAXjS
3kx9wPcqwWYIeOOCC1T7xY3TEkeuUz8aeRbBT9KwilxgGeQ103/SVGaYmDHms1KO
GchC6+eSXYL7HQeGTyIt65RQDu1a+mKUgyTDMD6J/+d6Syzm0z55k4IQPlvvarkl
R41ir4rV/aXJIzRm9+ae9cdYfPEqvbbfQt2GlV9g7GBu8pD6r37lyrC4WFEdRjNy
CNceJoV73HheCTsgp2i5ClrdambFD2Rd5jDsz087s9RIRMKsNQKVoN3Wfrok0ueP
sAabk9CaROwEAEGz7mHMjcmBx/ZmvF4UlcV6u5wQiDfHBxZSPfG+AcprcYPaUNOE
bAbVV/6m6DvPunA3IyuDdgl37pTosN709fSMGxRDgqoUWS5trOryVpYolFz+MU8C
unvpOAkIhvrrtiJ5ICEkNpEDMbNyGwLb5fSBU9chiWgBoUF/NV1HKVSqisNWtzWZ
UqwfUqkHXUNsiavCiPoOR9zBEjjRBITOZ96m+X/NXIBjF3k7pTQMdLwxf8mLkNgx
ZcZ1oFO1hGIMuSadOXouPUB3STZ2/k15nPgv19F/HXwCMnouNuR9+YXX2VFkarPB
Fc4fXJfmMPYDTepCVjRWFlVFXRR55+kkx40htLT7m+0lwK56Cbw1uQxAIgWUqFYr
AJY1KfmdIAM6863gNdUwnYNmUWYYZGfVxVWhiCCRuyTUO4Kls6sFUIKoLvtxpO++
HNPQkoW4HQ6OPXedY838GhaZ59EHi1YnEBNnUW0l8+nGLNAbt21BXgind5a+keru
NVsUId3XNh8PXGZ4RJ2EKryOVuVfLaHT0NquitDGk3cJ7Y/jSvt/Eul66uDpEY3y
N+qEf5bQhQIbfiQJQWj3ZhVWE/G6aYhBP25ew5PmIvRWrZvjlP1cVC2DOqYj1pk0
Mz6C+20Ey8tN4HKHvXO6+lx0JuEEVnyTHOs4HpFgWquwc9ilxdo4urIRYiTxYEAZ
njzvS1pDarkd80KAdj8BT6ekjVfC+mqgUyQCzvFq+rQfnl+kZXO1hlHTdO0jlmxc
tJLqgREKSEA9P0IuMCsLpR8n2ptEf1H47RbSQQZ5hhNnG+G/2J0VI86uG1ubsRXC
oQ+1xzH6k/e7+57M1iEV3pJRkCw817ET6XgQrzh5Qo6e/N7h7M79Rq75dy/qtFhz
u3KaXNmhhmWLkmLBMIhX/XF5OqnNutbDL823bC/KRCsPkozO9chpPxOtcm2FdAxi
8fmcuF27X2SWUD7v3iuJnN5myiuUtLiRecTaGkZvu8JRPRq7/xwvJzvN7+yxlb8J
jG3fsyNqExTO/MfBsSRB+cGf5mEkpoxiOrC2gGEzGg3dVraj39YIcdg2HfUWNhGH
POJS9m7cnR2yHgAllgyvWPHLP43aRDonKMFdf9SCS3ml52qMar1KdNKaLjHVoKxh
jNUfzLLdLUgILurUBZntqC/6qtAVhkNvDABunWSe1O8CoIJppNz9sAbUmQHwHq+D
juD+Fi9QE8Wvr0LJN5aD9prtBu1hZIx21vFoUhZonI8riRvuaTSUfu02zD3HZwKR
R9DziF2CDwaz0XSuELrDrY/QVCNZABZfyazoXXAA41FpnKLqLOBlmgQejvY+kcvK
fCaVJXctksIXO7L6KQxtwxOipHcxGxpTXvaEVWU6mJp15Bim0U+RoKeT0EnkAu43
8D/XindTinVMuV3Tf65EfAcxMjZAbtg2jp7wxqunXCAqCe4E+t9w+90G3ehd92BK
+NmWqYMkCN4MYZXwpB83tyvxXz3mw6Vo2W10gGB3zRoxpeNlaZb9EbFvjFF5Eof6
9ZF+zwIX9EK7DIH28RL179B76IlW364C4jrTfdK52ZCA2rZ8XZSwDmXe93DTrBbS
QUOpL63+EM7bzRgtShzRmCh6OIuxFlWOtBGvA58AAJ3B0dW3NxE/zpddFcbWC7Rw
bt1VRbFt3Q8AhuEmDRHwhCy7dheReGyiG0UIKueyUnfhJ0Gvu9RzCrjnZblMm0PN
yf7gQPUGUPCBCEFrbmPAU9Wk3R8WF4q/8gZA66yVM+NiiBjGwxuZGTr8sENqup4/
QIcgewtuOdf6/koOiliHJimNBiS08EcTO9VFwf0G1iDta8vIz+w0fZasbAT1VNXx
T83IVjliVcQ4MR0b+xL8+GMJzpw3SSGs1vHvxIhq+CaBwnVTGoDBmbjlLEKCbzf4
ip/wNgkbIJYJqW1fHYtps2VMbeOhFwk+SsnYo45yoSReMuTZ94ZTfjpVH8JFjLmL
F9u4D91pKn1is8pFnqzxo/1KqocpssWrYZ68UvtHlbxBy9UYZgFY/SqnfzxTaJgz
i9eyIFI9m9ZvEF2NhFKS9YOzSprRgyy23mwr8dk8o2obByYIgu7rt0FKtP7CYRRn
yFYG+xRmqiW3OqYnODRP+s1/ktrxBOHFBsnB/LY0ltfL5wzGuNnXfiwTSSuB87jG
rgawBI8exx0KE6wOznDfeX2qNknKimKn8NLPZ9FDrCBojGUv498hy6FmjnJGc4l6
n18BzvdK0fGwvxCoIIDHFqT8gDp1TfnTeVBf2b3gST97WS18xC5KyXszLZiR3x+2
HrvS1qq4DPJjRzA2YOMk146muf/00ZPzRyoQvR6/0ok0uKAYbcwMZnCfMMTe83tj
SOMgmJ6HaiiXRC7tbhCaRZOLanjBsJJGI8PiORQ8iVyS465W7bc4iYz/5fpZG0S0
WxqVJCFFpCyBon+xg/KcOjrRyYx5oXRU3IVfHjkgi7GNBx8waCi2d204ETzxyT0F
QsEkKsm0Qy3f2k5UJ0/Lv6vp6MiQ7htU/qYkx+9Z2m+IGFqjgUwQS+TXrTYZc2++
VzV9ZWelH052Dk3Tv6d3eP2CnOYt3HEVChN3hH2DxD+OSczxxTvGTxLLKnM6c/ku
LVQyNRK+wKd42lOQRsj0a2nsxGVyC7SiSjSM2djDPMhkKaba1l6DDL6HKLxoBsMg
C2bgg6RH9YPSEvVEAl59BfUqSnkWTs9fxY3DH+n/S8MbFHSvo40BCFv7XZN5zN47
HgMH/Eiu0IwGa1HscTnXW9dnWG9Wz3WXANxBxBwWmJvEy0FH/zC69PcYFcXsHzzs
DtfF9UnBZBFCZpGsKAilxt+NsOu39aufS9s+knNu67eiBJV8Yz4sm/xU/kLUf90Z
loJ3NQjdhV4ykn8py6baPCvWO0u2JjYks8uSlBgDIMwFEJ5L9I5JeXmloLfGfd1x
Tb7nCwBBsNqAdBuabK6jatVeDNnoVMPRN7HUQVrkNnbYP6RlgbX8X3ZeNhF7x+yW
glwc1ojGX6WdM8G/aX2D4BlptqAo+C0kWIONwyYzlwNeoAD56Yi7+hAnk721hUUR
7XNsny8tLnoz9yZkKZdHeSJ2TLRgkeev0rTpYo4EB/vZgSazrwgsBdgUxyeGiO7m
VsU1sCrB0WDwBUboSfIaTdzhKz+voCQ8ifZq21d3Eug4a3AQP7H2TCeE8g8zf6PM
B9/YNlvB9EdIyqZmyidwfKIFxQxDfi/+8BhJTpK9hOFL1PM0YF1b2r0wzPMBmm/k
MuOmLStBySU280QwmyudqOMfozoExxpbC3Fkwr/Zo/yUJZiiwfN18PqDwWWavJKo
QFBv/qcAxpbAjmViONHwBoJoMbQtTk+41R+FSu1UUblbYsXPpGdrFkAq7qJCU7BH
RT30GO4iFDEhcUeHIQULOxGI+OOeYxJ5KfxUqpGMNFcOSF4mMZNebmTVC5/2nuME
StKIIz7MWRCHmh6cxwx6E2pnNiu0lgbi33FVhPcz8wRtHnUOyTqPW85Nm7pkR2B6
0vclHaa0RB7nac7X96q2pt//s+XLFz0Br1EiLovJS72Fm+JSSzUDakme1PaltFRm
lZ0+IGhTl6jTEscuJJCDEOwt1LveqWDDgBuuJ8b1qOVhTqOcYmXdSR/Jkx1lelke
b5HQIMdnbGgIPrfUqJs7kCqua55NibM+vCVVPt8vGG/X1jH83LSIdNrEQnpNra3h
uvX+dYuglv3kXSt1koLqs1QJLSaZ5eEopBDp/ylSIDBDuFJCLSjTnWOPLUoWMQ8+
ebvAQbpUKa/o+4UEPd7YraGSkVD1mWPWl9YIJpVKvaKBSNEegNFbdUF1mwp7GrLG
Z2cCg/29DrRJnlKf1oEcDZdLPfkVIClxIDOc1RLsVmPYEiW5mmCV3unSuFSq8abj
M1mmCqHTJsJ3JCFTdo1uYx2IIjyROCWqYJmxsTI9g4prKo06tUhoqj1ewY5Pzyi0
FWOX4prZV1UhPSKhYxWbun/iIY6zAIpDX0Q0siMyaNQPrRY4Hd1YjlkpJTNqZA56
EM/lYVOQ7YinCjWPBopTh1PvdPVk02gTX/FgUHCvd0ByKbT7dlWZ/XMgW4WDWk9c
x05mHQcA79iL0HOPhwtnn9L8f5NqBFuFyFdyi66F4e5iLhntK3bbQDgJ0NPr+mBV
J0Ak39yHE5UZMTu7ms8oPp+5/0etxa/d64CrAWFbPDvJtw45TYye7qFyZqZ5LvP9
0nmiulgaZ3p80qphJ1MjYCZHmFEYVv6Zau0b5++1jbyY2u4OFg5DGiEqf5C8loBY
42CcoKjIho6IVjMGcmgHM6PFHgfsIUp4XCxmiNENDYkOEQsMHQwWxlAeH7j2yYjC
SUhvuzYnIUyShpcLnPCV1GWeJ61iio1mDvBK6T5qrRKaVmRkI/X/yaTmEMo1QsgW
re4I9Abq7EmKrBb2MHRBsWscIIZCDr3f/wQfLxwroOAFFWwcdLcZDJHQ0uqejGJI
YfjE08881xRF/jAL1Ln2qFZ8Xi9RzrnCZ4h7e3Q/CtJJ0lqrPWhzwirLBd4Dl5Tf
Pr4K6ZUBElhdq1XeF+9dkq4c6+nljDCX5uRTZXF7rbNeuQEqKvS3Q+AVcEqycSh3
am6edKoM/dwLk74xVnlHShDMEvrw+ITSiAJRUUR13tUZn/baRwG7J2ZqB3rh9F7W
nCZDDg1xFBWLEVFW1Ulf7bN7KtwNdvudY8DslWkwEYwssWvhYYPTSWAICYMsOKI2
g1bo3UGXRjVRRyQc1U90PHmCfWIRJ26XEOJKpdFKaO03cGsTn/D4uvDfsibP+0pQ
R5pCOnlKp+OukqZElsoEB0JsQbHJgz0mBXqhfRC15hJ5xIHkm0gNFFCa8mT4Azx1
ZUCwvm5G43EnXZLOL7EOFFD7SNFj8dEUGebX23N8Zq5dCBw9weivSiGrNpcZuOL6
G/qU8jRnZvK0p3i39+8ZoklaUEvow+PvbF7VIUvoUjL4bftfJqCMH7afQspy8O0u
8lTob7SEaQz4NWYapcnobkotDjMNX/4FMuJtITV0eAcmweDYQy0kzh4U69jA7hvM
lIaG16BA0l6Zi5jXEFP9/0UnFNsiHeFMoaEorXHJRBeRqG2D5pW0LipMJbrOtp1M
QoWSBBQIfi1YMhTJpMjHmeGl5N6EkmtZH5KgtBTADsBySAHTJ92nRBn9Rd+yYdms
uxa5aKn/LcjrhjWmY5QOISZJCecgFtLF6fGZJwTowz1sWBCNV2g/aUFttNST1dbP
ejHTnLxWUMRRqJNwIltb8AYkHr/Hll30uSd6qwU70hjKnFIa5btHOVs0W67ae6mP
GnGREb11JpH281uhbey7bYJYVxo6Oiz0Cnc+BrzV11XiZW6xYFI+xRmxpuBxtSMy
7Oph/huom1pkEGwPArcJgtZxZFaw/Y4K/3k2xOQZzq60ylv+1Suydi9dHlbbAXl0
MpnWN6L2m32+0EqyOUA03qJn3kqLhyiYW0A0WVP1sw+ovTxaaXxgs/Ql3TJuIcJY
Ho4glIlL9seK2tYcw31LPjgdzjXh/xvuxr/BQqX2PZGyOMsiwemJqxPbCfpmgJQV
KjKUFSu6yEWt4tLr1eWmxUazV9nzzVTBqSeVJ38pUbmFinAK+vbS88sgVFFtVIYC
ajZ9VJCGloPLhvnN3+3MEAgyC5C1f4FgPLVneVNMDU5WZ+rLArZ+9akWpxfIBWFu
Yk2h+tGvJdqYGeeUzcAQ7HY0VAEZcZJP/QC4gG6jbQTmNlsz9XY49PDisEDAq9W9
Hlw71dqclwMacfe/rrn2yNiLiQFiQkw4I3CHDJAn0OdtE8Fka3R7rWVnDDTzOeyL
+teD2y/LJnvnoMH9kK/nW1Nl7sEHZCuR8rhEsFKFdbpBT4y+4WmanWwkhGXh4Yml
ujaVfsHscW5r3bdYoCL8ez04Gm3FWtnSnpSoTkiOTK+NI6QrLWxTBlkdc+PoopX/
oXUK68gavEU++X7VE+fCBL5thNjzDdOR1YvKHZrYYcLJSbEDsCr0/zOB/ypUbHBs
SPWMB3F89G0J+IiPUuhRt1bn4yHbmSDNy7ti+WadcBUrwyH6tOviI3DdVefwAPu+
Qsq1vmKkCB9qy6QjOEnJ5q+Qt/rCXXCyRvDcjuEKNcv9aqVcWBvAZEZSSAudXqUE
HyDfer5ZxnwlTCAL9ON02BTwAdQXpkYNraLc7hD7ymnXe7Ck/bgSQYDtM+4ZTKHw
ge7cXXMiieTTgtGBpO4MnRsYMknu8C/0d4GGyK1xaobGBZHkhLLf9MUC/LNy1QBp
EHcVNwR7aYM5LM4HUgppNwz51jyqI4CbB38EMUlR+aWYqyZTxHCThfuEVAAowgOs
ofok5aw+0k5nrdFQu6P5sNxqIxapvRy7CBYNog0B9eRiyNceXbhrq5wq/QPcyIvG
Ca4DBpAfPRLirf5B8ezRG/rIuyUiEHB60tJI/LawOjfTeMQyMY03a9goBuYhc05S
hMdS4E8a9DkHU3+TVRLtS2K8oZH9Emni3WaqMK0TEz5Ek80GuUmK2FGfcwJHTHTZ
ra37UtY5LXHdQ3tksX8BAS0KTetjI8fZULyCqCRNbqpWooS0GJsNBbKIAPqh+Kwq
LMFHxyFryy7CBDtGfgGWBvkaPN74n/EPXcQaeMHZRHDqZEOdgZhk6AtVTWExpqcB
T9TaNkjDHENyfLaZla2tE4Knn5+6uLg103N4ohWloTf5ZO2kD78rUa3aMhrnaAPY
iUpciTisnFIVTsbykyRPGmD4EMqK5DOgqU7qPaeBg+ms7pXUum85LBiP4+q3NhqV
6tWfXks72fTPyUrGCmByD+0dFNsA2BiYwIg+uOiDiO/veGr0QO8yPdhS6/c7IZuZ
ot+/ksQEQJufTwTNBJtWwlhGt6zdFeYxHLw7Db/BizcWH3CYOfTKEIxEn/NeV/zW
C9wPI2nmMyvlZlG7FX4WwjZ4jMj0rFQe2g9DXY4kxpGD0LJuk7yjmF5wJGJaDLR0
mq2wJQZl2t8GWZjbcOC+3yMTvIM9+0uOIqHjlr+0j057kFblY6X3Mxd40eKIaEcl
Gn8V+pHT9DXNgqQWHDYa9xHVih0ESOwoYPc2yiNGqeFIZsm7Kh6DA0LmNd+hyNOt
Skl0FaNfQs+MtWs3fNTCXoPER+jPtkhyuDNKXb6fvm0Rbj19akuYL2DHDoxOj77w
Rf3UqULdk9skbSc8nDu50ODt6aIBxpV/wqSpP8GzzcFcCggHDDRIlAl6mcmSw8sD
3E5dQWAsJ84vpDGnrr/3dKTxzQiYxigIochsh/uiinnzAaNy12BeN8RaM3Z87H2R
dInH8NrZ/PXg4HsJbVs1MGsSYw3I1lF6MRz+pWGdOxmKHK3TtUcZtaypVYcFYNyA
1CcK+ftjXuIlTfQdXIOkHsVU9ju3nX8lNYdDBs1qIQY5VllBSY8p+K9aDJ5Bt8gw
4CslQyj7ySuGFk5H3kA7LqXCdQCHH7kiWCTWCUMClJq09KI8HDSZLq4z9slUmr3m
gFTql2dAeR1gsMQquv0rOk/iMq5EQw2KcPB5U+xuNcIrT57qjtx5Luwt5+Dlcsi2
uRkZL6cjzUg1srHEx0ZcPwtjGpOMOAAd56b2Xbjc+CvwQuC5wPhW4gYu91TjC2gd
PTFVM0aJOFLeQ7qYcpPrXz8aC0AFtc7J2q+MLo/74cELWH65VN7UwouWyf1YWKeR
S2is8YLIYk+vf+4qbfv2FKAIguW3ftfwPEvr3oFklVtI2AFN9BgfTkipSD7+wtcW
CO0I4klgF8Gar0QjYwithJ5WpVc9BXmaRhus0f46XNLSK+XRglvYXe3tYZG6Grlp
dM6UaF0w+P4rhSzbwkfAgckQBMweMTPbn8AKP1wj/ktSCthSDsu319EiJF8fJktj
mcCiOk57M9spDpb7Wm11bISc2Hss0AXhxrgT/krf2lEAAePQXQIVb8FffpOoI9YL
qZ+hFhVNn5IpAL/7M+4FiNam9FzxktbF/0Kc52NIVwRW8m9SCPMRVufm/5oUMnsu
ivU/VLw5b4VJ/c2DNipOyyrylI6cUvD5sRgiceLJWUMCpMns5DmGgfU23UozPLMC
eTW9H9OrWOAQV0+BjC8S6Kc1Y771iTGoGVI4j4RJ/yeRFQqZ5PYQGsqhpV7Yz5Af
N7S4CMUVlKTe7fDIIB/8dJYKHlJT7Sv+bP7yPx/JjxeJWLx9G4St+JnnwO/gCz3V
xQMAxCvjPfqtL6mrspt+M9/V/uG3UHisEuwtflUNxQjbky14zqW2uqCc0XavC7Tx
whvMRe5P8sQxGJVgOtMirKrkhAXBS+jo0EG1ZPFMy0IAfzNl/ypExkUIEibf3zFv
z2uzUmhzR6uqo5bHDj6kbFp/SCtzVZqxItLKcnR8s93u/AWE3mkr0IUVdDAGc3za
eGF8xRLEE026E8XBYx316p/RKqcCeljl6sTyNg+4n/XY+tePBPrkTeNcxwrYO4Cm
nnflpI+6kZscFom/Ra3sUa39qG+ydz2OzqeBMaFhHepISauriSCiTq4vi8AiSFr4
aX7Mp97m2b4riSPMD/UywbTg1Mrlvh1Nxmt/VmwNuIv8/RO9TIrHczVrIliyRpGp
w/nRh04O6ZdF1x7oQXoWas5HfS6rHMy8F4IN70iA7BLmC4WDU9mNphGiP+6BWys9
lm0F9r/x43JrxH6tRp9Nq88QyCeM+uLDYEZW36l6ikTjbBqAMUIF2TM06SAQlexV
FWCWsJvE4KOx3/6sh7TADX+82D/oC4ZHtHFkaR8iiGKOANziT6XSjXDOgxUxqmZ8
WAKG95BTVdePu8cht1pif6FP+nFZ4yxBtvLblDwUz5oxyk0B6PeIA5EBJ6yQ7ToW
l7cRkR9JITQyDsZgIQXt7I3Qcq4SWHLR/YAQWI3BV2FKv0DUGZ1Dk32cjJrmHdm+
0QgtXP9eKrohXo3/MgDXdCnKl+7P1NUbTOQxMLEVSic5z5Hq/hDo69NkpJblPxdn
SYZtGUlIeQxsyhFlQhzV9H+5Jjdr+X2bgr/WTADro+RIfPbmfqMHunFimb5ImnTx
8kKvo/q0vjnmkVu5koY3DoUYMSBuhHKELAaFRIaYiV15JOCaF7tW9AVbujMsjT5X
oeEorxIgG8QLikkRRMTKaZMxEBOup5yl7HkKFRv0lgj8xCuAk9OEDMrpUy7btvDO
EUeeSHcIDEtWOP5eeZd/5FFnQ/FnfrbU+iS2qNRVsd69UEDNAVCx4kglqVtFBdHG
q9MrAUwn/w+GKRogLg5JO+QtLijrKQnE4i7s6+uVyoFS1IGQwnPudvCKHI6jv0eE
ql04DUIbsePbdN1aDdTt4892WQMQYcsxwZ2b8ot0pUc/9akSTLw5+T4tFXABtvqP
ru8AiL4AyIAhVesOagpOUpaf8ZyplGufsF5SX9yjjFteS5JlwtRxSjN5GrnTO6u6
L7kjGOEaTCVEZet4lZIo+I6DezowQZI3cWnWrEr+f9eXEjGy1diJxVy1IN+zATot
1gQdoiUAvSS+gTVmCEDLaW5AIpdydU5sVLcmUtKUpdu3zRgCs/Q7sxPA+myY0jvg
SYqh7inFNOlWi5nIGkm0aGQS4RR6oIM+l5QmEEngTvoN/AgYx9YiLrbsAzZ4D2qY
IWW1lqJchP9wtKrIfy/p6WqsKWGtmosuqSy6vtUHwqDkIPD3QzD4IK5v4ZfhpeD5
AyBctXKaQAL5M2mQQynxOdVnEwMYhPa+MnUwPq6f7Tj8Oc1jfc7LKdgf8jepeiyB
gRSO4yXMt+WLmPttcZrdd0NJX7rwu0eNmMbViv7TTsg2rjX3cal29e3a+PosEhAo
I4n/ObcuO40ykW/y1r2janzW6sbhBdGeBz52uFdAA0iQQgfvSrwUk/ZRouM8AOjm
ZrevrZNbm25s0sPckrbbCKR5MTLFCv9XJaZcAYqqpAChEBmYwoJW+tNkU5NIR1Gb
ftuZU/mvz53Ar/8bJuu2YwuarIUgCYgWxQRqubVVm4acOpYOcj6HGs77IsStRpuj
Wfl3N7dycYjn8biMTmXrFc/RhvTDp1ig5zydjhZxzsFtj8Or7rJPlakwsUb4oomo
EZ4t6GD7OR6pn9sfJoT3PWYstnOmpJJ9SvsLiwWPB9vclVwIRV6/ErlT1D/tb/5Z
aiqLF5RRRqNZbaQVsERfeNADBSbsr7NNQEJ+Ub9WELq5k9hwMS5hga++C1lJBQXg
710T7bqr+JWV0lbJVbk8LaqgWhuKYf2/VWMQLg+/nB3pHAsJ9YbnHi/BXlzRfE5C
HgChtwYRVUMRInSJAXIe5MgiELf3FJbJbdWyLekbOGmQSD5rbMPvC6gosO1tnC20
nS1QHEvGjHJnn0IE3NPETpJN6mEITU51Un7HTnfALBivlQT7DGkdiPNimDfmwYBL
R5kkstHGg7jv3nKq5qMk2UA+syLyQZaQYITcPCpnrlwVLrDvjBTybGjOTF5h9Fv5
10PnJSFUyXluKqRYpXYKH55HuXYHSTG7z2omnk6yaDg7Ep+jR6Jup4Z7YvqH967p
EaIOWp9H0GWZvRWuFqFiF1Sd/5StdDqr410FrJWbLwM+BNW6IEKYzM1J0tG/c4Kv
uqkubAoPImX7uoINFEgjIkdUlPCkqpKbjqev7ACJFr0hWZ2US8/J6vxftFPwrzae
QL4RhIdRkLzkUP8Z/nB+sju2V11bHUHg95HezwD4dr3TWDsUd3qh+TaShdo4d6Ww
vzBYVsDcNtuIzEw1Nugllzq3o6QESB+UvFsan3gpuCOouhHqsPbryxNbQH1BfYX9
CHDA45PDlnvHxSY0pE7n+JZBeGvZvWTKbJE4dtZ2hpwxjMsxg0kAcPNOFqD7bHAX
6zWap1Hrj9wKcawdOGC5jFVCT602656Iyos23oVm3wmBowkXK1P2B+vyNOMrQ1Lq
kNo5Z7TL83nYzw19N8j4XPlUwM+PQ+RQyWCgrt4RifZWLvYmizEJdVZBsGK6mY4L
vOf+k5TXmZ6IN93XrfjrKixwMCH09xpvkIMGfVdBFG4d5/51lrArWvIRDMbd5N5Y
f+pkLLQDoKIgcDAMs76dyUKiMKDDZbCRsDvJOwTCQh8A7cCkkuRecO5GvdoFN24u
A6N2DChdFi1lngCZ5GhSv4yfnx+2YqlDDAifwJdXC9aMQg1gpMzfCnhkFZXKhinI
vGTe2S3Y+rgG53lcTKak0G9z0jW7bhuOnyD1vXYe3DmBHd9ydSMTPz2f0GOHwRZs
1M32FVYWNUaY7aY0nYf7EcFcfxxwtpekWAFVZXfxpk9FZhF/pIMJ+eQ44tBfvkOA
8qXpyv+yfMDVt9JC27nTkZM/HDJbuNe4guAfx1MrzIGJh8F3TSPOu4P6onLEZtLz
I6peiU4K2d7sUvmng0aor1+/+83UZrm4k9IPp3BVw0Nyuucfg618DRnpMLstkcOi
pLV1bnQsGTOI6FrOR5SFuvd/Xp0l46m6iim6mo/7FAQhIeEDKlgwhAkSU/xTwHIF
V2wdhw9iKmSx1nLIm34G8T3eumEG5C7kWsFP96OjUjtZNox207q/q+4bX7oGeq/h
QdVFY1ZiwKqQMz2+PL44vQRAXnsIAObULqj/lA33fw1MrqksQC09mJpdBc0YdUoR
BALN1WzgsLlndoP3O/cGWoMQAuXy6he18aHMXcVFm+Gxm3NmHx8rrqP0tyVIvvLD
SvKfNWbgYFPSQMd5c6NpsjfP0ZWm5gdHF15p5fy5hvg5KdZAnd5o1cx1Hudgd00N
xZn5xlOTEFMCKfgeS2btBT7Yv84+0pRI/xpTwUDn6MZZeb1FXgLcWvUF+5oQj5zY
1MwMbeTb1l5NiVb1qhr9MEunBbtl4lSRVLK4vuAPt2a+d5X1CqFCk9Cxg5P3Vg8d
zndQq4P5uC3u5xhm2KJZldj1O2nwp8AZUm5vLnNEIwA/r83jfx1M753RslW5mDGX
rmrAZapEjpWP+aisLvwOjIlx7OUG/qGjxPGuJtCgGrh29x2U1h7fLAkG3/KoeFHs
Qq0pXSIjG4FuXwQRM4rbRbWLhGAbCAC7E2LK4AebbwMcs+dYrWC9pcFsbuJVBh7A
KTq4Ex28q6FRDcyD9ZanNa/ZCTFqKIs9rF2KcAk1ua2vyTOPio63y3jkPibmT/OY
IpjE+zJEkARSHz4cihwoGbYb9p3kjrjv0YXnZV1C/BXrUsXnK8zwXtcIY+uhwkMx
eIBC4wXXrJj+5JcP/cu5MdxnhEPW3ply8ARIx0JY2S2eesT+AMN8OYK1tQFNzGWz
1/KDdjWBs9ZyqEimiWp6M9woh3x4VNf+pri1NDw3+KqgRzwl1CWoJow6QuT2MEc9
0nBzMVQKjrv/MpCx9cUrC77a8FruSTyidID8pD0H8aB7vK4cZuv5OqepSGvkAdKp
PqgeIvSd56dAX3672B20tYIXjle++xP30yCQofeB4roKBscDbf0bBGHQgyfFzHqd
7HO108hkM855qLi32T9yfHS6Jc7Kr9mcT9EvRvJPGt8UgAiBqbRlOJCqnYPHQzU5
MW7/BxVkOnyQ4vyZsj8Bf8I/WU3HGr5b1bsfXpB7bRMaL34Q/jZyRksNSFG1m6wb
By118nsRwa8q9ZiQb/68w59a9GcUGRDe6C41OVpVc/CwH1Hn8U1Cj/VNnoz8X9FS
EaptO/QjWVSQNT7IekvAGcEe05dLksV9AeXi2wQyqrnzXxbJe0tPQ6Z5aSi+ngc+
07M6DFKiWER+ADHOPj0DUNo2hRJ0/YweGqVKqRWfEfkrVNW7WpFIl/6HqhtmxpjB
PbRwsMMC/yJ/qgBOka3PfZ0D2FwvqfSmUMC9xIFz1B5y9PytzfBzm3HuIpdy+k1U
TTPcPRQeNV9qHzhwvtcEKM6GKFWamig1ADWDvALZbhyudqoBWjFE8908QWaHpHTI
oqM6YnnN6NrtJzYD6cKROblA3U/iiqUOd+aILdSfwxl5dnbfyGur+bZ9PHnvHzoF
39CWCooSU97N+Kzc01Oi/FOUjiBl3v27X86CR7gBAKVZGz97E/AvpJfp9p8k2PLT
LFlWbKfeL7r9eNfFcao7tvpSe/Yc8O/aJYepky3FDyk3Qi8ic4+jymxign5mjrK/
cL3TUgylgCa1tMIK39NsLpDOhK9hB/BKdXHbH/HBpLvPdbHZlPHzhfSQvccgJ8m8
Ee8zwROrbLdQNRWoaXKGjUJJcnb4eyCvheSYjpBWxHDkDOET6EaJwa2juy8jwdLO
bmnXrW51CNoa0TUmiHk1NcXeoSS6TlmBLWpfnwILFfz3wpZ/mtuuAp2sR3UhX/OP
EpLrf0sIrR9V+JzedN5wNWuxIWf67HIRvEhZaNtimUMgQ+y6OJIvwdrAHHqVlibS
V3eZd11MWC1OjQBBep5WZ3e1V7YABVYIWTdUvwFtfbUyyVBg1nyflXc97ZK/zybR
IlBdW528e7qUenLY335lKHyVMwJU6y2wpjjDu7gUFnyWjXtUP+Sy+BRnms0cp4Og
S9AvVLuuKvopht4WDy60QZyeSCjE78gD23Ibwg5blAl07y5zFfXqAQzVOGw2zW/W
VefbrMkHV+5wcQEKE/lVdkVluNZInIe7tHIvI2Zc6Tfwye0BMN6Jp4weOsEOZr9H
rMRGzYR1mjzZ/LI/9VIZHu4qneAU9fHkXBD5y/QQP40dXJDDeaDmaDyO8D823K/B
j5669wTSTKHeMyoRkswKwkDR8W7AlphFJzBV5v22bTEjgTnWFRIedxepUKAR+0n6
2JGrNogV9XXBokgCgHC1K0dnlcrwxvLIaNDRQ4J1RvQSSiPySYRkgRy11D2aNwOV
r3WByxTAFvIbLtK05lYOukM2UX2tAtRq0qAp/+QP4Sd4JcQJh1vF1V9RO3WetBjr
OGTv4ZcfdcyT7fdW78EBIKvMWaDimbV30ndJ7ERzULTkjd59Zibv3FLcPc6a8WH6
ufP0gT3xHz139VfPlLjuqSOgTXjTCxaW7rnD5Gmg/4q681oWI7OGmbm6MWt84qTc
2y/RCxrdHRtA3vsVMq2xzvJ3Ege++FG6r8QWi7jKTL23GSLhNtcSdVo1Fo4OtqD5
Rnq7dFQgaq0pEqqmJ1feqYu2cP0PN3URRZ2rEYkf06YFsdWHMccJ19jhEokONqoc
tWlm1wdp0HBVH6653qPh30GSTkY5KphOaFyPZN6SZVlq0Osrgm9dVsydCWXEPXcc
t3/8+IMigHbpucTUDQmB+9fffAk6vGwbvIuCgdvt8yPBFmdQB4DRGCvpna0snpL5
m3cXdL65n/1WpAFptmom2ZUxpsxstUo3GtXzpdplvMsymH72eoYoGQIq3QYIvvYo
7zvLLAs4egv/KYnhmh3Y33moqzIfoZvqxCuzHDi2+O9TG7VhGou+YSOesizPPEz1
EqYDxtMZbJwNKoYISeFKYpeK18JwkvUHPCPTvdQ3t4GOZCkSmmA5FxPQpxCkYaoe
B0/mxNBM+zT0qO8bELhl1qfPPLj8bxDQ03Z8oNmWiL2zTWIxiJyT6uAcWk/Q3G31
aAslIOM1hpogYuM5czmPdXW6oFBC+NRE4N3wYwLYIv0Bf5yH8VJS/vdjOAXH1Y35
LO99f/FGFoWnD5pRfPdGAouuUksGxKfEfd4xH3lppzU1gJPgIp4Ty2BPd9yEbO93
XMJVqayqUfGiJwmAQCcIzu4cU1vB6yabg+H7PbQH+YR73ibm58YjFpAYev2z3R4R
1cN3/TG6rw5tsPdtiMKsNJa56QjojLlhkgbWiNac644qcB+IfmFVuEP4+qgaCupo
YAoPWTYG/4Y9jWcOfvcC18ivBhNXAn+EIOWSuR6uEk1hAHzJ+5crDn1UUZEAzMP3
ldmm7D4kjWcat3YG/PPD4mueCGzepzeDvcVX74vvt+m/K45h1yBzmaKk+X8ro8Aq
F7QCiTqaWl7f4ydIOoakflUypcLG2MDi0TefmvM1ee1kythzaFkowQ2Q8W2RzWaC
FCZfpxcGJ42H4vM/WhUkgfKvvZ7/SkJFSiaWIxJRf913StvUT2O814YCyNU0Gtuf
3jwXCD2hRKWPPSD17sKVC8zsWTxjdehA/W1HpX7QL/2VkXPMR0eY7dcgFvO3BllO
7vZiRYlc+QUzmXI4iDabe568vpqi6Ak2Ia6BXqJvtABSi7xhlSm768PzNGUH+KA8
Nc15zZE/PjgKGb3RnKNW6bb47k7qzGg/TXgGheXdJ/mc5kxB0seQe/O3VjOvUvXr
qYJE93M6HKM4T3DHHKYSRPD0CpLfLLnFLGLnd5BFiOsttxb3RT3boYHwylh4jj4u
koDK4AgGtQTsrDIm7ubwVqO6kVgai71ZM9KuiNqQ48E44fbEnoHG6LqXj4WTBb1G
aeQsQbhB95iiiLg3QvgNVI+rJs6RF11NuxU2QWnUktl2hLYYAgUrAjGt60hmWvbq
yN4+h4ENBz5tsDyTkvz2qAF9hWUrl/93tiF0/z/A87kPp/7flFTdnR80koSJ2QiJ
+zPmpNVNI6IANZLHa5h1sW6vG+mTLdsURmtrGk068uOugSHJACtA+SZOlfQLZnhR
FK0fZik4sIdKE/XfRUPGSkVP05X5f2QLjlMeXPHoElSEJuULSv8B/A1+ttABX3Jr
MTrbcKpOL37nE2hFxzZ2RBwTjfPjouhIYWSrL4lb4JuAipcFtaatd2qswQfdKyBd
nHsSX/CU4gM2wltI+GgV+jo/dnw3PMDLmGcTRZFNQyL0ESRd3hnRTnOuGjzPranw
rSc26qjC4qJ5A2YhzXQxN0E9toWD8+/fmSboal5sOQkV1G5GgSPDwhPC3KSUAzSX
M1EXAyjGYgb0htPoFoyOnUwEAC4FeaoMh4ad7PJSX0vR54u/X21W/D2dkydnyr3z
PDA9NpuXRPTjOAFPWXajH6i3WSYuKa81N7p1azKNYhC9hEyjrmbHHwY+L7eS2UsF
a7MqU+8rmnJ2Q6LpxfmKOGhVu5Pb54oSryKoX8qggLYE2V/8OtJ2flkZkOOUZnrI
ccBxQhHbYhuva7HnhmR90OT1FJaGefv5l8/AfeiBPcJld5cs8IKflvSQvCseRrCu
k5YlqEex18OcKcEcPq5UkTuFipLel5aSchKObxGHTUyX6E5OYWzIkAbsdwBcaULV
/T0nWWyRu342dgzdGvngZL/SZ8UvUljrtE5IEj+PlAipFoNWuCC0QYnbITZSPNec
L6Urrh1/6dKfv6aVBrDptOx4m1A1P+jDCOVDd8s2PjISzCp07hKPUk5sUk/g/pUM
RKXWsmHIWJsd2WG/KWHcZw2tEdLlhMOBjAZ1tnL0Y0p1iiS0sPBoFk84G0YnL566
MCznXL3lPsVTFmyNY55V3kERS363qVWbBuSDg+ePWPru4YNCm/OG7+7BVk9rgCJK
l12CzGzpbTBdiRgjYJ04okKQWhVmBop8YJtQ9XR3Gpgf5pEMDbUilYqZK0MQRBkW
Dhp9/4rNYhI6kCpkF6YOdCuLcA4cv8BIgCqZY7M35DsET1mSdBK1DGdWQnSk3h7x
KWtmBlauSLalDdEaousxXDLMZO1hPedp3515JrVlKSWTpkg5vea3/12IGveXKh4t
0glWLEYD/DccQD0MCt6XiA+S3xJBmL+vrhWBrOCC7WIpc/kom7Hs+x5+HSh/tcmR
BbegLrr9lCAVGnS6GlDx2tx2F9/mcyXsGDSzrf5TaAxuCOdrPc3k+DZELBVXBIRd
eLULVv94USoDjTQUYQXyEQgiCG1QD2KFk/j73JP///+ZEbc2bHS20qsbR/GZ5szW
8uSj/zOQW86JjW43aQv2o1+YGuLCHlKChF5N+Vp4mADgk5ak2FgtGELmerWYJjgY
xlmBIs1LxLm1OKgBg0vD8x0o82RM3LRRhxsIut1MaOvhie8ukqhyqwLVkjAHpMw+
pQ/9/BcMuqNQ8MwcXOcQhEPBEKE6R+vyVOqndt7+Sq0mfv3m3r6HqQGaAjRnaVB5
fY/tBda+gFuS9c8ujiV8+Ml5/JVGSej9yNOHR51KWtcp0IeBPz8TpV1sqQMeXdRH
/8KZbYIDNUFTNR3lUOwgE4GjrlN+bkSUWokeMl57CN+Lui5jkZc2rnENy6alQVJi
Kx8H11KkzqV3VHZMp/spc/ltMZ08aMBWkxqodEUJVBZH6hHv+Cb8mTj9Bbx+dKcu
VIdgzikGmxyIigWwFC85WzNUouEWTsIFfjlOBSQAA809Br7evjr4uPNZIqRhON+5
D0Gtfx8t8nueqqT1LYKKgAuHiRFtGlj7hHiXbXRrzMT/8tkgybwe0szx++VOnETU
TNZcvU5nZVSsfwvRTA1xwEOlCwdb+n8G/4V7u4kvs3wm6nlMSJtu9dUapOMcGw3A
Bt81oKmrbvEOd08JRc3sWvK8nRVvqCQhWox+hE307EBYCZk+YR9zHEYJM7C0pdbo
OdebwsLGpaj3+atDkq48mrM0615iRYv8j3KYDjx0YZEJqLG+a3NwcpB8KnIkMr9C
4KXgkwEuMP/Zw/3e6xR2Jn70cjCAf//KGAkd6Z0FCcEkTh95fftxRB6E9uPnF/jK
PuFTu1ph35MMf7nBVSgoaW5sxn9Bx5gyMBb5B/3sdApEZ36GPIyJtF66AaLhXD2M
nnQYMtkUGPL25KHxMY8/0HUMZFWFYojaxBSSS0GaD2D81ohXKZNIK39VjHtL1ctG
BZ4tpoKyKSNGK+lTzGVRYaKDpdBS9CJ/iZfgckIarTL+QMdqx/SBuSV0OeCl1Pbh
f7rw2lqRc0YyQzuc6w+60mpOYgJtV5lZ6A9eZdMzje/vp5kFghOJ/Jc8LZpV/Z/7
WbuFUxt3fvmKRIYeOUziLP62jLo+gUp4iwDuuJYJj/z7OzJ5ou3fcy/w+1ww4dz5
2d6+nDH2FAp5Dsv9e5oNiUNnOiNWIMS3HiHPFQcB3t/YnOIxvihydO5dpjaglt5I
fJ4Eozm/EqfjuKk103VBvyQ3lQHnKXJmCQOcDRxbn9+7T1zSVodZ6ey5LBGceza2
kAJF9gJYJFghlIjDpucUIt3aIxsXZwbjWcc6nCcTfHPbrhUY8HbAJTMI+B4tEL2v
X7WqmfQRjRKDjskGcLpGfXrJL1v8S1MvqN2xwGPgFl65WUMbFYZgR2ThAMCnItCP
eOMgpd94RhkZYcBaV4u5K56rdme8XNY1BaWmj6r6zbVocV9xd4cbq7R9vP3zUz7B
SaSujO5ZZXK3zUkDcHogQKHulr8I8cJEVzf06F5USO1Dpa0VS+fpPVJLp+dMP5OH
6XgLIjDZnJq9MC63VJdBU6O3Vf0NxJqsCjX9+y9i3Q733mTbaCM36nHFiWUNPEIl
ozJyh3Mu3aU/0ClM8rpDYNqrzyM2Fmb6sxoX/KEa7AQb9JHwn4fEH7mRdUkSUkAa
OxIqdONeBKTG9bmC4bqSrRsl2QFkLlkt62XVAoouuo/Wua0Cz+dcHeCerxOoXTzj
Nw+me+XeJbnueVC6P8K4xvQU5fQGzIHx21SunX6HevTXpaOrPD6eHVvBQU0F/UYY
uZex2rR2dTZ3llf8A0MzktHbvBWLraqYhOGRpSd0w1S1FVOgptoPUdigJI9H2RX+
2ncp75j105F9DPPcOBtSTT0g3T3H/LxmMPo3pP0q4Qmx2ogvaG0Be4VZDYSCyHIL
tn2iM2WEYBoHPr4t0/9QZA/kgl8kjP9ilxkAMZL4sXVdbWqiQYVlnUOmUCAr+NK9
sbp+xpIpuDn+APlcXPISGRHVRmoUxH5Dvkdc36KlNrcebF9qMRUYYpybGKEcSHGo
h0/qxaQ82YzGNVGs5yAaLIwyR1RnsheQbQ0eRe4Bn0XfXLcIE3QBjee9Hl0aTdcw
jGB6WxYvutlz+QBabwtMd23BfOWGBWWxQnTYMcSHuIzACnrbOU//sBaUSDutGD1c
HU4OaR6F0lQv8V2aJZMtKMQBSq5+k9RVGvNNv87V/Q7iRPHxgWtJweE/uo1KRF2i
QDC/N96vPfhyRRRrnu2tkNDRTKs13oInlpQQ2HLAupMZ2+ZXWri3VPuyg+ekby3g
73f40vaZaXADT72cgBlVcOOfyltdB5lqBE0tLDn7T2QAMbqKfL3QA4SQbfwFM/CC
ObbYkwGiu2t3EB7NbDVBlB5Is0uMVW5N+LWI02zbieQwUNyXt+NvUHd8/4BElbSo
rP14vUJOEWcPSMzcRfyl79nJ42L38snH68gv48ygmrpEAGFf1fUsaul8ZRVZORb8
mvbkLir5Mqn3S5fbBHOt96kQO/3kjPJRI/Bw/uqqd/ygCYYnD6j0JqVEaPBz+Ogs
4aRMrxegQF/+OLb9sFhSa5k5QtL4KzPj2viXo0u2p2DXTfNbBuKpGio+GrdeNqUx
p2D/ahFAikBxF6S9ECEp1COl2Yggnoxg1IidUHCxsCT4gkC9OzqkTF5IBSutIQ7q
AgZGpwOHuew3kDWNYhfplcRetSHt7Vyx4K+E/bwALTOQ0jGvHBI15Zcxax+Xk0LL
mQr8UJVis97aQmGRb7QnRtuRRwlxI9cDBcdp/277CQCj7qdU28on85UlPZNsiwNF
DmsDGFZGMBqDRScPUPI4N34ZTTNrEm2IUlybwy0kuQJRKOe5oZWM+tLftMTMyBsA
2EJf1eJd5coDLvsme9x7PYQ3u9RMntwTjsBBOdtenygN0AeRCVtSbiF90LAxCJia
q+oXBTkRyiq3BF9f2sE69cpzBemUaEHC7wjMrRNb62tPA7L03jroOZrsnzV4v7qp
CbCaHeo+BVAdqize5uUQxa84BecE/fj29G0LkLj5rF8mS5pNXreCc85PBWxsNNUu
+WJfc4AoZp9etkVyvteq3qit/dna8/EnnOplJD+SLhfINiQK734dvrb7Ze5v90ma
Sp8H+6VYB6OyifCDRpiuieLYFLc2MM/bi20jKzaxB4WJ+j5c8+5gG407t1TJPHZZ
sfQStBeamoGtnMlg/dVT7ugp8DXBIl4o1QsovS+hbiPFdaFyD2oK5D++978p/9xl
L8xn+xuIVO7YjOsqtkGg7ZjbknqXtBLVZm3N+2Y7hpzYWdUbV4jDmmRG5gx/CGGV
6zLZBUzGs5TKMgaKQrhNc+10+5Cpvjz7qhC8V81NTx65G/aCk1/hvh9PErzx+7lz
2i8sHcrDR4N6jJ1uWnBMfqLI35bpCo5HeZNFK8UbqxuAZ5bzgezx+9dWGc+eJ1oz
KJftUviw8QzT7Tc4uhshzPY/+h14RDDG9AiZ3W4h220lZzNCdd6/hH5bBtmWvbJw
YgfHmnArALoaM3JeF9MmDcN/eNjo11O2ubQaAReKVsmk/5djz79BQXkkF9ZgRL8m
KleNW/06rE3PqcuMVID7w/Z0qdesN61VqsE8Wwb7UnPl++PKhl3gh+kIKVfg2F7r
tnzt7aQfqXc1srrh9T+pOi0uzC7HhStahVNh8sTtX7SwlLN+mYparFN8nsh7bvu+
nEpUnhaRDYzHl2g3wFJ5vqHCSzbrKTMUo5LLItSZ1wFBKX/nuJ3ru4EEB3fC6ibD
wqR+yhhQYwBOVFTFntzitZD8hPpkJY5FfQnA0toMZo2PXEz05wojkJi8vtjSq6L/
/kfS6J28Dow3TDno4VOOYaXLA/CAw6iL1cbs+eK4krcWV/3m78EeTIQ8n93FmDNc
Ja5TRP4ujo4wl6f+ibw9SZvSd4nYRUEHk9mSaH2SM/FRtF3A+hxWH1Kp0x8R6c8C
wkWaVZ0sXLq9st7obRqwHrasWISp5Xsvr7DMk04gxkVE2eLgs/t+RXZMf6CGvav0
TwbD4Co6jHLesaTjdL6MjipLYo8slSAoQ1ndh9crdbgPu0i9iFPyOCPgPAz41QwU
tPqSYo50f5eQ7oln+vbP4f82oP1SvQ5xSUzB3+FlyWHjwj3fDgIUVUfrWHbAjEuP
iDq9c/WfXYrJxE/oFdQjSo6055yGxc6RS2vpjuOeJe8AL6bI7t1iTj3x+Vw4YJno
THTCVCYCryh4SF6MIszke1ibmPAzu6X8yw3svbpvT1+zye0yLKxG9m0X/36yxCuh
ILO/6MS28q7ngll5Zn/tlnzmZODGOLrAd723AQHEpCdEEp+PalIS/fne+PbWy6+B
3j/cJxuk5vWu35ZziU9cn+W06NI1bgAe7D7nbGkFsY+2R+8xeX9Mk8Uu4RjGkSuY
+Dvk2I7FqHyTmOSvR/qj2kjwSZ4h4rQ3bb8XuDA6JE06Dj06BtCSXlTj7BO0jiIw
NmelKHATb400Sl58Nmxf/x4KdeOK+Ikjuz5JwohN/dX+YYA+pP2hz6EprzxaNZhN
XK2JYcZsHk7eqjtZd0fPYmyAHFo3mSDIFqokXv4xuQehhOrqNXBFvxa1Q4AXVOfP
0x5+KFDL16cUWQ15m05+hIbnDCTSZa07lnG/C15RUaoWFrQhGeP+oOKWN2moNpZB
fnREDUzXSzqlJ+uBy6MLEiaNMYtEbtFB/TYgGJWPcWOctZTOjG5MF+04KmjYpl9T
/yrFe1vp47J/6p7diTuYAIBSp3oYjbOOZnU1VwWPS5Aw429pYtLg23gb4AGavy96
HC6vTezbMiGkPv4RsdWcgNEdhV0UXE6BiEAX+N6qYVegGBsRYRqHzeFZNH15N5FS
EEht/ZpkC9UWegFs+epoPVPAAsL4ClbXvgiFTgFZ8RT7YsKAKNkI8q17FRjwWdyg
J+a2EohDXAEILkjKIucFZonF64hQZIp5E6IAoBlolFr+jNlDM0qZCZ//n1p6vtRa
OQgTba+J/yj2b97Em2lyQbtm3/vmMLz7AoKxFemuPFRC+DjxC8osfOcnPtExdskt
UI31cAcPi39MljFzCWMHI/frL/UFkQmnnFWeEYRKk8TiRVB6l90M6WlIHhvwkvtW
aY+bhnP2QxJ6Uqv2Unt476pSGhty3yYHg5B52UixsM5l0A5gckt3oCYx6wm79nOZ
06+SuGoii+K2XkYS4XK7JbCxNRI5ydWdiHqfQijThXQyNCtfzGxUzBAoRvWgkRLl
kFzS2ziR7aZNH9IVNMsezsqFeBk72jSoZBE57JSWdv4Y8swG/DuUTl6pLIfqyD3i
MtKHc1sl+FD8QSiYR9+zXhzFBnAMNnNu+tb8ehEx6XohS656faNC5SkYckV738H1
X/c4lRNHK0obax14iLvMDh1jjWZjefZvYLSDhCuRbJfj/NNKxRqqGCIJ2ln0fuyz
mJ5wILw6SKZBbXX+W7AbK17yviD7Bw31jzTm6iou8FZvin6PFM0QQhIWjuov2j9h
jjU/Y+8hDmQHWaPIBrcQINjqAclAeBZwFgvtb1iCuZDLwkml+TQc910+/w/zn7TU
pXAvq/VK5FmCtbGLGERCR+ZlZJBhHa53hqle2hN57f/4HjdG5VtjK+Hp3oC097xE
yo4XVEOysDaq1EuxNmiIkKxmsz7eet5bJ34Stf/HZTxOFMvIJGxnNrZWzXE7Ke+J
ioEc1vLnvHPChzfxX71FVcBhoe7JWQ9ItQu+cMOXNn+gKgXFiiDPxw8l39j+dKvA
e879p86Ykwny9ZSBnkcdBD6Ib1Uh/ZIVfOnf5k6roifJV0WDqBfH73UblSz8xzLK
JGwGh1RW7ETEzk03xS7sQZQdMsXXLiUI4zAVfE0U7DvuVqROq5CUSQA+eib5pSQR
hAwyoQ76HBorlHer6UUwN+xV0JTpHx8ZW185ja8LWcDQM8X2klIiSKveqFfmcgfC
5D6jrZSkzFbT9v1dDscUXXqjPdRhAvvnguWiLoI4zX+PLLlCsdavqvIfdmkrnrCn
v0Td8fTnTLDqelU8c148nC+SUNZAjPjz5YjLQuN7hxDNaVpjVm5yJrtXPPkW/ZWQ
Em4YlSyW/feYtJxT7fpDrui9QuaAqVzDFxVoOe5ahdRCZBnggjpfeJkhykcpk/hy
zhwA5JAuP22iEv3UdA1ssUA3nU40qct/kuIMTYAYkapQb3nrKeMrzA5RKQ4WIYpb
MMUbIPso9M3JXekxGHhO35op6T/NcSzB0J0jfchlqR1zymPuHlibmxx5AxH0FGRb
xLbxwQrqakp2xZEunPqDFdvV7lVaX4//Zr8H6KIH1EbrDCDHx3n07i905BUI8ahV
n96STUb+hNlM4csYWOYRRi1rwChkNCp5Tk5boa97dXccyQTm39uDfS7y108HkZj5
k1lT/vLpyNwVPBEdOjCnxEgITa47D7trrBzTIqvy99v2nf0lfMdB3mwsH6+xMcid
EJyLevdmriyYE4FQfA/i1LOdXxL3m6RiGG8Q6T3jjSTQYdCZO1gLESAiiffyMCy8
4c0fVA/lJ3UYab+BbPZRu9Wm72s+XNxqaVg9ahY99nNhgXbqBSfgkZqUrgwKtEeT
LxpITg5dO0sT+F+APsrQWSgnbMAtE/0DdpKCKBKVgAer6ey3cma60vHHmaODsYuF
OaJwPDJpsv5vH0upY4YOXW8hBqkO5eYBjr6QcsBuN3DpBkdgN013TA7dcHEALOxa
YVrP3Xj0sfIL0r/Odddt66TLzJUHht+R7joFxM8ixp8a5j+Wl8RwEwfPfCCtb9Gk
EqWNO9P1/gOXKN5phZ7EIU8rKU8yqYVo0Rfv2LfXpoIKpCdiFXvsbE0sPD0HNziG
r53jWHnyOIq5/2omWte/cMUoVTfKpnPMap3kmu9vI1vbrSFYrEXwzpc48+xSicS1
y6k47YVV64MagFOOuQJSlPvgsaLV+rdLmaGAs7ImC5+CAaNcqURvgAFmTBlJ4hPK
HRGj3994YKO1r+BEjw8KtrDFDzV8m7t6T4NRuZxJO8+XT8qAt4cYc7iW+aCbGzHa
w2Blm6NqQoxlEceYAs98baAKXduou/00PxMUmIo3EqW3N3kVmii/lyCazqZQQZMl
nGVwDNeoHZLG/DQ/rqRJP1ofcqjTt4oVFsIDSoaa/uxwJ3rxOiYknbb+75heB4n1
t3NNApQYUaSl9r2dRNz7fuEKcKn/nmM+3W6rFTRATdj3TJUftSgw3iJXJZLO81vX
dZG90BnuPI/gQvqVhmw/7SZRCeZqlttNoJ/Oypbl7/4c18tJX45/kHemZ+jufnzj
YwYbrNYi5JaWgXM/JqYGXGaVD2kyONEJ9DLOvl2UkfTPiaEsCzaRqmu8I53d0vAR
p+SU69DJRzLfUXsSPGQ92xfF95y6dA8eZDy/KL7CoGjVdqIe8KHY80ISLiQjebLo
geJgoUIpQk2UkPKHfWRG52c5kFvs66LDbxSeaTJq1i475uHYbjnLde6wFzoEBqA2
0K6xYuq9xsxUp5xYdTUKkdzj1hFHfQRixQ3/awLU+G0xA/uG05gQGR2eK0dtlam2
LNAm9PN+RmmK55QbtzrUnKVJ0aAytJuCgyID1dXNrFW4sfkOVhXcOBlN4PVi6XvE
qj8QrGSJbKpuzWPR/ZcnDub/NoPDHafCAbBRPS0bJYI7ghifjijYHczQ29HG2gU4
JZycDYhP/oN9PVFDkJCVm3w8tkBbQyVrS9bfjUo7Z7ET11sytK3zBhNlDI6RMLO+
HKMorsSDL4xMcP7NSdpOAdnne7u+ezlAvX+8aj8gmI9mJV0afXNJcjGaeoSgiCb4
4+F5Hnyf61IsAAghVGpyi46Z5opidoUeuNQKlnrx8cCVKABuf27BWj1NvdNj1fZO
snMMdIJgVhFX4HOT/PebF/JywQCh72EM4VLcRuZ1FZyAccS5RVsHx6l6m7SxVxsu
JdegCITiM9dLNGe9dbnUg+RN45/sT+ZAvIYvfSr4lxsPxsDshdoMTFAyvRXZzRB/
2t1YGKlEm25sfWgchCZN/7DnDbIVOKzdnjbjJ2/lIQxHXABHzSur/aYtoJE4lNlu
aglggvS90XKWWMNXQ3Ly7l5UG6y1uQvmm7hlMWDCeUjgb87kSZ/qHWsZrUmcEe8i
EH+ig4Uj3TTU+UOCIVlrzvKTCNci3iBRMK8lIhicT5HmOX0NEreTEsZADNRHK2xz
9WXoCu81+fvqnu7N1/KjfmH/uBBexBGSnHxG9LZbkXZq+pqUMKWWd2/heje+Wtql
2zlGhPhDQMEziwxYeb7d2jxYPFAo0YVv4YacOd8j9R8IDJl86E8TCSIbffMvAp+d
ZgyQifw1+jYiOeOrB0Llpb/Qv8QFumNu7J3kVwPSFbmXlswA6KPybrz9AwF9hGLU
n56XEmu8nOKV28W6RbTxNXnJHDhN7qXIx+aWCU/Sa+A3a30ilTbTPsxMqKb3/bd8
5e7rfmfm9esRtkXPgUDmEiAkUvoDxOB+Lp/JDMgmMsetxB+UHJRfMeRBvO2Rtju3
h+kEcEVZo/oyGXVJhRgeW5xpgFZgTK6nQE1Tr0511fBUGpxAIzIQ57DGhbFMFaSc
tHFc4V4dMKTnkS71Uk/AT+nv5PTrIZLGhGcrGT1jq2uoBQHVQ4hxEoVvgGZm3kSl
akNM92LPE6k6VFI96kb4McZgqMEvlLLc6smxYo1DAlaxex5ABmUwbkcQ+SF5JXqo
sS5gJ3mlccAxZxt6Bjuq71qOt0pvmAv801pvyn+aQ4MYER1QmCm/anQ0O66M55IO
lIcLd/CIZyzK2/KIu8op8CUVQoH+D/qRSSCKrOhKNU/LyDJh0VUliLsIsgRtoYq6
gA7IKTa84/Q12ubZqUPY1vv2Tee0KHcjjmoYUaI/XTUaCUM35OF4mcufDpokgivo
MxnVhGMcYqjp+rPUrrp622nL1uzpBr2ZIZRCThMLRMjAU9Re0GYOR3E4afIR3Ewt
QBWgmInWs152e/F5MLonjHVO47mIjWQqVzxeUe5t+pjN8we+xn7zcmXaWQ4VO3hi
3fi2XWNPFfxDe7jZzB+VZ8Wj0bFealX0GLFcRxKz3uixJO92g5eU7CkWUee+rgnI
gbmv2EXtKyEvl/93RmBo1fQhZ/gI9C0tBdFwTa5aCUI1ZTDD6bJByYBUkLjiwthz
v34z2UBTLHgGUMhL04zPWuSO/aJzuCeoiLMn5TiXQ0T9lhOlmTCU17IEjB5XRK0f
dp5PLSjyU82Awl07agY+McUC5/kb1A94TGcae2GGKP70JLoZB02qgB+obrUzuWtk
UvpUlApSa1t7CZJZu1GrJlb+muZeEQO7m+XNJXv3KDQChyAIbhcM+FFINdtGcp75
7ou5XGUh7jl2+yWEnvW6yhl8Z53BsmYeqmIBKa1f4nPH+XThbFYEeTkAZeekqdQQ
H8tU3Mmv9iaVfJfcowRYGd+U7qQuJ7d42QwqeSYhMT6oO4v2UZgzIX2+R1Uusudx
MdIWm8+94NjWA1UKLR7GyMyxRsCPT9BnF1PT88D81K/vvzop5rZQy2eXcB6Ofzox
CO5Vv7EMxAqW39A+7C9LUFIXIvfn5W1ev4zDVszXObWpVEI2kINselZP3xauQsfb
bI0cv2DLq9KHAq3dZV2qBD+Hxi7daGZuxQJ9D1fPuZo+bzQGR7oHfkNvQmiSQdlc
Xuj9RhffDeFt/M+QQj4ElkXy+8sqIl6y+SAGOtOqk6/CwAhXqtSPSwjHB8PPWJrR
7czeMwr2cOwsl+Kbxh9G7U3OIrCFnorruDseMFHpwGMQUhX7Et+ED37dSR0NGOIH
RJub6lTKKBJULHtL3JqKDoD6UF4gyduuvIMdVEvQsldIQK1VtuCCzacSgYgoZ64E
xfnO2CUK5IRaUuswAQ5O0l3Tt2VVeE24fvor4kqvn4E9wEmkdwx9Z08E7vi0y1Kp
z4vOoKsXQrHp7aQWiEKn399meERyojjpR+BgUIMbttIMqkquQSSD5qPoTknyqSC5
4CmaohWZdpIiyE7D+NLWSMBXXThHXIpsnjhk+JGoax4US2fSjJYG7MRrNdX8JSF/
ClrwCvjzRWJ8EHe+nC6+YKUqsthT70iJmjGBDAMS698r4a7cyKcnjLXY7Aixpkg1
67+A75Lb+1tI/j5F6CWz16vrv2AZTCD1btIfReboMV0zQDZdgr0vWauidxaWqhPf
544mIgyXCmLnIYFVQfC73vhbU5Yt6Do5Nj3uYXxJUCOTzRpkirm26xY/7lDptoS0
E0lB0CkEqRUHCIHhc67/wpZqKfWlw+ZJ//Wo1jWjttNmQNIca37GlNrT27DWv+Ve
ztpVZrdMbC8wCsAfe8GQ6gaPIgQk4s2KXa1vvwqQS7fnMo8C/in0B3v3t2Qjvkwa
m04HemXSFfl1jY8EAWQli1fhvA5FG6BKCRPnu7JzRVClXjJ/1X32BfJ1MGTin/P9
gQAwbME4reAYyIwUF4KB/M+Ii3XkyFbwV+2zuNZ3/aMXguMLFvYSn/EAwEVwp2VI
vgKJAsxfydKXfCzK8wJBygt+iWbhbCWoZoUeoLmB8E5PpspxJoiaTc9sO+1uZCKR
3UDcR+ZGSqrto8Iarf9i2vqRPRR4C7fApAPjrpSg+c0xrvl+0T1x3eFW8QL08g70
54dI61PDKcSqMy/JMK82UOU+uhdv0b2dP3K4cf5zx6DWiw+f4tFZe0hMrTDEpYCB
oxBLsGh4FB/hENvXyyufecns3gtb+10vwQOv5TzA1SpMcRi5P3kIRdnTjutLuYo1
3hsOLF9AR7O78Wexg9OGNFvjvGUHczlc5zHTFJp/2GywEZOvEtA5wwx/ZJSNUpVA
JETyEEZhbfItWlzffTw9WVJrbC30uHm8hNcdGHjruTossfWB+hY+j4hrgRia6IAg
X6IHATjbrlDgYZjxT9++afsSLtbJO+DAjRvebr4Xk9bY0kiwVCdDauGlX3/aUOi3
lrdVC3RNX59LeXFMfVMkyQY10G9mKVLe9F6imiafbyyv+p209q0kQN8Rgmw7QxWZ
QR5Eun0PXBnwtBMPbRBX+/gyG7N/kXNJJ6Uh9OyUaQRw9Bt0a0uy2Yo3SV/5igiQ
zi1KtKv+0fOZei5G6JNPWZZvE9LzIa8XGw0s/Ym9jBrGyKm8PxAeFlkZLviPtUz4
aHP/ae0rOeYfavakkB767bDhpe02j1KQMmJYb2MYfkb/82omVorCPoSgwK/HWsTL
Ek0tH/aCigUI6TU9I8d7Hi3hqtC9aZT/QoRhXIbpEaU1YYf/sgV8agyMv7yUzdDE
2TDK0ktT/GitIWUyUGtUbbWZT8WHPfFW87TRKy8/18XKmOHGJ9q87qOkDNp3A+dB
e0JaWXUCxZR9xNmyRF8oczDUMSG3X9pxWpQBKic4nA9FW5l4gKxKp5ILeXLCTaHa
fD/8ggngXjukbK7TJgFPF3dWk/wUzJ3/RRfVCJkB+oaSj+76ql0R3O7c0Kth0kOA
Gy859NYXhvG+0LVO4cbPFntWrKCvAk4Z/uR8PmDV7JOkW5Im+iHmHn53evGKVHwH
O6NA7OcL8G1x2sdrTI/Ivirog/mZ3oYJaAhIN548JcCE0Q5nRw3YmDYcaPI2oUKl
OO/m3w57sPQra7iz8T+bKGHVtIpMHQM9zeqUE5VPpmYreTLrtL9/CeOPWdQjcOim
qpuMSuCm1HDx/nzO60Pfi4kGHiaUdRfpqyMgfm7Rl9xYM9Q1HzWmXbDlMxY7cQnD
OcQueKfwGczSpNmOKApH2WBd6m+9UM43MiISrSA7ERp+Bfn9wXVCwnjH9O7jhAik
fDYp1lYsowT/QWHhhFv7XkEG1yz3hgcmtOUnZv4NODGmhLWzjTAUESp9mthRk2RM
mSqj9koi0+RF0LBrEpFbh24Vc6VvDurj9yTheJ1KfYo7HnTpzNW47fem2E7ukDdl
S+vMvq3TYnda56tDDEo0ibCXRP1mrZAQEc6fqZ+V7FIZdzOJ/YAJTG23flNfyYBn
qJIRKwJsHbXFM4bk6ZJKnBjq1LWZFsaqDHHh1EgPhq3Nw7yPlXQ3os0EiFLjCNTl
OfHrChwgDeTxpdapxSvrAdhZfiJXerh48wAIsTVhLBRxhJKtiMzY8rYYTo31uCGG
ITLLXYDNybG/VESZtpbhVnGbfdhzdDoAClzcyKAr9YPL1PUS1su72LSSkHm+DU02
Yg1OK1lCxGQZq5b+1GyJGO4wtxW4Ibe5GzbYxoaPEyf19RCqJF2U6jY8KGNAmsHd
FsZjxlY5GMK7dejQS6RQiKSmDhIG8dXPN133kYAKbOR2ASw6vD2lfdzC4pWrm36l
c1hkiju/c+vJvfAB47f3aBRxw0hHPuxOmI4TlPBnRJWHbd2DJvywJqVxs7eeTQ7V
pBzwccOi0YfWn4YLxt6zlblaOMlAPaQ+QH9UlrPhDZjsp8ITE01qHeKkoyl60mHK
oaj12CPMsyXIPrecoMvQWiAshNuabPRxEuE/ws3OjEseA+dk/9wMa6KCQ9mFZ3Hv
NDwABeHM/QWDGi0noqpaXvmT/FvXBiHlEMfuNw7zlnBeZ4FuGnKwRX2fpnqnlXrO
9cwRzRum0lhQvTPAQ9kGGaGBAcakosKZJhmBoG0pSl2XpNw7miBLEG+7RuuJVLgc
tCZdqm25LWqmerc5dvtFu7eMGRDsXgctRctzLq5EjO4fFm9Evia8amlJWntdiwL4
T9WT6D9EOBlTf03WUvG5xTE4ycHli61Y64jJCMdweahW5r97NMt6Pmlqc3OcAm2N
3SeQo0WQqQntt0A47Qs7BkSXJAFMZrRjjCZ4Id4lbcYcrADHqpkNifSDTHE1EVp1
7ofXK37D65Zyi3xh1RLfpx9jTS3i+SC4/B2bx33ft6gyeMczzLQ4dVZYMVHfOa9u
NEo5qM7v57xmCx3+0t1ACff7MdyOJZ6Ku7+EOQZWNx0VgG2aanC/pe+i7//R1enP
7wM7mhLYd285AkO3HNlXmzunwKjuT4x37HykAcfRRZfhlHg7GqGeQ3sUj3BCIDDy
p/9VufAP+yO+qC5fyf8tWcbS3kN8VXbUrSK6wQixgZsAQDDMwwhW9YHC7s3aB6t8
UCAInLazjPTzKAtbBUjy/p0qT6osa3RjNa7UwW94wu8B11pTa+5B9JEpgwnYxmMF
4xhrdwVyNqaOv7AHtoOOVefUsdQIlaTMLpQDzBHpT1H/vFB721bILDyXqTDhb2Le
F/VX+8Tddl6m8jHyP51sxtEzfU/X0jH4dmm3JEOhzQJxZLF1yGOHFn5t77GTTR0B
wb5W8pFyRRl1Yj3JXzm/K3vg/88e2+UJYbv/jH69DUzQwmD4MsnLqRcAUmwMEQee
+TUy/bSnBnI+pkiLEQilfqYFSeRpY0UAppLObpCC0jmD1vYDrdsLL6D1pMxS8g9Q
fUGQa9ogiIj3Y7SoFPZbUlAjQDovAj7owUWmGa9BuF7Lssnc9ov0pymcR1yg/hMd
5nTh+EcuysWQCvTXrU6v1bNClohd7occqm0YXmfChqLURHjAKXZ0+Ksgw+gVOqnT
Bq4JRd6+4b2ArjyphYTROfZbD+1RY3KPnx7yjQAjBNyWX6Jawwh12zbs8dGbh7zp
EWBWk4Tv0/Jo5VheninDq9AGTlsF0xr7OeyFJpj9oLMq2eSNNZL65TVs7bRPWe0V
uNZECo0E/z+RQXujvSVuei2b6KcCVYLoXaAXWw2qhR+Dk4YfAE+lkwy2dOxn/vTX
VBuMEprsaIzjAYtIsOMr3J10aeqREeejqKngGqbCsf1WQ6ihlw2O3f0GWwF7A48y
mud4CjiDNTn8t6imiD7AuNc4NyF60rUpK4Sndgl6UCoW2voo6SFl0x4FDlvjU0Z4
VlHdXpkXBR5hm1IJQwbLTf77TtJwGmK31JH6r2pvqJkdl4OCO7jAK/2VFH8hhknO
+gTxRmNmIwtTrWTBbdLSYkKYneXVylZXjXF6FLgeWOWJFGX2DmNCHXHNwiFGr5Ko
FiQvTrYDw2sb89R7bpr+kpSLmHaEN0rgda9UlegJkovLQiyutXqR20JGdPSPj/FB
5b3RN3uLSSZUDhI0p4aw71bTp/pnm/O6vtp7g97Yp8p/7+QTBdAL4d7v03He+clY
+GLH6ozfNRYfAcVkDvzu4eUm2PcH0kCsbBwscZIhxc6Z3nXU3VRHQT57IWZOX32g
vZ0Pbs5aaNUrInAjKL8UAJL6FE8lGHvXWEkEjJQvPqLLRa6ZjywD8V1I+Qkgp0f4
QX5GKvx9UqR2igSbazUvoQAdk01bGCZ+WuQLDIQdos0iDtMjas1DrQWM78saCuKR
VgvjJPsJuoRtz5gA5A5rYk0Im6zNTqL4z8UeaEmzegRurLfZsrL/rmVF0ngdoIVk
xJ6miu90yDvcQ0/jdcfEw06Qr2JxpfhV99rehH3OaB12CJ3Da9diH42RO8P2nvIb
rxmInpgOLIYdqR896pvy813QluamyDmjcQ7MolilOXYVtxPSrAUvFCYp18CCWA3Y
hHZO1No2rM7tRLmiRZ7VJsC+6ppPs79ybqoXIgJEjWerwh4J/4KNIMfUC8Zqlix2
zLVUGdgTMHHoeimBWNurZhmMz8BfDxwn+JIwMGJTnfWmsadPTAxvZLCg0yq2sXZP
6OXphL393IcZqFyKQhOThjkFNCyFbcOUP7snoxBnkQMt40AeKFqP2+UkQ+Nah5ne
DmPqMHrd5G4w1L1NGFlFy3LJvOoFJ+a/esbTWYcZk8eoQSKFq0uL3uV/a2C6HTR5
c6cCd4QSpQvT8G0VYDXr0nQhGdyhTZVlJGco8dSI6kRs7ZCB04ZFwVTtLhREcTTx
1iYN2vXsbTzgYwDEPoaJ3Zp/N/8tdCavpApBaR2c0164g8ZiufE7Ayo+jFQy6Zd+
PIds1dx9ldhSouHiXsLUfi61CAe380GJfqxFbwhvzpWsWiZv/mg20gUbz2ut4yjE
XTiJDs050QxC/0XzxReSY/Jc7kD2xjvyD7m66k4wpSjpw/MfF+FD7zR2SCEBGe6u
NMvKVCxs6OqlBop5Wtv1loyb3QiUQFCps89zd9dan4hC3AIsRpAyM1iUSidtytYm
YJ6UDdpOxGDude42jOiVZja4j8CaFGjJ471IdUj4G5z8wt8+HH/EG1UQnCmqgmtW
GDZiggI5RikSVMceJUDhlC+mgL/1dGCkZCrsZv8p/aMeY/bFLF0meamYfSSa3P3J
jYCR6oF1QpDsApDjSjRvWko/EL6X+HTIsN/UgsfAsqihRSkWBrmZshsZPAOJd/D3
0XN40xi2BK9RTVJIbbTkmKr1SKXfNcytpd6kFvAOuPepqYYDb9XF45LfDxpTxyfp
keUjRUSm0jy0fJCyB2dnOSQ7e6CO2WjnggGJ1Xdy0caUw8QcoRGY7k1rE9tEbUKx
N+ZZEYYPz8/Ln6iqaBUKKeME0XRf583RznmNXbM7OQmxZp8EXRFzlpN7XEQjw4et
rkI4ugl+DOPcHYiL1tNEZ9NlE9ZT+f9/r5fl9xTlSddEJOm/19d33mtGuQ8OID4F
XPmEWkxrw7OkMfBLki+F6BAxJz3fTH1UwTEEoDNUpC2MA8paqGL8Wdg6xrkUJYeW
zT7OH+xibi1kjFikSlLV5Xy2LyGXnLabeBA4se+xgZusyHCu0LVso30eg713ls//
ML7T+HJAFuiId8htNEazbGBJ1q9i8ShothBbKLcKQROHXiAZLXfwF4pF0qMaiAxg
dlt6Gapbc6CAHj5rVRZxRv+gdUZZ6yAQxir13WAqcSAcKpVb0tlVBkuhJFa2Usrw
d/bU0WJayqnzHz1QH5ha8dyUIwDUqKPVL51gMkzH73/OFwdE/jhUk9BFdVIifai1
J6l/4uvy0MQYkN9ohb5y1sW0yavSYlAvKc7LAP/Ca5SbsYhaqeK0WfT/Qf19yfq2
5GFS4B7I3Uvxn++TXGhGtz8lCY+g9fxEQWN9eGO7NJR/pq1WXBY8/0Es6PJvKj4i
P5jK+3mjTHBk3hSVKdlzEeqt2w9e1Oz6TtON50qNJWoSvUyJCHGNtT3AT6D7XId3
Imxia8X3NBO1wKvTdcflIB5X98HeRZLRK5lWlIHfJ8d0WRisTwh1ROz30aiOR+lH
ahhRKejai2FjIoLitqIH9hir3JGBXrKfhYLb/hb7DAOUeC9H4k9y6HJDtZNxp7PY
3VBtxS02wMMdgR4bXBWdP/WX6C1AhtPmtEHEVZiOWGWaqhGRC4W+YCuz3HP4d1Le
v/U4ukMDH6u68RgKhTvIQRt2RIxAvQ0EBcebecH6MZG6W+0LONCcmJ18p/DrUX+U
BNQ2XUM9t6UK8chfHacJSd09ZDSJWFAnK+ZN1iq9fE/dXyGbEe6mEyar1d02G1MP
AOimQeOv7Cv70VgNYaXyBAuMKKB3d3eeQWnH3oz/VMRtJxX3ulcG/IXfZZ32/S7O
t/9Py1RNqycsFaVnuBkKeb+B4z8BFWpZbtrJrrA1l9v6m9y68HYTXfaDOz2KBJ/y
9NrcTiJgQisKmWkeVNNh2n+N8Lf+BrN46yo9mGFqEGAIY/dIWfYa/4onw9TmMU8H
2LZDQ1ZILhxf/2N8SPu9l6/wL4eB/fCemGzxc144akRdWvF5elOSQJFLCtswjSwO
RBE7UK66sEmXfWeLbZp2ZtqzNML0HUnvcZNek7cdUX5B5gEDNtOzJHugL0y3lfqn
Lb49iDqNSIvTIWEh9KIBYRtWjAQg7grzfLnJNk3rkMXEqDfU7AOWSF+zpP8Fbv0b
mFYg4NXKJsEiBjJmrKthQTX+1O5oGkJhlmBlgLVaMHZq+un1y4QOiS89JspxG96s
VWg2Fx88aMZi2g+O6LoSt4co/mNMqR4mSOAarm+FOSKZrCOH4ra/XupUYlLM7g3g
1GMu5Rgp0tOa/i5T9SscXEWyCq5xMi+e3sP16RXM+dL3uRQ1qKMvdC6PPbsgwrb8
MaJqK9ey43FcSrL+UNUMTOzq+zbbzrQ0MGbo71wOazz3rxqpfuzczpwz2duaDmvL
KHOOJ0jGT0IG9YynoGHzZeQY3H5fB1re24Y5uI5FJzOBP62Pz9fOdTAw1x25G2G1
aGj1hDLZ2amB1lnTlFaDwFJ9/VCs0L8FWMxTwJU5tngjCbSqO/CJNE7UPHhF4bnf
CbNFHTG9tpRm+IF0oO9qrnUyoxi4ar+umVrHgySEum0zp9Eqcb6BDB0v64PBU9Yv
7w/M+qZi9F5/lvZKo74CaM594jHef1vgSw6cz/UN+h3ryteEan7fJJMAkpONBaMC
yBx5wZRw0mCPTT/f/261VUhlpNXE1GeuriKnd2qj6b/unvfIJe3XSXkE26O1ePkn
xI9TZbsz/lbgdh0Fxh4YEJRbpD3o+l++6PkUv2lHccG8dtnO67CZ+CY8IiilFuWC
QzVK5kJd0dCHeG5gyF8LWjNXHZ3cx11bVDb+pJPXpQ4WCpbYZGAKGUxhZRnp+0/z
eYs7O07LAjK/9qT1Zr15HeK4zII61y/7xmNsdbwNu9vmHKOXd1oYWOD/r5//a2EW
2RuxRPiOO16npRu850grRhpNbsH+ISIdFEYnBnufYt21tlj4UikGp/erWnKhgYCA
ZuyXbw8IVeeZQiaASeRDZ70v6k+ml7X+rnc9OFqVdLO4ZYJH2JFhJpe7vmin8z/1
pWvq6cWIXPDiSq8EOP6joDvQgbaOSvEGlF5Q9Ba6pgDU9PgJHCgWjBHy3AcMfsvd
eJq6G6OwVMY+lecgYPbDnJVqNpCz4odXO9tDvigMcfs4Y1ShQez+9xTFVZ8dAS8F
Jilbq8cY4OGklqTN3LgJJBHBtzH/6HOa5FgRq2EPk4hGGwhpzd6Tlck16De3nRJT
qrYRoLpy8RAQIxr9kMKLMGbJsmqkrsfnCdXGjmpHWMDEx79zBLxL7/1jk6pUpgqp
n4SP/91JqxNmJggOC66m+4J9i7S6ECpFb/dAoZxs8W+LlfwBxTG+7CVHdgVvXHns
T+vHLKBAVv+8fhKNKyEC6SzpSbA4B1oM8Ua99bkiYYrs78XZ81rpZzua6BcW4Zp1
KEzxsgGA1U+9PheEDjnM2QCFyhjRaPb4fN2puHpLqUoRIVufMbCXJhq0kJnI3YO4
OVhleqDW2ruVuCKE3IJp8tneS/EXv4sWVYxSvG/laAxWtuEZXKi8XIA/zCdiTDNy
s5vKZvmntEh6lGgCfIjmaHxTGc0o2k9C7GkgWTvDdErnoJU22h7DvnRz6ik253Nu
qbdOIklYQgdUyFPjhRLsmuFTvB6ogZzrZ3kp8tsnQJ8+QiZ60lpYrYU4Ll6yGi0d
0OjuOZWnZGl/alVQfpBjbIPWGMGck/BalIOIHgqcB1GhOvg6A15OVdmLk+ikJGS/
D85OYJRsfWRxzWkn6GJTZIDhPU7EtHc8jEDpa2K4iHbyMn9pTEJP2ccliLREeDRj
439fPJrm2Qy2q7wrEH88pF4amFCE4ILgZVfhpTTvJ6gEj+5FUjOwipuQ1Ip2K6F9
DdiWwXUSX/H6LD2t6fzfhdeLMHTb6irTQnxfYNrLOTjxenUpCGukj2WsAl1PEwlP
A0vp9CXpjI6ujdO+44ZnA8HGlTYFD1mKZ0EtYRlpTZPDT+pgCV2E3Uy7SActF9hK
NB7tZ1tUzBJqVQQFdqriCUAx3/A/+nfDm7J4l76iLzc58k6TvjRuzyrIdSErFkTV
mOHSXu/2oaCUkONWHd5zsLR3j++hGcUO4fLqD3fhNscgEoHweeuzggycxPW1pRwb
fSn6inYjqpVNZ9BurpzSvSljj+M7ciYau7TrrlOxTiWkcZrfrQdIadIvqa4TI7XH
zn0Q9RrrFf7aQOCWb1ujQblJv4v3b8DukIz0lKi4IB0ivO3EJXRvVibEq3sPgG2r
E+MEbgssp+G0JdqH29yFgJS8B5uXppVYY+IbkaJfkJ+4iS51YkuOsndkdoNGuvc9
ERfc3Sjf6apAsMfc153oc4wIInYc/UZc5PDF4ms/h9wyzyGlXObsKbRjE35V/25q
vl8vVfzmm44b877RyHI1jLaJPsr7+q1HXcZK0ZgBzRHlz4B1Nz7oQ2BGE99oIQI4
SrGapEf50NUfu6tU0NOCB3mPLqrP9s0WGaz0LONXZduUxgwj2rK+0NPqPZkSI7ro
3xukv6RE8Z27rfv91/5stOyf2XJUuxawVFBRIHhzyH8Qm3RggkERmqKwYglXPkiy
XX2JOuA/VKZeOcJUrL6y2AV1Awr2vr71V7XtZwwzESxyVv5CTmcggiarhsHqUnRu
NqRN/Lg0N28SySPMsuDrlsNFq6Lbe4wz39f8YuPGZNRAfePmthxGB3CG6ENXtjHU
+5liHpG0z/LCGXI2Lri9ywzlbVVvRq1R63LWtIN0YpyptpK45qm9IiNwaueWu4gX
CKFMdn38zMx8V1Aij+Vu5Pio2jpb3k5Kke+HbaA2YdOhvSkvMNaawrh5mV2kpvye
K9juQ5It0GqNtIrHhwa32CVa8UngeCH9EFS1qTp1/cdBunxPNPjinujG0umtzh3g
2qLgFY9KzKmLPwOLRdxRGaFwdM62qh8OKtmHgYT1tVNcz0ak7lxdvOIo1hLYb2K2
ewFJmrQAwV2LqqrPzejryaw3mahrmUPmQI3w7mSd0M4kOTSmMdENMRooeMQVaph/
n//nd/VeWF49OHMI34hBeemjNRoz5own8bhQFqE3BAnehNSf0kIYnxXgKkT+K7Ho
0qb9MdlKY+gUh/2Wkj7jBwfwqT/2lklLKiydG+uj+G4L+bQLcWPkElUEdEgivzZX
NHUdFKH8lljDjDLqfQXEaV6U/hfd9LMqvLEOi7wJN7uBLxjFF7ztZh8UcBVGfFjq
ajP0Yq527qbL9kkgztqRLtCTRgUvUpb+rNkpvEjv/oMNfBc+qC7eCFc6nSs0+Nag
q1v1tBQ9x+qF+XHEqMGCsfRcCoDZ4qtpZNz01y0JOlcwRPHVrDyTCdalx80N/SlV
xJSFAC6xb/ypjhDojU3D3WtPEntbJNfvy7NS28v8CGTIITwJmbl3ng6tlrp+p8t/
CjAMT229y492WXXAZDaJIWW4UD0/TyQpquj0g5tXPQqTFD+JYiaz0ppL6OYGW5gq
6TvbI92gvtpDcwWKq9xM5jsZ/wqeoZE9k9iH4FZkCVL4c6MzxmrszZ6Zt/15K++6
ux/NmFdRUix8jVGQMnSAutjJDFljBnlhFAIF1/4Mov5WeBC27aL0i1bV8jxreoWF
JawuX6WP4mRYLhU9PNWIen65BAsOvDzodtF3A/qqvv5n5sjuRZN6IGUtVda4KP08
K8DsgzVfyXqZ8jSIRBuWFJu2ipDTYNNR5itp+UVh76DTVuQeAHGr22nuVMdEF3A2
F75Iph8lsGIX+P7iKX+ENOYyU6K9ivLh2eN193gq4s5ZhXcZs+pR3ffsfMXda9gB
nfbFpEbazqTJMUwcZbee4m/+TaaUw6dx0zi4p0VdbahFyziB+nJyum/AVLsJIRV9
W0Fi8Nd6bGOAdKJfn6Sfvdm9eLPcZo6fjm2LKJEJqBeALLnw0hPN8z19hgQKdPCs
lHEW0hY3FgBuWPqpNc7DnrVRgbR75gicLreYgqqIyF5TJRABYHVml/+mVzrvPvi3
12OrHsoqxaOGpavP5AdksC8kkP5kPs+UUSH4aCNnpm7e8B6NYwy3lZY7K5QxyxrQ
UwoFkeAAU9uColbTXyTlxvD6laR6vm16yT6qGYdxjWEOUnkd43spJghHnliYDDre
8ysPqNxWS2QrYuA+DX+XK152Ks5u4lXnKo5Il0T9rqLx2lsJxkUZWB7mHipbFoqw
CixZbA/htzBsR4h8ERlFZ6vfBu94J9+sjClKUYwlWXyFYQh708QSWJxd60EmPDb9
8P1e75F8HO2dBhWgeY458bL78wdIGr2lyhSYVlF5qVnxmbEB1J4JIXPC0HTmZY9l
7MEHerj6ocWwa/0Z9qvaFO/6BJtK01RrEeWWuyC556lXJRNyZtjgY4x9CvLp304w
2LM5wH+SpFoCuEfAjNxjwcLfAOtjWSAsdD/El3+jL8Rf8uBqWf5RLthB9YVFlpH5
TBwET9QPfZqnTXPR78Co33upcE9/NiwHk6gvLm1kxTFxKUFOdP7l+Ff+pkDxqLtu
fmGmM2b/Vk9ylJRrJNfucTm4BltEI86E018acSVW5B+WqDNaXFPu/CrtiPurzQXz
po8mc0rpiFKohg9KYrZ6QBIbdjecievFOK8sx6iiqoycPO4DEkpPusVjsdkzkUgc
5PoVgEbeC7+lM9oaGv7yxOIiX9OBaTmGnITUgrZvHT5hnJY2fCPXTFjSC0uNtEzo
2bP2/09eMVYgloOUe0Qs4dmB03YMJ2UtF0wFfY7R+Ml6UaUBJH0QK5nj0J2gin2X
vdk7t/UIMuTVuqB8meOHJFjzYVN7aaJ15EmxLnAIyZ+MfrFLIU/fRQilZfBXbSuT
g8hQxykcGdtS20bdNsMQrVYb+Rqpe94JNMtfJMQExW0diHFXpM7JPj/9QI9044m9
dp5Ywxu1Cnjr9rJfIGviQ0x6tuxtJm1HHocY04cQ7zY/7vF0OCsRBOkV4+rAdanU
DSiX/h62SMR2Rh0cxXAOyeOgFdquTnh0KAx87HHGjwKj6x8VDeZr2gn44ulyWtDQ
a+KkIrWxkG1X6YZIe9olS72LbQn95AWHLFxS/jijKgWXvxWIrkdJZPe/rrz+ygJT
b8mu8kFi4UrtO+/njaVbGpbP07g6PFIqYeNuxW3VcqElEaVOtkJE3hxcB++YMO1N
5OjwSMgHs+8nB4gIe6qpblKXIctQqdNtlstwVR8G1m3AeqIwYetdbMzu8gy58Yke
P6iFSKZk8A3CODlBssXYcNb2mcuLjZdpxaGiZdG2n4iRppG0WHv5w0iAaOvj+Dnf
/bhQwT0YYKEDyJ16SDeXUponBuudN1beoqrxI5HJdsndAAa5yBj2qqIDMOD/3rUZ
ADFjgri47qDoCpvgJ55c0tvF1WkC75JwqCdazebM5j5cr+Nep3vjGdr7/0E7SNNn
wdJ3qPiiLF0Zh3tA6e5c6ZR2QO5GqYN29xev6iLUgPDpp62/S8YKJdQ2t4D6AdL/
vDiHWiG7oy7THIAH4bxQxpm8HVUE8OW0fSf4HIeiyE1qPN2yhyJuZrk49kXv1zM2
Ch2XGm98yEI2eSXddn28EwkZHW/Tel6GctYnL3Qgjv35+SmNJFQrRu49KDMVgQCa
p+khvNpphhFhuiidzuz9zj8wzqP3nxRqTAyeX2fYp+jGJPVT5iTIeJqGw4gw1xd3
hSKOIgJfGW6MdUjn3pHc5QrLZK49akbr/HYeeAKdmRQh6OHGOxMthkFGX00xF47V
JICHnRdsO+cpPTD9h/wr3E0c0JebpUZeNcyg7rKN/rmHz8zysIewDLYPma3S1LsC
EmTdf8tJfFVfx2SdUt86N/c7n0ypTI3rw+O+c9Apfouoa+PMDSWV8oxENMMIJzqa
+Upl7eNJGOmgH3NNm6N7bLqKWT+Ir61tAjGFx0KlhU9x301gXyqbYC5V9wJJCPhw
4Kd/rPNyv8/3HD1pdn7bfAANqobpYlxXuksTDw1c5xjlVfCQbTii3ephV2ferbyJ
Et91YYIII6EhjjWhPbMFrSNidVphPHarL4ulyrZjB8SfdOsZeY+tIiDVdVY/dxNT
tA6uLqANcnKWraylGI0zJpnX4SQeYisOAiDac9qIvnFeiufJMsoNsvir/bS1i8/C
U01PXCv1E6z+u23u66EIpJPvivH8iwzhrQMOHVnVxMKlU6bEnFfHX8u335GYzF2/
eWdwR2VXzeOg4RrrWS00BRe2G9G5j20VuMIMX1hgtbdtqjA3A0eSXuW3mHrvbA3Q
yijaYccxXmFTufGxEaPIVTbt4N/WtIeZ89XmE/GrhKCveGt4D6b7hm3bv94+NQNn
wFIbVEF7dGyE1Vrwkar6Q8uoUvqwQWGHpw29Q4/8wLJ+Z55n34W/2QPfOHJ8DkEE
RvAQOIegHrI+Ndi+8JHdUbvcqg/APRmavBN9rvuifSyermG5kKXPFpbn7kTXIPIm
uB+3xIE2ZQyL3HqcnAsnk8ZDemK9Ml5cibHMBsbcTCuqS+ifygvoMFHagN+UxMfp
RNeFXoiyZG3ngyXzrhPSiIpOoGVm5XlHyCZXN89qwZlleimpaE5fnMJ0USjUYOnd
jp9I7v69SUNn0aHbBVEcv/czfh/JEcwTdHqF747MPO8k4uDAafQHEr4A0UYVSWPq
lh7d4/xXz9p0785JR9Eyzbgh1GMr7J8sdidS0MyTNS1LjZo+PV+/VwBYCG4dafUi
bUeGv2oHqJ8v3EH6buicE1Ul1337UYkXC6/K3XbhhXRfU1q3ZoNV0cX/6R2IylYJ
0fdSV5xlbZoerXDacS2+sipx9YT9XRRkQS52l28YCoecPj68jWMb1w1sxXDc9Lbi
RcgwrSzkC09V17UT6zGjZVEj4RLws5M3FR8wbQnXAMSMQTYVxUKQlf2V55MGxU6m
icF+A2QZqgxwdpRcChQ0MLFSnbXRI1eoQI27xBCpUmdeSGPRatRB7q60B0kgOMed
KAGZlNMeGOSq9gAstFpD/53MrljuNDb2d5VmBzs/ZNE5AacmbVjSYYmky2o0LPAH
b67Q/HugzLnaDafU3wWFE6jCjsC2nPagc241zI8UAwUdmPcxckMGCs+vXSF+2o5f
r9X/KrhUjdMo2RluHPv3jgq/+ImufZmfrfNdpIYBfrcCT+7l4vN4af2327f7Wdi6
SqQZmJGFIN7wZB8ROHZoe+3iTWfxnyq/Sk5cRFQuYJIctQmmJeGTPM1yI2+lPaj2
UU1j8ltB7FCzVG92SC51DmKN4yGbvi/oQKA4yqCwsnBXFe808CXh9let1kAaC7wh
QK2srQSsNm4ALxR7cV+Si9x6DW34H/UTHhSULBD+AeGEYakZRIBMjtwmKYduYKdm
0vjDA+7ulJTFkJNB1wg4MVsFHqFj1ZUb1miO+RkzfcW9LrWmiXzokRoUAej97XQz
yL4fglOzEmOuMRodq7ePJqVwh9zEcQXKTKd4hVDSFLLXITbTXQW7xpWOKkm3MK4h
OgUH/NXJTBP+QcobzPeRdwsIHlPhvUXhM8JT0k0MgpfScxtJ1URHn7u7yp9pGzTM
UUCxjYKjXGWWuyDfGlz7UfYsA0XancQ2ACxLkkHFkfEG+2sKaJnc/po3jw3hs2i5
UDTRlqXtCPgQxH1GLWyikQH1qd56R3+FP0AdcYoYDlNCnIbIzTRCH0lorc71BRLP
ULNeduNEwHZJvLtxE7fXJt8BUXRLCjQ2b2qZ2X4dfoCqqlhsGg4CLqMsjr3VHMey
p5Cm5oBuksEhxZn55cTck6diSMagz9YSWEA2mv5r6UqQajZQK3G/5m4keBhMLhrX
ooxo7+q3Kpt2s8H/1ZUnC1BxoViBqACHByAQK5ik2zq2+6Lo4LoIRSqLE4Oibjv7
TQ8fmtP0SYmsz0RvUNPkS8usAq7ngewTF+sLXKDUUdRiLAuguNyAX/TKeyD8ibxy
d0pGWawzYhMpsFI83SX2eww7Y123e30MWwnMaalzgZfP5uBfMJoLaL7JkalqtE8a
xC3oxj8WKstSR+uilhV4DUQuxNfsOWnErPLB7cwB5LkRu9SH6LsGPcRfGyjiSx3R
eT0ZMJRlFYk+WWXXVZ2CCmu+Okms+GwIoqWN4cpGeHqS8s+k7dCayMv1ICAYWOzE
Smd6DHoW9fbxczvlRpAspVHroPs9MhHSJQe7j/07kE60hPvzcvUMWePtekDlgi34
mE3v3nHwTQwmz1pYPvzSgK4ugj6m9LgkBXONsYly/KOZ64Pt4tWL69IvVXh2OVsA
CtjP0bnPUuuT1vkPU2Aqx3s3WKm2UYuHGiFwsStGgcKeLfQoJovgbbiGFhdNzAPK
nmeqDPZgbANpXgf4qGMSPClGtG6pVayi/ZTx1XGQV9A0Hhv5A8nT7EGuxb5ZjRYB
D1bPjHLdJSoyWkJesv17Ph6H0uu5oJd5MyVcXEKdgQjYUA+Xma7bHOgPEerWUjPQ
7X/vMfBpV0/fLF2MwL+iMENDpJr59OYAfuQ3gEgBz5xMZ8TCXft5Q7Ieh1Oc0Fls
CqKwA0rNcn7thKm5GjjAD2lLBDkL+HloU4XUPbPjSyzy7En5MrBGSlgfhL1mxv3J
EVo7yxJyKHnEJK0XmZjy9AOQWW5wesZKgtffrD4tm8HxiLDEWZckica7BikHo0Xz
ndW2c1x2F191I+wdShig+YDudxQYhJ3CqivgeWeoMnwT3IGU38l/Hu+/w8LRGQgl
RNk21UA2kijISQbi4dZw9+cu6vPY7Yu4u3YEqY6SvsWgxBcxQMXUkkz2aONvZSKg
OgqjC/YHctWE0pbrjs4HTdeI/7yW1DFDxJdaio7LhgTYE4YqsGsl9fEJZN0g+4IT
tuXHBNCeEj06YbSjpu3j4GbthdPdWEyXfT96HpfxvRYnTFV8zM5QSOgwxIDDsi8o
RdTmvEBtVJGUXY4/BDgTNCPmbAmuP1hTGW78yN4Bmt7HrsuM2RlMHIPtVMB4YAkA
1r+yh0yO4SKwBaP6U02uzDk5BGKxfTicb1F5018CLI9sJ8ukTCvtMfCSJb+uTg/N
8s4xWeekuXIx4QaUdIywe9Rt/4Hr3vOqmbm8y+4Gm20XYOnHa4mVX4hgjwBETyVa
hXB1pC0N0lvnnZl+D1S4VmHkp+uiMlA6V2Bdrg/pkZ7bX35dFNu56Ds+Z33JCZbK
+1Tr88S6RwSbs1+FXV7eVR6aI8pvk7wB1/IkGPzk4z3cpu7BtypwOqPZltx4i+H5
r5hsmjnmqkjdfwbyTJxoTDt9aPHuUPDTD5BLdFDs/jNFKF/lzSKW7Ru7/2KRpOcO
X2e1VzNbVNXGpCLm9ayD4aGEumAkG3b3nvsHd3OOgc5Mae/B1enmlkDypT8856cN
Tg3nwRKsHghgwT72Zsu1kL0o7hIQhad0SWoplLirLpklFMH1FylfxQn+j1LA2y3l
qAziTMAUQ6ELOytg9tnhuzhvgojez4RXIueQYAJi1fVt9zxhogrs3Lor4ktrjW8+
G4d5ugIKP6vknq5AocdcRTWOyOwCAOIwVRen00thzFamRsDYqNrjhLVDgqMwBhWP
SENv7ip/xFn2VfiTnXvV75jQR1FBUXYnKJr6dsfTlNvaKPsVrBROh6KVsiKGj4bj
vhio3Fu7yZbBqnheQfGL8BPrLX1wtj/Zcvm8ex5NwMm0nYpfd4ZWEWyQJQugkwc+
vvn8xSJszmGvqJJZwTJpjy42RdBwU4FHiHOOxFAKSaq7ZalMIryYH57rxfjTuHzH
7luSzUmMkHkuNASQduzD34ar7xneN6VZUBSSEk7UVQeculj2dvNyMVUX9kxKD49u
kb85iqsiLozsQhr8iWirhxQ8+r4gHQ89n059mqUfID4G5RABoZ6kk9n8/MEMDwxa
g8Bq0VVckjzZevYEjDdMKR3qEwTr38jeac/NLvA5Rw6A/nvDTr8UwSVs77w639LH
hTkIDqNDRnoJPyLvgwfNYtbTauB8Si/KBRQ+clmbaNNlIoGnJVRi0dFD8AOaRahe
BV7SBrqwzjYTOLGRLjKxR1BdxQ4v8btHuuXtkkfX3/VGHC4bVZ8AG/hGIpov4G0H
aL2CanI1J7PJjCt9YdpkYCNZpTdeGPM6Qf0adlAvYivlK7vpDgOmcsWqs1zQBs8/
pxvSBzE8qkqPhV+SZHXMQn6QSativ2HWuU5AP99TdDJz4RyfLPNqO35aBCxwqxYp
3eTwoGjGiKtpyBroFp0EbNSwIhTFdDcKV1tZi+2cyj531UYvBufty9gcR9zjWUVr
mF7d2jKgOOX3xbUWzlmxaRNahJu8NWxiQD1aOKJszIGc6zvsdHAbP1B6/9rHzZtH
7OpkMlw7/B43OQro8gEyxJOwG0mWRdffT53BfyZDy7lMBmIvXZN0PM5EvbeBw9w2
I5oexQyL5j5/dTd1w2nc0h2a+NPEOi0B6lCC3Ywf340RYATCpYoTZYXIsfsu27M/
H2I24fZFgH81orggUAdLKCjN2HY1OOL5x/lMjlTrBQyfb3G2TW9zJCvWct2bScM9
tZYXbWil4tQbuYi/KYdFYjF0YWX/zHsGxg/JeL7nGUsr6Mi5zQRbJHP4BeTZVVzj
LNmPEjSkvX0UxyQeNuKxhClDNw/YlAAZ50uXg0ukxoZEZKCC7lZIjfZZXO8dOGvN
dHWX8JkONt30iCyqrTtP2+iyGb9O8gIT7MUHfhRqct/oCLm+iURcZ0uC1xRQpTkk
DnBK+SgfyFUXg5DSXAuVrWr+ylQk/nO0vSwJkTd4zH7H8+Q1uWRgJ2LqcZSjbaxU
en0Rh6n4mr0ETcjAlJ9FSy1ToVSXfcy/tlg7BZo8EUSDsJgZ4Ed8fwLkPp4heIU4
0z31pTeoNOwuIHY+pO/rYQgZWHh1UFgn/KHtq5WB+7cZOLvWULKwueb/fyPNofW5
BQtIzIMo3N+4Fv2dmitSQROE0ZYUGdqmiFWLwUf5+GiVHmVWkUWY9gK7uUq7RHg9
W//X90FSm7uEEw3r2veqn+dVq1MjjAyolBG3G/x8bS6ZG+K6iWMxeNkkYBEiuIYG
y0om46AY8D2C9JEn4b2UQ7lWwBaLPyDTjOPQZnN0CWMwPX2U53DX3KIzT3wbAE6a
sTJ++q03yWaJLJtb8SsGbaRStIqLfZyMF8/H2dGDkaIbhIhj0flx5GdqbbrB+PDc
GqgBOc+UNQin8Iwib90jEW1Tbx36R0Xh3+oZ71O40J3A3zAJP/ao2TKSyJOwFIJK
xYGrB950o//Kf/GV5gtVqmgrREECg00OC7Y4MpJ3wW2c8Ut3JzrpQbt+hh4WV+wE
cpxB5R6z5CUuxTonz6m0pEHjb/UuO8JG2e8x3FudI1eD4UWIcdGG9UYbsU5pVPLG
JQyulImNApK2UHMRkXDVsC+6T/fd+VB0RDlpgkryHwyL6KKTpoWEk928NqFclnsZ
AUNi5beJNyQ2hhW4Q7K/XQ6bwUPyodIe3gKXt2NnpbU3fi7XQ8ikFiV1bpgaFOL5
7QkURHtphbxckd5DA/rui7gJTLBP2CPnbqNhvQsugASyh9jnKd1FxyLGpLuX0WME
DvJZ+vfzERnFD5bgjujjIsS1jLbJLQbIL3CnxyZeUbHbIMTwetYQFFnzhi5ySQ0Z
VD2Lnt2/NWCf7Csp41udN6UHyRhwe6T0xQp9mJoCPS6HMu+c/aHaxCVhKT6NEsr7
cYWXv7TM6TOLuDnjX9SLIYcvgb5J59S4XsptMD4g6zzGj8AA4akCY9K/VMHAKG0/
Co/KfMblvrFdVUvmP3jQUW7EtAHIsTGDfnKRuMDcM8JidM19pSduVOXn0dLsxbTR
BoNFWe0irUrOd8O46LcFD6CPxJ83607BZVn96dYFiR8hNNcGcMJgUy4K3swm1Hia
53i7llYtegB9aitoeZ/SXujdW3bTkOBYVdC8i0LctmrDocWPjIITCbvuDGNJb9Vw
9rssJtgF/9yZLvXVKrqTyN8GJh4pDmeaLc5zLYKLR2GM0vWBX2/FJ+Y4PSDe6ume
Ole+xwvs4Kqu/0XAgngGQCAf2ssL5biwvvi2TZk6AnOahATQasb0AdhAoRVbYJSU
S29iSQinoCEFDCpGj5D0mJIJzVHbRSY4iCEo+KCvI/7UgeNWLh4ZaQt7WvVgYdZo
CRTyC4lYQouNPQLoCOfYd79XlUQhfI14l9kzOnwaodVrZbu39av2Pj5bXDhP8gMt
ITtK19bRg9tfPQg7auW4ieL1yYwxJfvNxtRDUrszPSgBsu7+3CbGVp4GZ6NXkamV
/CAm6F4pFl8JFSN5bhtV2pe6vZk5hXCSaGe7O0IUOkvU3HVpFAbflsF6p3vcSJY+
XEgBTI/YXbrQAQdIbgET0Op6562aNyGTt+pChIqGuVbOaY9UDhdLePthrChND294
E1dXm33vklGcvqMCVyk2amKf6TCe46RzEhdAPHn4PW+9oy8iRpF9TQ2xPsxjMBpB
/SqKngzx7X2imbHOaBeR09CXRmwvUC326nJ8t30xp56cSJ6cQDDLkOOtr+vzHiYn
hxqcbyH6w6+Q+0Hp1wkCwx35WnYMFpJwDgJlk8a9WFcwfo6yo+5E6mTqRvmlGIdx
xeO6vf99+kWB+NR4z6BYv0GWL1FIC29Aul1q9WqlInloIYgc0sWgm6mBIOwqXnkP
9mepuZ7ZsReSb/D89bYKQOdbaKd/i4yu6OUHLUuJSJGVXVif3uEEBe6SJcP10n9L
Txt6EyDHW+oWTRoo9o64ksUaUI9FnMf4lUcp5UH7zEdUNMtZ5c1Z59ZUVYEQYUaz
u5jrKK8a6+EWvPjYXehO5LhPLD/YGBBtwTEpgIux9YI1wLE/aqTBwZNUm9tswiob
VPZau1YiORBOu6vofF8jb18NundNocUgY1eaKr71e3fDLI1yboeiql24ml4KLnPq
SVi4zxuplTODlAE0WwXOOLQ6ttCzUSxn25ZvRjQ3vyF/ePQDhJ2cFgokEMPIv/yC
udxT2PM7Jbfh6uZZfjnpbtdZTtB8h8+JvvpxlwZN/sNyn6Ei6o2MEPwvYm35SFZi
6DC11Zn3vcAAtWtWrV4lfbvXZriW7plX5CMu/iF3Yros/bngcOxLYfeC/ammUgl1
xolDBT3JHrzzCWJdoRr0LPxDpwu7trLYyeMUSbEYr/mJYwZZdFwuO9zdyJNAYYSC
7OkS1voPMKz9Y6ocCNx/vewYlizuVq1ZZEusx6/fH6NWADUC0lIDfg13HzGxY7Ez
41/r1eTQnsohU72D/1Ppyxn/Xv6bV9fyZhNwOi8m2HXtsRPXBFFXrC0/vciDYdNe
Pq/amKiZLXEO0q8xpfJWV/6ERY9yYCuzGz2WL/9QB2ma4KuV35YCLMbhgv8ci2WW
wuxkLLkxjJ6/ZnPop+bFo1MXvQcYzTHmN9JTkHskNEA0sEwCpxsygroz/bSbRDJK
1NY8t4uS91ZYFZKm485SvzMZzeV2hVjqFc+BphA/4q97o9ZXakyeMHjZ/J4h2D3E
T5p4rwo6ZxnKFIBAtQLTv/m6XKBS1tO9Z0Kj68mTcLoMH2AQ5xDSuTpNQDmjpnEI
qV3s3S+0t357Q8cX1SQNViTV6GU4eajbK4CaK/+GSzS0HSgnxkA2jIfsPWusNHv3
JNqsm5LPE3lLhgzu+2PL1dhckG9J3ay+8zrBVEFKBvQXu3pK9zORYyeb+r8WK+WR
O723ui7a5ElpgJXjoJPViEkyy51LQjytdfFDYeyRkx4t6YSuld8VEGzmYtPuVYlw
XpgAZUdUdZT1tT6AoPKW2FbrmwP6HupiZwO/FG9r/E3r43QyjuESHnx70wB4z6uM
T3vv12QleosJpBeJZg4maMp9SS0Rwmz9FuSXCkb7OJEtYZJYrxPOu7KV5p4umR0o
jTWnulm+qe8vkBz9445SeYnngjgJteBxCx+tATxgOtt3aMsZ4mSdFPZGDK+7i9/M
SMjtHfT5IpE9t3hjt/RrxfpeP1rfRpvPpXc3GQmNtw13OLn6BiK8mjg0wNXfKzBm
4nWOIfBUc2Soj2skyDb9nbjdvYieVVWkHjkNVx6BS10aHv4REu0UTFJHEqzRekSV
oRgeMstsQD0APYbLeIYVFtJtANTdVeTECkx3gyP5NGM5s2GhljFtsIdqE5G/oNwZ
HUvr+wgYD0uxNy43tRk1I10Rv0ahtAo50GaKb44EH6A7aYPr6MPYqKPLqA+lq87g
nFvJlFjSJXU13DmQiGDbd/2Q5nsU9C9GiHFpSyrRLYPG542LUIW68uNeS9zJoA8U
eoUALFjWwrX9YcVWPvxPBN+BqMkPw2Tb81CHhtzwaIfx0/e2uOAJBTEDKiB5EUrJ
R+N40qNcxvvBnTyDk2YawdQxsrHDsslAjuyY/ciX4kuqZYiO5l8JYweRC9v0He8G
Nxj1dVfUYrL4r2iZuXYi26ZGevbBu7Tdz3j30sQ3BXWQlaGQdVO+Rd5S/v9V6fMf
wGH6PwO63SOdE5ly+aANKbQBhBJYqXaqb+DdEeLleTZz89hcDgrOk7evBRfPvOv9
3xRjPGo4v81OAibEk146lgPQcTT8Hl2l2B++uLBGnq4cgVGk4d0B1xwROgboGkbe
YrqHm8jycy+KtpjUz7j3TGhZKnNrrcbpqfgZALe3cOC8yoIgoxLutYIXbTm/WBqh
i97FMPLTgC1a8KVoGmMjfvgU46GOWA//W2+85b4U2RWR6L4+I7bxQtxd72yo/150
jS8C2OEBfIWKvUTzx4OR/srJHDp8pFSpoaGmy2fgnpHaLxcnmbxzwdvk57m3nOgh
es2tZJdFZx2q+yNK+9J1eQnE90+M7dDqOI+gPKb3vVkPQJFavjLQAzoA/q2usJSi
K+zPShpaucIplQiRzhGEHEwKgBGApYg2x+sl+/ZxiSwj7DKqkYL/RnXXSLQzcX8w
kBV2CP19nldtpHJgjPmzrCqmSLqp3CheoYWimAcJjsGa1UAVFw7ewSG3valkHIxS
9wcAM03hXPpYiOybIZ1QnKr4FqsIE/R/AnGq/dFhXHALnk4yA1JFWUdygtrqTpRO
7CuxLUveRL49qzO6EmqXrJhxZzyCTkBhOa73WxCks/K3MtAVJbNSmYtNgk1G0Mux
dwawyUxnsDBVcj99ZPRYt9OlghwlUgfrAJFQ+v3PW1Pv0jH4TCJAeF+seGm15YVY
ojMSFJsXE8bQXHWrLG0r4CRKBHBruZGTx9YnMMtxRxYrsxHsQJ9kboEY0ClrDyrL
LDIrvrfVgx0atsKdgklVkaF5Pz5ZNtMzv+vHwjyPdyIaOgRWyQg00e4PRyrwUt/R
7im9L0rXboPrA/OB/ESCKYFsgRxHek0XbfVuWKAnlRK3FTXPZJFklqflOy4RIr5s
4KWKC8lMyILxJOn/4HKLbkCV8ryrEpNF/oCDURvtIdyQHGdx4zX+xuYHyKa9Z4Kx
ZyldUh5vj/h0aLO1CUssdUpkQAOdtSyerSF59+LGOG9J8wRF6xGDXZYx+cxx3gVp
vFCkyj4F7lVrZWYF20GuLsfaxzQtcE5AVHfo4AMKRy8BwCYD70U6yxMZS+No/Eyk
ke+GjX5Jttw7iPNyCd7w1QbX5FNQwJUxBTQz733I2cd7+dMtDK0ulHXJjCvkqGLY
X8xMioM3ENhZmkNzNi43NPukfAMWMDqZ1pIPzOyiV6BpUZ251IL0WimHaCKT6dIG
U/ZCihGUJ6fuwL8TFXykJrXQ75nUmUkVl4re83wsNXvV3X9JmT6mVf6PZIxnBUqN
O1m5hZHIDNNJYa1j+Ur81dPY/FZYtraclpzWK6VKXqi8KkqsNSm+MI1KqFqqv4NX
RiO9eym8jPurjk8e/ZxdtB6i6hz4XHs7YZFLG29iSMALP7bdcA1oTeirI4WY/Pkd
003IeiHMdc1dQsGsDVAoOjUBWIk4zQ63FAFprz1g7PVqXPbZ0cCB1UaR6r3NC8ag
JqoUm2jvpY02JGe5NPvObUqj9NhClWytSVU+APV8GJi7oNIyVyhSFEH0u62k84cm
DD3lQFRs6dDpIie9j0ULYBemPUELJy10AW2Vgei0jEH7tzoje0YaTzmqpmWa8EwW
qfjfbS8uiqRrXdfifI4/vYZIvgdPgA96cvz9vbHUIH/vgXjB2pK9n7t76SprDSWN
hYkT8kXn977MqJ8ZkQqbfGeWVEDmKNFn4CYFUobAgeUyTYY4nbSYhDROofW18vB6
xnCiH2D8i2XQx+c7YEc9UhE9D7F6etU+2VKSHbOJRCi1U0hLq64CMYp0COLXzm8k
nAwUsv0O8s5B0iANgXaHDX0ja6Ia1RhLDpJzMwNhu5XUAiNB55kn/eWuXbmdpWZf
YHFSuGuVsTgs0LHeVDp9Z2OyxpNuhXZ7ucH4mjL6KP1WDBucL+BUGyXcYFV8X8su
p/2eHHeV7T9OGPg6EGUEus/PRmevgNQNt3TvHanbeBPrtUutxxhRQbKVcDg2hQa6
1PZk4WxbHMjL9l8A2UFDTy/euNlozuA79SpbaVhCNxO9sT7lSufq3T5Kg7iq74AU
Qq4BlnKuQjrRxfGpjAmcTqq3ZGGFF59h0cWmXPKDsFD/8A0Slp5fPhxPXyHGhOlL
+kDbfL4hwajJtO8hS+FrJQLQTwBwqWHNF2xvGqhaQkepy/fHWtf+w1j0qlYcIquX
JTt0Savsug3SWajcUjf5/maHbEQb0qaqa4t0SFXenBs5VgyGyJtZbX9nUbofMlxj
BUDPmZifcT7mJ6gjRlZN08VJ1uDy+4hCcZGHv6ZuXBGC0ahw/7b5RsaAFrJ7X2GB
TzweJuPFBdR/s7Yg71ezlQbJQ1mePCK00XgqUpdy7ZDicvstwvNU5dnOzGTinS86
CaiY8I+p4EC8pYkxNnQ93vd92kQHBuSZz2xwlXGI5gWzs9pJsIEE1/fvIdyUXYVl
QG5hk37da03yj8uj9G6NmPtgOd3UreveUGBCuvZtxZBDFNH9qz6rdUBef45OJ8nU
56rQEHu+69ZBXqn7bb1JQA0R1l9NUw7/S5y7Syxysjw/g1ET71to4/B7XIcaNBgO
y8yJ4x/jaqHJiLPS1GtMQsDAstFgaj0cxH2X/93oA012hl9BIH8jMfldkkUNNGoL
Q/FFU01zV5O62PkTNkzQEtLrRj8awBxEBIjjYZtn5+ZtIvutEvdjtEeMiVASwrBd
bo9ymZgSc228zStekY7W204lWwRxP4VudnwSIXZ3HSNErwdZc4BBZii5zxmtrkXA
Jhyr5KLDOWQvWHVwFPpYQcy0YrhPSMpke9YwSMQ7BadW2lcZhl0M4frKhcx75E5y
Hh2pFvyJQk5K6EbrPqxm+aYZe6KnM666e/FUSgshvItFE7B0c9bL+jTmTkEir9BQ
Wo3b8O/OrNKxaENdclsq1OITRQAYuqyXyYbGhJb2gzf3rTcTk3vEqG2S3w6tdhpK
IUZiWxnKvXNbgWD+DUumLED8ow8/okjcwgkXU5CpUkI0zuLti5nzimxE0yI27PZh
X3GwYwuaWqmoAM7u9ZLzzq4By491B7Ux6s/JSuTQpHewn+aYTMnmZbd3kspE5TJW
zPqz4Tw79QQ0BSUYcFReX8c8G18MvGgALXwQCDIX6OVE3ptytbzNrn6KEc+eSCPb
Y/AgTZSeZcDADCI1o1smuzBOoc5ST/Jylb8QKXO00yRWqQj9TM2Dur31cWIylKeb
b98kj7d30h6Q80X5JhdbwikufEE9KOKTIehehge1ZIoh5RqrmTvZMWgE92vpNGsv
iqX/OFcuIO7/6VSHoqqTmFMTJwoOaxAgTymp9qh/0SAzq9ipQ8007bwsyJACpqOY
Kif40lHC8ldchNlG1ZepzO5RyEWD2/o56VJCF5LZY3gnIHb1vyxambQKT5kITZeq
IrJ/ZHnUwh5VHNaUULid6RFxAyYJGq7bf26zWKiN2Vaw3ffVRFvPWbgebNOhV7Jl
L1fr/a2oVcObVb+54GkXY9FOpOPPbv0EwwrRRZ6RbVZYJboh9GhT5lt69vTFSc2W
hhTuLfc8d5KlPvR2aJZmscuW3JihplG8pFsJTyRTq1LH6N1NpMG4tLA0MzhgdKIH
nGBWRafE+RIX3pkHJ1W27kAYPnDxLzOtOVO7HXcFmsm8fZu5LAYbd7pIo3cM53SG
PdoHsEdSI3pyfF0XQ9u7BUQ4RE15v2TfwoQNGdLYkfkxW/61robF5uNBZdUHbx9t
Q6JnInYNvs6R/KrZYwj+Z1KuRP6fTWZsJjMYhB+xj6PVpjjBbcbCx+M12mijqZgz
Fbe65CXf5EoIJ0nscJbw6eOvlkZaHT4xPy4uS81Nz0EN9wEdJi40rXXK9l6jzXfh
U0JH8mP7WXn7CoZSv1M13n0rI4iQW8J0tchgs31Udq9e+KDQHSsyAfj6SdqVwfYO
yDd34tc4bADoG2P3fymoO7eliP5Es4Q1QbWAVS/60L26RdvFRvTRHHbQ+wknf5u7
A2ytS77w5B+v3gYqReBYiO7I8sLHeluRLdBUqwZEbm02mRoQSzlEPgeQgNg1YQ16
WcMOCaZby+Ufhetv6rHeyYDyY7iVQjhweGF+IzsxqQU/U2FnSGlO7kVtrWbJDlMV
LqIr/ml3VtMhGiduD//JaGINcO76rV78G5VUVNfoEatZ4EsJbOA2SmnKaM4VtZMH
HOtbRbnWy1xuq1c1Xh/MKHSClYUnKqnwsxIA95tFs7uu7tgJDSD4j9Ul7rhkqJX/
m0OOkqf30IQBWWPRFbQp7UG6qomyIC8jUJ2MN4fBXzNGnlZlcVWBXRNLuQcwv5fm
z2p/+uQDZJNnudHRWBBuYvdbyawm89IL0N0bt3LYTOnPaEUn3l1kbYLyEE7u9zsD
VklNwICJ00oo2YgacA7x8hsB55XKi7MknsLLetiSflbiiTTexVUqGrsMy0e516cZ
BVzuSpGWFrmiJi0hFFpx5HD6sTRX6ZKVu+XzD0tJX4vsoLbll+mTGS39tG9pzfrp
F3bR9N1oNsjbYJdvXp1m6iwViTlBrZjKsGM7AbbRSpyKHurkIPzJ0M/bdoxPJUq1
zI6M2rZAbL0lGzNAd+5/hjcDAKlTEwhgF+3DYaZk0Rf+aXVdkATus+8X1PnfSocR
qv/Qg7Ia3+J3Xc/WdGa0M6A2lWfprTkEGD9taw+nANNmzQUd860akAL/TNrVwqV/
mewkl1llZJKwRO0vt2iR/8WHTrRCIO4KosO0W152ea+q4o/HaHsBCsiQRYhWjzHp
qMoOJNUbPsoWkty3Ai59uIslkDEtWCmfWVJ/6gpp22hExbM9XujNBDn34iVwYg/L
+JeJEVOOtCoaSdV466hzONJuAqKccdE95x7bH6oAVoXeeaEOdHxhuhKuB7EYm4Ri
5w3sFf4R4NDIUrnVMGFjolKm5R9p40MoL1I+6s7yLJ5ClfaPCstYeCF5aKQQWaUt
pTtCdkvVR2ZrY2MOXmhvkPZ3ILG6pQRQbJcpIQB/6gF3D78c4R02ETzHQIr1z9nC
m5s+F+rD0Y6coNR4mohF+qSAH8TgjZMAhanobaghbfS09Rs1XuZmvoB7Jvhf21oi
JMZLt3VhmFKt9Iay0JolE+hQs9M4Js/ZWQj5KOOwqUeEHJAjzbkb8igbHPdXzGD2
8TbBqxdGua1e/VdMFU1t0wHmOM3DOQWbLDEZBQ6QmsWhcpm1fvjvOkNlppMGSIg0
ZihRJcUK9GLIXviSGQ3unfScT6bXzcxuhanxOm/0BVnSyEzP4kO9o+aa9QAimlNN
q0eHbnEX1ekbNyRrR/cPfiIyWGERHeyXgKvCuJAoScy7TAObAlzZDIysr+EGpm1B
IZaocnRcIh1l09Ky43yGRXhoCj/QzP2wFJbBCiBq0A4RepPNJeyAl3YOvC3hvUMZ
dWio890x8uWU59v3raMNwRdQW+JTzfwhfUU+00n8HKvlpDJmNXTnh2GVxdb8RFbO
XlMJLqk/pa8ajyrqIIJhLTHWFyy5485w6hq9Em6Q0Hp+iKZZtm94+1dwdQ86UhzW
1cQ3ivFCJfOkVgkU8Jw+C99y1AHmfLt4IkZJYyEYbWJHMK93eRYQoAE1nNd4GtGq
vU2s9iLrpKACaXTHYFqec1irEMbbEHC+qm+avGtZ2WUirUXCSkryJTZTRBC5SYby
nlR+ReYEyaT727ca218KoO/hdzkcGCaG60G1iwFMAyxUvYBoFU5PWauiXrE7inln
uumX96bW76QnbLu0XaqOr7il09TEKFbbW17UaogJESp01xH4mt9+ao4Kayk/GH/t
HwyLjPnaiymYTETY8dlb7wsixBAchtUOt+G2KiHYSsoKP2+ivCVTO7QCMGBxDD7m
xcWE8PCRrSy/i4tJyGtA2VcYUOBrVTJ6Kd/dy5T2Fkae5Uw+LFCXnUs+s6dBEwIN
ltE/jHT03uv7LhbSqvN8KMlp/mZLcrKUeNrcehVfVbNywauijZAYoRiNebV6jxso
xTp6LNYZF55awyrVVDzije0f7j7A3cAkAV+xwE1E5LeSl4hzQX19AER0JU+ZHleF
RcbJcSJBv0N53TToIoSdIAQPU4m4pDJajCh9j+4ptwcDbIctezBOT6UJwCiKM3+E
iwRe9HkFkelnQwl5YyjzUdCQ03BJiPfLaSRm6Q032zT9BurYfKBD2UgW2tQ2nZhO
j+Wv/xK4iKu1Xl8Jafqdt5tGPY696nqBQcmX+l8e9JMt7dXrwSTnlA1puGBfpuHj
aKzM2HrolwYHLSMkJVT78rCIgKTk99I8YpY787oH+1s3K+1sG3jPWN/riLsQ3FLu
eL6M0MqdRVfpdlJhvWGz85aWTgJ9HY1SKfuT/eCUmLBKPRcoWC+66JI3wAmBrcT1
Gu69Tk7bpdcqyajDz64SOAHfCtcSINGUOyJnOSjwHSxwjfTU7okMWuOB6FvIu8a1
dsYuCcCfSM729X2roWX2/ToYWmz1hVQkMhwtoo/4yhjxfAnBVum/uAoCYzeIiXfG
ycI+uKdDqIkF+6cCWUSEJ0QNsZxcx/x3aoLTBFjC4nDcX2br0+VHaitfKAXFOhF/
QEQl5l2ENrTDT1QWUZPFW1CzpGZaF0mm+X0wSOZ86gEw/6jvPad41EPdD8KSuu0v
qclDKz+62b5vhxRomz/BYWGFYtY0n4UXM4eoL8YFZYa42xcNI+v9kCNb+oPVcEva
Z+wXaMtfvhWLJm/g+ZthUwsAddePrvDQyHOPocGrQcyHrXBwy1Q+6/GIW2kR7rEL
sTV5B/YkRT7/VDUijUyi+vUtmLz+9kQA7YAVTjf2W+l+PZ/Wjx+nN+MGp/PQf2el
2Yt5ZicPIKaJMjGH0U7cfExRbdYGOwpbMa09VRBaZ1FRlJSV7dd8fIt26GXjbY/p
q3uv+6ZUgBBpY3GiP+z37FQQayUPw/6Ix9XJxLk3BPo619bIiD8PY0d9AJlMJE5Y
fqLmqeqWApuzl09FoLlxlMeWXLxDKMFtEoDBKxlyqmWJke6olHJJC4rXr0UQNkK8
ojDHZANLC4tm/ZU6wnN/LEeuQ4vTzWYwhiB/5b5tAFt1jM1qeEeI7xnKy6CVxv4H
9+sDBSJcRbZ/ugsgtAz6r7jYAcxWhl2StT0wULQPNG4OrFi6iT4PZ3lUbJTPOW27
NfXlgLVzmNWqYC5tsmxWnCOXFvEABQtKLatBhS795i/7Rav3G6Fr2d4bD0GYn4+I
E5k51fnvQVqXSXA0jtTbAxTL4SIAiUFc2Mc0W216M6vq6Yxkn7wKSiClYtHa/3g4
r73Q14J8CtuYOsMstSw1k6QJpkDlPtzJIN8Adh9NLVn2c1YX3WQ+fgu8ZwkviUdA
rUrD+92iQzblespIzL1V9wDWB4MwnZvbUcYgqPtANz3eVsovFwuVEOLsLX7t+76+
qBs9XjSPfkhAKrM8JaR/kWR2QdIQp8nfpVQsm/MhpvhU32P2xjZ6CBuZZiY7QqAM
sn/7igOHhgNiltxfWH83rCgKY2pXAYx24GQ0IyioQvcYeV1cjXq0Q/hatC5A+NDA
24O7P8IGDgEZ5xcx04X5CIHP6tYgpfkDawXXKkMx/mhnEyS3A6fzlGkT9jUaqcSf
oy8Rv/Np4M4hxMzAWixmdsYQ/hDdclh1VJtgdhkYjCdPMMtS+CZqLE5ea7bSQF90
XnUmp1GbxCK2SFRG60ndB8URMwDYiza+kKautY5Pxs2EsKuHAbPbXLLYHLpt8wV/
ZYgZv3IPROyq86K/RB184W+NgqV+Ci/JJZTYFhCiUbsLQ0TNUca8Yil6SkOykNlI
OpXzmwKtnpe7f5io8jC3LW1ZELkyZ/SJpv0rsf9RLeopU8kL6j2YAVYwrWB7Gr1Y
ZA9nDOtKyDfEGFjVddNRD5RKgaMg3JC+4a8xj16u4UBalkLqpnJphEM5jga+D43i
icR1d5acELHpOoedeYisFq8ZKntlzMWQ15OYdsdWaAVyWaTpSvp9Rv+MzaR0Qnx2
WpeHpd515jVf/QtCszqeONX5i9T5Z0lHb/ItBHLZJ0DSnQKGyijTsCgsu8hx6WZV
G8cmsGRP0/W+YPg7Jyo8JPMgb7A9FeYLn6psk6CWpVZHWAMKfo1ZqMdpubMz9Tl0
SSqKaPcKpBpT2Yjn5HfLg6H0YfuRyse7m5x8ijHSz3QeVH/X+COVJfDmLD83IAQ1
+EMbkm6zOoxCAhuAga+5JlvcgdC9ItPhMh4FcS4YV9On+n4U6DbZcZCF5iTSWq9c
WdkG1FgYjxAv5lusEOdwwktT1J0xHCFWgyPPzX0jV262YhGRO21BgdHe/e3gcfE2
GiMSycV1E+29SNFyDsSV+u8bTEjiWBK06YSBy7qhL9ohvbHLwytPDp2klF0/wH2N
H5zs4DVgneNKHhJeYMpa7aWXE9jeTQM0XmN1Yuew/rHzFWoL7dAqAtZh67HU41JY
5tBmRbeCi6h8+Xrz9jeWQc6QVYb2cvS6dDI5zTPmtTtSICav2bC0IxQdcM91RZxQ
UwyljlBYhubCtPTedalgNwW0gm68GBa9wTWknL6PFJkjwIxPWx7B8kf81JBndDJT
qxFa0Z/YNTjUkk4lxwYL4J7Y0F7ZtkMGSKuGLkBmRZLpgwX9q32t4GfTy6NTGn9d
WYSPvXDXbUBU81S2YmsK9PCQA9yr0pRRUPyLfNWcNyA+msVt6l1+A9Mr0rerFqXv
mZhd/guKjIRdBL5K+38kIVv0rsLtvQf1hzrKkj2BW0/wHRhxbuOj7iiTXVlkk4iB
ZZ37Iqy77D7k/u3y2psv5aRTSjZpXikoGOR+4jfLvcHBzlaCU76VqxlHOOCDfFFX
jbKS2Z/Tsmv9aM0BDxKhDy9L0s+UkyVe1DYdu1bpO/k4CpeTjTuSFUS4pdxouvJQ
dpewBDe9kYxuqS7x7i0Sb8V81noWRzYjg3S78W/O9689tKuUmaLvAsnjCaSK8HD/
HVpoid1P9fr3Zqmj6g0IuMleKCpahnZ5FMDzVOQQpj86qzzpuuMeLxdLai9iw/l5
jNDLufkv2EoueFUhkpUWe+P/bqizCWrp9ibWLeXYljbWuQg7VcMUtz+q0ltlFEIx
U28YImW6GdanjFdQB+IGOEkdPlptaZmB5GvAjaa2i8UQqWT5FukOoD7H5sOt/vuD
X6mbgbaEfUd6w3vNkz8XzSXYb+E4VAsSvUlaKiXTCv/oAsf+pKvR238LlZKlzrZX
+o70hWSdnXtrjMdIOydxSUJdOptG25VOXgUMBlgHy1QabrsVEBesaag2dmbWGAUx
5p/4DneOFHzv5xDxfkzV7qZqANnrIOs7UttaMd/f4SzV07rAmzzJ0psq3jGwfKFO
ZJe2v0CZwxyTwAlXwH5Px+JoZSIH9IAXYrphdsycTEutHQxsG6Jw1EUluiyTziwM
fo7PKDFE7DmZPPm1uvnREbznYahXEL2GRcDwQhlBJ9zr+29StJR78/Z0W0GcRUH5
S93n7ij/CMe+0TldJlSJECyHjhv2TufEXosF1nEQ/rfAX7OjvwLNiqG9okXLnnca
PHnJiZBWW/VGAl3KgU2PRspC1gZGFepDOMj5OZKxqzX4p5ZmpKnQ5lLQ9IXOEguX
kTgnsP3vUvBcucnEt2SfCtv8q70mIAI5qTO+ynOPmN4nEBnF9EumASXbRGl07F1G
R0UzIytyhbNba9QOZ0AMM2PghvG69N8Dd/Z0dhX8HPPp7hTtJw9PdNtXA0Acn3Gy
o9VOUrdsspOosNFcozgYQib3sPzGjgaLv8ggtnkmdH5/BzUeZFbLdmaomUnPdXpv
f9DvgW1on6zSSNRmR/3nGWGJ/aUTyGdGPPA9xF+igvjpWFAehsp/ZGKbaP5W1S6P
VAIJ/8LAolB4YGdKr+kGg51syXXpvwdzvoh9VHnQA/1il9DIRtYXEbKwZD+dTaFG
vQGOfklmSWrNgKhwCfZ6rb2Tm050goJVkgY8wLxAaOqxa5ugwaQ2hg5CMTSGkTci
imJMVPIivIACMuP+bhnin8k2kLYk0tBgB7On8OcaVv4SAchmzyhlyaeuXdRuBxsH
BHGCG3gnTzZUtLbKDJDkrCfuKUIuXYWBppcVdIB0gxyKpOLngGwmDZxflZa9z57Q
QMM2pYoybusNT/LRAj+R8MP399Gom/PN56ZL1Dej+cDyOFn7YezeljyMKo5oUC/Z
OBtpztVt16RIfx61yOFW27ayhPaQ6eOr5cIbV8w13le2RssEgGpCrnnPvftCBDz1
iKLu8QbP2OUkUk2/4mdxnAgB9gn1mAKu9mgc7uCefcdpcr7Dm2hboXgejMo495Ks
5gAvXB6Kit6VGwmoxo5wVBBC5KYI39L+IsXN55KbaJ/QGOapQdYaUv4+8kMCCGsX
pt0V83XBBlZfbcY6ioGscSv86Ng86g+zbkQQPRIqjnUTvT1+qVziJuu9GpbF3JYw
sKOjqRPGuWpx/a4b6Pf+m+Ndt+f9NI11g0eP8wgvnaO3jjAf89XViH3brWqT3Phl
ktjuKXb/3qR1+FWsRJndlvUksQcY649NYJJ55pK9MPxxRKfDqrt9lJ5LqGBd5qck
t9zAiZ8R6N0irWSkz+StbCK3P0g1wWDmn1oSrVu+iaHkSRbP204EDJ/F5QHsf+Fy
adXPXDxSDVmh3rc9bSMBidR214v9Py+8Hr3I8cF1Jb4hxNQizDB9hi+oUXp7c0+C
yF4zFQ+s+iDEQVDczfblFGZC/9EhUdR/hpGMJbemgNRS2ebSOPFkGIaIIi9QIpb+
H4/0pOeV1PW+CYlfKzVjiXsK8AlKoIyIML8ZqLhzCvPuv2biddedWhFHtOFuPOjN
YUudSFvlMZ9RRMze0ilRdgQ7dHOiRR8RQGEDwz3fDIzy1b1x04KV29PHgWjdzc63
VNJ/MP4TI3p33G/XbXdUkuKtW+DEY91TgaWlQpAGwy8jklx2rhYjGfB1p97Spf/t
CpEmRkDFIf759SvHzRjaECUU44JOoKotKPNX24tXcDw9NVcQvYR+cjsCN7CETBM4
OHkcpHBoIXzT9VBcDe+O9mJLHVcVwe3+wQlbelUXdHc0DElWAXKwtgJNWoQ1MN3w
BnwEYv0HeYxKPOM+Uj8KmKFPx/pEtFitp2DCAYdvTliY/J2BLiGL19bCi+WOPtC/
ko/fOz25mloAfipjvAAjScutmZRyjoCu8veljt4xesY7+WOy4t3kEsC53Z3iU0a9
cH9W8ZdD8tNmTbTzTLE0n5rusDOCyOt8R9k6C+gsybvVcsnXLLsjbkVXKOMl6xY4
XMYKH5k7Gm6BFMaFcySDIQ4u/ndLc8c7XzDSHCULyjAAt4Vl/ko6DnC6HZdtw+PF
YtkmGLFv8o/eo0luA1Cgcsz9Zweo6Q4TKWYwsw5XW3gCPHsFmTJwUkMPG/zZyBbd
g44dytnREa5liYJtsk3tEpzDuqmXiI+InmFpB5QXxzLu6dJN5MqToFZDfRcmPEtf
5/ZvGYlNLC0wk0Wz8kBg4M4cNe9F507UANVxKbVzQo9XzACVrPF4RML1u9uiNDtD
yxGpuKIHGeSDC9qc2Sbcsei5hO+RenqpJ7o1RxvSIhkjFfjIlvUUMwb5g5Piue12
OBefNhCLgSl8mVLxFFIZ3giEm0kPSQfLyG0ZpnG2TvZ/4n/wjhVTVMLq8LM9bXYN
551GOya0L6W64Kz28vlFiokoubR1hHY8EyXPHosmZQZJ/dQ6O1Yzqo8IsdMe/xcI
0KFDICmLr3R6Q3xCS+FlEAgLqBCXqBw+BNXH1xqmh4w0v1gcjb+ZPT1s5T1g9z23
XgXScGXTSCO4GQnPjvDkg5i7Qv1cqkbOqF82iPj8dSCytwA+yhnbVozI2VPa37I2
Xw8OrPeU6MpM3ZuJdlKZWU/KkXrze8oGdqCSFwH7SRNWU/7pu/DaFez+XdPWshZm
LhN1NwAEhYsYtddCdkHZ377FG2akAdtENpW2Fa4vj0q4sVIc7yfgyLBUyNW+TEYs
FnqycdQYlWl9hgOMlBwT/lrXpKGNIt9P01P38vpuxp5EWvsLXAm/8Ne+nPjdaRou
8GtHT8ulBNGVXuBIqYM8NnPZBniGfTvnHT6o7n0IiqWOjwXQcQ+Cr8mvcDEvE7tY
E0CLzeaQ1tHI81MDCwJupuKn0LTHmqZherlLLFZPIkESkAQVZzdcZ0kqpDB1ZNT2
rldOUcRlO6Sriekq3R4h2lnHc1vD2l65O/xIaXbmYBBT5jZCCsEt71M6+pePAna/
MBV+F0r2/M0UIRbcAeFeEn9soyVABUrPjSDAjAoSOmzo8BT0aHg2y/QDgxqdPqJd
jER5haQXDPhk2dpK+XF2oxftTx/Si+RD4NARgp1LRX7mE8a3Kb9UIBg/Jvy69pgn
5HQXUsJUabxFMZ3iJGh7cMt0SU2JG9hOTH4MHSL5+jsUkGEGY52IAZAd1aRnUa5a
ebkNyhhMi/Qa5X7E8Ze4ZSzFt71kGpUytw9vH3rxxHkZUxSV8H4wbFYdXocK1vuS
TG1DKTHFVtWtIQM5w/Mil4Z8AoztMeCOxSAUk8kSctmG0bgiT5LwZ2uxYJ+3nfwA
lPXjL6nJdrX78PfJMIqKX8XEK3Cud7HhZXlfocgM/0YT+645AgoDJKlSrQMeiT8F
E+PUKp/lDKZpnJRjC/kQiqNKX8lttSFgIqduouf/ZyaCuZCNGk748AYqmnrPeEve
d+U18UKYbhSYiFq4hjkwdhuaXvVMsiChrxY5gJAcOF5zs0Yf+AoeCPV+wDrj0YAN
F5mX/m65e0tZXsuOud+iDR39l5H9n8LTmyNqOe5wyMt8SoCYrJTHsbIf+Ab3t2tZ
JkbvXOYFnsiaBF4SB6HwPmnLj9nG6bf3Uz09HSksG+9l4lnXZwUV54IYrk/XYgHR
hvMt8oYb3xKXiQ3s/zh4wND8atzUwWQ9AXH5An9TIk9cBfaDMBpRK9JpEUyGCHQZ
67bfRMFRgvxXo9HPHQrT2USTbt4V0M64bzFT7XVeqtIfbF6XyDI61BgXqQicR9Vq
fid8wgFHQyDU+kv6aVdElhDCV6GUAJW8zpH6Hux9bAcpM9xr7X95IlfL63V/34O0
Bid14gW0k6y1/2HJkM6eAbTqKLFOk5Xc5WlrtzyG9ugnPVkTOcNnO/mROiBEQuMI
srIhPw3xU/wgafWBYT/p6JWRLUlbFEQOH4s3D5Z38TTVk+cL9ro+zgZVpjx5w76v
6DGBqdCvS7+xxZLlkYKIRnadamQ+mRNGZLb8D7AfQgviRNJGse5ldeM2a0XzZvpq
yisHNNlzZF3aOCI5u1rEbzFJb0GFTK6yCKfM2+mXpzUyR2kruqto2Ru+7NtgixXZ
CeXjvGeQGr7lqgS0F8FnilLPGdlMqkSPQ+yQuEFWYymG0kFyFqAISONGhOuCHQs1
Mb2CMwoOklyQXt31jUCLyVzkItTgXMZugsQqg3kvWVpDXZkdmAPIvRo8NKPcfgSK
ngUbEVQhuMFQSfsTrZlEMz2P3HGPYwyYIL2IkTGbpSEgTQolKTD1WSqrwPf8CFdi
rI3kmrHydjqAiX1zD2g9JJ/NOZARHMr5yQC0Y2IK0BJZ8Gf9yYwk0oH5ux1ORU7K
b5wpB6zpQR4V5ughVQ2e9UUmjOm7wR+htmdGEPPauEHM3zvQ5ZgvfHM8m+EJWTsZ
2HRwPqf+mQFIDZK3KWq9Gx0RfsXxGiYhLSovWlPfMhiAIfwSL5ZxCL4Q9hki/Soi
VnNKOWHNP368treENUliO7M7V7b500xfHrR+9H/6D2EDAB7a/joE+JWK+A9WGiE5
RCXvOQXXjosyF68MVlVukvsmizWwrPWcn3+ZdBTtcjmA4ZeUkyL0Zw8orG6CqfX0
FC7AMuoLyQgiVLpD5nfN2/zA9q2htEU9C3WC7+DE8jWp6yv7DbmwIzyA5K4trLpL
ek9O/2VDvfCw8qAQwignD6ryvFMbQtvbndAwDW88B0Nm9PToIKYvF42+o9XYrbwB
YN65YVYrcBl3QleDUNFq6WFi6EIcAiuV5UyfDMcjD9Cr3QQ9nYVbQjDwWRe+eoPD
LZXCWp/138AQuGJlLJkiLzbX41QoGukR8iD0iWyR7gwQm5BIMsqgVlJm/p6lhbh5
DEnTMzX3jxYMS4y+sRcliJqGipmn/2gC3J1u42J+dEmYaiYGPD1tF59MIFeu2bU5
2o2QeUUQkTBo8c6lbnI3c/3JZIwp8dvK9kgXSZdCj0+zMlK84KDVhGOqHnqUzmyW
/Ox4Sgg+UzT++Ml4s0cPzeXmDskS9bfMSE81AoMPDfxjEwmIM8B33NOcj/dFzq1H
5uwBMKa1nozzpqS3M9plaQnAgBvv7yEzhlaGJhvpXbtE1fhsq/b0UnPwIkDQcgQG
7FVbmdQ/aIdBn5/7oQBpoujmSfPd5f426PmZE8BvmlwccKg/Kq8NTv2PkTp3jv1F
ohwvbWJE+EMsRuxdU8vZsIFcbhtYeAGKCU98ZhiyhvcgLJDcg5OeLQjFkY9b6xX0
sFh+72aiRrP4YIq5d2iQXUSkyn+2rirU3XaUIpOxTUqdWZmKJAv2KFsR0xINrxPY
hWoJcEufedFPD2wwDJy4YQjpWCzBCStMMiIkrZXYl+uSxqsfiFjZqiRvVel+WSvu
QCZaugSwZAKilVi/0lL6Y2AUqGJTC/i23b3CyT6IqhFtkenRHhr/7buQajnQUuQt
Qd1Kr8vRkLD3L99lIUFNbkyl7qUU4VasQyWeglq36N087ccpX6m5j1lolDHaZVFZ
sik+bloxaaz7wajJqrvBhMT3SGCvRqGQs8S0AsR9cMmkkiLAe+PgM5JzpaP4s9wW
GCgwhI89ZwxRl6m1S6KAVG6Vsft0u+L7hfvgArUqY4vF6gkURZBzHdtAjUpcsPGW
rsTnmFthKrGyDaoeEjkDPjHuCIurrC6fS3O42fGSu5ljfkg38yT2b+y1zWBqi2Vo
1ufsFdKjPN8jjcxWYGASuy98E72JwELh+jJKtOV5cq6GHklSlNdfBsZL2EHHvi1e
aabqst6WVkLk5Y3Qw7t8VAfhysnJsohfWxsPyhvB3/eFOUumh5MBt77ERflI84jW
9Yts+fwYBzdn0kV3v8gZBu8P/OsjElxe7Tz+BViwov+1h+/PPRdebQhI8rZquZzY
ktNYQ4hIWFQW54cgd6V77sACLzzRAOPIvQ5bUNbpo9OOMrQdOusQT0z2XzQb4+WS
77UjQe2la/43JWIgGKtCDF636qc7ajh8UXuP85CX8XCYNNvOeXjXuGBi8whgqNAC
LkE7PB7rgnmBAREym/OLjDNGhy4ODHPueeDc029WygLBeM6XD9Fxi9Zo0/lw+c/U
wZGw8L8h7ixnpwrFLH5xNBZPjTfm5S0Op8fA0icdqH3D2ABvZWRBBQaokgIAf34c
cYQ/CqJ4qtRJaa5WLuCyOAyncaQHEckzcfvE961SZrLH8O/8LptKTMyVJquT0FqM
+XKymIxgRP3fzcMhErPcR8q+/P1Fy3B8b+Up9tPXf+IUIl266gs8eE0P9DOC9LoH
J913eGbhGA4/9nQVqitnIbv5lBOC+GyxmyPAUlWD4H8XdV/lH8hHFn7pXq4P/bAu
LBrh/XWqTojXm05Rkf0S8x3u+E4cpeRzxWmnOIzcLCT5fT0RcFM1zSt3AJU0g+M8
70wor6VSNQ7y87rZua18Ger0ejs35oa7SsmogszOcKnbOy1TV2ezI7SznUJDLp0W
QMz3u9cCZ4WRBH65vRapjSoTo7UeGH68FZ6V8CMW6zIiut/d0ubyoJkn3KBqPYyZ
v1h+pg5UbXYVUdgYb1/2Flc8NgXSmyv2lPxpTvX617ZN6BI0BAuoiFJ1dnm+ITns
WbCRfZ1VhkN2T7tBIt0qwUVuTT2uE0838hy1z60QuZyk+Av+V1sEnh64iCLXmkOQ
S6ibHpjp6uoL32/k6DhYrlEd7jc6sO+khirLHvqF06cRvqobveHtXKEagbmakfCg
iEmYit/DI9PrAKzuEBUzErhFvT9AJgQ3uYhwyiREemGEkZxX3kZHonce+fSUxAmi
xTGe4RfVhRNZzJl6fuqzgC8Ba9wWudVYIOH0PKkG1WuAlStswdC3OW7kN4AtX2bk
af1xB41LssJLmbYuaIeqboD4ccyvn07uIYS405Ni2Cqe9yB8YkYFhQuC3Ip3EF2u
uUhMhZbY20L9G2kp5KIH2cu4ovY/vaMoseFAAVtKXb6xKjFE7Q1ruUSUbKCUHQr3
05TvHhUC4gfsmgv+FZ2TfbIZSeXIZtVNx0CwvpwRwNXRF9E+k5j20hEjIriyr74f
9OpX6pNDedxMZKsKC9BoB0GB3FCjLiw/nz7W+jwF3yH0rhlf1ro+zXUj752+UVMd
X3ApgjTQvXA9uvJvYit3EP+jn8R0czmillUjPDl3EjMAX9hP4OJzK2sK3r/iU4hE
mVTI0JkDjnx4ilQh/YNmE18+dHGESvQ6/+alcRqMYmqRAuAlnz+9LFEMq7q7/CnQ
lcqVHuRVYsQ92VFtjH6/miWSY3URy7yUBtFvEW+Wtggx8L8izzxulc6xEbOughdN
XK751JXqhLprwB2iUiN5KGhc6hJKVPHgzsJ7sWyD7MpfKIqy9t1SwOAaP8ni3MEB
Pao9pkxB8OunSfJJwpwUkiNo2mT3exgZPmV5nPOPS/ian4LJ32vqHvOK+/Of0vqL
iztZ1q721ezxaRR3FlEwJTZB+WultNZZYXw4V9LK2pXnVLQFm52hkYHd7zJWW0wA
5buQCGSEZmVw+Yqld4f37HF1QWKlWKwYZVkiQ2R4Kqbsc2AXfnYXz0J5dSWXo+Ax
pZfcNj31Lhy7lUZIXZCmgrK4MOsHM1JUrUUrlibw4+OBd32vIOOPExwujHr3Gy3H
OnQhzY10QTWkUDOmbgrlKoW4d6ZpOddnJTFfNY/XMI5JaPcSQLfzOI0+sXBQ/vRH
0BPbfTwmTWpxFL88Vfqq+ic0ml3P9RggmxMY1MoKiRdwulGX7Cm7GOknuoe/LrlW
t4s6j89z208Y+XCDzVfR3aYjC1imLsEzLZgkl+NdTAuNfPa74HPRbZt9RvWELW3O
XXVmU07/i2p3L+M6shvmAEF4bxlesqSfb47ATzG2lRt2YZIyJ6DaYT3kEBYQbyoD
89Yp3bsT3dKSXFzUAWROUl+cg12jQUD4gNjzVhEiwngotyDEBphGS6rByeutmgQh
HKoeqUpOYc5YzLxRncztUIYcZltZXSbgOkDjDakrdieUjDyNYmSGi9BcZcuee6/W
AO4RuFczOVqsglA+P9T/RzMTDn5ITHCMrz1Lr39bu3G6SHCFnKPquMVrqk/sHGR2
MRV3ghFOHz5oHxFdBy6wx1rwEpXdBha744OonuvTFzT1K/J5jGDE8pDXzhecftGg
UekX+n7EEK4RMZV10d9GyHYwwRqhuBjejpq6BD4CqnHmj78V8sjaxGBAgfxVuE4x
GaauJtKYKYR6rajAC6g1Ne4mzLBvZy4IsD2j7L/0RkUJjfOsFJI3CZY5exH3b0lU
2fCPyXh3qigNujYzzVe9NU7TcYgsRsTnHh4MhPNt65lur6hT0F3gJsxSJKRLpsYn
DoueHqrGInQQVSPj95tKK4aZ3QyVERJAh82c3aeXn3j9Jk8JeJvugYOYgHZhMRXW
m2wz+wU50gJ1T9/p6s7CwgffPiAr+WIkKsERrvvOZsYSx6+d7OJGRdI63EcUWG6F
qETPyKjAYLe8u12c0nTf2PQEyU5KB3+VuWvgddit7Rpj8cjf0qphdMgwu/UIAXNb
gmEcIlAN3ApqjamRXv3g0uE9RmRMh0DPVi/PRQHGFngBUtnRUF9SNwOKMWBugRPL
Sfex7tY+XBQ64MS7sDUI4C2dduX3+9SkZ6+epWkhlw0r0ETN1rcnSrL3/vTIaHxz
0rXhnj+E3JxMyaERbFslokZ/PCg0ur3N3f0dbq+YZCGkPk8vfhvi7RBuyMKhxtJ8
LPbxUL/NaLvh02jMQh3EssuuMn1RH6omPQUsrnYt+KH9oCz3Y0hcj0/D3wG6unqU
RRHc560G19ZnlcW8Vr9Na/wiCP3y7Gg1j4HmiNbVhOQhrWeh8LrFk5ABBUmBLHjr
cpz1Os9ozWlOHhHYUrrOvjwNV/GKR0sypYk+lj0nPuiN5SWuXeGhbs9fUqCS5mcH
Hy9jI/06Msc+dXXPETTzJJn0+ER2JfO8T5ssf1vIW+ZKLkI4McEHdSCJv5U86XUo
4axLB8Wuuj5coMJ9S9oHofsmouN16RtZUwKR2XZF0oZrUP9XXsrQqmVNkGvL9Sbt
OIECrWLfMQK1pvIvQyrW2rlKm27fDMs3Q0VH7qntSObI29/o1DxvveqWydZd5H7J
iw3CtBCqjQqg9rrNdEBaFiLB5/loDfh/7JoaCqrQIF+QnBJVIKAINktxIw/AlKNK
HNZIUWnH1+JeJ/Z1Iuk8kouqsFp7z2S3HRahHSlunDYMYjI35YTepHJhX1B/xd5K
Hbd8mq5Vz0IyHzCeq8NC/MCZwElhdmivED8PZ5hcOt31kjD0xZiqeCRV2QSlvDwK
s+CH8LiqB/SKM1mKf5T33EYYfqMOfBRiCRx1idvhDDmZojiHwXwbMu7X2dDrUbqW
mAvcytRhmYpGfVF5XptmfjweC1DyeoplK4EFWubORe2uh6HchvUMueF/JGPP/ny+
KKPIVrx61vFq29yClioWoQBqDJpiTKp6dhmcL3zMGL1RfTL8FwntI3Dytn2K5bkI
lPIa+DLgKhaN0TwGM1ekDdZY809ADL5TI3NRZWdO+SJIjz1N+GbMgE80Y7QUUoEP
Zwu9mqOsQIObFXb8rTfRHY5w8IJxeyOHA4nqsADHe4YtrGNlSbISSPUHVflpTKKX
onlmYmZJZYSzq23BdHSmcV6gKGkBBf4IGnrAqyLMBfZ0WCESQU//dnILTpX6qAHS
E5eGWIhGkCfPANmfl3jwXUSQo3TUw7+eakMmD4akm92s0deT67ubRteoldgcdyBf
XPY0ZHQ59DJSVL5dYwRDfKH6WlB3upcn+pKkjpM5YOCu7TfwDKJl+Abz4Se2GQLK
aZpq7Eumi8zpKomZce5MxHAr/U+RjEIdI7jyXZvwaRfiSHKm7DDuTkG0nl8fstSt
xeZizCUg5ZQoVnLoatMC6JGArvOlGIK9TYphvMyQxHVF6fOX9rq/zsrs8RiJgKps
D9DhkV9d8PpDUAyWJSiPFUfRkMERXzsEiCXkcb9Uv6z6pjhywVzAa8UwdsaCy6mr
z9cNM44XnXEJklF0BUo7KsA92Qkiuyz08wPQSQIn0jlqGQA2uMEzs4mJn+rgOagq
fQ6fHQ+vr5a6eJGXb/dGSC7S6dCThFKrR7m6STKZPZ8s1QV+VYTwM95JreeA2S0C
GiDgvwRNDsf6erT9zDkhoD+4MX9LdVggQFYoN/KS9HsZ0pRq+mIjrUnZ3pXBiG0F
6WwCsTAQiDcpTetEcMZ9dtLg6dPAf0sxiBuhjOChCzfB7DOGTPlolib5xPfWfHar
OZ6gSLaSYre2yOhTQamwSIbsWXyt41UWLspYfCfdVLZTvyO+AcQ9cAoydNdMtznW
ST88C4oinqB6ngteB3oLbY/bS54M9bDrurqDD8FO6XMs8u/JA8PcYgHYGK78Mueu
fla1dZE9QpGNZqexmwihjsPWy1kkAcX2ul+rbwdmuz69jgYC/qCf/ortahxxrR49
l6pojc2jotS1LV0vDR5DwpVecGJAr307qqjRrdt61b9XBWD6TIHoSJMiuQLwDrJ0
cc1hDJffB1qIwEI3ybUmX88utZW4ryjf3u0yuvfR1TjmP649cHVejXPC8bYgQPoe
8EwOYph18nmUNZegy+IAec1+qI1JGkDyw/Ry/uZHfpQ45VR+6qkasnlO1K8aU/6P
wkmcqQJE7zzb44fqzMoWybdq8C6UJKd6Ud9Sjoy5Wo/lrJjXdVWj/IX89quOFoAh
nKi1yZhvDOyEW7GfVQ5iwg0Rn1hx/rk+BHE+n+zLPpqVfp+ptr6W/20AtzhaQ9wB
BUNIDI8WUuCHVjrawqryt1epZEl43du9QPQealTUDHAzwRyNsUuNBUKMSvPByOWK
bDENxjyUM45T/Op1zQX20l517kbXFVIBZmAnRhF8el46QkRe5fPk0MjYBR2Kogxb
UZCokEIWV7gQgu6/CgpP/ngev5vMwDTHYSvsW0P2XMl//PQtGcDo5tM41DvvAnfN
xFwOcXcJpJc7bTo9pInVoOaQdo42bXWcPvrjD9d0Rw1v9JtHbRWSDfxa7RjCduwS
d/vYFAa6iGRqFIA3hGMwBNoLDbf9hkkEESnfGoZ4wFh4USsqiVmCVX7Phkujl9jU
GK1UZDyYXj8ifNiywskIp4CXh/I5ZdulI6fofAbeJdvopP9iqYTA2Db9NOkcCBMt
f/m0T3TrNnkPiqRvLWmJ5lc7DeopPfJXtF43VwzTo+sFinZXw22/KdXPM7jNIQLW
L9lTp775Jk+e66d645tmOJPcsFU+cccyYlZWG9N0udvKS/nC+M0yh6n/2rAo+rcV
azCdKzwq8qVAYgVjrg9GLw9geIBInEPDFEVuh3T16yDLaChyVnGzg3BPWktlo1Ga
WOL3S3g5a6Xw/Wwek8UhAiAhAiT+JT58Zyp3y0K2yaRfzUtox2B65pnMXlkbQiRH
yeAXsYRZnHxF3fPeY47SSjSetLkR0HLt9p/YsgRgwrLXtT52jzahDf0b13tEiP/Z
WOE9sh7ZVctLFXJEH7VOq9MSYwUyGzKcdVo41JF4tCkqFcLpos404fpN/9q6aguZ
d49lxQXkO0mbGJLlQONiWwba9bbsjDjpZzzhnLgkh0B0gCK2HHpx+0ydJIH/q6lb
FBMuHY7TqTU7o3DsR5sleCe7i1pSHGVfSAd1Ff5zxZAtzR4MQFhCbVNGbeZhwPUi
wLjDTxqatQ0y3CcHIIguM4ZrXgqk2tTad5vgVn6YUi2Z7660pIUP6Kn0daD4+T6x
BxaDRn0ivMalvZ1BInjRJpxtMCYW9Je09eBML+nGBgGGHdQomEGRMI0eph42Rx6s
KYHXY3D7WYqyWP5z1N+dQkc9k5o6Mhn7CGiNYdV5kovYfOzB5FcvOYPTiwMDeE6m
K3M+er2u8LF4wzQlWuoGWODnGM/k5GXc5pjW6I6LArT3mYJEUz/W0yBOl3joZKAH
VO4oF1lg/azlp/82zq0GXYKUdec9bHg2y+xBrk2qLNbpz7vYm+bUVkKwzArqu5EC
lx7gp5FrRqFBsZcmV8MvYcKzONS8ZfXm/hYrElw9R3GRHhdqXqF3r5D6v9m6+LY2
vVaBOiwAlinEaLzgpeecpqlZN/xPxxmlHsWyrGhHDoIt6YJsxEYoG5g2lK3QESg4
5vp02OOwEm+1fxII1jRbskSsder7RPUD01fFBEl8R7T5l3TrF+gN9vm0ZmvyyaPX
xVpaCMY2NUyW0jtXHbx7qgG0bAcafUsMdZ/JOhVvn8tnAOqgXKLgA8eV+MxQVrf3
1Kzzx0kLcFI6YKUmybYafadi9vZhfYVdOea6r4q0e4m0uN++u+yWYAThMaEj1mcv
7Zfd8bo+8UYmiR9qSSoUXcR1OKagxSH9g/hZ5XiP26zuwWLHE5wGaVweb2T4Cs1K
R1+APsM6wo/vF36T1ZUfovXTWvMt6b05SXvXBxJNthvXaGQHNvi+5L7XR+4E+VwR
e2McyMwxZB/h5eTK79SgXTg6H/s5KVUzGayQX1If8NvpL7dt3phfYGiPUYrIbXmn
MXBHxmVrDpwe2vCbGZU6h3q4+nbQXqOD6UeoE/0kyFS04LfwOcocz71z/tWb9j/U
c22f/h+f74gau4gTBMAIqerAzC+IzK1kdzZp4amVLG75wlhp0wZaGZJx4tHepCZI
FLGwD5HN+iQMkKTNQYNOXabYRDmNVfAgTb3p7lVi2Ht7vNW7WCh95sKS8H2jH3wO
LR54fk3OhDfS9rxZfSois4zmj1nttfBE2/4jQQKT4KEXGkAzEHuaEr/RcuWaxODl
qf4vuDpQO6RITBhK9pv0omeVufXU33dvWR6pKSHtWQRCD+BQsrPNj0NC6jZ0PzVE
uP7R8l4iKNRAAJazjPD3qnTrV9MNnS5vI15HDmF+FJXsQ1mD6PIsKgLNIzG1+joc
vTIRAJMPuHPNMiR13AOJQHhhALlHbl8XilZ5tmlBzDtQAajRsKxpks9j3ZeGAq7k
SF10zIruUfMAD8jSJ6fC+FglOnDB5TUibQOxIk2QIlLpOM3XOk6ieJxlIOFUYMZJ
cr3m1gI895hJiqbIA2KkEoTKKRNiqf+wZ1XzhroyGuLZhYPy+RS78q8KoJcIKBRw
Z5xO2WA1gkAem40UpLbEM96jF+9hgFC6qFPeFU9JJkpDUKF38LLaliOZNMJJ/K7t
oMj6RlgAjBt/CLvwAM1ad1xhmXdI4Jhfhu3kkAxkLWtt4VzK5wXFc+Zzw4nW7fHF
mpKXNIKq/wJy/qBftX6nGjV+N9vaVqyQWEX1OiU18TDmTxk8hKGmoT+/JaApClR3
s83THF2IjGEtqdASvB0V1EVnr//DTgLJHpkP0suQlZkvO8xFIPbDaft9Vc+XhA/w
hBlEiU0xOAfiU+4v/D1tXGgP6s22cOqW4wikm20grytB6wx1yLwfS5hc/PZJfp0k
9jqcUKy1SlnuV+iYQiOCvUDWVw4seLwDDWput28iI3gJtJJiW9sG+p/jtGMVphAQ
rIMdPAGk4hP7OrcRft6ADo04DJCKKhsbHn/mpPZlEoG0ttkvcgRyDKgpOaPD7t3R
2+YQgvffWqLRp220QItAxTfoOGkVhPGassijICkA02Cy5WT5+7+BVHD5XrVsL3zD
OErJh1oN3fPMVAZfJsNZblL8ur6lc3WH3VNOC2LT0F6BGhVEW+97sO4nF7Y9gNjo
DWoHGF+CHswtORsQ+16zsyPV8+B3rDIO/SXvzIy7THPWsR4sgO9dUQ203hvK5Nxh
5uim/fC3elv7ik1zPXaZIyBItv/pGFJTEzE6LRedxl2BkOevFOg0nBxJ5RqNpBNX
YEghxSnylG2klJm2HZcZaQLnl01JYMW66ijuViyNCKo5l6GvTyw8pfiCjQS4oocd
kNLJbORuiqvmVzf16plQ3qw5Y/0T6+64jWjkcn0OSYgAb9PSAvi0BdbMvBQYsUOR
L/WR5eUic0aR85jd7AVm2/sASKEyGKnlsFT0TP/ODNyo2NqOIa6usGFYgDcMYk0s
7S6/NpKfBrbjlBgtKjyEldXgJf3MEKbLrlYDEkspGrZPAu1IKE26VRJ8EWFja/Og
PeHCI9o3jtJevq0cs/6qC0SkwDmdoL7wMbYvue9heN+KlKlBdErnU66n0gBXle5l
iZGMXYEPljXteGQAsaPIDsaRDfWp/JU+H8AXqGTv1fkJ5LTea8koP9DO4srDJX7v
svuFE1rImnZiTYiFmbmotPM/2eQCMRKeMXbNiEg7FS0/QteImtWK5Oa+RHMXOACW
gI87gtTKKyzpLCuJtObUNdLThZ5izcFu7FWXq79SD0QhWghLcSND0z/fi86zK9TO
4ftM/pMLleYPLhNYhknQ3kPugOoaUAajsAp+UTmygceDWZtJeWyGDdZ8w2e04MpN
EmmjKX8ir2pPomYCvvMqS+aqdIgG6PKcYj7m1v+qk4bNU910IXmggEVUXRpU7Wy8
7GkyBuWA7Sa4KLgdpfv2C5zBHClx2JkO5TPpMPu98WdmYUD/a/1jk1guaoFv2W7b
RawYc/3OXn9KLkPyTjv8uj38sEOcr71HeM/5NXtMLstj8KrMlnw9RUW+ZczrnQrQ
t9uOZZBerzonMbzhWf1y+M1gQRiC/94Xt+Cebp+81ZVa9ODv3JzhjQGe0OPrSM/a
dZ8dMCkC/Nysm12cc8MuvXaX/nFgJFFC55F0/y5TsTIB7ni0etJxxbfDycilG8ih
wmPAqTWbSSzjyxIHgdgYecqjZ45vc1tuBCM5j8VlOfgDbD45g5f2sr0ABLYd3jMN
phGPAVGKqafACYzshG+mcs53Yxwf78IH5U6Xmp4yKrMs5OGEpW89LrtFE2JFRLOX
HZMeVH26uvmvxxlQHRrOvyegsJhE5XwuAnu58oYU9T5UJ10nHamIyIRYwETMpWi/
NvbW/9UaTfZgLXp80bkzTJDUOQxu3WlnOm9BaqpyTbOc1je5t36CJK6+CtXJ5GYE
IUrHTl5OMN6gdKWm7GdSFbJz/M3dziForuuNcO29sG5y1LHyScLLqOY8aPxl4inp
TSwEZ0bZHGLS0se3ckfXbTUiny6vvb4WHJJYSbEqzsLceDB9UsCYUISNNSjbaQvn
R79XONpyJQ7WMEIThH2pWHLhejouIWsAcmuV+GmSte1Qo9zkE9+WrLZty6SnA5Yl
oQwOb6Yk6GaiMlJQPWWaPKKiLwl3UoHP0Sbxa3Vo9jJjsZQRj7EXS57DQ7Dg1S2l
y4gkpm8/1/a6YQjDXZjANtOqEPjg/XgDYChxe0YovUzwoFs4f6dh6GnxdzbzM9bx
gmvIJp0CvWBb1ZEOzqLfBoK9gbd42w5t2nCkTv51u1qetNXqoctnSy6ykhYg0gSk
fS1nSEFkw9KuZvTljiq3IgOWbrwLYa+eRFo8Aw8jgi4/kgCOSNYtVS+HQn5aboNV
CJfaJM/MBZoxCaifM9b/46IufAAFP2x8Ov6hWIOZSzZLVTmtSMuN3s6S6oYHC8Hx
15d30sV4tfzPJOX1o04AeNZ8nB+nW8ZG4dIUwdASbvJQBvYNB7Z3aiT4vytClyf2
nGI2pEA084bHKrpS5Sw+FoywYB8n2elFB0HEgEZ4uI8mLG4J+bs3X4Ef0ONSaClE
FFZXQuwjQi3l+cP8IytWmseFhceh8zE7/P+txuZSLRmlUkb+wiEySGh9HtLL2Qoq
/sCExp9MAG/uvIbD9TWwYHGf6WIeTLM1FnFh49XDU+Cf7o4gAn4zGbwbz76FWYVk
ujsMGfJH1lqnyISTKEAnq5ObMLrJYteaWV9Lv44kfK+BJtdTk3NoMBBZWqKwjmpb
JG0LQcbjYLMzWLhsYLlPWgmJIr/fPkYvcw74vvz+lQkQwNFFKWtFB5k3ySjZNCtz
/+fOKeKmYLf9Khbc/AEDfpOBXKig7A6WgXHne5VgJw0dz2h3sjTh1DR+Kxi451YU
NSuQ+NftYKJ1y4kIKATXkk66LZCiDnAfQYzelKzsF9wyaN5/yPJzslqGUPsM3dAk
bAbJl5zQaonzUAGguFKSY/dfknMYf37qu1go24eOr8uDgrLfVRh8Dy3PFllB509N
Dz9SKpoV6aKMjGqNY6j1DqGeFLkZ39Tf4HayUC1k4XSm4jEK7v0CX7h3r4e3tH39
2RA2BwDSSXmEodlYKbIZ1G5XJ7buoD+qZ1dx48ews0IWtqHe/P9sc9UuWv7n4QxM
OBp7o3685G76sioPuYMAwKw82TB9Tk5bMg0wQdReEboyIZjUTqE1XY3StjPwHN+1
sBgVX39mg4nWlw5MKd0smYjTfiMGH700S/blPMiPRgVoURtX1Mrnn5rqpSqHw/0s
yHw/38o4MuOp+YSA5XOCEmSmzTltVYPKMW4kEfL1cO8IVtN+9Ml00abnmmrskXds
MMMrgBJs3oCpmDniUWvMnBXBFCW8kPTOlPSdCZNav0Kp1XcSOtala0D032VSF2wV
wjkVDmX0opJLir/+wbMI8cdX2Zw3XJI0iBMQoJcPymEJ9Yh8M4IV8GhPpWjgjV4M
MufPa5zHiF23N0QoIlO7PdIvZWgkInnUSHdE1u0iFLUYVQsM9IMfPYRdXI9ltaT7
RbFtiPXoExhMUpVZnYA5q2DV7KjnWAGz8yQU1AFyXFsXz0uTvlDPJvN10VM088mh
h368EtAPLC1F8zPOzZPZosqMIBl3H+9xG2R07ogdDVicVrZFXhndg/sc4PNreZKq
/DKm83kU6T6VvZ7obyFnAHE8n3s6JPFgqejYQ7mrIj0N29VnDuIDpnEhQPIEt0ls
ztsq/+qYI5bh8gw+fa6J9aNewESL7qUcPH2VZ7hmGo4rrQkPSwwITygjrDp3fid/
rOGE49gXwNc+Iqg/AKnVPLY5TMdBzwtl78jZedy8AfnCGAxl8UZxr5iMyKGCyPzw
ZYB9tNy1r8ER4yj8rrB24JBd+amXKt1mvOaxrBo7AYc0OCw1g6D8Uw3MiihEcmhu
uvPZPFt+j7iKahgsXVEjhptokKF4Azu92yr7RBV5b9VwqjhXR4Xwlja1nVYBXxqz
Xfk2M0gO+hVgKLksM0YiORIH32bxjWZkameyQHuJR2GDp6lMNBNd8sq0tN3sw9vX
nUiTlaIeiSZpC1XNIM/RMF7mcqgy7DeBUeDLSTtePDEYVToCpxP7AaiL+dk+CWjM
lCo6Ell43fNDSrchdmxbuiqiUQTY3xORh4TbcFv9hnrE8pA8ADXB+e4liBIfS1Rn
vr/8RbEV6l5o8w8r7KVxBX4+PV4/2cd9cJWMIcG4wCCvB1d5kQR8dA8y4I+fLnjX
LpPf8gvwZrUx9IIIbvIDuEMoEoWIh0tlC9Xc5mYapN0/2wrX5Ed5k3X6+a1M5AvI
dOo+50wdG+pDMIBeDY1AhBdNPmjqUGFqC2IMtvEvqWtHff9uhD12P8yBs4/sNhzq
Dg6tlyRXmLy7R/l66RA6kFqLpwG24JUoeAm4oKpQag4Gchkr1ftpNv3wR82wbb3O
42KYpFEcnpUPjIiWglClQjkqK2s84Ey26d5LtWmlpgL1GUWFFqz4eiOcGSb8sF2y
rvfSip5uww/W/1JX/pD/n6pRJUTF0/doMVPui3XEG8xEqAsW3CE38mUIQBoB3TRz
bY3osF0pOoTx1LQy08CVMVB9KgksVvYv4J9e/pEZVa6Ilve3gLorQqIgPrzLRd8i
kguynwvv6Iw/ezWCLE0fdfaB567KmfYH9qz22XPKkO1ylG5RPezj/eXkm6qlg+0o
7LwGmZ27McDyexvyxUoN91riwKWJCCVOZ5Ini2bmDWUiB1owKaEKgblQCwBjYSnT
ouEoFBQ3mNsSETys6ovL4l7rvmk3D+fcywGLFpQ6wXQo/QnjuWY6fEp/zX9/KohJ
vxRcvK7tOq0y/k5KCnBB4tB6qW7oHsOvVLHJ2e5vAB09PR6cfhPEb7+w8TtMoph5
IrJzI5FEAt/8/8GVuuERLKdXqbGl30Km3BHrkmoeU+p3tNA/x3UcFIkYr8Yk/pT/
OxUecU1/qx4QpuKlclhVMMpvy4Abb+sJVBOo9PTkBqXb2MSs71EYJAOUqmKU45ul
hjYwfmI6yEHjINDE19egLoXSVfNzZPR21WqFbewx362OjPovCGG8xG6pYDD3Til9
bZ1R3JPYgOVR9ss/dnp1keEv+GYAG4rXgDBZvClcZ7hJJTtPyEtfM+gc0Xvw8CR9
X3x8uBlcI62amA5vXEBhZGGIBY6hQPDzJku9Lw/VY0JO7m6Qa6r+iHVyP2R20msx
8z2zsTa98CTdSlIDTn8uE7+An5IUyVRy6fOHbRXOrabWCa1QQ4az1mZAEMZMfH+R
YiT37nLSfzeKiyxxdLVGYBwb7n4nnkyDHoiQdTx9/qbtadkTu5cJUwV9DyFShHJX
pXViHGbQpacN2l4J2j7KVM5O2rPt7+4PiWxMtOW1525oXcjQlLhDRsLhytkw3HD6
SEh+pBeU1c8m44iituhBsjlG7noDUX9XM2CLwy9aizHA6dclnLp1l1UIYHtH575g
HGy9PFwRXPfEeTLfBFJCvIbGneDDgK8BlcCaNvo9fwlBI6GXrznJ8b8p0HPcUHFq
C2wMzQ1/T+MDEM2HyHhLncuewD0+qfDOt3SE0uHjoUhE9iI0fDjZIbzuwiH8ZAMr
FATBv8kh/xlXEu2yaU6BQDF0b8GyZkoYP8v0Xzu5DGfxmhQ1lpTmW7h44S73/KAc
SA2fM+gi4iye1S7Nze4JI1i964Aq0SlU4Ga56cHAQXN+C4vMopB4EBUi2GTTM3HG
MQV7bF+spNH+qMcb33PIt3EY2zgR8vuadYZSPRTwYSrU1bT2LpOJwa4A7GeBoJBB
lx5T2OVKSy4aq2oQqEBQq5cS+l1Mz/iI+U/gggYQdIF50r4crn1zYZ6Bnrb9znlo
CTZpQ3nhjgWGW8KvBrwP8jSs9Rfe/TbnIDyj+txcg/tcHdlK2sJyjPU30MCR4xI2
HipSeqOmXsutAaj4G7vPTJTy+Pldp7DJnO8sBhD5v2/9ENy9qeXcCHSFLulzh0L5
IYisuGRJa9otJMJwre99lDNB+SO3rw76iu5reUOMvitIrOhW2p+IYTbzNdZ8Q3yH
s9aXAiZr4ZyO047E+M7rOvxyeVwVeZMk7byHW+M+V6xz4Z3Y29xx/kWl0UPH7ldO
69LsEywZrepJloE+z89RnqWDmWU3S04gkWB1pWxHchm87EFiU2BwZtawtO3WX+s/
GKWTgJtwYWjoeMJB32RK+P88Bd3k6LD2s/1s/ZE2ihyEW3gisu3vB7VX5XrTNiQa
cYBYmrDnrO1kXXd8Os+rPP5nFxPEmcJ7934+L4IS8ZbOu8ssFSuXo7KRoslUENEO
B5+JwOdxAp+4TOXwv5bsVYZLitYIkScCQEeCl3xnyXoIL6RVXx+iig6BzfOp6RGG
7qelnmUpVxLXvRVMQkVpchywCbmqHJgQXyiM+AZnS1eOMOsNcRfkdBI1yMlR+6UT
vS3LY+LGzJLXiuBfGJARhal6u2emCigp/RFCzHr2c32Z7/w8He8TIhm91D2CGRfi
mLhS88+CkssBnhLRWDbYQJNoxs8GBKb5sDpk5mTQF5K3+roHI6TRq5Z/RJzPGF+x
8YKMngd+JzUmgKd0hnotj3SmV5eVu5BBadRf82F/f+Nl0G0ZNC/sdz3DbKpUCru/
E/bBxtZQw76dmhcA5nwqNhQx1iB48Ao775sXlJrGFF9WB0qi+ekY9PXqHLc0VcRq
rfWbxmn8X505rDkCr7ezmkCxbvklySL9hHi/kYde7pThyX2ZUo7qr6qqDt7obgY7
4s8AMGjCaEZZt/qBeUNRqSw4gJxmUdepdSo0FEtmTcSkVM+ct8YAdjkCBcwiMy5d
j9aTPd9Ic94pE+E3S9igPZh924JhnZqJozz+GS2DkjTh1zh/1ibj0b3/TafxGfql
hIWapkg6n+c7s0Kgm8lve4FsoQStlTX2ZiZlJGAlbVwUyGX5j71qSdpoqaGMgZF5
y/gkQFPM7m4iIKo6BXiSsCFXVz/4WnXBwOQlugLzsUXO5pQpGq718vyYBskX3gL/
HF3wByv8/v7hL/dewG+H5Ac3M1zDBv0hhgtk1Zk2L42x7tg/PtiU2eNOvL2CySJu
o5WxR6CtukDPjo2iDXVqsOO50eOsgrBh71k016P6GbpLktDJpNO8GYahhiqsq766
+BC7AtgOaewBRdYLD8Hp42eBSS3zFRRjlntXyLOstCsjAgXn0oFYeBySDmR7b+8q
zH0f9jqUduJVNsgZQ4HEbMqiM1ixAek8ti8TQLnjtiJN39HIavBszMrp68msmE9G
siiY2BVh3NGplbxV74Lt98K1HhYFIwZGen0xYAiQqbcr48d958rlF8u940a/fBuY
oaJidSsbpYPIIG33/6Hxd7e+MubO3TVhJ9ug2n5tyQX45fD/YTRbKOviW3kYMbEO
mN9EkN9CvZHS4e7g2F681ZP0G/7TYVR6Q50nPhX3MdULMl1LYAz67wmprbtjsREF
SS2FoUHkhVs9cRdVFc5Ys863psR5V8h1xuYjMY2mLk5Z4Tk5oAx4jITGaPZhAOoG
KvmhCrJFuxwlUeymiE1ugvUiTan4FG9UkekDGtzlE3myYjBEfnXNrzeJ+yl8byLO
WyAlWjiTWkC7+sGymsMfgoS+ZaFKm4C4dWRRgkfMZGnwwdUW2X8TAJsQpNrKid3T
l4LDtle+TPUrXzJ5eu95Ak1JpuwLfjdDbeBdlZzNwUICP03R47VCzZXW0rOWPkJv
juHjma3nYH3fw/PHSZhSCuvRKQyka4eVCkVpJ60NGcOhry1unOtOgFbGVzNjl+2D
Z7o5dipfUpngOeYdklsZzrEFwPJ3ZzUG3q+VoR6AzkvAhU6qapMLMNrvcTaMXKFl
W/7i1FdFbQ38q3PXyruZDrQOZMOAjPBIitqU9Q8jJ4LMVmhCdwA2BCRAKTf4moZl
1FpgZZ30ErQxJ6vqhhkxPXCKWNSjC/wMOJCxoj7KnwGPQhLrIPXsmDi8gf69OXKP
65/Sg908dbLgkbdcDhJUpPBzLwWWT0LhKF/6i7bo+N2TDq5RLXiRcn+X6Zy1UXEn
RTjHv7fsVbhw19F5AJ5K4+va6WCM8DHgh5jwyp4zrOO+iisXieqSdN2TAsn52fAt
ybJhqFNVFyVwfHdJM9IRr498v46ga/gyT6fiMMK+zfVJdBQLUFK4Al9hF5P6/0OX
sPuLqbOoHT/zZLJj0Sfy0AIluxHKWJb+kRS00JPVH/O/+iXNVWic83V/V8akOTwo
acrxQvqZXwtA8QgXH8pN1R6JrL/iZ/ojlipTM+1jXieScCiIeLGojjLliZLNZcJr
T1jZKqijsL+DEOCTNYD+oDGcpShYNdEvaSCYBhp3EUNGceZauSu3Vn7HB++c5YtN
8ctr1UKy/GE+AQcZUrpt79fApz3GlpfQdHsnCxTqKLRu8gwT6cqF42qvNoiGHbj7
ADmAiVhb8ceX7qi7JdDO7U0QJ6opV0Ssr2L5bW86lQIXyDKJnhMQD8A1FEABNn94
Cb/WB5kEkHblI6WEQCsnRHvnvMho6IoBKKk/zjxRK0fRlD+gVr80wZtVHDEw/JXd
NBZORWGtNB1TCuodv55Q+7P1a1JoXHmfqoEBDrF4xVMI8BVFV/9ID3qbeFLpGIN5
Y6KqgPghVoEFtudEq/ino+NpEwZYDZJPlsOrSZ8ID1iNzWlhK2vUDuge7Or6D9xR
xWwGOyfnBeQLLviFuMzrdERmyS91uvnKH5xFVmuTd24IB9bBP7MtSddOXHvVagVO
QUQg6J4opS1TCoxEsbQy7wvgO4oMHSCdejgM6H5qNnbKizyEdNBYFUJjHvCbO02e
C7tuRXb8vymPq2l3aIoIzV+vqC9XrsUD4v+cx0CKr8GdofyLQMmTHke78Wa556/X
cIvKEyFOXGRYHI8ZOh45nSvL7Yd+xl/BKR4D/QtwnJdxK3iTJrYVd+vp6w9gkhAb
pi+ze3FsgqwlqC7IPCsRtEJ6Pb3LIZZezXqVukpfdwwit4XQBvJWM2AKO7Kcs9t8
upKoS9HuH5QvxbkIKvwqh2sJYYEycxgPc/X5dfGRJLK5Q849XdCugwoBl+3mjBdn
5cmgpP3iPPX5WquoCdyWSajoPZQTnbVqq76CJJFX/6Z0hZqZE1N6SX013IdmJA75
/VsRS6UBvVeICMI/18xlKMHAAfpYB63GSjOU32pxFlmiiMce82Uqcq/cTcRNEtUr
Z6xcmMEIbiLw1MlzHzf7qnw+U7izn238SyQbdCtJh2i2Cvd9tZuBTMKaGzDKBsEh
gQiT52bAc6XQZqkVxbql+3HWEpbq/RBhoE+xJunh0Xi/TqB5Mgiu6oEbbI7Y/BvB
zzS9IJbS1zpVHNrBAKnTA+KjPybwqDy45VZXipAI1+2C4Qm5NPKOp0ZIJpIh8/A+
N3mLLr8RRna6eXmbv3ZDAW1JYiT1A/zA6Ww8DDsL4ctWeM7FMwnvRLd4PtkxEP64
pvNSlpwZpTyKxoCZx1WNQRc3MzfgzdMuzIwBxLmow1sFyw+T8xEvZpDAnJTHnME9
Rfi/iX+AXC4KzYfVXkwp7uL+99cc86gl0lSZ+wXQ8kvgzNeIIxdfF87W1o9QUpT9
KgzwSl6SEwSuEsgTYnvY7VZZh7VldbEmRx0NbltXeuo5gOehsM7N+t83031a5y4/
V697bNzi0JjGHDzULCP/T71zSCIOLbO3BGWC3MqFeRcL6dBH+qymP9dsr6TemQtV
TQ7Ylcoc9t/Dim4sUq9CyMNj7gobFDGbZ/9K0Jh2U66vOoYDGl1ZB3bjKTBIB1e9
/4W+Lmld0z7a3mR1DnhkEhULR7bDFY7E6Sg9TalEXAOtzY6a+xE4iKTITyXz6K3T
a6KOG+kABiT2LYk6CuWS2UScw8eOnqiZVH+7vxaEe07PdYt2oo739IVUhnWyxcR+
nfeRNkoYogFpeng5b+M7sYaqueRfLnt1dZg6TaTx5cVSO/57z7X97SbWFOcIhOUZ
ZJdCFTHxy0jxDgbNrD26w6ki2HAOQOLop2Pogm84faHaL+gMGOb1LfibRIVRmXqF
xn/qJmhmbjLHCkAhqUwhos8nh9pr4Yf82MD3NBGuayvT6hgoro7NZjyDUMF/97XN
hO0xv39Dz+iIBcUFT5akqG37CSNTAmqSzW0YJ8l49P3TL6ZkiSqeslSJ92Cmn+OI
TbovVONSi6gHDMwcjKD9vtme31NwHX2hIpyLZCETUl31ftIrFy4O2hSh7X0UG86V
ifaY/fD2cUTptYWNdJVT8ccAA6k1UK2z7ykdaLvv7V5psRNelFps5wbCxD4AGjSi
Rb1fthiOkvXT6uQzYzSGjVW4n3D4Meo+lVpbc3JlWG7/PV4JW+b0JjsDbz/z6dSv
lvDsNrqZqLUl+u4qAh6IhbXLkhCV0Vf2Txe2hxqUGbRbYQNdsJ5/uz93ZKxwhF0T
QUtthNcjktytkdYZIuojcww/lG74AFvk7F/DTml4wASmIeWorLwyzS/IyECKCjeF
CiKna5MGrzFCb3eeh6k2vjSmnH40abi3svMdObiimTmkurK4A9TaZsfDBNHR3LVu
6Sknro18AozPlPYHIqAqRCFb0m8Dz06ILchAA4ZuLhNAhA9v5eyC3d6tX7u2nVDE
wHJnt12CchqjgPLCJDsGw7fnkNbkTTMYfDcLJMErCAzfhPO7q7JV7RsOKcM9WJ67
B9qICbXhN1DhJ6+QV8enX3/0I4/DlnEA0bQ5J0O+rCPKsClrkQKYa2ut15Di3aD6
j3nDQu0Z2Y1df5Mz9uKfROXX3N7tu4hxU/PUQtaELujRbfj+o+hq4cgJlxwXsKXp
hSLOf89H0a7nOwazyWqlaQg6grNVz2Wup4zs4JHIFeoZbl6mZZPXLPwePeOYJtGv
5YZM5+TIWgzV18+xcPd4o294PpVO2Rk4oH3X7KM6DzktCMU9RpCdotlnO7Hez0Pr
H99laSDetDkElphfLzV+6NReNutRp5KezfTYhhkrrgspCpSrI+xgLoGc1cUhHSPe
YNu5hal6EfWuz/GIop03Zhh+sWlaAMhcv6pL5UvYXd+JTRVUT2Co/peHNh/LueaD
y9Q9fcMO5LLBOAzNw8rtc/0aiq7R8PZjHQCA/JgVcXcedf6ZUMyLKs7XVsIPGz4o
rnujJlhcZZtpWt1KiOWRYNlC/QEvXK75vamjm0KvBW5oLy/aijEt5zaszfBV7z0P
o0J0UVgR5/AbDcKzAZ67XVhP/lUzIhjyNBPdZaBrwaAXwE/Yk0S/FUWCeelSZkEC
gVck+YSA/0lZQUGHQqMgz1FT71Um+rRyYUeuqP2jMJrWHEqlmBp39apoigiwcQOr
LxbuXxY0gmJEqpG6L7Cq6ZfRDLwqMExKiYYuFlMgvnQlNhIo3GstfZW6nLtGQzAD
iFgVPmIFUhbEHjO2tNjXrYDdQXaW9rWIHJQVFwqpWPmTMWdZzFL+r94d52uLsOAK
MGj3kjhXfekSHz5FGTSh2ohsmi9H9YiW7osh8RM35+89EwNN02RDNmMTgvpk3D7i
/LN0/0YWhkJ268zQUSe4Ndxd/tkWDidr2o8N7+UAvfsixAWSTM9HwoojSOyik2jS
dx6yCizgtPwt//PlbmhZf/DPnLkQowUfLSNK4LPpH64IcDH6Ycg91M5DvL96VBFI
KmRBDhGWtIPJtA88irBgYlbUWhYhPv+AlLfqRTQhf9NKm2uhok5G5OKNIyoVlyQW
bVIpDPw4+qJuda6TG9S0XKkh/XPEcz5/D5oSoXO7f5ngdeQy9U7OLjAlzBZRlBGM
jO1M3yOZ9T0E8p3apzwFlgvE1N7NQOMqFRvEGiAJ9rClCtwlLwLTMjheeSNCjaRm
Yg6UpXSUzwOEzhEpX9x5LrIZty41OTrPzjwKCPM5UuiFexNV6kcCCl85MOAARKLD
7Gr50S6WPpdAei9Aj0sUvTxrbKDLqf62KVPBxSIWPu3PIFBHNoUdEtUwXXxg732o
WSVEE/HnFF768whe60vxEQaeyZ0UjAcd8T3zVooYmJM84DbnQgP1breV6nYrR7mj
1BfUvz5bVxSfblIPl9FHVecr7oensf2V6i6a4a0A/Kc1NaBIkG/2BaVC4j4lnIc7
ifmACzLQwIR9o/W8VGp0khQuuztjR8diaosJsUQKvnhy5wjx3Sp4xENXzaH0xI+9
e8hwqqS9rcVbQMQn9XhAC4uPT0tzkFVQ96X3JKgJJnG6WHGul9oOAWhQH9IoKXOA
2d72LxEZ0iqq+hmKtFnqJk6BbFA3CEOFfAKOHaCwqhDrJYsHWl0qAjiA+mQ7ue57
2uFNtQOnub2xrt8iyVcvTabwlBiUU7xwXVYV22oEsOR7DVJTN37sUpbaodWfEuQj
Qp2F0juYMJ/x1cHfkKkFFrEqr41Vpgvif+/brUHrCUMLXArowis7xDJvP1uENm31
IDWrVW9MOh9zEdF0oJKLlLKEUqIEGqBpSbQ6nm/a5zOHWCu/7kfc39LXGsERJPep
Y2fd+SuOLFDg0nLiqmzr73ignPPjSmvadUKs4KZmhpgamBBK2Sphtlj1iS2wfst2
z3JykEfHGJ4HEikJMXk9nj7sMJa9xUmGeJD6LlGw6kOoLx2PySnuAA0Rfaec4aNk
t404PFulsHnuEa8kKPvGRtqVUPEDUx5/ctM8cVXTEgmbe61ickwFFm0KOryfC53D
BH9K0gfW3uxZL1Wm0gM/5KCqHOG9aC8mKaJhEwvMWiY2mmlB2vRL4FANbZ0m459o
v/1CTHqFjfy1rFFofN66JiGiDgmCGmi2AmdLDgdfRYXba9EQmPbSiqOxIju2akfh
O3MxVOTprjF2Nu333qBxLwRwzr30d2m719nH/ni9RMm326DrNoBGEw/v9qFAjOYf
VDJ9BhR5z7VFgrBQRClOKjYycYWhYDY/biurZTGKitYvzBN7/MFIn6eMoU/w+2Tq
JOS/Yq/fP1YpWCvccyAyG5gtmWO71td0OfZJWHyuB9fCz7yqLJUQ27i9H13omFEs
UWpU2peh6SgDj2RceW3qNfsTuYz8Za0d/orgK+0MBhhsh2nGmz9cMeur14Ky5IVd
SmzbvFnKVeemN/ACuv2K4zpHZ52W6pim/Io94/qE/gZCtdW190mShXCb5Xeuogsn
IRarE1fhqc7+xWJRDLiXIX5fpl9Y0dW249/PKxaXI9R3Fz+MFTSf5AfFHPgA9+IB
f+drDLuOGVbHgTPMhoRQ2w6p9ihJgATIgU/EgWIy3yJtKaVA1DKnsvgJLuFfWIdm
sxAA9rBvi3xLww7IrbWXfsuN41e+5b7vvLI4CfAhPTcBTrvJXQxGyrbvdWmzvLoC
aSLdy7LfSqPKkEtRIZU0MAFppm/tUKCrKhUloxqSc5nLafWWbvm9k9LOjE1J5HWF
N2nlU9wGjnWj/aHBtaYFzvnu+mnUsV4QQ1pepjIUb7sKqLoZm5ZZrDPS4pn7dgjM
5iB5/95ocCMHE6pJ3LOVmdunjZ183LAORIZMCiU05B2UAJNGmHhxFmu2CogFw0nH
fPkAqMcX+WaQbNwld6HmAfocLFo2j33T0RRI5VZI4M1AmImIppOTexi4nGmesHrC
K15ZY5NmNW91ukjWwSztyyBCv2Xi1C2fHuKs4XaLxgRCILG3kxoFEe7j+MaJbTZC
d2SKQkMn/24iIj1eCcYo4UKZ68+Lgn87Zhyc64D+95C5vfIVdPLpfhhfYZIibQ5Y
hToBpulCjuriIVxcwFPOGeo6v1Z/cQstVqmbR0WOlYrW4dsqTImVtqw/7R4cnKPw
lDLB/CtC+8iSECp+9xScpL19HgVTkTKltcR7P3QoEhJhICFygeDNBOhzZFc7j9Zj
CPW7GPf9ijROqdCNp4Qg64h+k5nJ+kR+o+poLVMDzsTw2bBx74P5lmdLlWiEa02g
2hgN97ZtuMPg/6d3YPEivH8yrndkRnpygFojagpsuCoSrCixX44fWxvkEQTTVUhe
hfnx0az7r8JlgV/MpDy9Ei2C52wyxqcDFB8qFi4RPUJvWWTyul7Qd6E2UVlfqPyQ
Z9J8RNMlOEESvKY6S5SNkF6riMicqyweE/1+7lrqyXpSuR6TIIywEgTGntIORSJN
y0P25iA39jnBdParrhgLlEgXjUABfQlJZFin2tlfefMwuA/RCL84nXDoz/bMvEgh
KlodaGlO5yGH8Zzy/uDWlg6GeRtHIB61oL2CF+NCV6TPrt4NQzsaKlwqESGMm9SQ
kdW0dA4UJlMZ7x6QpZbkcTdM3B8I4pTM7zNYE8dsK6/9RWzV7aJmp2wR9glGAaCw
dEk+2eV/9FOKCcOSnUd1zhg2vf5Jnb2/cPbElG5DRernoQFSiyWNG387VgnJ55t9
WMu6bmZyskpl4Gs7DSb+xCwSCAAqptnQg9qRO3Cvt/l++X7YZJhcicQEIJ4x7UGT
DZo/GnSBZzsxevftgPC+Rtj11Dnyr0/FEaaJKltqtW1Oyfu7DFHAvze/fHFAqGs+
tI5tKX8PTOJJ9kXdrMLmVZ8W7Mvk0Ye26IOvFyn4qMBDn4PA/u0ExX2uzJbd3/Oa
TNK79a/FgwlaM+H24G9VRVqR24/uNioNrb/oE0F242QONGIMUumWX2UPkRDSBXMY
4T8FoReKmE2yr/LRf7DMSBRAMXw23BbDmRsAsg9kAamsj5aMny+ByDq9N7OHz9jj
LkNJD1gyq+WfVaV+v4PhPfHAWJRnajwpyza4LZQ/MG9EOFbLoLs6oaoQORrX8YEj
4gm/1ygO78fR9D+OIx4//nPjEa+n0A3cimpN19JWkZE=
`protect end_protected
