-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
f+ptWocOiAstPfOQEfDho/GUfCsLKNZSX460rrOhowsqMDKzV8QktY7TcbsJ7PVk
so+irtE87LH3ZffYAHtxFBmZeB8f9k2dQMhzxSryTqtd4fHN7EiGC4bv4mjUuPCP
RRseInVPSMrni5NR3FSaw2UCXodspPZNqJzyz44fWBs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9636)

`protect DATA_BLOCK
AUSHXq9JOR9DO7c+GJpdFgATTmy4FWg3jvoXvgHwOHywxIl9dcT40Z47EDjowOud
EA89DpMwdEDCokDQwl1mD4MdXrLNKl5SrrO7HrDtmw1XY8220AaqqW5+i6J+08TC
EtdgPolGwkhz0YM+utVMT2f/w43kn+6avBbTRJb3G1hulqALyT4Eyo7ShH1veo8u
A+0bKL9i5FWh/0A/cqRl0H8Bt7neUTpAFe8XXFtjmvMr6Hgjy3AJs9tg5Zgd4Utf
Nfq7l76Q4o+dzVV8wgrB9HqZdUmVpN7BgBbLX/RCrH6D4JrHxImqbcQg2DZyljOj
HZ3AWvsOpIURLQ7g5Hf/WvqjTLTdAw8hdYqAXMx2Ru4EusAnJrE/jOjclvE5kU9T
21g3p2dc/2dx94oQfXP2Tsh4iJqTDqIvnVKUyKy9hJMxe0Az7DkXDKPjkCz5Ir0u
Eb7beNsoNSmNtvMT99tl35FVji+6+VJx0ReazhiYd0OFfy/AYtex1NgQmFKr56aW
jLLUP1t6TnEBbh7A1rLfp/nEtm3hov7/LVbhHInfV/tFIISou8lRReqRVpGWVoQU
JdXqU2XnhTROTSNT34hNKkSoSEpHqCB17LBMYvKx+h0DfaBl8y24L03DSgisbJwI
WujFVFInvQpjnaEO2QIJRvXwyUKsUyD3OUDsz/niyoXZB/86YzeOGe0bXCD1OhRU
J7KFbtY+Xm/0E9gd7W6cGJkoZ+cgW9NaMXUYLoQge0kXSaWbVlRyBlduRkkvw0mX
A+zdLXaiWV8/T/Wlc56hZlYpjbQQjMhdOlCKcj9YieU8uA8C34nAE/jcvhd6CxCx
Kx4SY+XhZsv87NDRylbBao4Vwqcvv/NP75vHkgp1Jflhb8MAZ8lczfT442jugabk
/twYz7w0Js9cocj7qZRRszOmaCF4MAqM5lRW3DnPvEg8Tg3MULMyQZA57gV/h3nO
yQ5xggxj4172WEp1iaXjT7LlnkoBbfCOk+5F3Lx2iu04EkabdYcEvn16MG2jQ/s+
Jvyj3CIBjSYm1UeqoL/0ITFQNjkKFKLegyZz5zMar7ByGxcyobeWeahVVHNjSEl2
EJe4XpuZEkDTqYlMjMu4GKz/eoFoUWW9TupSisozy+23lZ+cNtpdc2ExIclI2wVP
DRDSidXEoM7/20fPRdtj/oTrVHn4CUB2KCRbafSn0mGdF44IdJ9rV/zw7kl8RFha
xtNJRBdBA4S0sXPi9SqFcxuopJ6EQ9pRWPI0p5JcsBoGlpsQzZ8KduMIYDOHwoMS
oFd/7y0QUWIeFXXtviA0/Ux6X0Z3zwPyH/atWK08LrwUcZGxQahqi+gd1dd5IZD0
tg8n7WNdkraSyNMwCZRoHz5D3mbOEHFhe1XBjCtmvDaqOBOAYVPavC/IFKF6ACCE
jK/p/2K6jC7TeyheP/euOAlBYT25xGY/BogTH9mMa/3YbketX7x9tqMjZIvG/sKp
r16EXtK6731Hda05riWPqYDz5aAcOVX0B3vxiiP46fyjSaO8h7DoLJOcvXFSJ4zM
AfaXhA52kcIWV5hAXpEaJTKvByH+DfI1YDc1E2Vm+e4CAwrBj6Z2dbXS3F6tfDbP
eCx2scJaBrB5xqWaSOOZlftacfZgZH3J7JF//iiaJJZhKI1THfj9yMxgPDeWc+r1
4S/p3LrmE5bZFz9IDCHV7t5u1suGzEny9tooAFPZAAWp3hIH/abHkZ2NO1UCHqaM
gzo+ezpxS8WnTLWfuGmUgurBUckVL6EDqm7rzPcVWPk2RfBdoEMYoGa44RBW5gdv
Yw66/nObaDQ9TRZAco/FN9Bn2Pb/HPJtce0D2KDqKf9O2r2sGSSl5O+XOMa+wZ9b
46KdxZrJQ/Th/y7wxAcOB42SFNFE4R+jRa9iQqC2KbzC8V4yMixREazHuNFap5Z6
mKTkLePRk7twt0Q2RcsM+HMt/yKFboAvUWN5d5iMFmw6JK+zt/uSEZxmuvbbkS9x
qHrsr2WPyBXk8mUVxFUbbfyubx4irFqlRf+Fcu3Laug8Is9hZbOJuEAVjVenWBiw
MhoI8ZjlT131RHJbiExgAnHapi2nJf/UBTVqjAGuz98SQ6kJ809/EF/pmnWYjlly
Xqcpt6sMH6ERzAMhdeVXRYvoy+gi7toFuikVnakazMrgepvzsyIMemLwHseZUkr3
viAys0WtsSKDfkCeTmP4CF7h8UiW10p/HGYgmpGskEVMeEOxUMZGhXzqnkV3xyCt
mZVWVrVi27jbREoyPXSir8tzDtqjkR3Ps+W21u3V7z62JEqtl2wejKIF6uZs3iJC
0jXb7zp/r3EyyqadUat5N49Xe+hejBp/e9B6coxCSVyQ0dEnITdoObGF0QyKjq37
kAMtW8zHWjrw8NLn7II2yQnnS03nHMd5UW7iVeWqmac1vjkV/dpViUMrnFIz4laY
jmzijWrMpGdIP1y1GSI7W1UAd//sGDkOFsv4Tj7Ev5VuIQ32p03kQ8FBKxbF57WB
kXtBfYKFgSrpAJJCXt5UP/ndRNLPdPgPmh/3klg0+X/g/E4oE4KD1c/G+iuPNfvS
LFM5Tb+YF2v+2Tb77Np0f6Ld7OutMgv67wzIxYjdJkM4R/wnuaVhxRfqdwkWGb6N
orf2AvbU7+0Pbkq82JqEi33lzDsbJEmweqmv5AHsBVj7msMr9HOTvaP1kDbT1hIx
muAn1mZOkkoyzpBMCQdDbrLqH61couurq1OuOytYZn8M/wffds5lvr8W5TU6SzaZ
MpSTXzc8uGhbt+aShv5HDTpn39VVQY5MulLP81hsbS+Wfdz5OHae5Tn1b1ssOaYe
2MX1yJGczjnwQwykmWo19ZXbrsuDWqn7VjeJIWqZVJuytA5wCzQFX1fftMtDB+2z
3wxGumD0E1rtfOQFiwUxpn9OFOS9KEc8eYx7qr1Vkvr+RYFcN10FfjTap9Y74erg
QSDISrgNMFy3+bP7j3PoDDi2DKgiT4m54UWvDW+rgMA2BnlHjUZUDCub+SAvRkiJ
8vy4ApJNn4ah0iNMSJ/ASPDS8PeHeIXc5N8ghz10EUIJdrTChaUb8PCZ0zJnqwxu
Xr1HzvpggyanWjP4CpKG/B9riARRfWdux1fLzC6blq7HGX8EtiQZnOtPGhKR98GA
/nW6W7pE9BWF4cQhvATDrX7bVT0fsHCO/WzRfttb7EE6cF6efqe9HP+xnB8lwv2t
l/HRIbWYb19DxT3Mwewa1u80ZOxkwId+0CY64CtUxpQEcomBDo1s0Ot1maqBIfLX
NV/tplko1JxJAZ32QI0W7JfbNqW6d2eQWQ4dKGTYMbenieFjkTNwdsXXcKMlHEB3
cBjV2hRFetOSjoZsWfaL4eL6sbt0YFWlcW+CN0kV7Fn+jcErtAM4MVbAWdghek/a
kTt5NYiRr5U8q2ATwo8/liEg+/2Q5OM0wF0LhrnjAOeseZ0DFjaQzpGYyIRItv52
d1X7eKOq/LzgFMjqoF84U0sROPisQ4kL9pGaiiQ16xhd6kGJvbRQR19NSCrzEcr6
LonaBXAq/EY9b0iGjdECYDuZYXwVNiZV4Mw76gvS4FzrKjyCYHxXG06jYUhWS2+V
cmkNC7ouBY+050h1RkuP2XvGsHaTBKfGTFghjzWwgRXuMoRN0q1cYvz7PyY8Z3rQ
+uzQ9qx8npN+n/Xz9FevS91uUq+h2tQQEIl5HCo7+MIL7J0qYXRDYVMn8xXJmcF2
tO4bu9xxe06pOoLPgCVFy6VALx15hj5UMErwmsBHmNd6qK6fWMCqK4Vmr7MbIlZP
mkAa0Nsk4L0KIkp1zR3AaFaT4YNVMAfAvinBnBplAAui1G/GkcdHVVJfYbDqN2J/
S43mfeBNvvT8wqlCs4vgc6T3oBw+e/L3KZYMrFB2S8PD9U8Pi81wY/FDamENLhW7
v1x6SXFBRt3hZURLfCavtOI45VrDYi91v3WnemOXkxH3dIZRtfspD5JAATzy7clI
h08+zR1Uj50ifDpyIoNvBWXbDJedub+4rNeFZuCNYO4WMp+oo6lfvlCNpneCP8or
Vq3ifBPxaeExqv99qv13eKcKEPK1uepmCmC1cfYILej9WGkgy5lWPYD8g0rLtPU3
8j0ku4cTCD0Ja0bM+fVlq/Y6pgQXIL34tdjWskfRPGNFS6mlsTs7M0Mq1aWQhyBD
TI1EED6berG5d4PMJR50W8pdDyQRbC/77pOpVxer5QZUnekUEh/LBQqOX++B6Ps7
l7XLMC0Dv/i4VJdbTRPqWcaGr61T0nnvmJTNUUgK6+mkK26Mr4RmNpN3jd5MjBDt
osWR/61eJpd7wRk3Br0n4s52TYoJtArwCxqGCLgp+LvxchRh5AdTjnuVId3hJueC
Dpg8EBQgm4XBiG34aXVLLiip5CmxBcBf7AGX6t74w+VmENgkjP0taSsPAD1OdODK
jZtfHWuhazqjTLza5Gd1JfQedzPE0k5zw2F/n4asx/CMA9uW+KlLoPBlakmoQFD+
aS2U+jQQHo3xfqEwggIG2Bw3YGWRAVHXk4tQzx57kG1AEvxbKa3dtIVDis6X7FRK
xZrjz7G0klZqkHa9UiOEgbsDRNz7HX8yhM0GpNbuQzpjF9FxZp0aluGhCdPp4uLx
Ruajy3ztVD3hbGSve7gYInNOa6JRlaYPZ6/5nsNHIVFnZ/k+a7MEjwS+XxefkjQf
B5GLanNfKGK6n7ip088XSnvoTD266o2yPSeWexEVjdCJdpSCXG7SLnnMrUqtJBas
qtEq9OmpXOfcdK40vivxgy/fM91S8v6kryF//dr8XJkQouvIvHtJgAX9JFpy0O2Z
4JTYHAYqK9WIAZRiTlfuENZOsth1RE+Q+KuBlHqZTan4paL2qNYZMkDvbKNBb47B
9w0IiSYwEnYPCF2zfmBpF/k4liQNw5khj2YCYo7FRYFxsBrH68Viv5BicWzvicyV
pS0+zTvAK89Z9xNxYD+gFvYFDm6zxoUiVqVHiE09+5cWd3xCpVlgvGXUjZ6swOd/
yem1/4pNbg4ebEkoGzMZL26jdLa2rjchsNoGCrk+8atIzaoOqX60nDvmpZhLVmEa
oJmJeWW9np9QzLLT++grBdwS9NQBC71Let3JrvZSY/U3BpgdCgANf3bU9mFpR+sV
Ign6PgLmJod4CKsoyOfA6XsE3f4yfykVDxMax/zyWfVUA+jPn26dYfBSPMw5npmh
To38zLyPi/OtuiRoQlpeg01v15NKAN3FmBswHJ6pdVfF+qjiJ0Y5lTu27bfwwkyo
1aAQQAg3ds+OboTZp79du5FF7T18V/rxNY+f7ypEHI/qDTDFEsz163o/XRCYcN1g
m6dUX92iZRqRp/ZS47VQsvJIHKvMb6vwugIBVhlpJy+JAm0mImH2cSMj1JNZWcS8
jNcSa0C/AHcd0qENXfb+DBIkPZCBQlbun69as+xMdisjPiqjQd2v+pVV8ueQ6Kb0
ItfYSFeOC6Wxyx+D5UylSohiRh7EowwZHdm5Gv+YARDrHLEvFNomFTfxaAucb4uc
RzyY6vs19Xt/1H1Frspw3egma3b3teWO00VLtZeTurGHxZdmisbx41v3aZvXfeIv
X/k/EEHm9vxRtqFFA55WOj5Y/kIysWg1q0JQJQa0RXdoFWIfH1TuwJheXOPux2bv
gta8r0ecRBKHZ3S4TEDDLSLbyXVXHjw09Pd8SzJKvdH81HJGyO7rqJ+23WzW1XNJ
MOmFrW0oqMBUizwc62wKM9czOntwxJ7ZFpbT1h0aIoDgNjVOIrfou/TCLLaQL3ae
DxhmVr8BNRYyGMb5ZWR3nFIrnV77qEJ1bBn0nlnig6cardY7WQXmbUrCL82+kz85
suoiw+HxEhoq9rvksgkb2qBSkkk/cEcwxYy9DmgEzXptEmevPozJ4KQcVyh5WwQI
/FbraCh0nKUWseZOawnfgJ6WXx39w7tgz+YnvH2axpvrAtrNAWVh5BQyKIISJAAZ
nBJHjj50rvCM4sNu+CoWhERS6CAPd0QcIsxMKbEQBwAI9cOSImZgUxsFNiF2+bKo
78U6C+YLRpszvYUc/W4DfWrAEeOn3UESMb51pTwhZuA+DZsV1q2FDwnRa12t/Q5W
W6YdefI5E/CyhwNwDpDcXxlwRSfB89xTfbKaSNUVfXIXm3xNCv2/QD+SQX2n0pVJ
UG4ojP937HjH2OEEBsxuSQtgLC/9VfLvXp+14SAWogvhUY/lBQ8eZdoiYe4Gqk4b
BvTYUvqonjoBzc5oS74uLw8qT6TDU71bgfH9GIlkkuTdCxG9UrcQVQb8I7w1kfcP
U6O0SlA3xI2usZaJVvUshbQAOpSbpuTt3/zK+tun1Uaxqn/XYy7jPCkSH/DCm8aD
77YAFnsWLFroCup0hPlF/KbT0P8qgNeK2HprgJVDP8/yMkX3ywK4akAnyU64zNZg
kcATAVsESLJOHqlee/4kkvdZzZk48z3AnnFKacC7Duktbp4r4BnbbG8tkdtpt4KF
gwJW4lRPjbYuhoT3Nw3tZIthOCCkFe5EqGQHltkYKoo3MoYsnU6v5EXYqRb0oVnk
lgMUIMBFKDpLwSRhiPodqh4sBJOm2FnHOcDiKcOzWkIhUMCKkfTXXwMtvV6Z+1/7
wcNVhg7mu2lv5NLJ3hGFQD7cUq9TY/9OqnD5IPxB0fpsVX0oHnqsH9LLPvK7qovu
DsWgGPEQCVQ/AFH8ua67+LTUl5h75PXJo/AYwLgia/UcFrUC/4JKX78MVe8yDnxn
FvQYzFO8KXE+ts/yewFGkAXSHTbFeYt/0gPwp9aCgwsJVig00wi6TqOSIqO8LhtL
9XJ9Ca/9RHRk+2WC/nmiOrQjB3yN/pqMg3fKTdLRRxIJqh2qR+VXGKfdNTerl7n3
SJOqLTTlHefgeD9bm6vdYi2pwOYmza+v+GOeFwzaP6UWyIJ9mdB7shXNdwqbMg4C
yNNcRuGAC+0HF1ZjxtX/LV3exlK9ulhC6HBJ5rKwewzN9d5XBkm4ZaziuoQH6LhY
U3srmebMgSmJe2f5pLCoVsuopT+EckamHvhQbwYV8qqtYe5Rlk4YbDOF/TB+AYGx
YXMco0lb36mN3T1AyxP/ZsLP+ExWjXYbgrr0Er270dHI6Vh3w/Q9y4BYZ0MesPNn
sTmyn3Jtu3wwOz9yq4zIqmqx3LVxRZUX8onKQ4Uj6Vh0LRDuc8ktOTIRMsA90Rsf
ONT4z/TNySNT/YtQ5EzVlwxpI7LzWHCoh3TPXuwo+4DO70bxNk/xlV9vt0Jm02eS
a1QowMDfgO/CauziFkFLUjOHnYZhzwL6SOmmYW3/Ad/kTV1Np3+CG7aRVMMjbDcM
hrCygVDBQZSGLJ6qNXNyyQhQt/DI1F9IWkOoP6Q2RoRnY3Er7TxidNJlSMft0JoL
T1uTSq0pshBZ1og1Nqdp/Pfd9xD9taD5PthGSHjSc1G1tXYJboSFvVbMGk2DqlSg
4lVoNBVUGujPrsY61PE0PBjEDqXdbSbNLykpEpstxxCn37ps527N+QWL4ZpqNbsc
QP1CiALLtNPOVPtM8VuQBIf0OeRSASBg47ir2M21K9DBE5oxN0sESOTYLtTVgKhE
DOszqc8+A7wmi/okAV30atuapu9YjHmuP4/hl51TKI1mjBWhO46mHFEaJdUDo9+k
ALPWlkmSt9DEdLBGQtYRLV7C8soCpsnQBbd/G61Bpa5BO91slx2uvD6psqdFYOt5
9lSniEkzUhGmoU2SJeFR5DVWmakWwS0upjBF+JbPZ0lXr5QX4gZokFJyUgKgaq0E
+VV27HVrinN5xRX00f0XJ4lmG8G5choT7QEpJHa/crczuORwbSy0t8Fpj05g1mOt
1aBEMJr/9A8sMfDl0q44P//233EJjnDbj4FdeaPMDTwec6jE3pxdQKnWdg8wt40y
4O4rJTKNPnYklRQAYaEV2EJNlnVKDI2H8xF0YqV49RnOVp/BLia/irbdWw5phyvG
IILlhObzkbq1jHNC8WjRN1E7BrH1qItFjJgYfBlYKn2TWfkQRu32/gmAzS4KiWlg
eHvKfh6EzZAUhW4a9AldD29orz6sbfcC/0+TnysGUBKNONtNxrLqCiI0Q28pPtYX
bcf2xe0bXv80WOcTg7KUd3QoenUx9qLcKiN1uJ9fqkWxcKt2vgfJgdBWEYr6D+RY
Mcmk4y1/qC+PtUNeGP9ELhTUEZjkS88vaft/EABGRfxfTt4Eypo3mqoyMa8Phvs4
t3CxAvzEhDnYHtLLqMvgHngzrEoFvn7c3C2IPsP6xw4M4InYLAfhE1RW0h8mZgcJ
MScx0E+kJBeFziPklbDU/eOZnhdA1hdc80dwAar687BpIB5ofZqMA7ji/d2D8q4a
XN178PpiMWH4Xly2J+jDFgJDWOzh8qhbFbVsXpj+lvy7LG9imOs0VXlDL7zmyLSm
uo7mMZKTobj9cJuAoVmKfXm/PN8wX+6wRyITSA19IVw2ycsKfzWii/1jH9ldu1H+
fw/ydpKB2VPJ2sZVzehP8zt3mmLSApGnWq7vObemf7vUZKVvZB63iTFG5SBIs4Pz
NgjV/YkwtwOrLSSKP27eNnHv9iSZigCtnC1EF9bD+fIvUNTQO6FOtb66w4M0Pk/w
aPy0//LOX8cbAAIkl26hT9xXfrIiSvmXbehVE2aF/pFsbimrxkDFq8SqyUczeBgC
8oiI1R0HA7pLkYhQgsMgN0LqbCPNU+SsfrEYsWWb3Ssoh3nxuVBdE4Z0CUo1a9mi
rQZJKwVVemkSZpDVhMElnFvJrGsGmXk/rjz+iGUIgwXxXchcFIHFAtChcv2tn5fN
T1R6FON8boLZCN7I3lgPb7rxGFTFrEFfPkxMNHbpQmyCtKh2kU70Phhd2z+wbKg1
izFEjnhtdEN4/S2rs1KNR07OUEianFDnMl+ucPrLV88p/+fRcdN61I9ThdqPGtII
L9j4iVIjgcnKQI28xyNwv4Ci8Xz5qCpUbTL8FmOmVSJHCJ4JZm2g+ApsNXhrAZj9
jlMH3x7MZ/QW+qmSk0BZhIxmY8b9th3S0Gz01YQtw5cUGtClyHKf9W6L8uqt0QRK
UsTpOhjLf0wG4zWilPl2xFVCnEj/ICJhysrXsu/jD+lnh8WO6aUd9/Akq1Bv1drC
MZbN2hBn/+32VZaxXrc9g6mOogySyTP/6mjPYVVg1Wk9VoAl5xyLGc+dzOjnUQ1s
vAS7zBMBtE4RW1P9/dTOBgauWMaAs2JPYjSIFy6mSnY4v6xv0d4MSRsa6Td4fI4i
PFKMCor7xCKuzYALc0qtzoR8fcHIofMFNQLAU5RE3y4VbDZzyUlQ7uMoqtOsrLz9
reHXy+Xa2sxmrblxOwybOp/YOahoSiP5zM0dXrsCvWjf2BErSMjdYS7j/bdrM+69
656cG/6dy6qbwkxijGnD68BhBEwrkRI8JBEZAcKu8qlyDULkAWVw8DiHqptM136q
FySK5OfUj/dDNPmdrJFWIpsv13qvZldBbjs2SeSJpRKrwraMarDwQ8+pc8jSUdlN
LiWENz1p8IMoZaCoC58bNr/tkUhsM9FR1RxP6QTEgkdao1GsNa8VGBL0Vcb9clV+
WyUGY56Os/Ar71RKcMQZYElUnA+iSG5omKVMV1zg8vKTBR3h5G7gM7nN5UTrBAZN
sPWMGXmF367mTmWqD/P1AhJ4s40YcNYgFyOahfEcGk5NEFefNLRZEieneV63adMj
m6+4ZvPv+2ItFy5L5WhLNoCfAl1uac5WvcMf1OdtTaJKDn8bUaIVce2UmFOknYrn
1bNM/Lin2H33/dpXj/FhqJZi9fmSj5Qdrz8ABYY6QCDzd7sJh5cliGSLnOJSehy9
fPQCk4rw1BMY/fXrKPNdIYJEJbdGbtKhjcAe6Zugf8/UTGLgsLE7miWp9RKz8DxE
AKBys+kpL0lMMx4Ybesd4MIqQr6UwQahBg2OYCaxgiN+iYbsgTmGnRS0viLGqaRh
1Tx2LsvEoerdnK2STSXXtJgg826QXBzBYsMle2T16b7NJAKG0iLqHUfz1oZveNQn
uGmnaIuVWrY2FME5skZRu77Xu9D/PnqNSFr2t6A1p79DMZzcMt/wmQgvOqmKKbNN
behzpIHG+v+OYpCp3CqZDxrxgiShCoApgPNprNm1xTvZ3M1B9UrL2UUjgit2d0EL
M/8mMUv6r2KM7MxH7XUzPBxmbE1d6QcTXoFrUjpWtDgVt5FEsfuVoKIW931m3S3V
PdSNTJkxGZCXjgDDmBCjinj3/LNt+0hc8IQfpena0tDmddrEDsAbwbZzBJHpWj2x
DmxMtv7eQC16yRmW81He8wzOIFbXR7YLVFS3cE7F99Mn7ctzP3Rd20EA9x2XS4Rm
KssSJeHCqyb8Aws+clm9EahhOWsU7p4GyIOFmsANJVccqKe5DhKnDKSyUCaxXmY1
/Q6r2xmUrtZ3FSGfDKtX6YEfCDpTJCSzKmyhJ4d7suD5l3KIQBauiA4mJfgxyEqn
UMJufYcY/v2m+qAZ1qWR3zgKP2wz7dC/HLraTIuPVE7G1aqmZlxCjfawoPS2S6gL
aQxvbbLWvMPXbVJhdAM0B2Of/20yRwQ8lQUPr7YAp6z/qSHmMsWqEw+6LFFjsgYV
5CQRgy6Oc4WvbDpaeiHNQ1o9jjpHFWMBuPa40rJXyTvIZn4AsQJIRAUvGlW/1QIM
HwzzzS+zF3bSOJ6xjO3waH2t/BMK/za0y7F0ZXKznVCmduhjDkk4YJtNvorgw4+9
VVV1GivBJURGMRsBr4wYkKd220sNuFqABcLzUTxR56J5+BAC//S76kYH66P19qco
HLDDIO+u1J8QE+fUEDR1icslo3P1QliRhtGR7EdxASTCez53Kok5H42kQHpBpG8i
z0+kBlgi/Zrsq5BW+zoZVtWzeXpV6WMqG/Kr7tH1LZpt/wDuvnc60cSvCaY3yA7v
A7526wtxYihLItHiGbg6f7jwZQxo3lVzBszq6wjoF5YZ8rsqpkYFEkK0YgIK7A0b
9XucNXQJk1iu953LDaJu327qBMmgUzXq7OGXmlI5mmE+hSnnIPEGF+MH4N6rMh6E
IHWCU16dwxGGWwDAha5ezKjZ7g9CKSD0q4nHcWelXtR29EW1FeaREzRssTE6+0Tg
+2WLh3apcbsJ+CE6F0MKHXJb56VJR0ns+Sx5mctmOkQKNPxm2h5SAOmjTUyzmmmq
DHrX/BqAfT9woB8/PcChYIjWxywCBHo22DTw6BxvsUGz0twzpBoSK7uA6UHkd34v
hD7i2FRHuwxLABJwMrB2K6KriZm1IDgjV2xMufZmExSwiceOlXqfZjJ35BsIwiOs
L1Gan6e6iJm7JiwqkowFCT39etMmp+kBEGF9lhSIAD+ZcNqNy4jEj4pNDDeEnWp7
L4iHZT+AD7k96dQ5z2uPqkAAcbKxxOxMdgxHMXF4Ysfjdhl9cCr1pttG8fWsZR4x
e23a8JgaD54bNDHNA70RqoqgERV9df5lTH8sM1NJ3YjacpPVUR0Iy99MrbrPDTuJ
13JSKRtQJFl8wWkoMTFft0wYQuwRdpbQNiSWfDH63B40gos3E0kk2qZJNoYJL22C
AQ0LwHk5sD/3H9Vr6PdI79w24iLFNuYClCYNZnUa1QcGkqnx38K6e6Z2fBYZ2TQJ
TZwJvgBcqCiK6uh31l/5xjKpSs944+uu4oFDS0xuI0HGbfYGsd7/ED0RS/Ick54V
kRXPMTw3r+X4uGE6miiS3ETeornt0hybGke2ckkUvdoNs/EILkyInatNPrKyQwH8
seLqWPKSxX7u3lrxZFvyXDa2fkcSnUy0ck5thqRePQ7mGOh0M/zJdu+M3SOgpUF6
PoqL/8zJp0ZSt0x1E8QI6azdLn/g5Yd0TIz+qtGBuINOcxvrW41hx0+DdxS9+au1
0GhEElNSFs4tfDsnT2S86IqIMW/JR09ahrOWTgYjFNxDuBh96xxjguEh66QlhjQx
wlgcQxucWML1JcLMGMp8sjiKimJTc9vZcsW+u2t3sqHm3cLiCQUpV5B9pDYcFcHf
JifF+nLVG82xeHx/cIbBHAMuFy2p8kw7z4bBouAPDmJ8MjAYRzAhDWT0JLHq0U5i
Tprn44KtgH7v6Fq/R2djIo1HJTyeOqc5b+oAn7tF71tnbUJqoL2tmAUJJT3XI0+l
zj+FUeMO7AfAN6tBrLR2ik2yPj7zVWVsJZmP/+sr8grNeNE9cg2QsDpsrfXiatqa
kR6oftRABXsF037uxKBE+msLpZ1x7N3PAyOY6IYtAsXsnizT3twXWREY00yG+oNU
AfKtwUTZNeqg+vBsqLF0UVv7PkKWJNNaxfbY64tZxcAIC3zdyqLdsaBEkesEvqi9
l6+8rhd9aYje5IbSJGMShCkYxf3aV88/OHOaAtez3VRIFv01A/4sMGA1YrMustql
gM8Ud9Pn0X8CzLDzlLDpiB3vwppDKECOaNgier5nWys8A+NIn5iBGGt14JedNY31
OZgApioo8ybB0y6k1SBV5RrzzW3B7u1ARpsyAjbcH0ch2AOSh84Vo+SY9DF4C2Bo
Cwfq+IssC/Eof8Hy8n6prjKEWsLJGRt9jn7Clz0zhebKR5qNBBj1ZvaxyiA2gaWF
AIASKpZxLX6ktmY6yLqnRYc14xL93C3awOR0sPCvj52WJys0JwZoNDsdOOcvUSeH
MEx7lqcmMgNqSMO7TUjF9wqnXubj+OQgjAygu0AOSRNmizsmG4N2IV4c05HVqWHr
Z4GRIggN7lLeREBTrbeqxl2P7mpTp3aFeBQwub1JFRo+CDyRP3+SALRzSa65CgBU
qDXw0ufEc6JBCLMbdf/22HGJBgwfhO1mLwxCOsFJE0Hf87yRl3BRMWFWiX/++JX8
2kg4QzUZF89pzYLzhSz7UGSFOOYw2+TmTCw4X+3KtuicEnOEk0SIdzOt4V4AgeZo
yqpuh0RIB8sjt3J5YU5GLQ==
`protect END_PROTECTED