-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
zpzAo8bRDJY1jiNVPx58TEZGVCDDO9FbYMovyyI2ik8RDc3guOdIZEUq4N4mdOIg
/+RVp3zUp7quk2jz4Pd1w/PPLFh4aTvjqpbv6kWfLDw2dkUAEbI62QRVEr2G5QG/
mlsgAhgL2JNRJ+awhCfCJiBkdSfzRDf2F3vikGspCy0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7344)
`protect data_block
amLf4j1iHQadijXbeIpjrBb8DDVcQQ6wZDVj84DDlREZFwyfP9oBEtpe48vq1NGc
94GEK/JBfhv6D9BzBzZMKE53TuASWebuLeI6JO27XHkIgsC5aBFugHvVxWBG+Zpu
pgktQJVdci2neY5LMFO52UX5roxghCAiH5TpeeF3tOsoux/Y6pPVW9AWZH69jDO1
LeB8tn3w+4G0MHeQ2sSQiytQwd4/gYys3/ir3chH/0TQr17b+bESRNBcXjnFE4Wt
RowR0FUSv6DDQGFfAXxAejclXpWMU3bRJexamuUxB4wqAfiyYf5bQkLy3dXG+ZCR
eE77jOaR2zAc4mKPSdHwc9aOoPs5MX9M8f1wXwCDz5Lcbpq2dFxWDB1RqcvdX4SA
LkBghZuXTK77T0BI3vQGHTEAx4l5+jLB/DyBNc1AX+edcrySIK6/UUIuhCUMBaP5
aXI0il6Lchc/esaYttF5BsteNQt/FAZte0jfYZkRLaC41yNzlBi5ckoGCbTTFNZX
Cx+PdmKPR+E16iajwVplRTH6yw3l/32qkgtnG4AUvvUE4NFuudXhrCY7RzTbQsVt
EF3yV80eRO9VfFfYc7zEVaROQ+FZKr4dswNUBUjmUqB1P3pQH8mEXXC/RTpgoiJl
6DnYTSWNpumzv2B191Dmdd3UZpomLvFWLdRuIE1SHATl568ZjyLpPClwg7PERG+U
z1tZfiC3blyyoP1Zqg4eObJ9/j5H2534KLKEO5yKq4px1Uv0a7HUGLVmi2qpBvQ1
UAb+Vxi1+ASWFRQH1HvYFZ/V6meZSXHepp9DPuXdsYgRG4xgaYXrI5ri1ZHtXcVX
Tl1MAc1ntewlt0JB5fMRmHiWmWZgWCConFJZGg44BBlN8FUsLhoQaQakj0S+8dV3
vERy4snnIxuSB2b6foDCu9WPFAJNAy4b/V1okqgVNkaBwgLHscttFRtGkySw90Iy
z47p/njOYajQNf2BrI6Mv4mI0bkV7zNQK5GgcSdc3bBb/x1o4kMnBs61QMQALsDQ
Cxwowr4SD0m8yLbwO4hKSyFWegnY4AKk3sMmH9CsppvAZzaYuOvpjQAsAp2A/jRa
ZDcE1FpqNqla788ZMRp/7l9ZO1TEJyOCulzKfLLNdQ7k7A0/jvNaUrewvUlnj3M0
Pyb7e05vUnm4k1JllqiennfZRZCa36tUuhMow/hlFVG8y+hz9EnrkcdpIXanRQxL
Iw+29sSIT3aSg52iQNF3uXxlV3wNJPHdrebcY8srF2rgjV8kQPzI6DTrwgPfdmE2
vLTxscyI2psTyDxPPt1gb62T5xwxSa89kKKIRx/Mb8jqT7skNqHyMPoVfhqufPEW
VSoEVc4arTFA282+mMhwPvqclFQfn6x0Qhf6fSw+nbCCAzmZRGKYXleUtxmmvsCA
dqWyE9L9i+0eF73h4p4opqo9bMvMLskVhVPVwseB7WM0F/BzSkyDVrFdP2f93Qoy
uigHFVH2mBOk9RQ3Fej+N8xtxrwDPPsWaYl3UhjPW9Dw16vYQFCl2iLBV8Y8ROs2
0PTNyJzysCo7Fo0H68D5ABaohVqGkFh3qWLKGAVWWn75REG4UyB2fwKoAHoEC2Rd
MVKnbHtYaCQauX47FKd9im6C1o14wAcwRYjnWExWuYojiUrFnyPb+TtbHteubwr+
99AER9eSxu88SHyh3QSjZNZKZrkjgdYaTA75hduVZcdhLrgqOfB46scsjqK/7HHZ
LE2lNoo4GsiXOIMdnyKgBvx95TYipOok81qhmxJsYjIMZr4S5+HpJKH0G1tUQDY1
Wh+VAezobjih+eeDLmNPsymb/5W4n3PMpCK/BarlwlAVMEFN3Dygj4WZgDCrKWxb
5nmlLN71utGSwvWsMA+9H+5N3PpV3MQ+3g39HheKNiRz5UBdBCCiBKZTcALAbm1a
pyBqIMzOv5rhrjEXjKe13jWGcGYMJu0VSMQ7OfNIEJ4daVEqFuwTVMBo+YhAZVx+
J3fPEo/OYCzBR3tdHN+SQcqW35xTyRCU0ogr6g83PzILKU0akxWX7i/zDVRQDWSb
QUTpXXl5CJXpWMb1cWD8PoPDJQA0pwZS8+ThxHa1f5JalHNzAcUUvqNgzgi3xbAs
6LHmWMjPjh1Ebg/LZVGQuZbt6Q4fXGc3YCv4O+v4Lnw7RmFalib38u/vCmI/ciJy
uEyqm2FEGMLWmNjC7eTxLOnkNaen47LsWJW7MNUzu83gVqch1vZAOG96gq5LORNn
MDAeqGf6SKb1E98RaKUclD+zV4chrahMUshAHAXnj0A2QlwwuPd6j1hcL2TQPfjT
uRZYML0dDbYdc2PNgtUetbP24d/YVJRffLPeHEN5/a01hmJRNdSZz/I+bPXdc4OT
U1ayZAoPmKrp9EtpgjwhOSX+iugNT9HQRLznPqro7WKiLEDVTJDpJIb69r0puvbH
mPW7s5a8Nss4eg0CQGeye0PvXXJ86QAkWYqnK4BMvipndjrTMLSFnv3yjmoMdwKo
l5+ARf1FMsRW+ETAN9e/i3oCThzM0wgoAxdtWtUTMJtnSVRVwyS+N+xZPqcI53Wv
GdAL/N0dVRzR/JS5k3ASWXpv0reJoFWXtLiZRiaqMmR+sr8JxtotmHRbMdjPNmiY
nJWmZq4UJOAIMmv/GJq6dpGJlUt05IQvPo0Csf2RUIusA1+MQEJ5k0zbzlAvWeS2
aZOqHqtbKFgxK/UdTSmhyf2jGjHLsJG0P19qdrHp/tb1lbtGbhHvpxv6okjH4pGS
f0M7upc3LXIES/5Cvg6KdN6Qx2E4sJhNp+NnL0Z6/ebUfMyjoefPQMcVn7y2nnsA
nci7DUgHatkqNcuK+qYetqP2lYWYq9zqcRK6wVHpWcwMkXvoZrkPkvahb1lWsAbX
M7aawQ+TjXx4wMfXjbbZM9BuLO3YIx3TK7gUgrhbXlHqKEsN31chcCWkLu6PVhZm
SwFlG8Xti2ZME6vDFNMpgCbC6KTBsv3/pIWLa2fsouRNK9ihpGwfyhW86EbkCIZd
A8Ndg9LSOHPZVoGKv3l38wWoqSbx/hQjshqtMqTEJb/cO7oPgiS794pQW6bovua7
JeK10OqwwO+rvLbCdCm3Mu0FpZEqz7oObo+R0pVjelyr7xVcjQkfYeZj21uYtCgb
8LOrLlAuwkoEDTJSGcrgbInNx5pDM/iCCW5HM5JOQMpVI0sYZ4JXj5yO2Cv2nUe3
+Y8C8/bed9+SO2+SPWaHnp+hErfnOCgMqoQdV9fcCWE47B919sXhggO1Wj2HXYnt
ugxRGEvywhxtFfpfJYy5szlsIul1mc6qFgUXcVbMRSQydobfKl9LXOgu/zVf40lO
WP7AoptWxRcIvpEmw4BW5uMMp1ssgtV1h2YP7zUuRNn7j9AYTqOTFBjdknbjbd1a
x15KgZiEMZvPRaZDTjvkXBVvRIiEzOpUvRiNQmwzOZ8iruz37HNa7Mjrj4PHGL8+
8lecC6pr4SBAvyUVnfuq1cJgt8LR8oEb5wg0OO/RDjivGjwzlBgEfrJiUJKMos6u
QvO7Y09fc3isArZoyN3zIpvun2LcDRbFWxYkA95THrOfq8s9HjSxcGMKQr+85HXG
xmQgmow9YIkWunb1PPmYLYEPiYrY7AbETJccL8zlvntuYmvYYXBXlmM0E+qFfXnu
6mt61Gy42JeeeGCdjNSuCwUQwRxUZq16LpyQY8LRhwXMqv+RJfxwPRFeXi9bV94A
0alGc3piSyOr7g3EtD3Se3Osvs3ldWu2GXlsCD3kjrsJwsgi1HzbfS7jx46oPbSR
b4VXb++saenjmMK4+P44JHudu0MJZDdFk6DsAoZ3lVeoVJ/s+EmAFUf63iAEH9gM
3FdqHkFfTzN6uTL1Q9j+tyahxzS4A2oti67ClAgkaisVOp7SEWOC6elPxNGZnVRw
LF8EVjFUrpPZ8w31zKJ2KdfJMWBP1oR9JttI+nH01EVzvowAMU4O16HNClgw1rNS
SFelRbKa0th5gL/5dbSGso17aDTlriUsBUUlNDOBqYtak4yDFuq369wDd3Kx+vGo
m7k9+iQhAGPlDNDV4s0TWaWMx5lk7BnLNlyNbUoCy+mukNhwoKzA+0b5WlJbtH4c
6Drr1//eKicBLjm7/E+JRzWBtMlZbzng1eVnjgvks/skG1ZvZmRFzTZgdfE1fXhU
MhkTpP72VmxftTosvnZE6zRlVhDy39LaCM3VGvFPFy9JLZ1CRUn/qjiMf/d/XW60
Dxr79Kp3ELXUugxpksk0QXcnuC++d4k7bDNo4uHy0LkTTW49z4kK2H6Ro1uPUGVT
PkFBH1N/fvuQG6vsW/WUjTZTDC4C5hPHb7dIxu9Ct1O6vnUPxPnKY9mh7lpMSnsk
MIY6Doicg31Vt+RBD3EBsvAGgZgKw+LIeEy5hUruLyVhbh0OY+A8c+saLdDZ7Ops
LHw67dZ3YqAiAqP03Uqj6ZQaCvfXDiLiQ+6NAqLHIbnInr6ONkb4u32wiTrXVJLX
s9SMogNqmsPHoQY9zT682ZFLLa/tsVXR29ediz8fPONxqt5b489w0mX9LzOEuaCD
NfcSSLKphIX8Br2gGgFA8UWxwHZt7ti921/SXam5jcO4SZOVJ4KibMFk0IkBfLZ7
w1gkSDOwlmNwI3eP/3RfwsAw8T5Gd0cZwYT9oewraBo4A4O/2RBYZs6sYECIBRhS
AXn8saeI5Mcv02tD10VXFG9t2mmQXDv6JfycVQf8i06Tj/I45mkLFCv8CInBwlpL
LFnVCMcz7diCqQtVD4876BGyusDzeg7mz+sWFLiD3hWEUnwLgSCD0uNz/g5SB7Mz
am0CALkFxh+05hJpEA0bfAoX4enyyKHf4JymzxUzx/sZLGz9gs2gvePxvghy2okk
pQ5GXjdAgWHprH6eqowFYr1nioLCJEB0UAs8wijykMGkXlv5ZvUvsWqGuBwVako5
wYUirHxP0aDWySy8H0wcZQ5uTqAYaVbCjlmyU7kKYCAjt7g350EnYuZBLKnsjY2V
PmBvuNsBJs44CbRHxDu4Mn0oAomM7OOiQ0vkFdkK6kM64mGSsbDdwCHtUm0F6HM/
OY9+biLvfL1gJtroLBQgxVZQCunh2/5ct8RUUwXv5Ep2HbAc+4f3MDyRIZxdQj4J
DPQ+p62SqQeqrE3s+zZ5SjEgE1NgWNQQMhJGZoYnCOaJUa3Sn9bK6K/jUi1RgJm1
pOErEpfD/VH70Voo7SK/uvhHmeVFpWT8aTxcrcY1jTjvq6/DuJ8vFqHoai1m41sY
0GCT+Ndb//BEf4m83SJC6MabIYjpNiAvJ1Qi1CHywqvUM8KfCTslSQ0ZcrsN8kE0
yk0cz5NknIrGmZtujexPY2SV8lVTf9bzfTH6EffuXX/A+YlAZ4+XZy/ujShkCPAN
TjHogIpr1Ux4odfhbAbO3MabjpeKh4MniCxMxNHFYEGsEE0AT58cGUAnUuT82BFA
bEvObTDvLwmGLm4mGR9Px8wXtNXF2vxA8Y1LJPoI83r89MA0XDjKzEgO//i2apSa
kDJWZ1od5im6XMVRHb1Y3LWyXXG4wUdQ75NhYw2L0iXnPsrWWt8PIjazTLcHalhe
5BtYV9xJslQM4zOwAS4nIvkXxxuYlEPjlMU4zwHYxnoJbHu5yEqng47AvzYnvZw8
n9NjAKsqrMM623SV2v92ViAfbP4a/v4rAmcghtuLyiUTXGFulJA8SfA9o87M2Jj5
QvPVBJaGqcCBqSoSoT61zLSWhWICkKZ51bflshKc3dl8KsDMEc3UVjL+1Qhva0aU
egqH+F2q49ZgfZuMH7qH/wd+N0VlsUmvB21lA+RITGHkeWIyUzqruOUT8w1qUKvS
dUtZCRSjcIcyCbf7JL/HHPAW6MEFCZbN3Cy665DuEmE84Hvw/7/4qe1hiWj7C9qw
etzS4LA5M0EnBeBesOKewqIW7OQuzdPRSwE/RqMZMnvNYZ7FmX+S3xb6cAzVKiWr
/WyXTUpEUsa61aEhGUozg9AO1XWcrmV0q4YE5+gWYj5RaFy7xWspjiNr2BLBbwy3
PL1BoqX2h3LifVL6z0u0QPhTHj2PCri8Dr7JNqwDT/VPMep85CK8KT2fUmgw/o0v
vfZJmGulijIOuaU6Vx41Mh2zTK16tYa+XAhrvezC6ozMCpOIDzdRbZqkJ7qRZieK
Wd/Aj9WmZ4Sm2stVLgPCx4zho+SqA7WryJ0HI42KzUQBiF8xXobhYQknijDTJ+VO
nW0tiAhFncTOmhM8BLKGiPCQvJ7HDMcMHtuobBwHXGob6983ItGWeXPCZfHvbVUh
maNHzX3lBLES85rRpA77Su8lM8+EzemeckRkM0jqv7l8t8+exblveOMMMQ9P3+Q6
Obqx7OXjcGbcKGz98HaRmGivnf4+ef0ENk3p3N7+P9IhTHvJuBNMgXfRcTotzAQC
su3n56flmAOO1TwwekGJUy0bGRdZqGTAENOEY44yjjW/XHq2jFdEKaC7xqo0m30R
4IYTCMGHqKpnu8PjIQBL134JM9VVSNW6LXufgjyeoFzPgK5PvZxFhgDXjNzVuAX2
P6P1/7neZdoUmxz45eEZ3f1FIwB/WX4YzVYMglfvEu9uTr6+c9TEIkKvzeu1sYsq
Cu0px/uXsx5geL+Li+tKJtCiZd4zbGQC36SSFKEswJaLY3iWt4ObAcI/h2px3S+o
c7PX51mcjWikgWRzgNZ7poPN8x0urjBH9H5mFlYHpw5b1qJ25OCy1uFHNhad8+1N
5cMQSt7GGWkePL9MmqXTVkhP6LBvggaHfRV1e9nsNFGUs0L9SDFPqc2QFE/tbARt
+OcpoNBmAEjdDg5a6A0rxmHAVKbHc2gK3F3owb5GvmkOxeHrC2a/xmsMIoQZAOvy
xrHR0GlxG/4muJ/Cl86U8SnGO8y5SGCa6SsE70IpHHo2Bq0zVaeUKb66NVGy0gqn
CDmNywPtw6b627kEULs/3+TlzDbIvxXRC0xL4Bevxj2nMKFpdbRzRbQ83AOiDUeB
0JJxTN11Wh8A1mUkgT/QsNOvMO39XIbygslRpN+GNn5l9JoOhBtL5sWAAMZZYxwH
LUET3np1rX7QlpdrxWPmNWp8sp4t1WOxADmFcjePIuGNmnbDvqF3B67tpPSLDd69
L50Upx6ayn8KYoP3xCqFSKasB0twdowdwoTmu+iljKarLLyqOt3GikNOr2DCOEIE
k6kSTMAr0En/PYjEgCIWunp1HWeLo/bdfTb8HMbIVihA6xIiPD7F3bUTRqbbKeyJ
YOs/musXBVz57jjZJRxz9maZWYQ1WIeKCy7KgWQmognEnWilEFc9j4YgcEpZyz7p
xoOF7CRHPfFPRwYuV8JLtDfB/h1iwrFFmK4LGp4n1NePCeemYFod4pqfJA7IzCw7
MqxkILTNQoWpHxI1ylq0ZuJVCU08sZeFydY5jWm3mtG49ecBgKjHt0anCwNhGGyG
IqxNkFEyH43LsOTnhiCxKpDr8bKw17PmB2avTOWxpLE+awVcHngVP785AV+BmvjR
kJHwiQWU/vuLtWtfXi51bzL4KsIo6WOM9kK04yPnApLzpktb3eiRph2BqPZ2ga9o
2Okk30YXm4LEv0LQXttoineI2kXqJs87LA9cE1DZZHd8AOMrCwmaBksZTj+JZ+Tk
PTqlpvKwK0RcrUV/7dJF4pIMajwp7s9CS1N/PFhNO9zdm+MwqGIuc1i6hT/DA/WW
dhtmpHrddbJcfiF7TPrHMirJeS4odswuhn7xbq7FmeIq2EbDpLaCV0LJ0No0Zr1z
ftxygVWKHSg5BsT3jJTSW+JvxuWK7m/tfwTSt7qbciz3a0NKR4aq8lnOgbVROnxt
Dwi199ALelKYO/QIsiPrU9VLZ9TmFIIQNOSkRcCSV0T+p37b2X5VrfbrgyzEvtEx
LZMmZYX7Ih2FrkrTe48lfQHUww8XwQWJS3qb/OQDN/abw8fzV3v6hOC7r9T0MPmx
CZdCdLg/jNXGX5oK65eWbcylZL2ep5LNW42kUmt79bIsW977NUOxInBn2vblZTNr
BA2HWIYVZ56eskeE1hyezieRmYX9HQ2bbm/KQwxPgjKSziu2g2VSOqxkgKoZ74hm
HkmoC92YW0XlLUmBcBS4f55FoLznNy6YFok/xmtV/YierRkk1iUUWPzWmVFeZw0T
ND1lsjG7YtYygi423GphLI2fSIXhoFSjf16cXjpDmewQh1a4QMNxCFO9Z5ESEmr7
GLpGeF1hlJWurCsP2lOiEQTnklrW/40sKmyc2Q95hT8df+e58JjhX96JUIBK34wm
k7QvwUEQm3/v2UYKptO+LJKBla7fla4pw7XDMHGN5hV2dSEpvy5DU4Be+jltGEec
B5YZ5+i/Vxb/zRxGHxxmozr6lo7mui93n9668O4tjRR/LNXU29L3e3DxstFEf9hc
U8H3h8X5fvaU+1dDjrOguFgrrK/SLIcGtm0jsOZ6r3qOujtRPrPmsonxQqGGhfLv
qH20upnPbE9372MeZyedVOuWWplgjW9ZmpL4YjehkOjFpC7X/zdc7qQkSP/1whK3
zUs3yZMwkk+sO7VGFBXl12Uo3cFNbWl9+Z1jxx197l4fBprZjB7wEgPHGVb9EP5Q
N7u3KbJGnCETgedinddm42ge+C3FrKQVML2DtCVR6RTZ6HUjGOjuw6wQH7r2ho3g
nu50vlTTqGIm1h2VKERxTPuj/GjLdlWWf/3cbG7U7lMTK+tPfw1M1FfWQdyS1htk
fSxtgBRM/Gmfp/ELL7cjlt6KpVEfDoseg7APdMeOWRJQAHPtm1AJdPpRby6+r52e
wpeINi/nkz0p0P3T87RQ/NQNAL4ZxQB0Rhudt54TUsEJkxM17wuYl5T3RWCfMnuf
uD9HAf4+Wkd2D0qIfhildCef7ZrlCobq9eIRCj1paIC2h75VZRJPp3kEacJOmVZc
1qzLxJUGXeiYSfO0gP1Y9M5EEaqWIZ9Nq4my4v9wacrQxnpu09DwmlGKYD/6DD0f
JSKQITbGZqCy2lGuHMMx2leL1nFeZM5YhGVZ1pcLHcwAoWOJu85sDX8vOotEY+tD
P4eAb5DHBG5fpRh15ZPyXwPmZLMBwdUiKQGHDbkNaLFFNVowUZ+sGbYqHJvjudes
EAdxPngPt59SxVuG0pD5/UDhLFCjMK9+nvb7uO7xXgieqF95WWthpI01ZLW0BUDi
V5x9DFGg/a5Z+tvdmBFZHzOe2m+ZKI5ufact01Ry0RTX3SuiX05lu3c3vvCNar7t
gc5dcqWkIFa8FIrv4bHnszHRQLIo2KkRV+xB/DxnIWc/K58Qm0S7s7L5wsfyZXxF
/ljOtJjJ8hKq6m05U9LRTTRu2SLZth72sdJYcsd2BcM3OMbQraqtRTMhBHfZvDW5
Nx7YCiqncGRmrFGHfNvQ2iwMv8WjH1SF83T5l4/15ebwBSFQDTnoJ+ogRMb0lZJx
rKfQewwlD1AKTZbB1zdjFAL/v9M6wDobC7g2LssRpDBO9+ASQoq6LWDwahs2b7G+
/G1/yY0qbiFh8uX/5hVgVgCUtXe0ZZtkkkJ/uOc0HwI990DFk4kWqIrpBYqGvkLX
x3a6QIdf27jGIgasyLXFWKTO7CURey/g1pN+62K/Evem+l/woSqk6EHD8+J2lcXT
YaxGb2GQWGDul5lu3d2lYOGV7s7dkrub2ewbbpLMmTAfd9FpVcTr9jIiyKvMLUHQ
eCzb8C7I0CaQsJWr/qnHCIiDFhbV0t+rrKNuBzPl32/JMrIqCa82iMlm7bQmULzB
rH9aWXJZBuGPEuqfCBU4CuAtP+foV17IbagT0dNoTjlfAwNN6VxShGc98yVW148v
`protect end_protected
