-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
IRizdhGd+LB/xNA3Fs+Ks8yTw3IccG7XWwUqy3BomqKyrx9WACwL/0uWJbsrCy2r
L1mVgwbApCmSMQPuxVbsYuRFNLWTZdwB4g8W0oNg8soiYVtEimQX7rQYTXWTznHo
E9U38gOD9lQt5VRg/M+MidFyCnmfF+fe1UHUWY0IrPs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 52288)
`protect data_block
TAz6UtUO4Cs9R3XvMQyzKak4c7VFCZGlLDst9jwKcpx2wPsAAff22Fn/GJn+PBfE
8Yv1UohqfITfQTNr/NWYJeLftPzI+66JUh0Eyiky4Pz4EtNvRzcU7LC4tuol9duD
Nq6UVhTfX4QPVywvbS2gvuYAZp9/kUJiNiL3EwbikfypRZ5EPbR6zygv2fHMWKLM
uZTWylvwxHmr8w3Og2sm4fZ499CMJC8/yUJ+kyrbzf5WcWXV/ZstTpSwSh7ynbbd
fEzT/k7iIe0KoYraz4+9dN+TNARW6aIV+wTqiRbIkGqy/Ao6X1hScwS5FVmQZQIe
/J5MoVCNJVfxQLBGSK/XOZMpfuKE9x11sfqv0zCILo6/rfNYH3NYUGKEOw6Ck9wb
y3FzqhJxr5TtW4ydsVKUWlo/VXN0q7pylC2hNzfWTlsDx+VnD9h7RlE9KqKsc8TU
Xawbzbe4Sad9WZo51pJa1nRwRXa6pJhEB49RWCGccEPkfxlbzMkz6jraBBklLkDs
3wWlhu8PEAG9Csuj10dAb3WqVpFDtWaB2ljcTRYtKB/pYxhd+PegtP3BwMCt1V84
JwNoFbJNswGTNwksuKM5Oai4pGM3kIxsId0FBBJyduVK+9yceBnju5QCXnV7k3S0
N2KQc+VSAYWxiEEmdpBVtbRXEF/C2DEJA+66gau600Z4/O7Zh9gWdYqVmjJi6Sdu
bmRrdrwdZuetG/ixgEZcupZrgNUDzxkmv87hgA+7fALp1JpOi3Y7kJTweV5tUzfT
ih3ZMO83HV6umD7kJpCF3EgLNb1fDzOErT3+FmHip7gNNViGx0N5DMvR7p9EojqY
Rtnfqh7wP/jxIKXIBfwEWO7+TTOX8l4dMDA3zbUubMO+kXl9IEsnoYokcOabBU1z
2MgQBDdLk6k4ZtOwyXWzU6nWH983tqoCjYzVNk7ReivR/kitfAEknowaBjlLfAP6
kD/PdU9s5h0SOgu6mkHKluumrHmhpOWDhbDu3cQA6IgouxjSASMGr7UAwIeMBMX0
r2+LIw0XIxPfGXfzB8uRLcbhGlHO3Y8XqKksPu9bXC1hpUp9Zkdf9U5AuxXjToKl
9ootf9GlioVKk5uOgfBcyD+XMCi8qPd+f7Q+qHdh3G8QA7UI/kPa0IlanC+y4kuz
8pePRsUNF69wkhD3ohSK9B8xN7sH4ghN80tLC7g/cyNgTO6OPGqDa/vlYgEMCZrP
S3i+zdnS+AauxGdABwf4P+dgWNRMwYlkVIqCvHggW1q++Er+SJLB5V036Lp6Aowr
k86L3xnF/W28Gb778HVkv4fDNBd6sYKiT8MTeZ/wmdMJx0t3cSi3rpy6LHFbu2o2
8zuYqC21NlNysnrkm68TA1xZQvx+1f8nWAAa8vIblyjF5/TnbTGqW/2XdFqSAuvQ
vaVhCIbVNnPG7yc44+7hLjHDj6WQAGg/DJ/Rzz5WZ5sgo0l71AWG92g2Zysyeg1V
SzQFPo6TG4ZzGiRz89aNYdkT9I6J19TrOk3vd6MRc5Z3hYLT35MWcFFOk0kHOF+b
BdgA5rQ/WgnTC197y/6KwaSDKPBdsg1j5ppZmJyhSwZOgrUw69dYcWzrhyeDft8w
vcX9asAFWPaWwoGUBYQ8no7HyNQKE9sGUveCuVEjDYPCxvZ5R34yQBLdCfqfCYiQ
yWKWqqE3kBZcYK2PoQi0TQEmRB0h9aIr9vcfOn6PIhfZBJS+qWDDk2ROOWhZp5uO
jjvtYD0k+RvBoM4Jxy0SdGB63dnwCkgk7JliH2XHkEzmMAdgGEYVYW34srbHFlsQ
omrBma9VKeq0DrzZIIkx+MTIfVG4eLYSaozcK571gAHVPaadQatxwccOT6Ks5eGT
RlHXDb29Ow+uHZsTJpBbfoUau/NSsg3nWZp240WsJ2cE7Ru63+00PwTUuz9CUW16
OvOzbEjAoUae+1/hr2erLc9NW7+PNZivCNsXsB+AOLd5bgo7QMuNBB+XkocDEPFC
hCSgOfSBxJJypuD4fwMj/WZB3uzsIsFPgAaWd8AJ0mZmvnWowLyvwXq8kcfOZvLE
WZw+wJb+sltB3h+35PLXzh8OM1xUQzxlpDI7rSeNFrmtme4g5XE3HRdIt086OMnt
6FbXURNEC6XkCizL+VXII5AzKakt30O2JSExmswImwzX2fxeovOesAsh+QL5edah
snr6tNCwd6NJp5UIxtiQGNz0+wax6cvQbfp4c3YMl8T6iaO0sU06D57YAl6NV7hA
ZTHBp/iRVwXa9MGHomfWnRph7OZUKc0fARuhEFDyZ0nujOWj/h7d/hxZyXyYlXPu
hZpnpeJtABbVlIH5+tjC+IL9HyawXwbSoyuLm1pfPGGWLOF7wFs3a2rc0oUon1lu
rKRrUdW04X5t2uev5e3GINvfTidKbat+CtkCdSap41VnK/97REJqlRVNwcJNg2cC
+aDaomCuuvz6uDV3nYkslHce/GZW0u2Q1lxT5fZ0LOS45OH2U3J214nvvmHgKwY4
nhQqURPw7KV47EaRo+W1zniOSO5qr40x+fD74XgSDTKoZT5ktObsniACEkgEKedF
no5flbY8n5eZpQi5T8q6uD1NAW3zJJtkwJ4JJU/vZDRmYSqNZ4dYeVE2GdkjKfdo
m57MK7gTlUy3riCDdvTdjHL0M9cdH7bKHqsPgdmxYPDzofEcBfFMXamtzu0Sy7uO
HgDJKwZARKCL23MLQl0gdgUYxtTI4+s6ZBpGMLxTUCtNAhC+GMIO4x47a7vS4bpG
VnOPWvkOdgs8k0o/i5ysWV52A6hOaREwGkgtpdZvOUfPvvDhlWEoqp4mfua09stQ
6RWu6GC1ukBqEJiD0u2QfOJjGAphXcbCBoTJQGlexNa3q6Pf9v4+OKDdo3SPQL4n
yo/s0BXV1ftm92HpNr84yuCZLIBZlXLqYXENyPT2XXVkV0EeN1iNVQ6zQOXUMTn5
VjlqqJoVP3HyGmFiq3nf1utnSsIMKMlK6Q2ovXDq97dGsbCAh0f+aYJNpfaCNuFs
VN4rbR+7Lh0OppKmM5XeV6duQs4Ou7oj1XQ33QjEFrKMy4at480jI8GLNfzJuq90
Tf2Jy1mkIZXCci/683mnrfomIVwbvoK3BKdjvKHpwMgwDXWH5yW5uhBBXQRFHvDy
R/n6O8hE3NhbaYNf22Dn9JGSwjXSNgchGJZ0KF8P+uI8/0Gz8PWPnVnmGHXfOSuD
WMAvAqIzlrMtN8D0up1+5Q/BNgqEEiyw7ua/klipXM8dBOVFVXIScPiLxg4q/miz
Z+gqNg+NKZh4ZhMK4sWPduWkG6hwka4di8Sw3OtSu/Kl7+uRT5EMw1U9l84dNSW/
rlUAC02MeaSYWfjbJZBNIwxFVFSEr1Fr+Mb1osr+Fgw2uHE9cCuNCrgNvp51TPLU
g7jdOQ3On8IAfIV3PrDXHIbp5rwYajSwF8GKYn/j7FIy4Zh8FC3J66IsXHHoJmHp
hIIG2PzVZpoQiB/OH1h/2zPpu2D4pn+f2WyvbeP4bzHjY3HWLFdfso3fbQuYJyhL
RQTtyWhx9jFlZa9xZ2lWv0tvndVH3nKBtchBo8mJzKxxlC7KLFA5f/+Fhyl2iauX
ns2PASJu95iQ3nU6fdDsG45m6Q+y+pb7IfKXWGy5MuSD2SArRHOKV4vtROxX4Tnk
YeidoLLfNjP+9QvWBusqJyQrJXUeONvv9DEbqRjZVDleGClIPjc2DV/gdjsmrwQy
BtGf6Da8U5MDXdQo34NPKCOG79+Pk2zGrzd2WbahBgTU43VcnUSfvEnCERCtW4kk
+EnzFkX9Jr+lIT7vidEF9Ar5MbBy0XPg5h88amQD3ijxBlyedzFp7R51e9jTaMbk
1C3uXlrRtFi53bF1faBYFQcTeEpn902YGIf88pz4DZ3GT+eGFdSwl5nVxAKxLhcm
83MRRTULiHUzp3QYvq/qw8/gVzbCxORjNWJe4oXsgw9NiWoLZmy7yGk3A9Z6M0G1
g1Yvc6mV58AQ7NyDF9j7/5GPQgE+Ydw2y/fMKWxsdUveEWG6BhAIqTM+yBVBFLeN
dWS1PNrXA39XRg6+B+Rx7ycI9N2NN3soUPMXTU1lKMkgqLVE3jJEE4EqJ2UkFJSP
DdbSt4H2j5nUQ8bA9l5sxJCvPgPKwKcJ7LQbRf85lJ1Q+qit3LjJha/bMlnctNLw
xNUuj25E/LC+yfXaTYC78LSmik+tO1rZ8E640HBDo75awFOAOvOo3dhZN2hoND/+
f0QI2O3IkO9YLiJrEiqya+j+Pku5JrhfejkVkNhzrBy2jhhttpDkfltfcCIMkA2+
MRfaGWo4RDREuTBE4drmZ6VCPH3Mc2DNpjc2MauBjo+qiYMUNsEhIAD8VpkT/XUw
l1yMfEG4AoHGsU76yKqgTfa4oFLT72y8aS17DVUU+HzZQEnfPw/5h4tf49Ai7r1+
ZX/APYwvQ/nBqZnHNAGsNXcapiAwofDOxSQQZRJA5/IAWPoHPo4JZihlewqEw1lD
rysj1+yPUmGmLSWYG+eCXIaVEfxPOfCndDocW9CSAUXQoF/NC+CqO+B/PyqK4izy
uvt1ygyB43MALMQqEyQYvjliKimTXttrlB+wi4QLE0y+czwTcZzOq4PcMknOvIvG
I92xUVRyHqH5PAlP9Lgt+UWMNft5HCajLaCezlBQBgcdMp/ceJVhoMFzZikv2DC8
jJHBPINpABdZ1uHiPym8GwIWPMWtCwFolfX5rOvbm9jvRYZwzJ0oGWbJNpBPcvZl
uvy3EhQoIptgmDiYilEmjsUBQHGLqcfsxhbOjIBTUpDtt2bXHR/YMF027C0uhH17
QgjpqSI8dVmTvA2RiPXphX9aTankqZKoG5fs1Vi+P0f8GdDVQc0f46UW/6Q66g3i
GvN1bCREk4M7+MFbMDOSd2yKAr91pRUJQXcqeaFd1FDN7AWm879fxi03xMwh9g2t
eySe5+RRaz/WLzcdFusHqOn9bXB8nMUHMnAaDzBX9QCL2VHj3X2wDsyB6bmx95JT
4MjA4AV6miu3nJIXWpM40yfVfDa+qI7JqeAKqdQ/67dFp83+RwpU4wK09SLPK4om
mgttVWKNoQQgV9hLQPxsjEy7lLLoopbMhHyE1iiUHbYX58GZNyLo8XnEan0LuoTq
Ca9m7UsW4Bu2x3l++eRTgCX9ou2Yq7mkZ8g7k/FK/7ZYBz7qaJUiW1sFHzw5kCM0
He6cxLkNG/mW/m0OyNSsttHUX2N33GWsUn+/btg+jf07TqfQS0sMZsyCzqygPLM5
SRs6NwJz/SaG5JKP+faPkg+jpLoPWTnBlTmAixDbkEeGf8qgzn2w6EZE9YiJVa2B
MAurzZ83K6cn87Q1l3eyn/xfHDixI+pJmSPHBI7rmeoWgW0MdgQYxzvCZcM+yKCg
zjKN2PdQcge0xmpnNzuV+pb0O+h7oTVZNrw/PAxPbt9dCMujgdECIsEpMg4bYpr3
4laE/RHY8J/fHQklOk2t0C5/HDEEQqNC0xLTYI0fuMeXFqjYIUtMMtjtum5tuJ6n
9jtyaOH7s+2tKni0QzO2dBrEfpbi26G/gF+kfC4mezuNpCQNvnI3VbVlNpfreYMv
zS4SUTl+Y/dnfz9lkZhAZ8RmIrmkTDphZgsube1i120Cllf+U3ntG3ARjYfDofG3
NeHtZtWgHSJCHlZ4aFTMUXvxJ8AJOBBYBY2pGc/Uf8DdnxeM9bVFCcXb7wJVH9yJ
/WsQgpGMWEfBvFU/yZPmSCFnwpcKPHC5pWxhQ9u0NDX60LyuzRdfnSiE26XwF8Nb
h51q02d5wNrO0QLH2VSE/eJelUO9tR9+vGhFFiyUIzgcd7aZQotSuIiXJcr3rfLG
+tTWVP2YRuCyzA5y7Mblkza2W/Hh75I3d6utxiLfQqdlBLlbwk4rR+WH0bO6l5gf
jK/M4Knh2OpI7Igvq/ntNLY0aT+PkurLocrL0XmBW1yb3Nrqx/BVHR+Hj2eW7OZZ
jmo0dYNysvtTnysVi/2AYUEFb53A/HYz33vCqAPnJA/8Cv+gEaaTpN6cNPrUKyru
nJzal0nmaneb2RrKvVquY8XNBkb7AEPE8AaJ056nj+Fn18IsByTmjioT1UBRFTEp
EbJA0Y5aU+hKI+AgYaFcEYm2lsnq8S8tKl+bYUgbhK1Cwct09Q6Kiw4Nlhzu1MZy
RgRuUZPnkamsCg58mdiic/HDpfP5huvSuFxguqBClfY/trH2k7e/ftwbFzmqj0Mp
YTHvfp+TW2b/fCZu/CvP8LDPviMGzzoww3BnwNTB06RW+e4OO0NVNReTkSuSv/t2
heeaHfZhj3uECHgsiymcZ7elEruMRM77I7qf14nsL587zulIhNslwwZcWWwPG5OL
DPb7JlBBj0VCJQ71wJbJ9we/jLiL6kQ92Ae4Dcea8Zjf3wEL9liDcyUQr9MpYJvr
zoQ+XNhT17KXiA9IjnjnhYdWWvLjflJ2B/obsOE2+/gKHvjjdyR10+OLDiSfCDQP
7ZYXabTWnrqXjlsHfTcTKGva47SGder6WTqPlZx53hSLaLPVrOwwPmhCRo5xoMKj
13dyZYkRfNDosEC9VwZ5rWpJxjkgcWVIXjHjxKlULCHzguJux/PprJ2y+cFlLssQ
JZVir/g75VSLK/4CAfINzkVoUFfti1uReYhCq2mDjb+vB+jMlTCAhCnqVWg0Uosy
oS1b6QjKWTV1QH0W7e9fmU6+210FhEvA6XPddvc/ungPSzhjKGaueKjVtPYTzUXm
5gOIHy4l0gy152YMOUvEmMfKQ6huywDh0S/vp6wRgWlqUqFHCTGWQFT+qKsVI5La
HusiRwgh9pCqADvKvSpzyG7WwlZmcCdlodIiMqV7Ej2icL1zfci2cNaoSLeMKjmj
xtHfRZR2HyV4M8XVM7XHhJtSB7JdQjSk2wj7McahZu6Fj1n4Y8nROffqUBsW+U5x
ornKxlxkoT3nFRAWRjNCISZi/OSyg3NUhqDpJkkfOYoKOqeF+dZUQI8unyMwpkRt
2N5o601wCVxuaA8uEGOENZ2xrLoUT5DRdIZasFrwH8upzDg9komAxBdX80WmT2kD
yr8o4/rzCVNKOFTYznp5Rlk0nbdvh6bkHP7IOUFgbq1B+BfgUbqL6jSFTQUKmhiX
0j8P1Oz958X6DpgBq/XCrZHLXoblGth6VdObiRgAUnZDsV9b4RrooJCU25sHaWz5
HHBdPfeIzJBIqH1Xj3EwiVHYT2iowoerYoySGHdGT3msJWQQnKsZmEJuPvLJKGcR
p4yDnM5NaWKfKt6XGmOj+qjj/0TQ1VOhHeeZIT6GajzAd1qOEevrgNXtzSX/Pml2
H9H8sqIxVEqZsYCwrDfHMHf111J090p2Gb2bHX5HuY6dNnA2MNHAlvvCD480Svti
NTjKZjNEsNCoL/HjpAeYS6+R/uDSJdKQKSG1lzD6Yz2IgDMiauYCmMCCcbdWYuJK
fw8osrqUfwsD0SXke9GGeyMPQZjWhKi38JC//myz6i4T/bbBw5YXg4l4Jh2akIv3
P4UPqMaorQkO1S172XfKK2we+x+XDkbnoz9ILXW+2K6VrO8Gy5lVwbikDzPDWS4F
78zh/hl7Ra0qdp0s9+i3FgB/uXKo9lA7DF4uzoH+se5KkLWZhbqnvw+yqmJPLwpr
UTK8en1BXYHPFntgeBkpIvGlPuKAlBl7DiQ4GzzxKn1ymUo0acKUUdHW32LhWnyG
mh5EPJsjUHoU5MbiCKcKDRHsEOe6Ddc2/nscM5Jck/e74cA/HN8MtsdRnkSBFb9i
LTm4Wk8pjyGIz0uFCB5dhAUvq4yTifWonJaNbg7znXQR4frOZgujDvXNsqBxxdqf
FxSRe19TU/TV1D1fooTBkQowKfyaFNUCZ7YEdWX6RJ0MMA6dC6Kir6WJK3aVgYj4
jshkxsrK1LDad+qgxaDDYFtrxWSn1ae4ehrfP7FUr3WFiVLRPDBjjL2enCv2LME2
VDd1WIoVbxr20/DDQ1Q03fnw0FCRk1HYD86o1hymfeaqpT9Qlflg5H+Cysvw/GDW
7rMzfiMrLbTeq1KwNY6vdYDnAp2rFwBn4xfSnMI9OcDPI8urjv3VumCFKXPpVVXn
MyHoWRsXWLFYWKypOXJWvteUePGWoYrrexHwPt/bcZ2J5yknqT2X7sBrHfvk5k+9
eavtq4/w9IzVuk8YlyCljK4KclLt/oTCXmJOXN7gcQl21zVWEOsvcVuAT/tqP0ig
bGS3fL+kbb4nINNJ5COWdbGz+ria2s0I283Bbl2jNNL3BwqUWelhG0v+D7vg0miZ
JG2tVY6KdHKh5I5qARohJt3ybmsahZWfOfFhxn08Eg5bZ5o5PNkGGMHxqO3E8oqj
tVn41cuDUA44Upzmqi7hM83JhoxA/FPWTa1xi9Luk+i6AJAyfYkfJ0/EVizUS/mA
VlKhqBd1gEX0WAAZ80PniMPKPjNo14+S26Fve/6Rx2+ZoqM8kMkvIhXMDsoPLuUl
he5xo0MvQYKWbIOwFvglDcfnri276ehV0TXkYDfPzbayCOgNqUHSrcV4N4yv86ri
TjZFdNgakfNJKUgTEpLXmM4A5Wck9wuwqOCqEpvweNBT+3X83solRT9GU3FwEq42
Hp3InJVcVtKCn2kTsVCLRJAEebw7LDFrRq/zAHXijJwbnWLQKpeDnRNyD8+G8X3Y
R10ZmCjwMry2XJ1drAZnrjFNokZvcstcpKO8nzgU7Ue/KtQJhfaCAr0y9tcJqrvs
JMZNJ/VxuuLwY5DMdj91QD9oxvYCVUZdW59c3vg7u7GPnPecsTKTkh+6zhWC1ly+
nEN2ms5alVGGAndaqlmHrAm+gHSUdstMIBtzwTsTUd5OGwd0jFd9PPSBkyL0mBlm
xUm7Q23Qk1Hrph21PZ2AmYTHQ1ii7swjfa+H5xXKNKGN68kjRu3fDhupcEU/CQgL
SKxydxZsfV7IZBIhw4KAdcwrPz0/lLzFsAC5RSGh1S++YecorZLa5TO/pDX9LHmS
kY3f5FMuyuCOvuiz2+JEDcZDLWNjIF2zLUayBP6dSahHg2EGqXlW5mxXYlqaN8Kb
W74lzrfvfP3rTYmSMwZgU4LsGpmVyngwRei5PVmP7vjT0fIbPojTV9XxjGmYj6oy
Cb9yBH1Y9MXF0cYd5H/BxPXpaGrhlYNux5n4b1hth0pRkoxGeFiQix8eAdtmes4x
1Bg8ILLtGM2sVLoLOHfcNldjve2JxrFZajILppleNQUrhe7+6lHVlTyoGRKWJO3x
BhlDx3OuhVfIDeZajn0a1p81/5YJZqDCmDggykdPG9hTbQDm2kIXcHNmmmdEPh04
V8e8LtkfhPoaDgEK6yvdnK6/b6W/AP8SXzFgbJuwcfuFc5VYdP8UtfCzSdxDal2g
JDA7P4iO5oT0FUM3WEVuD+KW6uX4LvS1hKKoxReGihcK+qDjBqIp3yCeD48i0ia2
g09kegPo95HZNl1/qWm7ROzmYMuSfdtMraCaONlBiqHAo8z256+6nAebaGXzzkFS
v04tHA/u8ID1DFYHyGKebob7qjJyUxRKIWXK1HCmozPfI8jjp4FTuohxjUrDEhd4
DJ0knIngx76gl0TbTlAEB8GZeE7/2GQRhj1Wnfxv43IwRlhetPrmEh2q4JOMZz27
mGG189WQmceclZl+cwjAjwB1P8LcFui9QHSPNSZiauNQ5GoQz+Wfs6PFwyXz0Gp4
wIKfhdqfupgjGseN1GugdQuezKHBKrgc/49DqtySlZAhXYgzpmnAiNbhf9QM92GP
hveKNfiWyens8EsYqFEe2pMTnV54V12KCqE5nkYjw+zPWsHu38G/DtuR+u0CtKlF
yLc3fvZDcktB8+WRftLLws3ZVvTLZPQft3mjZhfHXAIQHIbFu4d2cEzT153378ui
3nbcq/gruWbmMheqpDVsOitsS+jkWyKXkX+8HeDh5av/GfPX0yppon6k6DQUQlAp
1B9qC7z/MlQ2wd46axbPw5XNDwXNVsz7GpSbSX9TQPzpIkPBQyvYQDCQJ/ugJmtW
cQmEuKWp8sl3GZ7DRzGRb+995CUseOp5M7Z/L7wxQt4cZ+i0+qbJDJ/HI8CzOGL7
+JeR4NaU2EG1rVPZaE8zBRmvfEpUg/w1H6eYexGDawIFVkIPzuPtIeaqP7m8Gi+i
ykxRRWSO9yX0ptjHV0X83AugyuruQaG7mOK+IizLZRkNFah3xbQ+0KarFyuiT9Fc
O4jK4oxETRiZ4bwVLbOEEMgYkAaHYq1ZY423oGGiYEDFDMpJNwFhLm4BcVGlUWB/
3bY6BKm3Qj/3FWYMK/JRzJ6wcWC4Sd4Z7/oc6357tL2r8zkk2Kubb5TnrothZO89
VMl4I19jm9czJVCHZK4jhwJLx/MWv7PixeYBay8YTqpks9HEFg6R1QiDLdOv/yu/
8aN96r5I88A7wZLu2ci+F7QVGEtOZJZHV6Fq2sV41xRPE/Jexj9G9i5UKIQEnno7
s1hTDwfAAsJoLeo3ppAaPkIN+cHPZuc5SvZXlM25iRs1bWuluE2+uLOOgDNcaI4a
zS5ckAbZCMzEpttv7zCPSdH5CPGgPcMsI9ZoFmhS58Q05i1N7PhzQS+WfpDjUNfM
p1UqTkGnvmjDaZ2PuH6k0Xi0XLcTEU4Xi4qObALo0nkSEvGFSJvjp8VVUq2/EMIH
uXGlTz1tEIgWW1B8G41xLJEsZ3zQo6kLhTdNojifoYg3AXT2VrZdIULgon1xkUoV
9Whul0z5p6S9r0aHtO7n5MvbVI0OMttqB6wzC0HgRBGGPVCoySyujtdVHnupdjfs
m2aCq2iCAOg7yS8DwZQkX4yE3PZaLxMm3aKp4RSZWwybKSCO50icqoTDOaAEcHYA
pBiUl2Jge1buDWYuQtK/pFvLeWJvxjuA1Fl6H/Q7gVuy4Z/CCua7ieeOdarb8uJ5
veoupalPZiRYCIlwYjeaUGAB655jq2UxVueKNmeBBYABryDahLLucdOvD2+bpEju
1QS4WjJ27GZ++y9lwwitvVogjLUt/mKXzje0iNHgbcczDWfRRiUEovu7ldfRCJgu
z1FMwQByum3nH1WGr7/kU7yngYjhj2on4c2nmXI8l97ahz+u+svoJSi9pbxgm+Zw
C17K8YunvWyD2FK7FhxNOoUYdXd6Zu2anhweeWsbVNO+UptoHaNdFFpiNQ+izSeZ
zgZEAvbXQ1c/GagX3tgXj82ryi0JEWyppN+I1tgXQY0jfn/05R3LLaqJHe5MiKGA
MsGcQEIAdeme1W+RTEymR+znCxVeaF7H5MlTnSVtwqSCP7KHwCuInSZRm1SWkobY
DtWx+GdhDFJTfPg2jQVMfRAovQwPK8hZnHy2e+tcOimImVdXFLNE6q8rjdEZQnqE
TL19eXnHmKDJIl+1rNnVBFKFmi8BOIQ+Ch5ASUJ5EKLwZiNUEFtKucmDyk2OPrS+
dnDkU+ltnA1y5MobuI8h8DUi8bVWXR+iVSYVWF9CxcGBeu9ywcNY4EDZdwJaX5bE
UA8s64j5h5OSRU9SCnMMXmZ3C+aBXCkwuDhjOpjwGBplXrXAVByyYIvikQtNzMPY
v7B0IuYWqzoS2xAi2wv6fqtRoImD9mGhNoCMoXWTLNvmajHlDV5E/24AEmTTuDXV
eTCh3BCXS+uNIl8LQgpqfezPrbLK+cuEbkMgWnGhsFPLS0gNY/lvUEbIkLg/G+Rg
rI+zA5V8B2xN7Wz1mZKNRsBUZiGKWuu1cmhSYF0Ryb069uxgxk4yXr5GqVRwdwj4
ZJQzhP4o93kj1TcJ2VJI90nuabGhgmodnddIa2mcRBYbmvZPPVVpR/TKXqAlJVZ2
sKKRSA4C8OYqZNAk735ydoz7X26RC9Pk5qDR/OwbnqBKYQdyhTpdbE9h8NGVC5nV
1SfG3GShKuah8U9x5/WDeDjKanVoSCIOdn+/mrUz+oyD96/cadH0/52YggLNdq6t
h68qhgxRe/D62whDHzvVvRcL1fvBbPnaaMUkEhM2rVR4h892sDYKvgrHv2NGxnuH
6HjjO4zrGrmJsdSGLc88pasP8d1md4q4hJ8fJLCskqs27/oxOXaBiESMiZDH3A2g
riKnpThXOsRH+dS+CfSyDmyIrAXrNApvv44hzJ0WsAgExKZ2XO8kNNn5J1G5a8v8
s2S5zt+tPAFcCj1YrelOhfN7XeJkhNjxsZGyKCtD5lf3ufJRSm5D493Yo3TvBBJy
Ck0GmEV4R9cimzym1xrSPOFZ0BcD06SdZ/kUzDwKLG+au63+5Rr6i8gTWFB9UC62
d0VhePCj7wMsTv+ni1rX428d9T4USZ4HgOjKzEHCxL0aXi2j/1rIEm/lweJDEPGQ
4qYP3osqMot3YdoAzqCwlTk8hbuRq4QwbnXZwLSAKMDSrYFTtFCsWOoQ2wWLis9h
w4LIP/qp544J/xLRkWhB8p8uaiLkutmc50cEOEoWMTW3xxLLtkDrgWw7xMHFwiaU
fdu61BSePh6ev5jrES1N+MAG6aeXnBkLeYdYt+Sk/Nh5nf+LHpTXMw01KXvjTZq2
AEBskflkqigHVl6xII01bk/HmRqMbxsWwu5QDkjm6sEi2lelqJG0PAmrrCGU0Bw9
+o9TfVGBn5aoPwdQJhCAAr21UH1KX4qEvm9+7xsw9Ho+k+f94ncphmGFx03FjBj6
4/zE+SgJMWzi6jMeOF51yOfQ3KzbIJ1HM5Shb5ttkfj65OUyXZsd8Y/uQM/LMxFH
Bawj+Mnf3t8S6YSxGnBxwNJ6ywx8a8wrU79vAuSPTqTuycsRurFRWyG0Tzs2UOJw
SWAraaz2Uzdf4WfhorO3TSf+sImshwhK4GdYS4LIhQlgjW70JUdACsA1WJuWqGpO
s6VXDThxST65SSb+c/ilGP8mWAijYtJdJbeH9kcjp1X+V75tUh2+5sHtqHKLjkdq
DQmJ5f5UOJmJc9Divk0cCQMGtnRloLj3/ryn2ryBC4q2hNyaW91tck905JyiPIAK
RF25mWGE9P/NUNnkr1SJYAjfhLDY3A8ufw9JIoJatK3b0YibVbigy6IieOo6BcPa
fYF89OtUoTfWXXZ7eJ49RAMX+si00GWzTeP8nsGQuVWVH3UvV5IvouyeFONajOfg
kfXNRFQ4QapC8NHd9LtHA6QLFxl8jJhcL+usMSs30cvZBxzchJo4JjclRs5u3xFi
zlQGoIpHgzFnbu64Q2qgxQWF2qgUYAd2SdYHhyof47ArF/GzMQ/WWxNWTcxrG4DZ
5ew/3jZdnSxtcToL7htKo3vOLmtXWpCdwBUypIJtYYAP0lQe7D2UrfTalEd2D3Tf
dWAOtFFaJpbuHqiJX9FNZnnS3x0kQSQttEx8vqJwtAgujIzrv6ZVv1lVBQMSuMRK
oW5z4+7vcab3vbjuA+0uQFb8ixL5NbHm/xwL5ZWThhMcxd9ZMKXMaMKhmlsJTV9m
0+5UhC3MQQmrp/0sQeR9BKRzuExTi5I2MEMwN61UKBQDH/0AJVVFe8UVIEGyJE1U
C6NVvPydcBRmdK4t/mm2Yj4cdHtf4FHp0PIiciWR/3C8Xolk3Uj46HPSEcDwkEZK
Vn7w4EEhlEQCirdbJTjo2mNNkyVxV37YDcU90/ZsYydPDKZY7eyR9+ZQhMdFdKuG
K3t7lp/NA1gS28dU0H5tn0iqJaFQ44Ut0nuL95rN/N1orc+f1PiwZxgZFN+6I0kO
uZWzfKHN5qaikw5hMfnhItb4TJjYAcD9eqeWNq3C9CWKgv3OZ9Dbf5XTzAdzGDDg
e9tjmnUyRSnAV+oIUN/IY+GllN5NCrPzQJfVLu8Pwiou3pIWFaMHeKy83cpmdiZR
8PecYq2pWUUc/KafwTRUijHyZ1YUuU4BRqqy+6hmTx2Yh1/0AvuIaQzdIu3KPF1y
ie82joAIBbJXFvXFj4IcyzwYyItLLVqiwGCGzHmvxtcWh9VCt5FYwWPVUJk7OjQn
nadAjvo/x0FEepeRDTI5E0bJ8j//yjOuT1LNyoFincvrdbaaNUabCiKsScJdKwdz
We93vsrbNWbIseA8BuNXthG2KfxYLnW51lN5JiNpGK2FmqgIXFJxyIKzw6w+WEFJ
ms3bWlnHTi9DwqUKQ00VL3G/uVAgUgCdZBVlvEHYHXbncJ63UyEDNHcObbAedpxN
ZoqJA/0YCmi7BYtJ3UQor03UGWTfzW4aOcGu5H7HYpua7T6ADBZIZoBf0OsC7l3C
Y/YIQDy/Zc+U0W2vW9Mm/qEg5b8+YMORUD9b+5IB8/pXAU42kotWi26iqIeAxWSZ
1pgRZASpVafl2wCQ9yRpqYOjNCXQ+9wTDGnEqCalDLwylcUjYs+hDrcWFN7ZkfI1
yyyZbtv/s6Jmv6rnvFh/lnoqSWSC4C3jd3JBMkyrSQv5YzejlQRU0czyuSmhFLYp
eoUUaB3hWwO268JFikVel+SYUVnlEwOvhp7aeU/iOVDpxhnkIcjUJqPP/jIoKF/q
BZ+hlfBCPimH564xGFFSQ4cNEo4mIzb9CMIdRN7znI7iv1iaJPHfDT1KhOCxbTFg
xCRYQK5LIvQQNDHDATMuKpZVXn51ivJkjo6Io+j5sdGwnNvm9mBWSoyO95j9KLzx
eo23xobqb2QVBRNKtqD1VDrgPghhiK7AQY6w/QunL0lbGELsNCiBPYhe779OLK+e
707bYKMfTo5bXwyLYE8nvA3jtQ7Wo8pzs52zuC5OpiWpYp0eMCr7cjVZ+ToICm+C
0qjIM+zeztrJVjo8JoDGr2HIsA5xkbE1OMHjqAUyKYBC8RQq5ezc/THc7OEAa+xF
FvAbhWuX+1KNbhUN7NKDhESPGQNjXQVrMfPq9b9YzCu/GSbeH6yrjBZ+B/DInzG4
V7wf+T0g/XFomjQF6XTrBR9PzXFNLrEcKTaPropKo20wtIE/W8b9ubAQG6GVxjTK
l1mgHvzljdW4LD1Fu7P0D2RGhUyFpDTE8JoTPpehlrL4NhUx22N8N0CB6+efa4cA
xMOsnZ/8qQBsbULmh5XA6+0PVg3Lb1pHowwPjzR2Ii7/ul4unRJIYVu1aRlgbUjY
3K8A4/h8nRKB9ZUuWaLKAtii+DkIkTST7+Zzd+IpWAmPVDYewJBNciIKeYGhgZAl
45Jztb8DBRVypUgbZ58aFm3/glSEIcVgoEJxCLn7hAmb6hbTjj+28bmomirZozys
YDze7qk6FeEWnfFsDt/0ESYtBM71LseAeaxGqxMVKz9R3YRt0p7hnUC89dXEJp1A
GgbzIx89LZm6zjbhlobKAvdFqlOLMVGnP6CsjL7/+sfagtRY0EkGMED4c2IsY+aQ
BhM00acOdRF9JYxAUQdVBlwG1saQwKTYeV4LJ3XnDPasOUQzZVGDKYCz8I8P6VhW
c4KYjLjNZaouMxa06Z8G1izO/Um3kVzaS9ftfktpTR/p4GQBTNk6l+cDVdynL0HW
FB1pW3yireQoA0goksERMNpa2YYxLMystxJCp4d1nXrF9H9R+B4vyUE96Fvp7iEb
Et7BW79fr9+9zkvn3SrhvUhmb2yATyCm00atMwnJV+uT4ymm/4GHA5Y56Py6eDrg
w9A1Y7BtlrJyQGGrZXKPt7mlQbL8eUTC3QziQ4lBqmKXn4Dn/m5tY4L4NQw5bV3c
3yojH2eK/iT+ZrTz+LGVQFVSyvhgHOVaWggLJ2IvC2inZa01lZzKirVqZJhOYbTM
HgzkgM69vBxzBVvSRre/nam9lDETJJ8DbSse2IT5b07BxKdfCJlYq5LJ6PEFlLsc
waJ38qMruku9kpUjGGsoIbdJVhw/GOGhQIC2EIcSGCEEyZIihcPrXsbeL1oh3fQq
bg5X6lTvTRn6ADDJFnJr1Gsv+wN6AVDb/lGkXMYpQUnxsG18A+SB4hgtkGD0StSh
pRM6GzrvGBeETIomh0nDfnkG79kJGQIoJoJhDTfyHWS7SOrAx7X5iwVnRakA3n8u
waMTZqg8sDYK3MFJ3XJrJOcNpf2QB+97504NXcwwTlSULGFX5zTw1tx+iYDEl5+6
7E6SS5p1uAu97v/QQLFVB2qlqbdfBZbT+zMcXqdG/v0oc9KlHdSj4FLits1LGlhr
VnjJ39h0pGMdMWs0ZZttFvSTRcRLmv+zna8TC+NapOQ/26olewSdtHliVeZzmHqt
faDdUPQGRvx/T7dM9L2/Ql6r39obos82mEhe3hBCBvPARz1RuSzbAMpTWsLbMKZx
CVA2426Yi7v6HAXxa/oyo3VNjdSPxrhlZ82Y4hcq0osso1d31IabKq/MmHOjgt4R
e0l68Ra/I7yMVWg8jZ6IdGD5VjQGaPr98svyksQQR/9p34GwBm6rtezvmQc9BT5p
Itu/5G5x74TfcX9mhWE1O2DvIAuxJwrhxMvHNlcFscwdySFdFIbUlFo2kjxu77Te
lp2NVARyFMvLM+JFuY/iFEeh7E/ISDpCJv5kZlpRbAphKyle4f5YeNX93PsGWCW8
+VXA4VM41bVz8kTyaGDgTpJJrZJVAJFdRvkClZMGguGfcxnc3rOumKS77yxTtUT6
AkbFi1654L6a7TA2N0EVY/voqO9SY5v0Bg3xPrQRd3WvZZAXMO7WIWyWsS0pyBLt
Goruu9BJj4WG4FLhUqfcqybtXe+ZRk6RfHRPWMtRTfsyAysgB27VAsRY045h8J3K
Gy1ve2mcIo/jywZdW8Y84QS/2iksT5W0SNduTdWYVE+ogDfPLf1Abp92hWiKB4vs
4xPnvWCjkdyaFjGL2E89oP2h7Z/eOMOl8t8F++6scJGc7yXisFDugmi/bcODW6Ry
w/SkXQEkfMnk4HLowDgLfRXJWxJBN43ycsG6wcJZ61ht4jOI0cUgyxwK3qHEA7m6
1DP6f4Ay/RIcLOAfMVT7qrBhsAUUTlqphqO1kTIUc+d4/rzY9GVd5EwDwh2KuDHQ
M5SgxtYrH5O/DT4Pc9yP6wYE6ArCl2uxnVvAh5OEXAgNQupFq6uA8bq7ZVtScx1r
91Gf4+f4xjPoY0x/4cIuWXW/SaUCfaemma8m0u2w0FBVarv7iBlKT3bwiG05mZ2a
1CQRKzNIXjWFK8s6rzLbq+XMbSxAIvOgqA6n+EHOp4NBZFCB18rEbI5ITrV0jgaX
HUw7MjQBUbqv6wub4EHFNA1peP8mWsFhDNWO1Kk7BmLq5lFnb/ca3hwxmLP0ZTeL
XUYuoTD1Y4681NBN0OXIlEAXoBa0lvj1ODhavHFSeYz8OPPP1iqDUivrj3sAbqv9
2mrlxCjd6rk7sufr4Ey/YUMCoItHqVB1xuLFnccROZg/b/lquXRcbiGuUscfEyfA
HDIdwvhK8IMmBDmPEdN3H3j8lVzupVUVdIKXNQU1f+ocd6JQ1pArs2NbYt/cUmZm
TpZTDAbwIfFCSUhUj09vLiGPUDcPkQfhPXoJmDdw7KnSPsUHYVkIdxgV4R+jtaK2
7kmkIMuBSM/BtLm3exIfUEflfdmpA9iaSmsdDOW+1GpG1xdtYqpRBfLt9BMHVVge
qZhfJM9JpiRfmj0OHPlCwgyhLi5/c6hJMdXrg46zZ4BB6aKldjRkcWr5iA39eqyW
Ce05ncL3OtRf+FE5q/PWnteCrpcLrds3hgzCNDUHHXXKlP7C6gkz60W/b9hZJdEh
cGnPpyT8u1+ruaVcZQmv1T2tIuEVpLwBxohaHXDjE6I+VKja9AQzPg5DjyC8+dAP
drZ25NJVTYc4tDGm4EZpChwbyysNNRDqMzybblEaVcCTKyOyu1XpVqVQ8TsTiONv
rN+lNBRSFJ+iYc4Dexjp+ipk6qPgvcKUMyKSZBJxS7v/uk/Ys4lWlURvIGAJP7kR
rYLuG2SwsaIpGs/SrxMU7D9N6ZUIhT9kefoNNZsOHpUgzJJKBHRMq7MAktwF5zKM
sodSOF/lbSjW0sq3qbNc4RbmZHRmZRR7bTMdxuKoUu6mMNqz1DEBLKxirMSZvmh4
S9F3GDYZ7wPPGxPcl/MAurQxmw++HcJaB3AuIt+oXDCHZiw18ulFWQ/uricGYCdU
slqWL5Ed4AKq2VjQmftF+DA9QDz/1yoyo3XCcFt4Pltedv9C/H7WJIR/XfB4PJlO
Xy1heYWnFYLDS6mlE1sDiYFdQb+YaO1ujBrEEDqfuZGkrr6Nx9JuWxTRAMIjSuG/
1M6jBs+8RDlcT6AHBwE2zBy/J9xvPGOcKG4QXIC+CNudz0w9071uckrK4k9z2Vmq
ZjodmfhgaPKXPGY/x5I/zYfi6bIuEyzBJcZqnW09C3oxHau/uv5NyvJ/QOVci2TF
ZhApB7iMNG4siUAp3PwG+l4ytfxL5cyA00JJY0aOxq44FDs7qLzL5g2t4GPj34Ok
nA92PDYV01e3OXx6eUK0aucg86+psz6FwQ3RFjYvkgsntREvL2CSvPuLoOjJ+AU8
j/67YVUs/yDXTgF4+pMt8mw4Fz7LCLFs2oPc8uS572+B0/xByAqdaXataRbMBBoK
yCPEWyCO6wLe4zTp0/UASZ8Ome3vAKzJeImhNrxFbWIoF3dFwj2OXwJNIr2NwfYH
nSHbuYfScWolkqBRz+e3i4skvBt0azlYaGhxq64mYXreUyrddfGuJLyRqrQGBbjC
93ZF3DIYRXwGt9468TmpPkDhzlbin+97g+PqmvvP4oWFJoLq/OgkPj2MTcP5sMes
5cC9aupZ9k85lmq6VPa95hUDvqluyaPx/elWfWXsNhWQ7F1laowxk4NwnqUnGAMw
vhYcStUlsECJkUCeDkbMY1WPFTSwiSXnug7SdYkbNcr1Jemsn5dfxCoErfT3YH/I
kdUp9fs3rOQUulqsmJxSLJhLQ1v11qzzlpgwjTZFpfj98z1jmiF4mGDeR4brGfER
eHIRK9MVvBBhrQXhO+qUxR2Wd3EX6VGfV4Ef9OGIDVBSLmZ+KVI7gBD0I/PXehfS
jUub7wGTiAoaNrStw+RyvL2HXMAHlzdV3MWDAqLV1899ybkJWRdkYnNIqpwl1UXY
atfDvMUfQncQ8d7+UQdKV17PHvvrwN9XHZ8/sW5cxXLgOLRVnOwweYXsU0XLluSx
ebXdst8B+b23qN3+/lbLp2shPmlBonzNvB38EoclcUB+Hz1cK0Iuo/xv8AlWC/G9
K8rVfS768a8FAEPmtiJONDLUXV5VZ967W9DdjyJrRqfdhU9j+cv6pwE6/pmcan+z
SMPIzJSVPvgZNV5eCaPDnDTXIMNXgkpwTD1PkrHtJmGx6n2GGxAbPL0upGHwt7Sv
CSpr5BBOuHWsYTX8xCd+ott8HcsNd3TnUsBGhoQF7Pp9YWKKAnfINed/QxdGoud4
T2BElYufaYGdWBlrC9tFnkYDMyExIqLQx7ojtJULviYSH7ZaMuZwFnZvHu6UxIO0
+kot3LPr49qWvqzoC+oyyPhvHastxpMc7l9BWM6KXMsRlBZhNkeEqRzzFoaypYzw
SI/++bjEhv2VDuCvc2KMPCGZrAHV5h6K+a1I4njAU+7u/rZTXhmyxjLFwaPi46o2
Si0Yl2oRcXSnc2Sxmlf8uM8DDqDDTDrtEKb2kPC8PEl8/Eurm5fQFUSEa2WBGJtF
2Z7Kf0uy7R1sPQA+9daRfW8KoSuv3NETu74lVwkOrJw5xekGh+dEogO2HYrFngQs
oGLT5aQP/BoJKq0VoQd9ZTRKgq4aohr9EZPL+xETi7oVfMffymXdoY8Q8KEk0oaG
Jbn7OMsPO11FHDq4tY1aT5QOjnv8KEM14BKM/HYPbCFPTlPOPAlMcq5DIkZok8uG
V7/EmzL0qLxAO7QYUJYf0zxuGspgSLn10SncAjNvx7rsaYGd9QihLN36gbBpn7y7
BJv6rSQaBXj1Ne+5MG+98lb7ub1n2WoMC+SFbQzO2XIFIciQ8xinpopjvCDcakcY
S2mhAl4h9UhqQv6efsGRieJFUFlvYUCf/xb93j+aNMtMe829eUW3OBwei8cYTGGb
zmMHc4MV42+ySZDN+hKjm5vjKYn/x2admbi00zeEfyV4hGD0i4UqKCEfC3Nm/i4H
ZbJ/PfR4oNeyg3IQ5opt1lSszZnnOdIyYZlP7U0kQqjGT4devWgb1Kl2/1WXc1gA
muw/rkNhd15FnPx6fUS0D1YRUHYVe6LTpmXfGWJjDdyjg2QeayZEsduNPUObFib1
nETgB/CIaIXlROwt6DscW7dXbqQndtcbdbPaI3W6TaeaW3knGTpNlFCTd8e079kM
LLvlsWfjt97DWNHgqh10+683LL1THQVxeaypaVMx91JtFXqER1gAcKUh26oGw2JI
GHoFF/Rkf6yq2AE1MUOtFSrhRHkaCp7pNysf8zQehjDYC+xXrmfNiEex4tJ9Mzyl
gWJnsQcJzJKOJ676+3aRzZPN8FLymOsTTJCLZuD3N3P+yL71nrB+Ve7W5yaMnLQT
7uhRjw+X1KZz9/KaSVN/Ozevn0hqiyH6QMjzYRiGHaZyOyvY/MpLH2nTmWlLXPt6
41tcoOs0aRk5+hvUEMRHLbNrG6dW9GssYlV0OmHOOF9ntul6iItL8/jKoIRQgT3I
1HFs/8rLqbjeyOhlD91/3AkisZwxlyW6XgJqVVFMY752Trx4q9bzhC0qW63sV4OU
RXI5EpCO5DIarWWSffEzd6BYzD6TvVCr38nENwbIvhhZ6eIbOPDs6aRywsjvf+kk
4H+9S1fx6iN5dqeqQehuyuRo25bCvpKdfWrKipBn8TopcN770Fw9jsDXMffFKB+6
qRuT8GjZhR3KsDYlNMirPmhiN0g9BlAKqpnOWkSR7dK6E6BatYNbB8oYzSzKHepL
dXRYCo0W80Dx5hAQHJTPeJaCZjaxA8p//JtqqyuTiLG3hMv8B/sxOpuFBK+PMuG2
SOg1Hzghij6VDm8oY7RvVU36SmoYuBYCpslQI66hYcnLzdtLaPPjXvMpm3jFQVbt
C+zIysxxlo6k5YTM7gFaP2b0CEGosY4xEp+g4CuuXYogkVA1TIa2HJ9UxG4vqTaS
clVuWphkJA6JLGtOWJlp0aLqVuzi9a5wRokW/SIUxhMZTCatRHR86BsdvWbIo2Hu
QQdKnZi/6A/yBW2OANlBaNjjolfu2VZM7bMoiVERHVwpBt4sByXBlIp6Q8UmZc+p
Xfy+SBn2vpECF0lkUCOX9GHawk2j3cZqBE2ty4rgVEKWtJ9LVknLOxRmjaRLTzGx
XzA0b8LnWIYkWvzd5IEy4XORS7oRNvt6Qiiyyk3svkLC1haEDJ33yxhOQ4KSQYc2
vPZdLXvYTv6CeBFhr61MRbHUTpi2GykDmLeHh4BcCRdeqQFBKhTZl+XVz2llD3cv
LOPoM4G2qkpBDw5k+x8RlnDIioQEyzXeL9LhG/hh0koZ3231eEUY3+U9WlpyLUYM
6zG6Ij+7nRh5eDPtiHFJcTrtMRCPXU9DdHxA/3yOY75P80UhceKV3EM1CA9Oc5Bf
p8/YyXKB/n19oj/blYFQt46UaIySYNtt9oGEzTtQyjET/pLuWnYmzBn3KgC5GKYu
saCZ3wPmXibbmlJd+hqeuj9LNemnoY2k/LYb56/GOROAwrbAylZXRJQTr20sqPaS
MlvACNGk75kJHzDOZW+cdrtlIpnj39e+v0uzwe4ondWbrNj+J1YUT3/GkRXb1vh2
dzHwcxf9AabDZRlHIY6M8duFXCvYCr/f7jfpSFrJhUvksL5o805eD54EwTAJ+uBS
IFpQgQlwvTk07o/WqvTNfaskTyidhHq9daD1mqT7zv+VAo/cIs8EOJYZJLRbRtv9
qTlX8A0qjc/W8VBwDl/IGUbcdsYrxm1xmedt2v0sJhNJ/Lu00KShe4iaAmEyxi8P
R5AGWZ9r2Lid6jnluuI1NC0gj0v83pA3e2HjOkDjheDh2yPlB7bUCckjxzl0EhTe
BJq9jMJANGy6nL/4UYWeMsnPBn1ShcJOVKa/UpDC3WBsOA8nswMkH8TuAojsXu2Z
3pNXZFIm9SBphNmPGzJWgrMH9G7L3v4OhnBH0CWkNP0U8cMtY67KbDnJ5xibYv6D
/mbWBn/3hEnC0uylWjE0Uy2iaIdliZ+BmMVbaY8zllhcr0VVStUXK12gXycFBTS3
MjiOp/57+GRtUBveS4EEuVWUBOnY0emnDOURx1pAkFUM4NHQ/nBWlPtRgDIUYUeV
NcqgHExdopsOqi6PmAlbPbbLddynpaW+HfNNjQGiLVTaTgnlSrbxHlGFzmEP6aqI
+OS+cb+XRIRVtwOmYJ9wS3U2l/ANCaJORAncJR5EYQ8nWHEh2tjpYnz96/Pe7KGs
nP9/nY30mi3PFXWgcc88uC0IAmhYqcvbkkLM+OiQ9o3hVyqNpMqfCwyw6vT2Mzbk
WCs8RVOBfjckYGtHfBAut8B64QXBKGY2OQnNAfqPdR+PoO3+faR87fU7lYikHJB7
oe/+vrYDKmNafI6n+B2KoEZunn0hjfgi8wNmcyOz+uxwhMYJvmlyXVzMOFYUf17u
ieD2+zZy647j07W9C2EGhlS94Bu8nGTl2VhkkNYVBddFDFG5uTZQ4d6XvjmdiokT
Fhd2Mv2+ey6aNSe5X0oL7O1uHVtyO84G7GiPUo+zExqQ77ccj8cQrzkQaA2oT2QB
zfUvZ9ucsmxhBRzTT40vcTrjQMaOUASqceL16MlCRYN48VkmX0nyxbM6VMxuOPaz
WWdb6i1Cs+WQ2SzWfdc7hI1214rHgpYxIlK7DaqV8jTxJm2NTGOdgruWMSQMPiz7
HRUavw4KDg5ftKZgal4aUluWQ/0QHR8HGXlk+ONipR9/WtvE1cE+17wV8VhNsJfi
DR3AWrwjhOugD425zPQdpQ0PaxU9pVE4AJCO8cVpY7KeMaKxLdmX/EgiV/FnObBU
9QH2nJlLyRfBnwMYnaYOetchHrXw4LOhgv426RxX+cW49iUTlX4k+XUvu5En/K6/
1qpNd+4u8qWOmTp+5wNfULkpQ6hT0U+ad5ZLQJf8NcWzBO0Jq1IvFkLcIz8Ip0kf
wEqQZCWUUhtm0mIna8wzu1Ydyg9cNawsG3B5loEQJ2har80UL3a+lXKQ8LNbWRvg
pcvivouaqRnUnj/Uimjwu50ff+yo3R1MnBegFCB4SVBx+9rxAwZM/TmC7k4QSNoy
U5tKGCGTOzmAA5DQzkJx+5ARNYClKeExmgOCUrl6Mg3FA9gIzlFK4mgDeU9pu8Kx
bORAT76tlLsta51+daULHqqNRPegxWG16qzCXzfhvLSv+2CG5T8oeAnj4CL2O7u7
TpiY7CiFHex3N7gp2FsK1Qy57VcV36OqfO4EB+UYvPdd3Amr7iuG35tovCPDI/Fp
Jl0pvf0Zh+ivzb3TtGxCINeg4KxC7bMsX7XsBi/W0DN1QmSLfB5iRi7lN9ZS/Ih/
eduUFDU/up5HITUfaCc1HOLeUy63x3TJR8gHpn6iwLnbHxG7JI6o99I+pztltuuA
WFWlUQ9gVKHZ1K+FshpdNBEYgR0N7F57hmVponRsTcMKWNTjoIM8yH6kllpqKSqb
RnxwYg9KpokbN6SNfAwIOhazvD8bUTOyzDlyw4c80tBtY3HtVt9r0RgWA3giwfzk
3IMtsg+naA4AOKPBF5BOdMRwY/lW7Ez2V3qn9nuLCKJT7lYktdfVRACp5F7+ftUP
jQP1+11tpeZwUlujt3pfjsKoDT5a9sQoU8x5hN0vmx+QhVhdTf56+xQeJLVpZCl6
WOo9EyKZw6FoV/KVXunC4+xOn73ZVtah7oZsqJbkB4KUwImd2YdoQOCRLXXSVecx
MLM8Zk2DgYp0T41tAFc0V5btUN6l2vLov9dae6VtvwqpneXKKH2lMmuTXexIzEhe
O0qKQeLl8FC5vlL2dDBrywG2ttWXeBZR5BLtwZiEKrdYDvM4cOO/JFvGTwWlo2fm
iRBoM7sDjLVw9FbGCb758VVgrS72OWjoGN+WY+MhXNkF2DET4njg3G75Vpuros5l
WmAXCowYk3ESi6ZY8FfTH8T9ta+3tp0o8wFF0Ojhg5NNvmpEkahRGgIx7gtq6Elj
1ZdULT6IbjDXzrdZolDWORvb1mgsCAc/7QT60Zxy4c2+JfmQmrm5QeB+OG35j/OC
684Biwo70cA/hm+LcbHRIY+fIz3u3Ks5oGN3K0ksLNOSDZhmkWmkYVFk+ciECuSy
xVzZp1C44LggvjbIiLy7hA/YNNeLgD4toCWIlXzNR1/VLl9/lE2UZQD28AzYCfyC
jcm8t7hwP2zn88ci61pBn9I3hnwzlCmRIxUpj/Jaw8xKZLaDG9Wis1hzrHUYpCZJ
1O4PUfeN8OfZYN6LABdBA5DR2v8picy4ZRnCCIdBFfj+40k5H0pPxj+j1JssATDM
VVy7vjTdC038r8b+gqVuoKuxQMdRjl/ZYOJsDPaQ5CeH7ENuUwtqc7/1viIa8Upn
vd79s3YJXoho+7lhd8A9buZiiQLuqLzdrB/OfnVWAE9KDS2HEODT7hy7BO8uFbss
SCQLwn5NJKjJtwewvjKGGxQ/5xCLfbZ4yGtCPvfas8RNoliOEwF490zJWW1XbOiR
v+kd1RTrT8JV95XCHlnrh3SWiL4iN1uaknnAU/FUU77XFAwAT4EQbjTpfE2qCI0h
7yMJWLUdtcWFOmKSL15TIw0QhIbWqlm2ncS1mxCB79AisaFYfql/iJZ4IKTKOV4S
CFSqDBRPglSNgNV/cxXcNhz8h07tknVZN7/fcXkLskDiz4z+5AYO9GOtcoP0cluA
cThwd16SYy82tZyHKVSDFqMaiYyKg8UPQNemYEMw2Qy6ICiKKaGl5cLIS++Zhl+J
JFvPwTuNVN1Dj0VtpPyyeXaJdZD2U2QEmFYpBinzIvIwAIdkyc7bGlWweUMf6yE1
AM/c3dxfcWepov0CJXAfMrdavPG0S58d8I4LCt7IdZ5MzVqLgsRSfBbU3D3/SAUC
mmSIYAtYKbw7sJKyR1/TNEeY7spnGLJEVCBp5teUbZHQUiDZNFRYMMZnZsV29Ig/
fdUyvE77mtPbeYV8HfyooUfVFsl7lQlhhzN59APMbjoyQY20/FUzzR57jHhTooNa
9Dw2YOMT5JrukN+kfRut2TpuDSfPF8yWnI1iH0UWD/wzN4fIq5Gww8Vic9mwq+/h
7xg2BoEZ83XSquif+W6lYStkk3lAbmDAowinnlzyOR4h7kaGG27KxfoLtTfN/mEE
WzJD3G0Jyi3mzS1/xPBZb7FKhs0l1jO2CMekwI1jTPyV/9TYHyF13+baw0g4zOs2
hP/08krHEGMAFul0ropvYOI5Az8CxpG6jDziDq5SSbqWSGQNz47BeLfjHhDhWjaY
1e51udFH1OC80MCqPFjAmnBpjuTeg7MaaekKX1MK9HjOq6J1Qe2mCBi2A7iL6uMY
+iv2JdxAStA+2AvO427MHxnEi2C+FaGmoMt0C41CWlaFp3gKdqqR3rWKV1xuvlX1
2cy3BmSphTJkIwWHuCyeXF0CNkOie6snRh8IpIwMGBHEixNHCORi//AjESRsTheh
q/HgnbIpoBYLWHeZPKrYGo5BruUzsWYGy1uLDiHIalN+PWADGuL/mkbDy9RDYLw6
wYSvcjwlOKHJFJrlXeaGHqIO3UsqNynOuwYouZoesl9DNf7ZoBcXnVlHgmTAh5W2
vpcAaM7GFnni9knlNepl7Bnoj9+iBJireAFTG/OlA7AI+mZIQpvu9WLHzsKapuBB
bLAZZ0cdQ9pt76zZfngstlsSrJBzW97GQHtZKfA9d4qr6lXOoyBC5qCbjrJsCHfI
0ItVEG2H/e5Shb9XsTxJTSdY9ArELBPa/PjwqGoa+O+8QpRxu9xRbryucPwKkcue
7dtEiUMpudWsdsOHzZXsLqP3BCZJhNrcPRH2ya8VNmc6ovjl+saFSiZ4bQa5Lgk/
aprylQLSw2PXsdS0/jzQxGPtOK7HipBX9174nG+JR2LMvuSrt27lJV1vrXGPRZpg
HMgiiyvNPBXKQPOHNbit5PEvcmLQUc1YU866OHIpasEQcUK6RPQ7A+GR+iSp/40t
mjJQJu1xwTFq/B2sJr0SmGUmflLZy9GnZecYUt29dZX0xajGwYxLzwZWOA2UyJie
WfeCZ5ezd4gFkkRclRPtgG9Hx7XeFECefE1xi5TxIo/yzUivEzl0eDKKpmmUc70v
Fic5Bi844ItlPEk/y4ELiyCGFV+QVQqS8NmT25HZxO8qCaFJYOh30LPO7bWzH9lo
FCsHeObTlaePTNkZV8Geq2eW4X93khhyffpfaAVk9o6clrGwNfHezO0+x4Kgp5YB
LdbTRa+tC35r/6RKWCxoZaEJzP6IWCCJZ18nxGpgSYgB855qhYTldmjVK3v/p+Uj
V4D/OIWtsYjd4CHjVQ33UixR0kotU4u9wqyOnqo5K3LY5IZL+huQOzk/vM6+iCjg
U+JDIhkg7Egc8vdCRDbjtS6WvSP2zhXJJhFakwubadQNTYB9Wl+dM63VWzJ1GIOi
hblff8L06/+VY0slkqGphwSPPylwS+c3grryXzxIEzWlYW69s/6gJqdwrR1jlzIf
oinZ8V+qCOnJCBk8XX+R+4FLBvvQ9oWIR1J2fXwWiZirB4VXQ3xckQi9MNOIzJGF
74uJ717SiycWIwdk32EmjpXQVWZRJEB4SZHmcG/z1y3420/D7qzlWbJhtllHKhVU
FmvP4zFrp5rBwgfPtim/6fic1xQ6tF7XHKj9eIpszbeJ+ZgiboDMgAsj1w7glWJc
rkwUx53CK0+8fTBBV0DpnuU5ngavcmW/pKVGizh/VepLzck9QazA3rRm839hxT5D
jsROJ12w6GhujC6Ae5TqVXkfV5PoxSNnOEvmrhoG8kB86cGGQtjwran71IZJg1fa
Nb73Xwe7jsP2Zyd8IAtzb36VgObv1bPRGfiskOkgC3rxio1Ihzx0tyeY5wUAdOJx
86FSSlSO0LXY2C1gp6ekv37wGcrUjwJoPgFheHPBQF239S2y0zlgr1BdzQiWvs6T
HRPBu3gaCcuQjxQjYA7Rij9X2/JWxFp7EryamKXgBpv04nH+swe2GBzKoFxhbInW
WgptnJuKK1zgKhiR36+0zjvPFDj9Kbid33i8Jux2Dt3ho9YvNrSo4YOgCjX8V5rO
6K3B6qtvBHVqqhHgFy1/Phw6uRbbBERUMHJKNxtTW75q+0pwcnZMR2w9kGcdSA5i
ry5/Zm7eYcOG2Kg66lmGjUOb1J6Ad5doyWb7tLFI8p9Dfi6ei2zyATvpmyw8haIy
tDZN2/CjVJPbD6+7JUfic39WcmfhKXgLDj0tWZx0LbQ5sYq3h03SNJM1sashMwPt
l5IIqQNwwNUQ4/LtHMrQTdZLqvPGGsrP6s1+RUVntD4Zeb7DICbEkTnaoS6umwps
YY3KcyOyyNUfJ63p4xBPiJMyCVOoaeCbG1IwKtbk86AnEMirIa6apxMhOwX+qhsM
3dog+j+Z+Y9CmcU9WrU2QGQNvwEkuX1uSWOkvnpMRfXmtYJgvBk9PeqQA0gq0fW0
/Nm5GK9oea5ADtQSSaCl9AUff7npfQD5gTP+nQcXglm4e13c2x1ta5BkR6xTXi4P
JJNQ7sDBz608su/CPKTwZpEntF/LkKM8dKlKCH8NcNJ7+lmqB+IUVKQStaYeKJbB
JYPVhM7BXqiefBlxo4fLJTwOJTTcOB+y33rX8QXzU63k+taORSCteFUYwY6rC3hy
7GZBAVYAN8D824gNVejdGsrGh3991StnEmPGIFBjLF1E5y+M80Zle3+SCseMoCgP
a72bYkpMrWJzPHHBNkKjBD9/OEm83RM8U7PA9qJ2T3VaBQ1efOqnr2EQfDefPRO0
tbe8gyD8SKr07y4TrdkAnaAuiKw+GKTCb6kkDZs2ZV9F0M/Q5tkgYjPPg/wMgSMv
jFxn8REkdkSVjbrTTcmdttz30f1JYS08jqsLkjGqH8R5O2/Sk50dMMkigLRBSm+K
CifSSEWKAPf43Bcuz2OtJPvWRKS5p71NqcY3B/dgCwrLNyxvQ7TJRy38BLt/BA/W
QEwbBzfN7TjzxvyPnBpoS8LPuKZ+fiqGH7Q6TrV89Ia3mp4qJfgbBPsxsWfffSlI
Uf3paLQPUacCkTYSn3Xkhw1nqJY1/HDAZKg6+tbgZGo2SEHsJYJ+FM3H5eFe6t/Q
x3O5HId2JFo8iIuyKJOIeGMpSjdF4T0mFGqyrOu6x7NwBjyDOZ5FWTAIJuUf+9ps
ko2juQnaOLvTAOZJCu1BOV3qpzuwh3OVtyuH3w/pyKxpC61MW5E6BgGKFcmwP1kK
TthbKdVHhrS9BZ2w86Gi04+ee2gQO+1NJaQ9CcWCTG5SqMq84gbHVIr5pKRZln7u
Mi7eFmNvW1hTei0zcltDyh9eQieBnxk2aUPnBp74JWAJVZ2Qm12myXAHelbd5QHz
DWn8tzsHcTSXZlrAUFW4iNUZimSbb0/cxN61QzX0/wbdJYfZi+clS/QhOtZ2K4jA
IDO0KZt2hiBAHfjtoIW0h1Sfo5jBAWp7eObeJC5mJXYEiUgaNta8TozDr/dDDBNy
QQN1509ojnJALRTUGTsA+Hy515L81mIpxnJybyF5Wp5C7wFHlmqNznZFi/U2LA9Z
2yYvIYpToEjJWPwlaVsqbxjG5HcYZxsOIVAAXrR4bXfQY68PJqUhbZgs4va97ti3
ti4X4dg6grS/g4REUrXBKzTV+CoJOJNZ7MhVhVzyYuzXPl1w2pTd+bSaM4vO2PNA
iwqOl6PJImS1qFKP6gMDTEcGY9VTTOT/ch7X7x+T5FwJDZwAMDU3VSqK1RLUTOjG
hQ1CWzoew50YbRT8JwmDOYdioamK5SBhgwWL58QSrAOEXlYiBZPcEPpuKDS7L1qE
iPFUCcmd6jAcjAA2Vt6fRDzJ65yCTAxc8OTgEMqPG9xhajUUmfKTpp7iEMmkib4N
La+mnXwPrvodH9l01M2CA1d62zBFo1xUrNhmZP8o1kLJHBAt4SW4cYk6QjMa1R2X
HRVgi8KApEMaMBebtmH6tj28Ynx6N/tDVEoT1mTk/95BkBQ+882Si2ivxnwD/6Cz
EhmwQ3wY9VmREu8VxW8jUbaCNe+5NTOUsJOGV06+LzlEFS81vAV+znXpgfvhSyeI
kCSMzI9Pm0J01ZTpovzU+1R5ZFBTkC9lPxyzyfYA5qAG6GSGwAL9+DF9zhhYQQqg
KXNUWDn6RfZTIkUmkmLwt/Y6RnoDNJXt0KkHBo7F4q9D6U3+7G7qu8ZfruT+KhoN
7HN4u5eXKisYGVxM0DV2lQcGckFWAbtYlCWKoP9zJqqlnUfQIUBm6llJZd47u9JM
QO8byR3nlhCs0TUwu67TVeROT0c+LyZ4fOUz06TbHv1h6apl3ZYxY62ZbGOlKmfc
eDeiXMJslDafkxLPbvibg9fgZY0oEXANy/XTKX6miqenBaYrNKg8uu0aCvXNJEBS
m+WWjCy7sn7LMFjHWzvA/4P8WIZmHHRU0D3a/q+I1DvARPdFVz6q+4Evc5lyp5bw
xmslEiCU/mutMoG2D9cmYk8JVbhr0B2ByQ5mZGErJILmyGDqq6azhpINSaWZm1Oy
rSmM+geSBnf4n36pEr9L7+pTaQXE3c5STvn3aPJfZRWS3bXKAY0gP27r7Zte7cN6
pLBCfkther4dlBdDzU8sVE01E3fZ4lYKOrvRRZ4+VP+JL3Y5kRzzELwjkb8S86gN
Ri8hUj52Lbm6hgii2jhA1rw6rUZkQmauGWyJiTkpjnbeCEupqVZGMwH/gcKQZXZn
DPoXQE3tX51+kbI8jbVpGXi3Q36K6nLvTywWN2fpAkswU6+aknmhAYfsTIMoviT/
k2wxGhKDtnXtHlDDp9+4A8FwwL1vNYsGJtyTxLktT4/wJsdMeiEiFxQRE5UUbH/B
VdO78o3vIOdfyxpG88tJZWx4TovedYf+w2w9aOXD4Sm3QjMBeRbZStUdJli4BiTa
Mzz/hj5xpp1HFD2nJ9YFK+4r23Xu/H+hOaI+gWTatw3BfPr5LKVHIBO9kgANNljs
ORT93i/BUoXl3CPoK/wNq/ziGTKMIfqaEaMBzraVZ4p6KKpVyPIgwQqVGPEmOBXV
VfuAB3y/Nui1c6IOSbAME0UGT9fzYjLeTaN+pR6Tzh+Xn7FOSgJs4tfiqvHdAoJS
SEygHxnt+5iP+eXvrefDZCYC/nAxbe54n+OR2wHYUe7XDSml00D/w+qgqfOeDorS
8Lq5qHwf6glXCFvs3FuhorYGcEBtPYVhtH3HJslPCZ8YqOi16M4Kgi/UfMR2EB79
jLHqtcwXhNyqA5ULiTvkBzy6E++QrCAuB8/3TGBHS2XU92PV709ALipmY2RwAp90
nJovyT4LXdO/De3lUlv7GJBIqX7Q4cvOSmAnJPLtwpgLojo62qE4hFey463adzMV
ym1vmmbGJWivU0XfDXicCatwSk2uUVL29KN1yCCQ716M4WZhoipTN6ml4p9ZzoLW
zQEZW5ynk3WOWyA8I0rgR2mhHqouJI22z9TJ2xcv9VoTLh9V76Z3XnVwvU9EYI71
3MNcBvTzKPZ5sfcLGwHusxgoMNAuNrKEG7+6/sh92MCaP7/Bu3inFiwWLeaVmHFY
56dKAHHlihrxbK0ddfRkqp567883bJ1Bj6QkhlfFuQooRq48eFR5AHJYeLAhb1Fb
lOfivAJEGfTApO2Rz+pQP55q3iWn2tGH+5x5KqAHqimtkTrIlLXr4SzIvbU7u7Qw
fCZeQpAmIglBr7XadwlTIH4xvp9LriApm/9wu8p3mM8yClhzeCPtfOTgnvdhmu/o
pCF+T79qbgLbpYBeG628po4gziS8HPI2IPCf6i69Sp8bMqOA6ij+gYd3hlcO101q
vTaDS1RscJ8EniWbd+0OVkw2VhMwjWswn2s6ej47tGEaiXDMLif7m2AVOW/tVlIf
2dngcZnoK2fLp0hwsVkGW+WGtn/E2ddIaltENTTUT0ddtLXFI9aDnyyFW9r1EGpg
qsgxtMgFQcKqlLPoBet8AU/GGz/qqiHbpC/UAHJzemSgiD23HWWCMXgpi9z7MV6v
xMyBxQNIj1EpkV+fZcMax65yy+bfwmyMy/1B8qQgk3b86yKkwjbWOkGW9i/NjLsG
qPtGqmU1YpJonIPEkP9WS0M33ur7/fgfoarK0nvpo7Lt5v9brS3L5BEuGLymZBzo
SBf8nBeIiiz4lm3qOKQEHEwpnlE8QdPEapxydWjEV+6RqSiQZo0DVDOAIIU1Jw8K
5X3WRmnIpWoS+NGuIXKjjSErnfSrVVWqU8kMGKvylNPj4Hu+RUxeiwMGfFdNPSRP
Pt883rFH467+84w5L/tIJYS8IBbLvp4Ohq3DBcbdWXFndVx6aIWhy2aBolyd8Pbm
igzQ6zFHocCgeH8TPwvDT3V2+2UQWqG0+PVojPJP+FWol16Ob/5ehJ+kw70TUp5W
jbT5ly2oaz2Xg4I/wnIJFNpiRdim3BMmiOeGy313Dk46loBNG3U71iVXfy7Ma0jd
kaxHvzQ40NeWnIQiYrVvwv3ugFlyd6Y6WJdwRWkW4joCsFVPGos9riSqDqRdp2io
WcIelpHcMXfyxUmP2+bg3aYvFNqe/KAiv/z/hY9isGhiz2lJIBT//gjw3/TU02eT
9vFr2OFbrRDft4qvkJjNjNKVToSxl/padzZ7Azj1iuABRBOvne88oBeAtgzZ90Ir
/h2SLRQJxEhYV0vgq/0Oh+kJfxYaQSKJSz9tZUtK/FNiqy5trfOCjqUx+nW5c7wO
rTmSg5NqPTe3bQHrvDXuvW/hGl5Q8NAqOEsS1ao8aJ48+LBoQZDVy7GrD7CtJveo
/LpgPmB+GuXqEsBhgR9UtaThgAiftnD9OvmdVc5G/mXDQbeVUDjlGume8K8PgxFE
JiCsed1y7yGIWUA+Z4Lc4VTzGmRa68OqL76TaEn6B/3Y1czpP1LPXb7jJ38EDt4i
D4mvdzNaQ24dv6y5MPIu9qHydlGl3EMHSFwILknLAEPeJf8ASq/SP13QhDr/AZGY
IDEdvdXoWFr7YRp8MY+o17kqzZrcrRbaoEuMeyZMMq6nmFCCrvQjdaOhmCehWdv5
snWAIMHVcQ5JvqYD2ySLsuMmT7Jcj2Mg7bZA/ZMcq4vFfwgAGDkaC7gHsR4yEx+Y
9hn4RRmpXv/8xRuF98WkQpIcjtrBs2NzadnAnjHzulIDtRErEe/HlGkhTrm2e+g/
yPYZhOw8mGoH+7EDsNDamCFYb2F60qS7MgwcE4KUh7N1vJuEsrlohKBfRJl85tc9
IrOCuU3+Do+ayn3w+K4CENLdjMWvcjQXxkmzGjXnbUvSLyWT2cAZjv1DhDD2ZYgg
cjyPZCF4vBlqu6QHOci0q7xEKtO+sukDtEswvvHOXsmHZiRMFdBCe+sK3Lh6v+BK
aCyq95yghH0f3H+Ana62aoBaBRpwfMmGHJR/BoPhDbw+bab5CY/gLcbG5EuxY0MT
SEq52LJIDNVCxyUigJAq2De79aZsoI5JlVUaFS4pCroQ40+YiNC31HpNS/h26sWU
JeiSuB0f/aUa9bRhss+s6SMYXqombZrW5xUZZkX6L+joU1Wu+lYGKNONW4l8IjUa
Pto95w5isHtCeyRjIsGVo9aLPl1UZj8+5PBf9SdDDrCml9MjWwY2WUY5IcEOBz7F
UzHsOvrKjbzyHT8IfAEzNxqYN5SC8XKCx0j1u23Fr5O256H6IdphkwzZednwdFVP
M4hjfYxUEHTgxahOQbnOlksmqgXvvgTDF1SGBGNweqxjQxSqfrgdeWS6k1L8Y1H+
5HGUjGEehPkKfQcnfs5chi6IrTT+OuOPV3F1XKpS0oobBKKjVIpM9yprnPUdoqC/
UhLXwHICGoJY1+ypHZ1PP7oI81O8YAdMBoLH06A540cgP5IKPw8nSAYKNnTQusSL
rN93hXprtGlyLjWcs+WyauZp5VsLLYXfniHCKylWkKnHYFjl9woI9WnjuNDkAH5W
Ba/+MpNYNghgO4DTApLefq0r0f7P9/MAOafDZWcyoucLlaPyCk0iHRn9EF0qGN70
NBHg9vupgJCza9fOixgTSmFhTHaPywj7qL3Ia8C7loSGi2BUan6ZDuYK5gyuD5PF
hdeoUQ5x2x02F5XtuP4XE3q9xxwAKoICZuWyeY+sr09RGofpbDVIuiKaV6NMTH8k
R1BrV/Q/zBtKb6TkgOCdBRay2mr9wmZqA9WPXlpsSavsyIHte09Q+e09FJ7t77Rc
P3w/4AFuraZ1c8At9ofnEJogkqldkukwzsOcmtglGDQ9Axr8p0FWS7ZJoeq0fMoA
Jwi5wFNfl/vhmqpkAIIRAQltQo/apxD9fo2qmqGtjDtTFMDsZPHV03nUO6wbmZMN
bYzw03n8THdk9Ukh2qO3TgWylrEINkTGEgLt5y6BtoOyaNsOosBTLp6HmE2QbDfY
1F+XFYB/MPloa4K4tbV06NpoxRt8ohyFVmFwYZmbX/iIfe4ja2CStPlPt8bln3C6
fnEy9fIYTWM/TtQ+GAjnnjCKUvX6Cbx+21USzsu/R1cGcFhqdO8XZmy9QD5+vIFH
+BvzyVi/mOilp0xPc2ZnZz8BH7eeEhnj3Zr/khRTiocINgHsJFyKPj6w1kVrAWlY
vbmp7HN9OvNg5R7Dkmu+EeYnVY18oB+e52MLkXALX1QM/Zfv/cN7mUNQoOVLK36I
Pj0aPoUAbhuIHQKpgNdj5IYEq0b8h+PkCM2pBP/L3Qg3+gPKqov5ChhvQOtQvSy2
KmSQRqvREXekns9oekoq1Z4pUHWWJlDNa7VKPX5TwWF69OCzMuB1QvW6jLvbMWap
FtbXuzFh9o+T70auJBaz3KaFjcL0LVk2LYOwbaGZIkJhzNIpniO7GezyBTkNGkLv
9XrCqaGdD7KIQOs/vYbfosuKPNBVtEBoBfycKwjOCgBLpsNrOg1VrW4mxK7Uxo/U
KqcCj40hEJQi9TzTfejF0VqVlWMID09LDe9JYTs3Vl06a0xT9y5gbIAKZnZvWdmS
a5X9f+jDuRbjse2XfV/8CAOiyYUkZMaPDc6WuM0Fp80V+84FTVnyUxwS+z7Cfy4H
MZNTSAw6gZSIODcoHmw9WBK97LcOEDdW70k1Q+ePTAuD+ZKnhyekDUaokymKMtTd
e3cJ0ecbBjxBn9IhekFfpCPaeFNuGDyRFexezJpGG2B39zUstSUdnpdU64Rk2B8M
G6YVOO5Jbt4kEVn0ilB7JX7C/aAHpTbJ6mMwZIkp5rkOXKXajj1c5YrIGNuX9b4I
/A8sL650YPCqA9PnQpgPKZpsAD+cnfmmSJkLDy+hkaWkySTPl6t2q7TMY6Fuhfld
J0QCPalJ6VPh/ifjWr72XIX1o9UT+jbwJKhA0GT3B5QMPjlVy7QliP1Qiv7n7TEG
L5zEPrvajwJlHt4M5miOnUwhYidPz3lb4E8ASNnmXSxmWEGT0GhWCgCFa1vRpSdY
dV8Os5ac5RTG1DxU1WYHzQjT4yNYaIe8lv85LsRBa8pImy2fTUNHJKdo7/eDpMRs
g1pab/KOC59HNCOxcjdoysx+pOapUy4SkfGXDOU+YsYIEntcRXZEgHaBQec3twWV
4OgvZ9L6TEwUyb4nPZ9RAsXg5/e/SiJev/j8rSRRyHDgGyB0L9m/iIilVjRf3mZo
xTYltl0zy+Nb1v125cnTrPGnAXAJraHU1AWkHu5pTQQOOsXwBBa3P4C6IzCbW5MF
QpdZVZ8KzlU1UV0JwAFUE1h1G+ooZtnjkWhVpafD95gJOD6HwJe9gpfUr8c1ysgF
TfJgZrY3BZY9iRjhH1NiwqgnZa3Dj6Mst9ICZkHvAstXwkh28I7M9ssBvutXtNRY
Cnwhti9JzEEimurpWlctDxO+w5lGFH7iBT7+3mzN3KVAWsL92V6Ap1YiEra3X7oJ
fGxDZfAIKXBhXvCoR8GShGUHAt1U44y6RDbSKYDI/t1ywDtN85bgHrXpAbN2B1ov
+xpEYYICBL4sdE+I4z0X2Ep1pbB2gXehLb8W+94ynAAA41JQka15izJUpTLWpKOM
JHBuD653TFDcc40IHj6WfQKskR2gTF2Xo075nQzca01umx1+4H9k4axKTno1Q5j4
4q+XP7bnoFxFNDDFcIB5UZ3fzkc0BNqL1D/xh5s3Oan9dyrEVJhYjEVe5eOegNgt
xukjtHMvd9wtGBR2yh86DQkWX7+wiYdeQUw+ytTbZfX0mjiWQ8acezIQZDF4UuOE
Mj7lyzQ/XpeBDuCCMArIbE2Lkg9NY1Uw2sC8TLwzSCLAaWzssdKN8XY/RbPBJ6PJ
E6BaA/KBcakks0Y0geU3v8lDk5tI/CRxQm1bFHFZoSyUyDCx7iIQXuvwtl17D2C8
xcju5bdVjvsDVS7IrIPPiZjVknTQSOTwXtgxvrtByMM6PviVQT9pZy6/s2KTKUW7
fDPGxm3PkZIC7IR9omj3XkYa54zo3V0hewbBymKFHb4tA6U5S5RDu96lgZFQynES
tNdpZ2ue94yWU/gGxQKhtFROSBHfayxgfY+EhGbo1bGicxMXOr+/VQCDKphGIm2H
zQ46NwRNXGCRYD4srRtd9cZKKmtJbfwJ4pVT6rbXWuOMG63CrXRRdobkRNrchFDJ
5vH5ZcGlcNtIQFDJPzLq6RMufWntMrBzhD6dyGOrFFo7nbwHPVFb/0hraFdCAZ/U
1LL4+x41708kzbHgzKCsH4SOROTPojx8z+o9XJJxRxJkwUmfwv2rqN9L/Y6+lzD+
6/2m6SkD5N0FOoRaPvskfuPyKYlr4GwUuN+Mp0Q9A8el5mNqxw3ZMgQ6JYoC1HTG
O3GbHZHTD/MJrDzVWDgGSZIIlk/NZERKeMFNdGCXNhruKw854Nw/KGIQWzs5GLU2
KiLmxLrTHk1wsfITSLduLnjjGocT/VNW96RvoL2DlRC34M3C5GN2E1/FZoUklMC0
0lXHf12VInBFAFyyLvTRU09t0TdFUjJ5oMgxcL4TilTS4A5pxJ/7IhFk+t5lVsLT
wDzw7+N5D5Z8mpnDzl9IJeMD/5ep2gCkc0uJQrE/zbso72YNQc0ppOOkizgPSDy3
rm0sjYNWSQ3yRQ2N4uyZVRYX47SB0WzT5o3wTrNgFgNO7EZ+DWEfUnqL6+AEuUXU
iIGNOprGJHqqXa6f7RaP/HM6MEyxCA0Chb051D0M8mHMT0jCIDl2FX2hCkHNpo1E
KmKGhWfqV2eB6B5fPnHuE6AoRU57AU5+T8OpoeAbURRv4Wb3448f+tihLd+tiUfZ
O/du0qkIxdzxUyBsVK6HPMyUTdWAs6uj3LqQd6G91fUaR0gJhYt8MZm8eKuXHROk
Hu1NrJI61AfCtFOiIWmtjsImd+Eh+lJu22A1oEcvTRzbGp3/eCSkyTauPEo0yxL3
OlSb1gQMCPmuyWYCMf25qsdgb8Qvq5Q7NchpbjycTJByG9cjrX67qG3jijE7WYyh
lgJ+n1EDscgDEnvd0qrHM9uDI6guisjgPQ/xTW+OwSDiZou90IL8UN2s+/q3IBR2
PRyn6lbc41BJTGqNh/veNVPzO81MaSGPPfmE977WWjDbY1ctQ4TfIAz3uwTm9vm9
j4Rudg5rWWFFC4+Kq0ZC/3XZSetwkn26jyPGrFFljChPK+pmkXnUNANZFWrm5M7m
EpJX7HHf5RasUekxqFGc1z0ekkEr+ED1fa/eX7FuKCyIRG5K81ZeyWhLnOsqraRF
XhtRJQumfmPWHmqo1eImm8Ll1Qz0oVh9UB0lr1sxFq5OWTYiKDVwTmWz3ZZqcDYw
mo28ZDs4RW4pkCwHS8PH9KfJ9ih+CesEFkNeyiOggCpq77uz3UagQQpqhigAa9GH
T0ioytm0r9EYtk2dWqFt/vX8aXN3SQ5Yq7Rbv1SvsKYtuAyCHJ5cmu/Yb3thgmmr
Hn+mfRy7gTEErU6hf1bRGGyfAYTCIyWAk8b2SA2zfhedVSFfITjBVjhUf0tOm7RD
V2NrvT8z3WRWl2D/zjFJT103V6ZBPtyDLpKd/g5Pyh0+TpLS6AI7Typ+Ds8RIPKY
yUNKSbWL9m2fNMCYqT43bGlSaau+2YQHieOqxM3pyc6L46A1AMylKCElfuT0nDO4
9ybNyj9HUocNRYcLEXByx4e6mjwN2wKtllVa2VDbzwE+TtJOZh8qNTwIRqSeyt2v
B/niqybL7mr863JylXGpXt5UbkgRaDnJYrvqgns08YnsX/yRL9Wxdvl+pvk9Eg4e
2LIDVgBqVucRDfI0+aGHfTS5ODntV1cDetyYTXgaL61dA6copLTjmyZbo6eTLcGM
DstlAkUW30X799yT6F4/6rLrxkpgkJUfFair5RkC+x7drHUm0E9NX1y8ElMQ7eyo
jrCimL8dNoE8Whv5t6PE/Y2vwk88lPRQsjyZQWuulhUKy0RLi4tFmzt+W1sBnS2V
DeUOIaJ6Q1pTXhM9t7gMU50xp1FlpKrm8h+kRPuZnbjXqhCXRMY7N1meBIEjRKrE
omyr9xUWg/WQkfMJF+BKyVkLxA+q/tLbTvlknzwDSZCuwpxxmfYOJxTqONLMZkbC
hYUW/0fjo0tcFMyok8TMccyvr5oXExhZP2RCvio1VsHARGzLUa08LCAoZexj8lIx
7oM8CCQ14W+sN3A+W4Ho3qqctz4MsbtCFw+BEPwmIhH7Wi1sCrNcz/ZDH87nIDWh
ri6AKe/kT+/A/keCF4anwZCch8JD2CFLK8OczJkfNYh8qtUDRnkgD+9vLAfVWadX
PE8e/tk4i6sPqJtLfe1krpnRWllFOHj6cJgGzu5Xw4SitL9t8nTDVZxKrt0H60Bw
bfD1TG5YI/3+6PpHyp5iXKSIZXPH5HUcbJw2NeZy1IJhDskY2tFoGdlp7KTxeHun
fxR5BijJT3dImpOaOxDp3PhSktV+INuhYCasDbUL8dqQFwLr8gb02Tijur4b5Hf0
VZQAB1I0uKdijDhjY5dQ6X1/3iP0ZXxTZjfMjZg/3Y1avDepnB3wk3kUeCctyeKN
XbBEwdbT21ICE8waYoRnhfrxCyERy+wfMIRB3wuqoID+G5SNnqjCMOa8rrN1XAcF
gqrYYb8dvWQR0syxOFlWdMiFbfWNpGPQkaGQiO+F0wKMEToiYZh1LabUQMxG6xq9
R5v3kSvb+tuX5u+UPQ3rYgNzzc52ms9XmiIc13JFzgwMOrK3RNI6uVpbqvZkB6ZQ
YXXCj2FvoUEZ4j2Huiajo1fD4jNlFWAEKNX+TeTJVka/o0Y41oDfl13IiOCOThAY
Ctyo7vVCEinI8DMDaJVCstL62lA3OFo9bpekFnFC32SSice2jzsQ+UInZ4Oeimgo
nWRWtP+eKoWjWrAviZiRBS8WJfSoax4zY1qTUjaaVRwkOpXI6V39SZta31edpp5s
jpaD4S2OigV66q4BtNyeL6oCk02glF5qd0GW40CpfoY/NNHeCZQMDdQn/00RlC4Y
MiS34602Lr4pWVNiZCU/wo29pMvYLxfMQNbnOP+db9usp2vG373HVD9IuIvcqStd
XgwOqdbiZsM3dUCQjNTr3xcReTkwStQqVFVjoZTvQ08qHfAwQ+CBZ1qwmDXNCX+V
EJ8aZBmFReEGLRfK0d0fAjmjvBSl0EbKQ2Tug6LLZ5fhaES9905RT2FMQIzmuDhV
zXRZz02MS51hxWvG+ICxvjGuJ4+KuF244Fis/V6HazHUq0aYweYPm+EyQW2mayYf
Sq8Vc0TLDXbBieL8XqZ1XK6PVPLqyj5XqswQNbbY82YUgGHJVC0WFAvVLPalZxvZ
7gaSO/Rf9FHsBsWx7NJmtOFXc+XINpu8JAD+XZPjsNh73FX607E/fueKAdmaIdZK
fzukdvK4GPoSYzcEU45BWzL8vZOQBO2X3pYF7/N7pt3G0NyAC9XOhqcFWrXRB1Vs
AI7iby40LZ0eVDU7Yh6LVkQkmTgj45PhqaY+UQLHSIQucLckhfVDoJHCUkPqEZG2
OqV1+ycM1zN9mMyiwG14CKaCJODWkjcsJHy2bwmTPm/2Zp3jbaiOapkn2M/kY+Ni
dipxSW7xp2jCD94o/f4yRPlg7b9oy8PVM+w91R5313FHGh+ITlLBalODQuJ/d7W1
Kt0FpPIImyOtstjeAghDrfIiy3PRo83fMAJsFvml1CJ54lYFt0nuGPPH2nOuKTsO
RrZNpM89xg9JC2EXDM/7A0zOkILgmCAP7Wz9FS4JzFyjY/6uIIoepqskp2GBtZj5
x+gBP8qTanKj8wDOmKFgQIdnJQ25h654SWTQw7bhL6QMv7Zj8a/KV8MrvSedRryP
H24h5gE+8FonFZ1UYdyfRT71hnz+9ZCFSB5Jpkv/uUSfqiIuA7lZNht9nMKXUcr+
u7kvb4+sh5Mjo0OOYbQ/AojaypU7LFEW635KsOthyoj1rdtNMgBigTNJ2YkIj5n5
x/ZokittZVjp+JUFjpm/k2hf5DO3TF6+nRp10ItnMxRtMz1leGHwhaeQtELf3AZw
GNyTjw9yikirbQbsCDOXQnvoR0j3oB0S6pX3iTo7mpbIJDoRrWWCvi7gZlrv0MW+
Hzv7rJb5ZhY52C80TzCFIVTAKZeB10SSgReR1sPQX83+5BSbKFvVuT88D8QevJkD
i/GW8jY+kB+4zx7w73ZF4E4nUpQ7p/rtrf6rDybrol+QH9br/YSs/0PH37x16Uqz
FcYG+OPQcLYgAFGi4z8bdN5UGZ5HKaYtZ5osq8iow4EJ6i58XvIdvwz/LE6K9Kz7
B6LjQR+hX3jmVbo6LnBh98GcdjLJdmGJ1YZfEREUITq3WicLVZpthOdnRU3FEBSD
S0Ehz2TXV2gMbkUj+X2TN01uK2AWdEkuWYtPq+Mk6UGMQHZZ3fBco448ZMzfqDdu
QmJJRyU+qZqGH/SWwiRVosc1Or8HszadBzONJGqHFlXORzflUKj8eFCajM5eRsD/
lBrX+PJr1R/W3lhYMOw+gMi04MxrtZ5Fp5lb4StxLAsfRFwSZtRUCw/o3hTsED4N
sFmKSnGjlALZt8hdxRj14LBUel31TY6M0urSuw40gJWZCruHee84UtfoSXtqw48I
m30GPWQq945OqmKb1C6v5i6RkTQwcjS3Yqw6yRxzy90zCkIWtMMw0dk41cdg/F22
3kClnlImVbc9t7VgI4mBaeLAk5Ye5lxE2gOZ5KTiX4z55YKoqXOEAWtTaBKUzNu4
WLOEd5u9DhNYWeLeljnpBy35Ytve9gQSxZYfPFV+OPcKy819df8uGqRnO0Wv6mYT
BBLkg8WBn2WKHFawUIT8z2doQyEKfR2qJWjpuhycQ1UDzcr7HSflCzyF8/XJmJae
PFnK3xc7MKp2OB+etb+l8PglHuqkkINWwJvTzV8P7lLg9IKLLkgYBGXbNn1WH20X
rWPpWd8P5H8ko4Uqy8UC0WbAuJ0EQLDPLc9I6I7onaIOAvCYsHubQIT4OL5kOQVk
DoGfy2cVwd3qsrdJCvhOAl0wyuvb/6SMtyfTAJMr/6UCU+eaad1YKvsEYmPnr7EB
jcUY27D4+ssa0q/jeeWzVjyVe/SsUpssSCYQLpn2OaSCKo4GCTPbbPGGUtPk14d2
CSXSj4y6JwvB7LCG2MOZbpNM3vuXohTA2J6nX/GOTqNk6/yMef4BTYAd1nyRvtHH
WUZjJzlrw98g5AK6fVzeE7VNEub4dtN0L01SjxJmMklPNw3yE8z7RxX9eahLZLwe
Rrg83gUei8qzj0gf6JwBXMxT7RJ1wSrFBj7n/USlZj4J1WegP40A5CJ/tu9j6AXJ
f1zRHDeCSKKU/Bj2iYC0HeE7RBmN1aq/8zlL+ZaHuJyKBPpFbamergMO2VsuBrzM
v3ytxHdpD/ga5UAtzUb51yOB9cZupSrlL8Nc1OZn6PsQqUwasZgN7PdJ9Ek6lIP4
jZ7HyIjqSS3oChyCsUL5r5vaBlMKKqYCiDCvqRamfXNfLaI0sCJ1SUIKSwGRCF/o
hCT8p7HZvGdPvkfmyfC3h4kcvp4nbg34SFKYC7tELw0ULDJznjkFcNej7gU2BXVA
YhbzjDgHGra1VfLu9EffqpBqeDE9wZzmZgyHd/ek5eA6i209bNujLZ9tpWZHhY1k
tZCzx4EM5PdREc4dX30Y0YE1toP0gm5cL+BmnAO8nr7FYGarVYv3VfZbJ6T4TN+/
taIBwUFSW42nb4SV1yZcqnHutfEbkX1lSpbGdkBGXHEP8KLP89i1WYntWnsQYDqg
xQKBEqq8lFwGGXeWpsdeLvtD1fnrKweyQY86BVOKLGsJcp7ekXosJXr9LD8/v8el
nImG7axVbWpPGiiaR1Ni4EUyTau7g76+CRa7rAylcXJGK5cNJSBRDNKTDp0/RpZq
h4DHTi5kT5+WEK7w+Qv8Z40szizyz8vG+Y0rFp6SB5j9NUFcIKQVROUxZHzxv3TS
W7PPdkNxVGLOyb4MspUy7Xz3kfFL2mHwHsIIHAkt4Vtx5YSPEWfle0c0XP3xURWw
UQ7e8Gpjp9Y84gQrPcUhmWXO/JnkVxpXYkQXnGZ9C2Ha0sxlo6nTSOS7XCCAxw87
NvLXg1K9QQXhdAgV6vnesbenE6wp0Cn0YU1urQNvQSHuz89JN2BumEao46UzM2jT
/2Dtc9z0qHiCA3zGha+KGq7wA58gqCyZch99UPx81GFaKUZC7CSkLF/eoLa4J4pZ
jfmzrU7s0PQUxan/hTxn+FVatUbCZpdhqD7Hc3m64p26AUPcLXJmld8cNHpFR2vG
VSAqdUHO7gzni9Fc9OCXalRaIuy/sVV7ooKN8SJV2oq5PTd4p3HEaVa4Oclh0oLb
weH3iQSKlJZ97lJwF1Q0qcSqHAxBUiFv5VlOW2tB3MElTjWcyfbmeTdsmFWzAPpP
HCcVe5ndd/r/pWljP1iZXkF7OcvcUHee1QBZ0rWKjgXYpKKwnwFwa3PCzcTX+92E
6hlHO/FW7rLHBfm0SNybSd2vvzgz6U+b+52dJ+kZsY+vruqVEWgLzPeB3ULpvtLP
vQmI4vI1ADH0uk+kSUoA9jPFjV0Q6IWouYZLKlr2ZwsJliO8Zo+tjQGQv1GPpvii
mGyqvqh0/vIjOC9A7qG23+rfq+9QrMoaIJDdhgNef5FIN/9gC7ca+H66P8GeLi+U
FtCpLOp9Rynvut6OFg/b48TQJERW7SuvgRSg1GxF2ypWfMkkXzbsi7+kF/dgWL3H
hSfU71y/U0JJdN/1Dy1KUkXVRM1c7YBb4UuASBfwBPPf3tATfDj7FaAUSshHcTAl
rX9tZGOo/eoUQaal/j7uKFSa7YYF0Z9T3v2FuqgfyeuFQ/WVf6hL1PPOHW83vX6W
ComuKOs/HPa2qjJz0s3LCHOAZcIwx1IiNQL9UDj9rhJx/a6ylSfft0YNdMU1skaI
UarfwULb/s9xaBIV99stgcYgSSK0yeZsVV1t/yaxmrgYDgFn/9PLG47QsY5DVmpM
lpjczmC0zw+0q8K9K25CXc/GfNxLu3uxtXwPSxurPYIsfKREBIMp/N44G46PHT8d
Wl8CXYj49wOICHUmLNl6GBjCXghbD7Zq+3Zr5dscB5DPMIsUkMUiip4TlYbYiEBk
gZncyngscpE/EqegJNbMs/K+Y99/Si1yIWn2AP4/KwIKXohsFYYy0NUfIPXryVtm
Hr+cXr6OFSTCzOciLmr1fYUm5RxzDMbeRGIJzZtJsykmP+wh0tR4VpAEA/3qXnCw
ir15Ju7frLdmfrsoLaMJHTyiTuCad9OzEwnhhXFLDxoudSBfD26WtC5qlMX044Tq
WRxeJxPOXoroZ7qZV/F2OxdaxUzJhHWVIxCPdULrfPogHacGsYI0UgSyPW+sWJB8
+slcc8lZ6d8dgiM42C1YYbZJWJPLomBIa3gupZXRjI2k3rmVW9d9bnt9PXLfL4s8
+XRWOR814R+i5Aosu0XWk3vhUTjwH5RNFDB+IbNxs/subYksofUAqXMVVVayqxHa
NwzcwMNVys8GFZxacufyuuHVa+d4n77zj0Ta7POYoijVzMcq1bpqTo7eBcK91V0r
QZvBSgVgHVhwfkARrIq/1tISCqU2GKvOTmTEStd3XDl3Y9fJfFYp7PBmRoxw5xuo
vEsp16n4UQ8lFywI3fv87lNLxo5rXAIh0LWjPt069JWcTuJXOJOQEVdDKSJjPzr0
Mvy2ZHn74A7pGLsRXsGZD+VdnnoUlxSgvM0d5KkcP/OLcCTs7GVeB5Wd/OQ6wXqh
LpdahuPwrIxr1Ts+7RIDR/zmYwfMqBTUi/lydMoCiFGcIET2JBOsktndnUlKxJzo
esz854Mhbkf9Ah4QaNaHxi0T4PoxpurSvqG9LAXqrjk7mVwDQBmWWw/gP37prsnJ
FaQOinsckT2s+tLoaYQCKSePtlWRWpE4sCwmG1NeA4csrGwH2AYUdDa2BoTrRkyB
wcA78j+vSUzR+9O6BZ97JJ8HXyKnMYD7H/5XtqX86eEcKSZH1x3SjqvzRcPubi1S
SO/xtYMBb0kSK2TkRlv/d+OZ7+8AK9nob76wTLvWD8OKI3WszqSTIfvkaFl5aUC1
Eppxm5n6i6QFW4M9ckaEAwLKPO02Qb2mdZBAyljrDQpq2TejCgHiFaFI+cl0DLgi
tyZeUXykz2ISjjd3JqbfbiAjm58R2PITaQdk9jaTNBNN1tJaPscZi0QymzkMB/ks
72G36XXFmyLrrkdEiUNvdTjX0FMqhtGu3J+O2NagmuWTLHSPJY/cM0B2V0oygKre
4f1S+jJLvFdWVwDX95bsgU5frCPKVCOyTD+ReHL6X0BDwsvz9hr6eg1vWNCmNBmj
v9Zmia1De9S9G1y1nGVvMh3BJk8KX+LapKltGMTozDBW3eECVFq3MsohCn2nVJnD
rd6kw/SBGRt7sGgqgI+rbkApHG4u/h979lDkNKnbyl4WRAOaU5Ld/q595IERVuMt
dhvk/uEjycfvoWl6fTM6DNne/JsYy56CE6dpPxUVq6q+fCVbBbTarX9qZRNTOncW
bOJEm4IrHoc4dK6+niwcvnTg2iaEGqZLkoRDcWgDqUIvMU+rmIhP90yERkCw0iAO
j58053Ttx33c69C5+Nj+1ddWrt2Ttxoc2W0HECJNOo3JKzTSXCQma9FN5a+fp3vM
T0sdt4PoxXCeQVaRuDQlJHoJXHQuuRykIcGwWB70ptUNcDTyGegRopH73fJlJG8v
7yF9v3I0LTgKUS4cGMbnh4JdYZTGb07wA88ZNt0ieKFxQC2rfF8tqTV1M0j+IUsh
U8Hs+O6peQ0i/l2JI3ScmtYYVWG/9Ux7E6WpAwAQD5DWMPyZzEDwZSPRJU+GCusG
pxNPK2QPz2AUk524dI0uSRJpJP6U3yTpkfqRul9dLEYXK96MJuldNlFh423Ymyi7
RkQZSAO21+5j8qTC4SzFeVG7RxlTein7cQ1cmBHnHUcIdEx4Mj559EqKacORonbW
H+DTSmwZz+HEE/bJtBeJr90k40lgV7b3QFuOj0ynaS5BX7YK20v1gwzibx4A5h+i
G+1pB9NkdFSgCmn86MtXBrQvDhtIRsMw12EC0KUbjf/3g/s9Ly7vAoNi2xdLd9Jh
QGWyS/yMt7UmupjCHnuaSn+OKoBREqdNer2aCGYqARpo/TaEls9FNDVwmAdepCi2
sgx7K2FidxIJFgeBZkWhboAqQ647yLJhscBNVCYyB8bu0T4NRXdGs1HU6+6UNxmw
26Zfm/B8WZ9cPFAhdTfcA4NJmdlVuGBTco+4bnBOVxYYXYZoNNhd9yrIauP5OS22
26+r8cfH3Q6gC6Wma9b3kCj+seFt7XIxgFP/6yjwvybms+BA9oMvXzBdYS4/o0L1
xE6XbO1D2cpBTghQdhJAYdZ5LleLOFjXcBjtwjwd67Oo1SWae73YqeKamPHNj4bU
zMXtkYneZq7nogLR3JgzgZjF/cgMlrpki8TD+P05rtOa3dTPNbzw8SNRuH6xSnNW
F+LK+jEcZrYteGFY0AhdvV0ptcWvDKFGNnt2rIkkPb7hSHGYCKt1qYLl6mR8ucQN
uWScB2a+sOx6VePxYCBswJhI3Yfi31uiuVPIAdLUgpazyHG8g3DxvA0Yks38omDE
YgFGa/HuELgOADIbf1cKcojfrpWuIIiYyN5XthcNJtbzBK7f3WxZZwfywpSRT8d4
sbUHxIKFbmsR4l9DbjUru5OOMH91KqPbhTmbgtHdXgPJi5hHz8jYY46K1QhgUbPc
53oEVnGRSotMbndThTiapr+ZVlzcPvMCoRJmdCIMd2jSOL3XuTQh79uwF/0XitLP
xhPdo9vTr7XxqaYJhXNvVx7KhXq3ulgBbyCS2rK24cR2MHwSku0yZgdU90K9Lil6
E4DBdndzICLkjlIcbmMIax0Aowb+NF14Q3DXWiP5CAW4i57+rBqwrFM0jDz+TwvM
Do9JJszTnyaSPt+YThE/Fv+jsIdKt7AYtPEV0ZEk8ZR2esqYH+sEBvPIUrvglJEA
XxdrszfHOpvtIb+WscZg6acMPYo7z/By0lk0mjiBQaDRivRNe26nht10yXv7mZp/
lIqsm7uifAtQXW6uvKQlKEYaeSXL5pT/Gvd/5wKEluEqeYKVGoEXLFMEVKiRqThj
LJr1ZBNLsucyTt63qNmrlEwUMXrHnJ0+W6aBBFjOh5ld905ybXKEcUSs4WBscMfz
PIGe2g3IRYVigDhA49T0fHXFwqbfKlzH8DFhvx3lKGM4DvEmfufh5evYoB3+mwld
nfaUe7QrHjMQMj8in0iIvVL8UnyzNZzXhfPDF3IIiHD9qdc3foNwm6aQDtjsYbtt
J2gS+7lrwLrFSDi0prVJEuILo6NsCnn1j+ZmBryNQrmb4/84XbreVPoZ0J/hVVxs
qzEes9F5QrE7kuThNuXRM72UEhx5UMK/+8cYTj3Qqq1ebQMHqyji4n+ykRQspkNz
CL3/6KDanK1HlMya6LWQSuJdRsEToV176cPEnch8h63gigIOF0Qcl93cF42UuxbI
KqhmxY/pcQ+icOd+EIxmEL0jloJuLG8jRkjtB6EXA8NvYNEXlMPcS71V8BvmggCN
zhJDZZcBsLqQHCxcAEEh6UZQGdU2sK5WTHZN1xv/iKrk5A44hHHbwnzsYOsDMoUd
zKxgshYaQXFxLbb/Qgnzi7KCK57IgXMslAaY5t3sWSL0uNN+m+NH87gyXvM0BHeB
4E/VTVa8MwwuZgc3RTxYnOjVBi5XTGVtlZaKFtdDmWmWrbFFcu7NtRkphzu7qHCe
18/ogYXTJio6HyAER43ZMAX7Mqw8f3QmFx3sNGIOKBs88sfU9h0xtaye3DlJkSos
jVIKT4iso99tGU8HC+K2hCujG+74PBjlJqp5NlK9Kkxoy28fVpK+XGgTgpsz33YQ
txw4G4WolU6Y0w2xHswVqfe/XKPkyaniPx9prYW/3r+hn3o1fBhH8TVwaTyvQjt2
PTCuHlhCLAAH4eQ9BY4jsbtoKXeuO+A81sXdI+pER9bJH9M8GayaCEH/TUkX4l9u
Lq4jw6Ea/zsfX8hQpVvite0rYOP0fsSfmKknz3Fy/rqeuzuN7+ZDhOuVe6Qx0t5q
xQ0hHcE8XLAV9ecI84A6vJpjyNuXbpuu4v4qeS4LbPoJoZJx+xpM+H8p3uYjUUGZ
8otwcyqdKtaMa3WYXBhy4/Q9/FcYXKY7//ASbCt6aS4S7TD2XkkPvA0cHGP4fDTD
fdcRG9+LLhqtPMnwCXNoieLcNSdgW4XfEmnLAjkOa7G20eabcEeGCsoLtmmXDxZH
JyIwym9RW27Nt+ObJa0mteCNFowF0RZZm2Z69i4upYHsy5hQ3qdXC+yGMT54KrfC
F77MsRceazLjbn+8cGvZ+mdzz4BZHm/3d/DRUXKX2PVlhBhEGKFcR7lFsZMPzWhA
yQTN8UbEWOfZtqtn4Y7WPtHKigJ4CWtwNXPYBvbYulJ5CsWsYjkxvFjXcCYDa4FL
olZZigYpQ6luUI7qTjZLzPCfIOQrG3aGwKYm6R3dD3Ck04ljIBYcl+Xc+CFzsAtr
tQ6GKJS0tXOczJRpYZPWfwNwGgSO/TcL8Xx1lqOJ9EzSCND0pjR+KyJd+ldj/6np
WzyLfv8KvKd91a6giiPMmkbrGVwvFnM88UYhvodcSmkfHtPwi0oBOrcCDgQti7N6
8D6A1tEPW97qwz11WMm65gB//4VFCAYT/tRtUxcQAmLVQMFaDOyCPK92o1iipmv9
nuUcjCK6I79L9f2+1tj3jjxmKhFT/zb3sFINoy7WgKL3JvaxiQhtBC1L6hdFOMps
+sH9Pe3OBC4V3DpPc9byhYYxWXVhA47zfMVvi2/uGiQzImsY+DG3B32klrYXJbih
N58GTt1la9vLEhUy6ZMoguJCMol+WAirvNvhzgmWRbKQKiw4qnMO7Y9uHPShSlRn
TMYHXbW9MNE9+sR5PO54QjF/AXPReFS2nVnAY09ZEgO9P44YZnEIiqrblWyuf8KM
L95EJjDBjnyPV0QeW7Dp87fo+meR/qJIcINXdLQTuEJwWfdakOPfcntipeBoIdvJ
vdjDZrRq1QKoxQ+sbU17fdD+HFAIVWLoHrZXQgqXXLdTdlMAJgJFqp4ltREBTwmV
3PnCCiOm6F4ciuTEhbZMOxfVwyKkSemkZlVdl7N4HEjY9xrw1qbE+rM3nMpwtHC8
7/bLeuF63uQe6U83IpupxcoGPfxPoIP5uL31j2KOIWEzmDu943Um/len/qR0ORrz
C4fLHYbjP3aWdzl4piIKNspKw6V+Z3RFIQtqiiljOGFb+2oeMC7WxbL+pNK/QKTq
R5bWMAsUKMlQ6JGV8v5F6X7REjZO1xgjuE+I6Q75wNUwnS4mfj4JI5qz1VH1strG
H0BIEAnn1esoQTliPS0Lbogu+ifM6PE3cPrUQgUXoenDAysVuX2dXPGcOadXdRLY
RInnd8DG8xaREI6iamqvQRLcxGL/bejfpGH8Y1KJosY7WASsvqMl8pH93fi2WG7H
yhV1hEdyiQItDxwgvZE2m/0ELk2UI6kaxkw6TWHMI7V+I7WFRxcxDQ1sJdg3WK+x
9/aS9SHCN1OaxC3cxLGphxYNhiQIKDONeaBNILx2nzHJW1Xa6LDmEM51Ey0Q/zXU
oSszEo5PEK4yz8uedM7tM7jh1DVKhh1x4nKghok08BMeRCMXa8ranWXbyYg9/tRc
pi5cB6Ks6Ynv0yKLpqWZn4fe0SqYC/6cG/1UJZ8vkHDfAXG9jlgBEjAKHy+INDFW
4yzUnDC+KdXJVyD+rF3/o7vIGx+Mt+4rgqKjMGuCIy0VUvc7FZtKaOKyzG/75uFG
D4a40XmlLQirPQAxKaRWCFb7+JgqodfHodSJCy9tMn/FBs/i54GPjbDFrEKwmHO2
3NrHBmN6AEc3I/Vfq8nW94hFHGKGc2sIKCUh6Zo+A9YePDvCqHzmL+T69JvIGEOS
jy9bZEqE4uWN9CMYKwj5TYViJ4WhHncVObgqnJv9RYKH+aR5+A2DHB8wxpl/jbMx
WZQ7FwprhBEqOYo43ZN+mx3l3BvXXuVidVzlG1dCa3RB+XvsrLOUUP+BPD4SlAoq
wYjsvE2GGejrCK3kwlTcWsTBnDNcxLw+mR3jPKHtVwPlZ+UF7YPW7VbX/kLo7beU
9msiANn9m1KnUgSYE6WlZl3t3NT2bL52fJITSSpoeMYLNA6VDRKGaNxC/XJOU2g+
1gJoPEYE74E1wCnZ226/pRUPWsItn24gAABdsnIFrNdUPkRtiyPMfCGDGsINAv62
aDpx0gFOdNLYa53Ni18vm5jIAp8eY2Q76fUXF/QFUTAJVaBybnTzDoGStmkxVIqu
9o+zvnqVaGESQ4r87HD43Tg+DlTJhVydiaWbm7T0c/yKH0j+QHP4DK0Wpk3Dri9L
0liZg3VLMsJR1TX3lJ7Hc3qSrqD5RjNEKhDDnpQ5k0pdiEgdJzahp0OG4FFlBAD1
7JFiU4b5VymKBxL76pIndwOKMEihCWMpt0tV9bCQYIyBOE547fqlKoaMLLsa3Yo+
7el9/Ud+yZTPQUKUPaoA/rj4C26o+qgy7Bktf15aHu42Lwv6HNoVNAUBckSkNDpl
RRrKryd1qeU/0XWTZyFZASeCZ/tCgcU+u0XA/Ww7yjUIpkJ6kjJOZptRoyZYJfxO
C8lQ9lJF/D1NuS4uWWjHm1mpQqWE1V0sGCc02nwI7VtUkbTBb6qAG9rnDVzphgcr
7TUYVFAivs5R1hPd8lnMI2/Lw6E6f7EWLSPKU8fQ+xm8po9IV10YTDWylCJ7Bn+Y
EVH9qIm44ksauZvyFn+VHRYVCSpC7sPGtFiMXmkkifi0x699A7GYNZXCSYTGPG2g
HygGJNLJlRAlghOOJ1a8ZWv1lp/Jjs1WEFq9NDV56i6VBwTePFnHF6cwW6mZ4YwU
cMNgIKXbzz9wDmPFffFaDuRX6r/OZGcC8B9uZwRIcTMioi2IwSmIyGQpGZF9Gemt
8N+swi45o2ndc8BqyxF945gxkKAzhaSihFZs3GQRE7wfFmnMW+zae2aQhi8Qo/D/
Itt5urZxX1PyH76tgX6KKdYYP3yP9xdq4cLjNW78rb+JDNN2s7g7DDqlkM9IbNlt
j7PqKfvQo7AdRRfemLxs/3kD6Sot0I5mGn/JkCBoJxsiT3QlgyFGkJi1xNjDGQRL
K7GFPfX/IfZ8nXPPGD2wDmwhy7kqyrbdq6yiIfViXO13whtp+m/OVlwZE6k1H2q2
duks1wmi74dXWLtHiOjhE2usigAfjgSyxX7V1dMS64HZw9RPEMLfz4xad5RE2ycj
xkgBenfHqwZRvF3cX+lRheOM9n3bb+r1BxVZGqEZ06ti83iU3APuU25dvgnk36dx
pNrbaqfeGYcZCZ0SfsY2NOpv3/UKYRBk8C6r5bD2nj7zLj26sRbYZ0xCgeKssBQK
jXOX3/3RufiMYGb/OTjU4Ju1eb/GDWJgCI3AdmHg5dx0L3arfmLd0gaWv+/jBubj
r8w4y7aunH/n3L7jpLT92YblApfmfHryhpd3sg3sN6RkxD7202DvegoalnWsliI7
t3XPSJTsOXQipmDNeCnJH7H+JiXQK5DP4r4dXqS7B6ejSqFTbz6SY44Z5hc30uHD
XxQpWmQqI9QkHRl0RhhP74Kg4BYez1r9P2AvN79jV+GOttXAa0TYdBA7SMxeXMbR
91IfwxqT9lDOvbM2vdUBOOEkutyCucc2eLP13c1iNXwaW1qYxKTuGqXiW8GmJq6T
ThcULFv7yrHcVTPdKB4mSzdTXDj902VR6QdZXJx09VVT8TJ9vkHWDPAqIkh+kZjc
BwSvNcYXZj9N42KdBBbfm7QN+evK0fvo4R9ghI0Su7rNQa3Ayn731e6L/fio7E/q
ChnDrnGm7TxBZOH4U22AWxFRFCzrDTtOTMKAeyZ0OK9s4LelUlUtv2Bl6ep1DBi/
nr2Pi7HhYszbNWAzhcs24XtY1fwYj77y2Qp1oXsiw/VA7zS7/oD/o8Po3n8uMHda
1bVLir9BHhaOrPilie4+PEFV8HF74sOtWEZMBAt8b7ZUJN9PqnDmiKLh2plprcUK
aWOyL3exHMiV7LNJ2/HHBC4AIc3jNMowHhLq+5OPKi0DX83qFUrNyN9jpuAqTtbh
48ORYp3uF+xgt9+eWtZoU8uVWFz/ZIH2o2ew8eoPJljTwhINGdIx9yo5inUFMWIp
AyZYfU/1nscpZd1mo8mzGM48Y87EQN55NkkH3qNWKmBxAycl5pvfs7WPkuWOnU8z
6d9Wy4bg4gHXMijgca2jsIhJpf6BCT24IkPdT0tGBPBtbmsNDOQUua3qi8uSJHCX
oequevCeqjvKJBYdAMGEpWPJgq784wEwNUpenLrnWARTmo8Vl3VBWrZZfwHJZMY+
bElTV+WWo5eOJkexZrpqlOiDGVx/CeOz/y8Ti550FAkU5wB/+zR5bsvgrQF4O0nE
J5nxaLHluM/mEtC1DM+DE3eaPwIs3AePuFf83kEhcvLs7prPrBuEmRf8nzaAXZnF
3LH4MXrHTK/NfOfAjaDSiZ3qO+cobcUz1FyNCouT1Rviy9uujlIevLlsxEhTsAu/
rUjl1kw/9gB3rkcQtkVQ5BsXrBt2j6/aOD7a0XZMWKPOmFBFI4T60wS21Une6TIz
t791sptTGsTld4Ni4RXV2QdZdG68Cgn7EKgZHYKtYbZAWjDb2Y7LVNpeZ3R95RPr
L7LlUXj4d8o0ww1py+VCLFMJbj5dcOm8EeQ52R5nORYjx+hboi4pV2WtlTXKuPgs
0kPdQbqcI6TuN0E074N0lneZv/qjhRs5UpwIlCW1sI5/k16Uf1lXDr21pobDe4nu
75sAFjVGdIGwEhrduD3TvOvR3D0xzE+f2/EjkhI8LVauAN4G/dfFzCDizn/fcyyZ
I/KSvupagbDSL2Tg0I8fKgopJViza8J51BYkH2cIV96aTkqSqmNvln2upoFr3gH4
kxOrkugWQGoRHLnI++5wqqfSKNMYRPawtBwIzN4ykLREfH/qsA2MoVQ0K05qNzYX
0JnbuEC5NKkL7e7y6yYht/YCVec9HVdGys2WtFb1zs7aSD4cxtMmpRZRZHHGIMP1
N9uvwzBYY1rs7k30ex/yCT5d/tP0igx7kNkIqnL0JxT1MPhP0ljQw7YeX7/4XoLy
nvbo94+ksCtap1EBubm055cbZFm84JpvJgF7MRo2tuzLmMzGwWSthKNeEk43KNJd
LPCceJ2o6BAhytNTqUFuC00APOLG6IgYbQkvMZzcK+s52RaKf35KmoFBCLGq4onA
2DvKOoDzytJ1NgYbcZEorjMl6jxcb5LKwfWbqDy0rZ1XhDP0WGE37QY3BRmF54ms
7ICPdmAw92jDZZbI0wnGCB93NnodmLzNBHWs6ug1abIh2XrUSYekYC23o2Wzvoaw
xCq/sfjWw3QwzlAGcGgPSU4eg7W7ryFF7OR/B/m0qlyKxHg3SLDvKs9GXfcTE1En
s6AJGxwuW4vZ+wevqFkRV5ZzSJ8Uwu3Z9bQ2yUJ2q/4LiVNfGE7sEEY12/OHXUY3
dIXlhb+kzb/0IEb2V2zB7pLYmD/bZ2/RTEtOMES+qY/fmO6BHvBQgeCGkBC2O43G
yOrRIkG1+rrSv+/ETniRyKEvtYBwig1mU2TanptxLG2eNU6yjXDHBXWc1NFj89Z1
t2/orbLH29OMjAemPDdyi+o4VmAB5e+wJo94sbtlF+zLDF099lEtvdVHeUpngQsy
yuZD3hZRgQxzsTRIBubthsU4lov8xoHKkVzFOPlotMeJXbMPLGlmf9BSbgU3qdv+
mC6qv0dou03rdY4EQ2GHWEwmOtuM0RRfihiXQhKOIZXngwEcVjXsDQwOXDZdgL+y
dNR/uZFEN85vQNaDlTZre3IWMLn78ZQp4ewrFJ1t+3AKjrvKt8Rb+rxSH4bRPx/w
2zXXn0U2PMntM426J39ejI6sRMR/hK4sjPI0XBOJPKVDoc/c5vdPSUxRVLbEbtuI
jqUEEl/s2ofP4C9Z0LR5Zoapx6m96Zkuvx/9y1Wq2AwIFhdD+UA9+1sbPys3302d
pQxkUsDvDZD+4jKBRe8PcK+JMPi149NosInHGVhmESG6oazSA3giuJQtah2UM8zw
pmGUBNKjdOCdIFndciSaLdyN9KwOld9xoWhcjFToVHlenjqipnhInd9TxvYJxjvk
ZJBERzYI+Yj2h4rrW4ZsY68HMgDOtVhRi5ZL8ABFqZPHP5aRmtt+Vej6fs/tn8sD
k+bdtKCg1WUeUDpxbKZF9DHxSaPSeoIpc09AE+08iIAZrJfAfVdOPyPeHqn9Wawb
eUmvktrUjl5ztg1kOYWjbYLPGPhlhL2mbDmShCUIul0nFqCK3AJGqOVZ8WkGprdL
GsKbBsc5tPYS0hgqXhEyVVFwGST5OHtr4hoND7NERqPffSOF9Qklrm3Kyr1oW6jN
XH24izxLu5xjQJ+sS15ZhGMnTTguI+CYb8IcDYJGnHXX2TTja2luMx5haeUASz0R
WyhR+8pyGQpwrL46Af+FTPF0z8b5YXdBkPEBIEQ4Rgt+qo1B/8Rt6/EPT72/0u42
IPg2tqFxDyOgJsaATKczYi7TuYSqlGp60N6lDQVemwqnHLulL9ynGA33Yo9CVFC6
3o6t2QgZ7icpF0gAvpcZEAuZq2AUuE4GCUWdmxJQbaBgtTSqgwzS6x+uGe7N69e/
VtMmUWfxApqYIeLJVe5I8e7EkbZutY1ItUjcI8o4nVYbuIZQ+xA0lbtLkiXr1PtZ
fvplrj7+ZMxZqIfWnUAsGpauYDT9qokjgOav5+KkAPyrHsPzeJU+P8Xa2JwTkAji
+xyyfEal7fqlLNkd04uNyB2bd1NLhH5JS1uZZ78BcSvsVcs5j5Zm9vWFWMNsfYC+
aCMnituqOc5lxYT+HXtQwv+wGCbYc2/XAj2TSPNO/sRM4naSiSsAt9UuLpUwNNqh
+y4MeEVANoVmr1wuvltXl4hVETz/17M3/CKbIBiwxTySGc5/ZbcAkJC0uGpQFrVv
W+fhdv20L0oQ+ynfewhF2qozNBwE8+bx2AsDD7fgxeSy6lWDQGVfiQLB0+Zh3pN8
o1AxqQVg9A6jXAnyrEJDvdOxJvxFC8Czq1115bjB5yVBsD5eJEKFdpAOygDsaxGU
rfEFDhaU385ksB1ioJT0O8aXYfqm/UBl0+lsCYXyKrQ6DICq9Cu3KXHX2OGZf80i
nU2cUsd/TKG2qR87Gl/q8FHz5DWrMQbMUYmQ7r5CMAiWSAfvjjTEbYfIdpZv87K3
22ITKgEUr2FlVzipUDhYNAO4mSI3DrAeURc46vIyIRj5rxm8ON3pmB1r8v00V1ZS
HVTRrAhdiNL9tXXWFodZTBP9JfwEYjZU24WEKVnRgtjgMZFdmcoGCQgL6oSd9q0q
6txHLnEti6DtunJxsQfje9O0N3UuQoMsy431wa1QbO+6NmX0kHyvdTcadceFuSHG
uU2rnw8C3a7SxhsRHTE40bchiWJEbUvafhGfmNTXy8altRlQrCsskq+9Hckgc3bY
kzFU2SwVKE6m1/FxWXjJEdGAhd3WTVNI0Q54hAyL+sAvYY0l7GtESPjnUFx5UF3h
OhnPp9RRyeJJTTmYaujJg05NoNYfwhKTvuO+GTu/XVBCOQkttXeJPSulh7zrP7Ch
QDX5f4112YQfqWTLxTru0axNUqQr4oXG+SHCHQBxOpYe2lPJRpjhlQNAnLdKfiPo
7re/odVNYO5p+yV+AN9C4p21Jx9nbg3DHwMxj03pSSp+P+goGEKJTKG66OQk4ti9
+LRIyY2UyVkNlpHX9KwXNPSsuUOSQMZJoH4xwYqOz/D5kdX90QVOxBxiQtdrls6u
v3/mScx9vNmLyyCykKyOzlzaP02bJv7Ijy7oGJLZ698zL9rw/YtpZcz+SwhfCnZH
yUag+qSg7wb+HeO6zfA6id/RGeyKj0pUVjCFG1WXmzjNe+Tq+pwR5c4fcfviTniJ
9iEZd6ZZxLEptn/fIHRVVqIOiJUooXeHm1AuCrMzu/HHAOo1B76D7/LVnobd/SJc
V6MsLJF0/SS1N6VCs+EE/uaNkIsczo2S1C00qFg2OWhZHA8+oJMluvE6LkOxM/7W
UNkNLHfXySvnfQUPxW7B6tChLYpxSdwvb/0KIdxfbsTpGX1hpdvPmHpWagGjVvZE
LPsWp9kGv9V1t16bin87ISS6D+CPRfddJRnKe9dSARa9/rH31ESKsBxc1h7hZcL7
rrTbYN78D+ai8QZ4at62a0/l7vgXj++Hg6bhU3RuBwCOZPyefyg1UP/cdR+qLubG
p9ocQSoa7rDi6U9xOb7YK75sierd4fnOm6LFntYRMIjyBqJR1zr01rN3CaLqMzvY
tw2aZStsi4mu6F/HJ4s0GmYFFMdm9Bvwj6QfLJtZjSHrvwG1ziIzNW6XfpP6+BAX
NLXvIdPr1J1NTKXMsrT4PcMeyUElga8k06gXXLS5QW1EvY2RXpUVOyXVc0nh8sgx
G5koh6UJwepH8maXmkUsXC2+Shr/zzFnBhw29C7IxZjG9ddTEi9s5rNpAcGAQvPq
S+SBP1gGgON1wBqQuKp9gTI+bYfb1RPwWq5PXhhxfJ54/3t42oY7NS1Hb7NSCjqL
Dr57Bdl9t/ES4pQkD0ECcpsdNQjEpIpZvRwZaRQbQHI8pw6J9vl0cT/jJG/pHGrQ
bDkw3BHdMBaazo/esAOB84VSEUi2w6SrOzppl48d0m/EJczILDeIIxqARjWbB4nn
V01JAFoB/KAP6968Kr/84d0hd+iWVxL9lAHmCSiuaTu+PwyE0Hi3NXt21zAzle2r
Vrft6K8XDLp208w86kK1AqGLBr4cJpN1/Zmtml2wMxwyX2WRZ1rgz5XZmQ2ymRXa
ZzOPWazJg/1931hH4UUcKpQV8tIApw4H57WWVCL6prnba3qBSSCWl8F91boo4V53
F8/4J0oejivLRCIlzrVQSlfzpKELpSX9s2BIUeKVfpdesHbkBhbfJy7pqzfb5EyD
XpVagSAE7nowO7xiv1rbCJnz2l2LvyiyIJnRZvB6/Q0Bph8IDzvvsUxhYskNedIM
NBObUvoYbOInudU0lo+PaDuQ0MKRs+WKp2y8YTFOzYIaUaf5ynlhGv/8JPslkDCg
dXbZplGPKqLqwa7+VyFdn7p69r4SS2BwqP64lUAxp0joC08BNkKpZZ2TbL0H7WB7
CSNsRBEiOC9iOo+HItzGn3CdexU3XjzzZWQ+sfF6XF29rfPpPHmy05zD/QpbH+nt
Sk7/Krz7YIDlLj/cKgwmi4ALf2jnkOU1jLJficWpnNz0M+0VI5DXm5EC8Est5NFo
B/IsBDewkO3081PLFWO3w1/J1YMPVO5AtHWEHsXyYFY4tPUrksWENqzRwv4bon9/
B/hbGBH+DxzfrnNdvROkKrXurwDCGn1P2AyscCEf9rfA4U28LRt8liy3Fb1QiYtg
dyQmql+0afN8F0bUVmbF+AMryFer4kaaVgewbDhQWpgjuJ9Whc2wnCEURoIYUyOv
ThKOApDg4/0SDd8qc6tCO1Qc8pV2vaUpWGMM2pqNs5GvMUTeQ4Z5afnvQMaREnDr
OBkGFP0qGJBwkNYhaJqKjD2BonnhhZ891FFtvyOp4iDyQwx8MoxGCSVQGS+jp+nX
67OyNtQIGOpYRKqvSHBEdBzDYvbFA5Q343RXKtTYgi4LODPiWb/Xe1jcZS5qAWhL
SW9u2JtydAUqg3DtmwXBV6YJ4OR/6X0OAdBvAvAhQP+vwdYE6Hvx9j06LgSfRAi3
FpSQWXefEWK/s7ln0nSjpRthz8RovnLDK4lG9/CyqBYyvt7+7TtS43Ak/l12w2vv
mZw7XhcrSNm0hg85pW+GU2YobPkul+LVlUumkb6OiKtGyjSiKH2hJmyMaFJCoFBD
B271fxomRNBlaip8Z8+J9URUGPmOgBru5oW7msBvPkZKYQF7VYrHNtF9SNrnBrho
y7ZT2G0I55RaMSmoIvVCOEtb0tVC2AwZ4/IsUJH6QDkK8kB+275SefYL+C+o1lMb
ar+rBtZH+WFKGUSoX7cXKFdhoXDYUY9vaRKO8o3TKmYBW8mVP9hpt0IpQYcHbdQa
7VSKrvkntGCQp1AusggUCSSsoer5KqO/HPOaeVxx7ejxwTlVfe60ABo/Cx+9djoH
4dnE9687ozoVNwFTp1yoQ1Iyx2sx40RmZhSSKmEtUmF2/s/MYHe9pywAX7SSnQzl
ZO6LaKaud+aMbSXKkLP7n6mNXS+89zxcUsbrNqvli0DX8Q5Hw2C3fISRBzt18vWk
pchqsCU4hrMh1ErZErGTutpki3mBjt/0wp3anfLJW2NY8yUiD8KxTy5ZOMVHEGc5
BDLRaDrJx/QgMcJpvSE4guKXVRnTfVT48WZlYKRRlc6OyvRqM6wXDyZdNymPovME
WBA2Vuueqqi06YwqfZlmuKOr/ZMMEAvWqpgX2/szHWkcoNzfNrEq71oj7WRxQCoh
GS+1q8spkn1aNp7H3Axoh4q5fj+PufKHe9/keV1P4yQLwN8g2jl0ajKgLIQ2l+Y9
tvaPRZKsflXW2IbHpqrYI4pDp44/EwzUr/mgoecxVMmVhlxmkk7zImDMDrXtB1nA
0MZ6kwojvbe882BRY9WoZbxSIdnZIJXi6SEkaaoheG0k+KqacQjwSekWeV/7rAQB
n9dt4c0jhabyXO6A/+ZsEldnCLyqB4eNmCnxKTpRbtyKljh/eKLATJSxD9WndlfA
KqCvNeIBMpS4jLr3FlPd7xiqrSmY9FtMpWvqx8XdH2jmHL21v35v3wDrJ3A/Jlso
Mhhgwu3kiHV3kkgOlGwswiGvktl71x2M2tMkryrnc3jHwOQTJb/J1Ws8XjO+xbeJ
8/o17s1nJ8lb5l9+QiC2iCS3yEDhADhbJbAAhvtKK9VWAnUWA2EsnbcvSCJxbNVk
qLL5XpBtsJevxXr7Sc7SDJmNQjK5hAGgsKAWikrp+d1YKiCMTGE2BYEZrFL0WyrI
n1WVNbv6Z3kU9iLjjMYcQB0rHR2GztsoFucSiVxPW4qOtCS87h9ownKzt4EyylFz
uvo7Hd3DwDvKpn6/i1R+E9kFAy74DUrBQSt3ElTN3zL4NxSCdPDz5BUW3/L/5jOC
80oN9wtRkdMlmwU+0lhsR9IKXkhSzMOT/vt43VfNvD3Pf/l1AW3Ky1yx/ELj3EbI
06poNjpRRcjukfQowL0HJDZy9K8nu1+H/SmXVzdpJUc/xagMfXEiJ2OyQ1uKaCAK
7ur66hcriR/WkV4D8Oe7wFpi5/9vSpbBfArMpkSNngJqURlwMzu/DUWd4SUtA7PM
XnKO3jUU1ak2xpZhTpaOX/WE/xAnQO9zuHV2ruXfZ68llc5zA7LUecvLPy27D54l
lmAJimaYk9bBCckxDOT6FbMaAc83fndAtvZhrcAtKbr85XIcwf4Ts0DClwd7UMTJ
63w88HX+6o40szqi827mw9x/NtGgepQGO5nts93EghbTclf6bGW9z6FwuMNw53An
oUUtbBcYPoXuuPbYGscJ8CXEdLuBGj0hx1KFybiJWsrtXFc9m4fSApZSZqlTivYh
2asYoxIJcR90DJcyMGScWA354Sl2fWmVIbcx8qkpm7pMv1lw6usXSgt+CFkCJxM6
2fwa+60DNUTiGaN00F9K48vPWmwgWdDOzk4Vd5VFUNmwgtbhWwDhlTxfYS35o6jA
ZkycML+XgNp4i9gVY8I89wxZF7sakRAyb7xyy9hhJh2+iJ0POCAD+0zlcJt0n/8F
5zfZXzAHWPPm0YIHVXrDBc35SvS0r14VB7GETrZKCZkm/PqwEFQ1flF+/JRSvnJB
+ip/2KBdZSeQgGB9wWbQOBddV/CYz4FBbIsWyDRDRSHJoUfv9rbeiMgwQRLUh1iO
PRCJe3owRmy06Qq5dibU+qtrJfvRpnUEZAvfYHjXjAxhKSd/rnWiMb47EoNXb7ME
GAJom6pIj7c8V2KitQdtc+J++flwcM97Oprk9tyCG/iM6grHTQ2m4WkbALU2MAhb
4TZNFaQqsFXuWVnHR+SyxTOX8bzAvCIA+U0ba/Yd77Hj4Mi6+krQ8ASnhGVi3VJz
G9m0XZtTy57MIAfS8/7NAs8EwZpZ72eyHicewr2FqtpQQVgfYrhFkBSdPw3p+Zb0
3wjZOybDDEjwbPdGItnAj1kuN0whFLnOBNbb+ZMwzmrwlxmu+e37ebnDBIDs6ko1
BSMV5doynUOrFUZH5Z3O+r9gHLxyTWiq2C1CeS4t1Ey9D4Tqbn7CaPowifitII42
R2BbLmU0tEaPXmdLQVMTDbvj0d+Hbcyhm5pn/OANrfYdwLTpcCQsk1MmGJhs64up
hafSvhkOi7t4IU4oQZMnXeXYursy8Cc2+wYdHVjar5qHqECgb02kJODRvDcF5gEb
BkJhuvTGDvooyJJ+EbqBIhqt8ghzHrp3U5BSmkxmpu9r9K6Y83QYkrNqkgm2Zk02
5xbn8KjSMadb/rlWfLfP4AglEv5rsdKQdBvrhzh7CiP9Jlg8CnOOr4teJpL22HeO
IsocvgetlmhryVQmwjMsOi19rztFriLYmUKrdHiVD4mRRX+0L+xYlJgkTHAY3FKE
2N3X63/Q2SIW46/L8ZRHFojCiBXw62jOqTf2fHkruusobOs5CNkx/iSwSYR+vk04
Sy/YHF2WlmqtD1AqirmsMjrJDFK8SO0qkHeeoOKb0zY+FimW+xTM7PgGyffcZb5t
rWwFkMrAThBiAOjxl2DX17EfB+TkpWHEKDSHSV3YlCjG4ceeqt1g88vKSy9l4r7X
ap3EylnwAk7x6UmHItlew1EJ6dDZEtfUucC5Lu8MnlaBAA2qYl7YXScKDe4DFr6b
fooXerGI1EsvAQRQ6DbsdVR1zG10nlDo0Vsskk8AupdMuBcd6zfY3Y2zqfKO7eeM
fsdDeFumipSapZSAEmK0jiAbs2BWAunY/KCaAMGPt8jBdWc7w03KCck1A7QT/geu
9+gcgVfid6op6SKwJAS0D4FcQvFfi5bQlc/JPWz0Ug3eS/VraM6RBl5BSAoN6R2R
bFC89NYcnU9cC6aeYqDkmS9lMrV5T0WICqWurS/7AQ7S84/K9KPefMT6PTNkbit+
gIlBgGYbiJVS1DNJHWm5yabUoh30j4MiDJAorqnB4KBJC9rN7stLhTIeC3Ov/Bd8
JgrrKlQich85UXoFKBAh2GZpCX8w9zOhKkC/umvJZJD6QGmoh8VyP4kPacUJ0Sn1
SvP8W/hHTxn3nC13miZ+yq4IkB3oRi/r00nVexu887XbOCjJVBmpqWjbbWqkJp1z
ihNlLagjGh/+gX0i8ads+wJxLcKVh82JWlCknkK+3dD7qEddlc/Il6839F+uMB/6
EkOMtJ4TOHkwQIATzBJfolVKBBk5esSRMPc7aTFZ16Hf92eAjh1UeuDemLpsOWpK
b9idw4ukiXYhdYBSQfbW4c/siHLJyQ4+AbxlCiECwJxJ2Lukg8Yjk43u0r87oOmo
vF1PuPv5x4oO6kPFvotvFhxfTLoLXKdY+Cvc73JB7JE43Jue7awSL68/kmrs/9/8
qxm5zi5V8iagh2/lIjeDuCGvmo0h8qinFSbCrXvF9ckDTn7jvUq9s0JKeZ+BLnfI
53M4YFq/O38FJAuMJQRL+e3FDoVA/uvmGrV5EmTOtCYO+kUgUpf4m1aPHsLVrcve
JTexBCJCsSJW/Pmq/zTdKrOUOlZeiINBany29cegUx2dTNVYN+aScMo9x0KbjYfr
Z9L8Q0N+nLVqp01/tjR7Z9rrKeNPOxUwqeQCVVaetl4Z0+48OfKFuAc1az3Mro/n
bcy5BYYCE7LqeaeKKIgTrD/8twDetPXgFfaSs5YNGZAGIhwW9q9C5dA/kIAnoF1+
MtS0FNV4cjAjgolghBrJvoFpr5bfYPCQpzqkk7Xogb7VjYiDmrl7/owSz+RE2UTI
hMGgJramSCHqsH9vEvyEWqAe55eomihhhgRUdmkRQYvfViA5QlBKCh0x6SE8REzC
epgZnglyx2ObtirogMKI8/YAcg/grqAr92TN6Hif2xMTlx0I0hDl04jVfIYUidTw
FNYPj7JIxN6Wxod00xvvKoYWG+69rDEKpg7FIfBuAA8Od4dAxkxFyoejaheEm8Or
fIKBrKjvyFy0HEoOdN3u9lA5jIT17iRDlUbK+4Ul44zgXaKaVIOavsInfhHGHASN
m6kuNSKG6RF9JgCPolmUNrThlFHao6fWpLWl+7eY99XrmAGsUJt9kekKM7fNBA24
qZj2SnOzcmLkNuEzV2Sbr0stuijizqQ+hV8gMxR9t1yoUvi71Yz/DKwUXNzIRRCc
0HfiW9PDiQnKxhp/ubgpSve83w9fh82ERHKxZ0QZNBTDrA5Kk8+GK3T5g+4h6wgU
98v0egQAukdqpBPxe1wwOX/AB61H/KeZuL0f62a1P5HWccdAYKdINH7/rXqUsxy3
Rg7o4G/tEB5mORK4GmtVFcfb4gzeDZoykqtRsWSUCDaN+8BQJA5TFFQzANdNaQVF
8xfjZkIbCXx0ol2DpphUeDA6XqaMxgBpl9uyG7Ix+IjbLrgJRyodBvBmRndpla5F
c8+FOMX1x4YyyqwhjCGFGlYbTiekduLfBj5rE4k/gr5tls4xRLtIl+NSKJzgJpsp
ccTklN/DN7iWPcLkfB4Bm7rCTsU0PyhNLzBPgLnhACtqePbazLlY0jm+Z/LYiZGA
K+Ti0KuOwlmVSY0tXPXuYyEshAKDhCoW+tCW50PDhoqWObnPMo3CxH3wkPkIpXf4
iDu7XkkLDCTAGSZcKygAjxNzwinjyhoRCP2twWjPx8qcqwoI7nrwyffj/+d26h6H
ApIsvYzI/UgdhwF6RuiV2d7snp3xgRXmywqPWvRCizIjdvQVsrPYYzBdwhXSF6yq
1Qj/hQ0b8zS62DF0bda7YmXz51bUUY0A/l6a5e57Q+C6wI2I9dJ3c+K64ibjA1Hp
rYTjbh/plXT2D1v4u+FhkO1t3+YdJlrt//HvpQOb8M+ESH4OlXq8e6uOGCh1qI/k
niyHBsLpvRxyv0WYs90gkIfjxDbcTC5zpaB5IXsg9U9x0al6+kklGfDZikBtgcKZ
e9s2AX967MJXzZ2VETxkYXkBmLBvxp4OkPkOJidi7Jn5OPoGG+GyCd/eccvVLl7D
Um69Fvgf98V1KJBjh5y3ucYBvuRRzxh8YFVbksQOcfHWRwS/P8gE5HeMNPcOtzHs
vTzsMZ75ZLidrc8tUe3hPxZT+ai4TIxgxuO1f2hjZhSZkD5nR+4GeS4kYLIiTGB9
+dakRWkSlxjr8UZsJb/EvYLLIzI/CrL7nEjXAXD37R/DB/+iSH0Gwf61y482eJFa
XEoMr7DaldxpojNUWuXCeQcOfskFWx52ut4+OjIX1OJKOsIUPrjb5CXKh+1+Cvsi
OcgIB2+kl5eS7DFBxcerzyUt8jXZ7hOxnJJSk5XM0XowIf1oosclGxAGpqTN9ILF
/gJIy8x4B5yBYXUvsfKih1er+Yln/VViqVQQ2F215PpVMGgct0uLjMDM5X96oAio
yVKuhO/f+vwUszGehs1mSa2/yqyfhStk7eRi8Z8LlMJS6ZVIFl1zQAprGb8fE9jL
SENL0z0c14GmQ74tfE8JwGzpeZ7Vt7e4FSgadgEdo9viG3zzrMYZ8XRZPD0DQ/r5
Jl8envpyIt3F8ISkZv4mmizUFNLFt8H6klfyhnUPLxn7qGj4ao0ySk7iN+WJja7G
hN0ajHaVMv/pmvLSB7ZrsL+LqYgQRVdLSmre2hY6GOKyCJI1rt1HYuvY0PEMPy6i
nPRQ4iao4RK0aWRxfcu6bXqTufEJIu4AGoj8Zgyt26yt90HxzHmD9/HFj6O8h0VE
7Y4+04tikRm4uANDDE+xThm+TuPVhwj2p+IvmR7U39DwGY0qAi2EyYIqTGKZM9Gm
jFjkDMbhWo6fXlLcCaWuHFHFMlsjV14Ge/QsecOJkvcL0MPjtprB8zXU8TKbtrY2
3R62ea9fRHz+vMHfVJTZTuLfuATJ6PjInMIXoZUoAjaSQdB8QQPKJ9PA8K4S7kFs
Cdl3VJBnCnA+Fifaa3fobrhKmCrPv0fuEq7trdrcupFLy6AyIFZ4EHxE5/a05vRM
f+m7g8W1C0J0VEVtLORRGG8JMwr62B4aQMye9u21Lq8+HL9yEEktmL2EPKw8WtAI
i6k1igbQQw8NkPbStbSsDUB/bAwwYsNcV5AOryfynYldTysaxteiy/JdIpoYa3u3
fWoSNJYBfvsYtVPBvpeyDvC2Y2sDer3Amp7mahLxy7Z3Uolz/yCzsFEbupi2REUb
YCpAf/rVCVlZmHuMxow/QvkI2jAn7hP8hS49hHie0ZScyRgkRbTvcs9uA2453xjo
3Zdj5gskIKhlzIIYQ28RrfGM3LjHT75Ww0k/v3kQqqdlhV00th0Kaw2gShzcSkCW
FwFN90lTIhcOKI1RtAx9Gza9qN2BuSpXVl4Eki8r68OKRbjgqIPGv08kCFwFxyaM
hTB483jPfwJwRvXXjFp3Cm5UARPdeqsl7DrsHTMgnkcH4uJeqVzX3jk/3JfUdIkU
EALR5JpPJGD/sHWbfajl2xy+MvZZKQtAn4f6cpuWWUKpDhotMRytazPGQk3++Q6G
TQ9/JDZ6Hmv3Gnmj0J88nFsdGdr7vo5A6SxquYc2ut3HF7UaIZ07ghiqqYGsUsj7
a8F/PJ5UhbTXtt0OHhsRoiqwPkoZBPatPXS8frSqoGR7drbWTaBj6Ldp+m83T65T
Fo5fzjpJnAq8XQVz7u+x6hfkFGweE3X4UiDRy0ff2+t63lByUlB+xwQ6j20O0VOt
I6E9Je0dx3jug3+e098+4i+EGjCstMTnhpjiiJIOnq3ePPjT3MbbyckgwrN0uWh3
uWj3ziWCaTghMZMX/C6q3qOM+HY/8u7lcHgTe4CvOfbBw69Vg0XVnFKs3ZSzUqWj
+NYSRV2k0RWReh8UJtaeFl5cjM+xnFC32RVER/uklMtZoe5VXNApwJ5YCIglx3Gl
DCVig4AthWziuQmzGp3IY+3TPuD/AecbTqgc8ZjkYJUTS3VRoqaGNw1qa/GSagwp
MEly0b4s/Q8Z7nOkwEVCzSpUWD/n42bp/MpWlOIpVyBc1uoZhag6KshB0SUMUihk
PpqYk3OOBI16QpTBimH7Tu5D5sqoHQowuYdenvkMgVYPc9CP/UJWvFht1WmiFx0G
2XHRMMKHD+jhHrVnfhLaIh9mUUSD225ydOY+XAEP2aVT0ahTuljFRpgIlRvh3KWK
VSSJjN+uaIjmXIyx07WEzTqeIhu9slmaX/chAoqc8zt49KYV0lmr8SGxsTBQYnRW
ocWstglDYICQ178f+KtnF4w2kVo/0YLBWRWugCjprksujW4IspFjaBWdIbCofPfS
FUnmPThbx4IG9HijPkho/clmxFHrpeRqirdYOBiHcInxDsInDv2TDyBMewaPkg3I
oj3GcRFeDUJYf/Vb/XjCGZ5EFIwPXATP2g7lDJ+wEyt2mDx00W9T+Fly4vwfhaSl
8TKNLq+B0efxRNDVtt0u5KQtnNeI1izS+oARLU3LYR6gANYa0GhhflO0A8nBfTrZ
xxX/FUvP+FZoXpJG4a9I41gMo8GUqNTE5LkTM3I7pfJ3CwV+tPuoZh01UBk+Uw7W
06ZFyL6qiPTUPA5jB5cgXM8JIVgDua2gibYEuAUL/7Z+nkEcxVTG/TguUM/5xw2T
UW9Zd9sh8Btdu5F5yEbaSIz8i/GvmUDqpxSDbsYeKMEIsjBExbw3JmzLzjJbvmWD
tKv/s6iA8GQJZLn4vBa3UoYXYldYdW6Lh/hWhzvmopyEMxEcpYltZQdpwmiDCtcR
cdcg9O7CAmbbiZcw8j/tqMYCLBmkUvd35pS/DyyZYUG0wDwUXbEHJCC449AiinSn
VF4zQkHJBAW5HvKTIBbcg0f3AWGCNrv4BbCA5/UA1NH06yxm8hegUCJBiS1JxXRt
RO9A1LutQ5B9IcVoljPdqnbDoRvA2aBKYsKWPG3tlTBI4Ie63ShqcJZy2uMICT8/
2bx5g90CuRkI8/decKFqpzPe3QMZkDWjLN2uZeqldXzIHkIGurYm1rXXo7hqiEhX
XXs+o1ovAmw3Y+5AxnixRdZ52ONVD1pu+GlSBqkL0OhQUo5nB1qvCTNk/sYQYAxP
DQaw00ACIs298BPTGifWCiRh0QI+QHR1sp+oE8fdeMUnacNbJ1QfVgFqPuOWJKRS
EhjHM+MWYra5CnHED9BAWqG68PmDNFpNAHIIg9o5+CIU2D/ki0K/Igghvq72sd7/
EevzJMr3I4uiZfvdFfa5htRti7shOJqb8voLmd3nsvxU7QYf01RwYI0Id83yXCxp
nbteMzZUAFMsVK5kU3i3JiFi7jsL2bE0k2SpSylzkeNdSY6r9Gg6NdCMYApmaFN4
RTc69p5WTS+z+cTuE2Isa2+95IJppl8k9v/r6/LEfMjMqqYL+iBLRVRLTchaB8o6
nPk8XLHjjzWv/K1T0NgF1D7+YsrvvmCj6OuNK6idzAObyCxu1yVovV5S8j2x6tws
2QmQD7mG/OV1mfZXwTTrPnQBe9dNfZF6uLTEbDVO0H4oPvZMP7aFlaTXQE423coo
Ew07zuYaFis9zS9EtFOEpH6hBoIh7RX6lOcexjQB+9cZ90kUSQpX33ZIRYTPIQ53
YA1ldZXEhWPkCaI1VLPj2iyz+WwvbQLclr+Pln3p09CzjGgrFyHxHJD0M7eWPRgr
BYMTHE2ycqW6jpR5CG+XU6sysFm9FM8urUy7tkdo07i5/uCTHS/15QaJWB5DlmtD
L937ilzLInZFoU/vpKGkg0inKVj8jMYr8Eg52O1OvdMygq41OutMlSWdLy4IVDNX
0cq61GqXDyG2bsYdpq21V+Pw4RJEbyuWK36iCD/LDwzZIzzobHHSN8+VkY8stdqz
ps3gxfIXWOb+XfKwHqY6yyEHwTjVxdcuZjUiqRG5VLh6VXUetiWffG5w3fAYCWfk
5J42F5QXXDjibTUA6Usq695kmsTwGr6CUPuknGuOm7HT/D7Ig7VibsW4dbpZ56V2
mAT3ufLzR3sWR0ItEKUMzoUA5HmoUbssV7FJvRE8Xlg7IPOAk00mBWvW2Iap/En7
5xfUxqtfv2l3nCQUwiHp9JSni0N7PORBsKIb32mNmqr7EVtbt12cTem3c6G/IiCY
cAmRgXkhQNBip6FZRbnYtICfU7fw5c/j49ygIu4hQ2I5UaGSoH1yLKNf7ZjJgC2q
1oKiaVm3JclD0j8ol2Bb9GPMN5RV9jD2+vlMcDARsJepkZ0QVw7U95lysGsqk5Z/
cJGCIroofKL9snN+GZibC1hIGBwQZwct9+Ol02I4T39788WFmU4LkzatgJMG7ANM
UY2DX5WDiuWJEvkqI+f3HaMhOFD62o1ccSuj2Js2LhxmUIaHDCVqTr7fcJqDtbjx
FOlAR6eTHPaYaPNV9cUl3EeRl3Yn1YqB5tIP3egXhvmFp96peLfDQLPJVPnxpS6f
O0bRK4R0OKt5ixO2nu5aN6iFf0WDbquJCChm7k7AchT8Oq9Z3NDeWY6AtG4Ci0Lp
SdnvoMgbF1IK+liu2MsFTVCUFxaMeAUHfHZWKUVYtnKLkFohuqooXTGgmlMtuy7A
lxKYZmQC+Z1e/w4/rpHLiNKhQPHiKiWOfzj2ubaSALcLwG/EuOpcQ0G740aKpdAb
pUdJUkDPTLT6dC9eSonx1VxGw2usQxrEtlc18TUpTJc2CEzZG0U3YIJ0oFYZWuoF
rMVFbewejlMQ029f6KDMFSgYIMzZuGhl2wIGf0s1O5Ixfni3NnohrjdUXvyFgCWC
3DtMbjpt0BFwhqROMi7NNFRPVF0upTjvrR4KNiN8b4yD/RhQlPBFnwCLX65MZoff
dB62h4XLG2L6E1E6iLON/Rf0LE2NZJ0WhkA6nHak7NVplMc6chbPsvsFbLoKoZC6
/F1sZoDAeVYOXrVrVJKG5xwVC73/7gn4rzOrLCD1qpETqrjCZKz+9HXrB4YZDwGR
C7siXIEgywoybzxYD57o+1i+vFZ+57k4iTeKuOGdgjZx6SoybrzHZvtCSdV8jSR0
KGXSkTziencCsu5KNc2VT7moqjKGvvYsPmq7cjkE2whlG8dttjlEEzNwkGwqiPFf
a7XUkqb6fpTBDwWtT5RV8bQ60u/69PjC1koeRsqORG1tuPCgKI5rQStFr5x+QeiN
qvlEQadLuP0skyq3BNgS2cxp0/XqIHkBy1d4iud+/cTCcNV2M/erUWsbW9po8GYZ
Kt4X1sQrKHiuXfBKX8ADdyizV32syHTHSQZVDV0KrBenC20MwF5ICkok2DlfQhqz
jHh7jG0RXmqI1ZbT7qUCDOLKgo/X9/Vni8UBDZnog6qzA6Ad+1D13EZ78QoSDHjk
7yolqvspsq1nLC3pd3GDCKNyVP1BJvlNVW4QWLv3DvXPbhf4DIcOO147l4zfShYp
BRVk3fGrnvt5n2kbQ7pnzIbKg6n1TrcE/b/N1ntUnkIIZkB9jD9yhZ0dBD/yk8Eg
PRRL4jG/P6b+E3g+YH/j+VduW1VL9boMWpGkYVydGWAEPZXgj0CBGPHj9QWvxSTk
JlnyB8P/x5arrOnQLQLdZ/J/FBKIFwxCEOwPouuAW2MXl1UBm/Gp4GKISeFWkOSX
8oO5VE7zh2V/Q6EOHXB/rF0vYruf99dsWzSywDE68h0qVHMMR3dzKtXgXmhDASjY
TClzzC7iPBF7MK9UcHj4JBsQJwIj2ZjtW+D1TXX2LIjitKZtv/YzC7liUwAaxRtE
tldRvQglDiwqHZSYMn174DN6BPTUG1ZmbvtNXH0ROq8SbXk6f+xXde9IrZIwGoVV
a/WTFwjwKLaqT0z3eqvvlisDAzcIC593Mt/jOm/S7XfPVRN/OXSv34Kc0KkXNZUw
312etQ2Sxj//1R5qPZqRLKTVYp9LrFa/0/3tmB11hC/yLwAqeeMC5qcsxPajNRLi
I5Lsw2MwZV0am8V2STfIlYHaGNsaqtep6suXMZ+6vvaMQ4wKlLwFpwqJ9xcdc4Gj
RPKT2a4bmMH+yR3FHwg+M8iD3sDzhH+NebCubGk0IuIMRHp1m0j3z3Vsp44grr5W
ggT3vLMBDnB9aOpxC6QYv8sCIC0LR+jeovOuarucqahg3euyaQtO+o50sm9RIyjJ
NzT9akWdpq5vLJVOxUDuFC+KkMOsGd8eEPNq80Q2t8JWPmVqwhJW6POc8Xfe2YbK
SiQTSLReZo9xOWzmUMNaGUg1bzdkhEHn+9TnDMGU93FcwgDBUjri4g4u9hBe5ATG
ezKU7IoBDvByBHtJIXbi4t3xD6/a55DyzZk453ybCMwV7hGahEBy4Ubb/1zzQOjJ
e11dA4AV5cU8u5s+lQj275oiG0DqOqOBQd/6TCJBd2GH+467ubD0iHK6Uwf5CT5Q
eCffl09G9PBVpiFoaGm2l20kO0/gO0yN9HwLDMX4xsjwHxYVn43IT6Jpaj2kTrVH
crFWWBAt8+qqM47oxqwA6+hGwEtCnljOROM04zqYPUNPM9BFw0DcBuLA+hlfp2UE
Q6uUN4P7088/DReJJwZYcxOmbDNr1PHI3xqPKXx1LI2CoRrWcx3VGJQAOcmqdytd
EmVvE5zZCSiq8bQlsO9SkJBlBM1uW8TywLLdgKnNjM2DZ3gpd0Zqip0BDrqaOeGE
9yteRDBSaEAVwf156HvHEuqEEnnT+DLApqZBCik5S15Yq6FmkY+VUWKPHPmuG4ub
qZXkzklrXUVqHboEg5bTs8N2aJZUrTevKgswTMvqlBTN/JTa1iboui2gTfY0Y+RD
GTF0wH5+KV41Sm8pKmNm7wIRv3cfq8wxFtuYJdlgfPJMB9AhVVDO5YrT84/1EI6J
vQemy6Gi/zwbGSutdJD0ZJeE/vICmTsFLSBfFywAZrFRu7rJuD0vgTDjC53b9GZr
pyU0NeaajS+7DRmnPnSOzQk7KhkZ+ZqBQx5zG9mp+5dYSgUWXagxV0jFkrAUrtTg
kG842Bi09DpWCz+4gBSNhgNtKStITzhjhuUMHSOpHYM6+vN5yC7BCYSUaDdOWK08
C5ZG5CDdEllPWHTKULhBAM1WdJTZ6nXTyNNLkaAeYfECi7dJdsu4KSNeTu6eyKLa
Tw1otiwIaFCPj0QvPgQfgXBZFpzuuIK4u2JwswlzBmsIJUVLVjmL1PZAus2kRbYv
zxukvUU9QKc2v9I1D+tzEElJbNXosmGTGkxrslDh2Q9dckolZ3Xj7Kf9PIw8nhLl
iqw2X++K6DhnmtjD6rahKgSe4S7pC4tLuHYSNANtkw2oUUh1EQiv4mY/OfbeqfPR
NCFbHup/twLk4HZdLsN0C5KwMrxuqmo3hSSAsEEuZZF+9b7v2jF38FpICnBzBWmg
cRV+hz9uhh/BWSes9D+Q97YVS/G/29bBfbzYaNORLIuecAoNc4Pzs4/DOKDm3sIJ
vHEnqeR/Xu6jqOV8FIjYyNDKlFshfAxDUADBNLF9llfrJqpX2+AB2XXMmf3MVCRY
JE10RbJWFuzim9I8esApiTsxc/VafWurzb/0pJr+bqYhLkgP/oc1ATcZfjvs5ywb
/gaLTv3mXoNwMdWEc1pTL4VuYvvUUIrQmlzvf2MvhfypEeACfm0IxhBwtkkVeHEv
IL4uz4gOcwERqECd8f2Bt3jExUSjT/HkjNCu62MGNdL8aYzYFVDqyj9OdRN7E4+W
dznh2N2J1V1e0DCAjJyQ+TBizjcj8BScGLCYYs6fGBkes9v1jMcQ0Ck0J84ozrX8
QSa8O2CFP+1hk6lfzQHmNANY9Y+zyppOjNV8vJ9eocp/f4S8H2tEfjBLQZa9an4F
D7LDXjDqA2VxbyLGEww3zmZw0Aue9lPPWSIZfacwu71fXM8fVi2Af0EO1m0dMva3
MxYHL/+kLnrBfPEkvsANABM1rZ/FafDyrLL1HBb40z2r0fkiCbrVuCo6mP2v6Gzx
Vbe0cQKnxrkzaYr1IbBz0J6UYBg52JM1JL3er4vplXZPakoPZ2zFj6ewQtiO2nAW
opSlwyfonYIFdvvx09fyQFyQOOmv3N6Xri9r6ojWQPQvEosienf5l33rb4Cut89S
Flu/YI8C4KAQPH5+BJ+Eod7zGkotyUAEJDj9gMujK1uVmHpeKQzVHM13S6VoHc6S
9hE3mcAqyHa91uzYmOg6+fp1OttWxt0FZYvwijUVWgdHCjtbLxfmHH2yh48Tny/K
O0NOjSfZ+x1j3BIPl3jw7eoIVite+b5yc1YG0uRsRCNgCWDi5x59gBm/JrxhmH3d
cOtK+APDiYMX1EeTkUnQuUKEuxaaMAfxV3WRof79WMXUFxWm6WlvTc4c0FNbrMn7
jU7FXqxTbjE8h0W7V44aSMN386ZlGLUWxKIvlj+BJCjASTVeeZmq18D20DZ4aatl
P9C+pbf2/9OuORxldoKuzg+qlhjWf2HoWCzrXdNuQ5uVFaVyIKYuvmvFwoD4f+2g
wXWy0d7pjUxR+QKMEu+SbPtV40YloJ39JtKcju6ZCsBRhaDJ13jG1Dml6eOCxwsc
lpXXehcHyXYQLamT45i3iw==
`protect end_protected
