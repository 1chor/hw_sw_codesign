-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
d6RBKqGQIr0Ja/GTgNvCkCcR5IiK5Yfj0PRbScc23E2Raa2vXTdlhGXqIql3TpDV
SCauGeclLpES0KPQL4ezT5qw/mn27IyR0WmKeLzRfpxE4MErWI5Sp4xQhsoKsIS7
qKEY0D0trg01ygIWqVRLq+4usghOAcCYcUAyqTSsKxg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 2656)
`protect data_block
IqrUj70F/ivPFSeiYEOe1eRSqv+ucpwUMD8hX7hff4tHpDgliLiXZam2m+Idu6G/
2c04tCjB1llOEJ5vDk6BzlQziAgZIvKHQ0MWCxpAKKU57JLKZwkGASobaX+0XfBX
37yCdBgZqTJ7uTNpcPg5kBPohRH4bMaA1M0pw3K7j4pN4FQzPSt/NAJebcMB9kgY
FubQqWkoFi3+tqu8U9V0W1wUEb3C1FgacVFIzdtKg0NDluGiVPeiwb3SFhONnVck
jLVPKEDpJ96GcT0yfzKvzZMIE6EnDoWsxacGdPPu3LUydrBKS46QUt289LxFcHk1
CuynqQ2xRRPCbpvAlArJFF87EGasdxpkpsDYH2stEk8x6UBjvxx/31f0dY/TG4Wt
SGMdCdJy3csvig2Vqt0Fl3hgcXppVfn+GtFxaCSssO0qIULGCl9HY5l75husLIwh
uimpHfQRzYz22nsVxk+ECvRQkyFoLB8fwy3RUPeI2DADWFz+SqIqU4TkXgUiOXsL
ngu5TOZQdLFamKPaolc6N4gpuQrUMWZZrY7To2Gv0qFx6y+REc+NShAq+DoyBwcv
0RZCMGfbd+GYbtpT4a/iCh+C7UpMl17Nxc+0EPesvbLYl/TYMGM7D1mOiMve7c3i
pi+yb66aiPr4Y2RUP8TcoSt8uRaejMRD+0dVDr/QnSevaiL3QRjqJrK1B8+6Zr9x
tv8+WZocS2HmeVqllUqJ0qeacV1XMv8LRUeVIzDF51DCEwtl7ki5ay2BgnCC+33T
lB9o+fdfE94XfdPDbK09nrMONYBXCKskurEoGBzA8KicrE9c+1p0Xb6jk+F2ZhGs
ScL1G9rvhEyZN6+0hXrcd4x8MVxjkSYaIOLKmoc//bnNV82JNLCuswiHgaBuouhZ
hMnEvr0MtXRhIrPjQ+e0iHOracYJFHZZss+6hvhzKj6VvZuBKD8KV9MH6xbc136G
iyM+5R+v8J1RAmRCW4Y5FY2LRiRFXRYfN+H/Z68rs11pixU2L83GdZqO64vmhu4j
tee2ZfX6cEzH+0Dt7LCZrbjjGmLatfk96cfM0SbY71leOgVQvIIUzoNkEotqGNWp
OemnV86RRMn9Y40GSwqS/0ZhlEeUcaKSU3O/dH3ebLCXml62dF2OQwwQWkNoicw6
VTlpnGBUMMddxYMLKcqPQM3TF+PPSemfLg5YeKp3TxsLWy3SHSXw49xtjnmZ+H64
QyCf9CD1EWGnObg6sk+SMLRVCEYQ8aF7RXqRpHJnfeTS0Wzsn6SBcxnjMQ5GdmIz
+9LpyaQ6zOywxyIwv0zjfO6HSRxAX2hCEhOSlfrsigJsuHiwpWWziE1QAtIGzW6p
4elNE1uhxwdAZV1gcO9g/OMKIyycd0uSvNfeeu6hV8lmuxt4gKxgYpABq/XuBJHP
cVUVSMGEnlpr5rBnBRjafil6aoGwmnEh90wdisF+Fyp14gpnp0I+dg3I2iTJcpNX
zaWU0nGmc6BqtKIbYNNqY/9EnAT5R5q0ez5lphc1juLASSJJACN362K2vg0dzm91
IOXrxb46aL8t4YsK2Gqnu9WTY405YSqXv/pIOPx6r4/wv301Ejyy/0L9m4snVfrn
P4oIVvsujY1xQsmdw11gfSwCTdlmnxGwLErDIi2+W4qGsrM6ZXuLO82224C3cFc3
q+/GykU6/ozKtffpxs3v1a2kNQJeMBb4KNd7M2xqxBGQ6L816GuTRLokg6MeYUV8
9qERZgmrDqwqWMT0CJfA6VmL4dttw/Z7IkIYemYRj1gEqKmvfGfo7edNVeKvOST0
D9f5e15+mVCS/JUWehJCSl41Lsjdvn+O+RM66B0Oz7xTONHjVkgc8K5yaFFfW7RO
z5D++8t3T0ulghlltz/iHHUTnANUdAbQcXy0TJ0dSwEIz2bivEomkvoIM2KGRdZ3
S7LdDqcv2hdmzFxTWrQAK2DMCnwxnTARYGmKb4FAtXEbg69ak7g3dBnXLDsn2ywX
qz2DkyQ86rOzmB65gMhEXTPSP/yeRbLtA5EHjTAmguibdcP84Ng9XOMZ5Zu5MRL/
jrI6pOktQTcOdObPGal77jA5upPJN1mWRq8TGxt0g5PJTkqmhB0axvXe9ksuzUUx
ErsrLdRSk3xGgFCu1vWv+CC5+ZMvLqwlcRPpjH7B+r5TkHR/7qF2U6NtfXYogrZJ
z+t4xaPztKTkVr/4S+25Owi8C0ASZROkZ9mUr4dM0RdflIrnVixyCj1GLhbFaAw3
qPBToIY9aer18HDSwQWuXllEPyod5q3WDeyvUZaTQZzv26hd/ZxRdE7IQ3AlGjDU
RznniaIPf0PcrArruVkZIs6l1GLKwZsXKJ07Zyc2/KVATPKwSwGUWhaTOILIQaE+
FEKiAsJErafIUvmmWfxtMqjMQaotYARZrAYPGUSMMYDCfaymn9SZRof2DKZtXM+3
szxWBTFbC6xTq/nqHuBzUwVcQcYjpdL8TH80VyJ60iOvRnaQf8Jzp00blPV2gupr
ip2kdR/D6QQN1Jn45fSDEZQNfarGqvg7ZM6aqTo8FYBu/WSivTlvzy9/1ujxSM2f
5720tYdS6kt0FiBkDeDDXjQ8aRU2dha7JlJDmka0us8e3PXclwY6qeRiCidmlWPf
p8ztZCgZjUIC0TkUHGqbalLmmUNqxFnFfMbUv5CEitcGixKm2z41q6+EOdX0cvQk
0Q9c9VDipqvSy0DZfjF2ylfGoxJzqDmdQmHHnXBLM1Z7RMIYEzAaczS2rPPcxPne
RVUoxrEsQouTN3+M0Pux+vO8olZs4aoOPxawd+St4gvqAE/79NRSFsJmUF6y4QVV
f6GHUHHSBwe8mXzkV04EFrsoE0iLm0TfzoO7AQXDRfPk6nO7JmsKddMgIhQz7CtZ
qojzv9qHEdAGocNkT6sKv0z4+y4eZGsJTirhaOC/HScpyd224tRDgtEFn9ynin0M
r0Qgyb1x2UZ8pTpXKtVA2VkgyQLIIEaDGqcZV2njTPuTbWgUtQQ1svPfC06k84eR
stVGLWf/fyMJiDuz3LvsFPmly5V7TOq2/A4D+6Nloxxq39CjKBkShfR0rQWUq5Fj
BJi36LtXYqS6dRE9wJfLrn4PKUOjb1iyArUfyyj/V0JGIH0Vb7iyiCFcckzDEM6q
fb/0xEIGIb/fjK5P4N+pHlVc3wg4hWssnN5Gh9YQSnmQ2V4oX9KbI5oBBz1x2Qox
vb71YALSdQnMkModEEuQfH14kzNRsj+AXfpSE95OkwzmUXlBcTI6kGS+jI5JAwbw
H2OzPyRRP3HwSguo7TR/tfGg+YDxbwpbrnaPss1CxECrvpHrLcBgPcLpE6lokYs3
ucTjSIXX1CaianKkdu0ZZ7oSBT65DPM4p/RzODQaPIKgwxwMJo6vU5IO8rOAuaTh
Ll0ywv7jEL6QmalGdspMVsn8CVzCMxHliBEyrm37ZxUpiMFzBGUqGhSDIHFjvvcO
nVncQwg4y3kCsmLLuvO6KSd1NCZ9R6DUnxOQqIZCCx26HxFKOqbnjsV584UGCD5U
/yslrOuKX2MypLR/xsGVcg==
`protect end_protected
