-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
csUkcsi0IHsf2aCgGdVP1NAroYpD8RAewGiioAC/Mfw0OMkxkcul3M88oa5U9Gf7
/pWtp0vgkRGyX9EBwFXQJQrYRPnJqerVYIo5PL1/4G3MJZ7sMBNqwsnBt4uDuipW
Mnj1ysDQWykLc6U9nPuZTKCBUOCxajcTKejWAQzOUYc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9408)
`protect data_block
wwHQ7QoMqwYo9UkGSe+jSmQigClBfsZZZby+kDfyLW9XOUy4uX2spIithUOqqYpY
QaWFNl0eProQvJZUCGUA06D0mwBHcbOL9LxtNMNnLQLqYg9voZ0GpXHiROxLxSRw
IA0HPwhgkDTNob+LZ45sWYsJCPg8E/pMVCkqpEA9GYDrxkth9XwMI0sjVlpWWlDa
SBK3V2/shDDgCbqJIpfip/2niZF4IMqWiS3ThtLCv7D/mN+Z+ruuClLv3IbzMufQ
u16EDEKzY+8AgUs6LFsZXQkyNbcu1thi4GgF5FgoMJi9hFOOsWa5kTmSfOjYFaQy
aMcVG3THIr36NmxEPGEb+ndQYRNeqqL4GpwSzo2eveoyZAkYrp1V6viCGNK7v/cJ
GKM34OOQwjTo18j1giDITPQdTBV1EQxAQO6vzhGLyvROh0r5OiqahUV8eb/R6T/v
bw4YRr5ljWc5wzAJVOT3VDlosB9YarwVnVqyTiRjAwvaASslw5HaXSrShZNobtmp
slipa1uFb+f63DFK8mldFUB2SiLERKB4bk4L1g4C3yjNG1BpLQ354K5NZ7fVWzC0
E9Pb+JTWtt7qY7pZP1dc3BhsPZwxo508AYtqk/2BNzjiyps1IA7YpS5f8aeb8Dtr
JUquImcrrewdnEaCr1PnvnLVK6dHK7JhtoZEAloSP9foAut6oIo9WQRaQ+QQVAKW
oc+XgvWMj2GfA/rkEpWKYktAEFiRRt0IxFR5tJ3gkqjasQG1WmTHCSVTxDwqiUS/
zwDjvmFeoXCgzUCgt8lOvlcR7DAUtGaaO42aaw35KtLXdkriTeBokHQk2JErTC6E
kvBcRBG7sjAKPL17tTTpOQJaFp22ECZxryrqfFRyikMITGlbXnekoOhcMcnWOUOS
pcqEaRMq8mUaNS2hFacU2jriD7+Vok3pPYhKqsVTYagPf0tgIhrjkQeeSYNEQ0UC
/Dkz1YEF4MJvp8PM/iynyuAQ/31VIO/4WBLlS1oej06FFO24txjdq2Fl5eUQ3mGU
0uF/+/GO0tIrFuiRP46WM14CEvQscBBo60In4h57Xdlx8+uZ0TccTYbziBhq9Dlr
u8G3lZK+nxEBvRhzez7R5+DB5aml62m3yIoSxvY7ZTR2Zqo+StYLYekuGkl43eTL
B07sEc3usDFXy3Q6OIt0buihK3s6E1yXjP1tSN6bKTSEQgvelm0xxbss2TX5RyYy
+VKUgAIW51HePH88rJaIEDXpywfjtczckgfcJ3QO+rFWS9YR/vxgRS/yQP1ImZGH
8afwqbsC2/qEODN0Pv6dMxpiQpxA4qr/GJ6d75ea80raZw774OfNZlYYlAqDEaKA
aRiYy6lBsUlOiURbKlJyPXQxx+K+X4GlXzBFKEUOZzLU0yigLCQQkDnJvg1sqaGB
4mjBo7TA+QLHEAY4PamUuDmwlxgwpIQbqS7J3368Rc/9E4ITfwtfmYWg65lYCEfd
9FLaBRp2ftaPqrC/15FNPxJ3DKNAaHTqYuisLurND3R1lDkxg3jnGO1m+lRZ1L9O
0Gkaym910rAbFqaq+Z3ObHiP6/RjzRS5NI1ieF/V3ehL8u1gknL8VA5JtAEbaH0R
nTRHFV0SjvsnzAaSR9XNVxYRehFM6FAKSi4hEx97RAYe3kJvHp/JxywmbX0oVpoW
T7WWv3Cl3K7renBT9048/z1NG7HSaY8Y6gOH6HkLmjQu49ula3H58ApzXhTRtA+D
AA8kcyDDKg4XzBBANemEokqgQhKGXXIOKp0HCuhateKiy1vgR1aE1reF3jIwY8Ah
5KJE0LugloPa+cH8p+R9NgKRPXEoOcxRnbWGaBlsyZD0qeF9QIZEVacpjPSHYKjP
YV+WXTv5wYunhig5LJhxE6zRyar+1xjtgv54PrrcK9qEC0pCuqvnf21surOA+WOX
CoXcxJ6RigbF7v+cS+w2K5or9sn64TFV2ZG5ULHoMZXX1vVRkuVHwH7UHCAEHA0B
zH9V2KtFI+/JUFbpGjoZwy0l66WbbZkDKi7LnKfWfcaIPYoZ0q2FZ9J4QyyfhTk7
D51niAV9gxeJiHmvTfymF+uTZ2gp6AwKwChR/VroCKnnQk+o2db0B1WQdkjPpPHT
2YWirbf1/bkAgbPYlfU/xxdgZGKJQBIKVdG6nMW1zVF14OoMkEA59NZt3AMST9Iu
OVHHVSY7N8DVptU4DwPu+BR3i7c5rsOlY9NAl0AQjsT8HGGKpC03TWTIfj6IEn7n
u8sOfNKApeRY4g0KL7LFJVal70UjXV0ADnZBPaTytkKfdv8x7YVbLk3QIXCH+uD/
mM8F8phzsGrNGELynQ2zvoy6A1/oGYfSrsRxOgimu82sbypnSls78oj3f6QtfChB
Ea9zbfPjLORJoM+95ppLVMNPSnlNHiyL50am6sEptPTf7/nehnuNe277Yp8WT74F
oopw/bdp0j6VSQ8UKz3b3DZYKcAB+cA75xEdTWvA3x9G/Es4q+0mGl5mF5DdORVu
3iG7T0Ab5U5A1mqgcjdor/Z3zUpP8FcqBS8qE9ur5/En58ALXslhzDML9Kcwdnd/
Frw/Mx/b7RDGAS33VnuaJRXYWv5A9+wse1FHrCex40cnrE9IZGQQaGQiKuCDgYSX
6IPlVD8i3/newpPk4QMj8cXGTg9wWRib5Ivb73q7dFSIL+X9YLUSf/BnYazSAylA
8t8Z+IU8Ax4H8zxvp8LcVtyCQC5pBiUdsq8Y7fUoELxvZhVvAta5aOq2khP2sW5U
GsQbm2QCtznsnG9u0Px9PrQTH7StgRhWLOSnekVu7xShC7lZYDM2BSLF3cJWRTcP
gP0+zIAfrg1PiB+vv86ma1sv7r/kSROXwPkvbXEXgCAdj4Id293olq6PYP3Jq04y
sns6g6SpBsKQTDtuKT802WfSDMQNIFt+tWR70Xu9h4tBzZYXEOQqduKtYRYD3Z/s
nuwqmruwcBow1Bw6H5caOoPNyieDsQ7CkiC3yj/+jBpxvTsPpdYdJ2DgqSYr5/T0
OTqy2nCOvlGQ7B+okfu7I99tyQnDnqL6TJwaKLAcdSwh1qH8GKiTIfFloZmFirEl
ksOMBLKOmPFn5ABv8yuRA+HnBeV/oGt6zAaXp2dUgdw9j1WcA/r5HjmEcjtD5bm7
+w8Ti0XJ754FWhpD1W9XJMZQDK4FC6heHZGlZHJQwVPpFWCRVDOjzc41nxw+hHrc
KOXn6Ud+i7eJ1WAI38v7ifnCwZmFyRdaYO+q6JMwVdfpcmdSysLLUiISaaUnGsuG
k887cWn4Rv3Mh54gT+QFO8BYjilelJoK+F9+7toOroTzU89TZw7QlZNqM3cCCqLW
shLNrVmkCOgJLXRUtv19Dag7bSEu+PbJDQcBntgsvbzvs461lWliUhb6+KxiPhbd
o8rPEKYHZRe38gPhHGthrCYmJR5U+jEMhXc+d7mnRyfyvgV9Q9Oy8iH62EBaH8Zx
8R0fBNt2M+ITabYMQ2YXG6f/3l+sUemmUw1sU+77Cg++Qjn1mHF0qdLzAdajxhE0
cQhaEn848Hq14bNPFt5/oSdjWUTPeL2e0IGOc/JSfjygmmzih5oiqZhDoa+W+/Ko
HbEmLMU1qSWKWiM46bxuVxGtexTRpatm1rQZIU5aIFYOKiJXJjFpBrKuEwTEFxc3
Zk6UsNpOJ7sPEGUsBF1+5p0zTgZqSTbEYBXSdbkvLAK4o9gEytCiSUBzSm4Ognfx
H+g1/S5hIf+aN+Q6/16pn1CqxBvVVHIc6ITi5MTUUg5vLlo8UmdE6Nwgalj2xktk
FAtpv+K4fSJzjUM2FDRQR+vZlAx9UGewwcbvlUoc5lv66x3RmVjvHeDZYoWISxzN
t8qQr9rLrNrF5S3f9cPm03dcjS8V39JMoh8veiGayi5cDkUW5i/Z60SyjgJBuFfz
9r7r1yVJc+4gU0HU+dWl98UJa817RIN7rxdOGaP5ctI0zMdszxNMo9sUbRcxoaep
I251IA3kLMnxDtRPm+QEZeeBkjTpZbQcQgPZS/ZvVFIVDJP2Q/JjlJGhqblGnCjK
HhKHrBjxPXzv+vidU+Ac7nOchcaM9IDBGYlJOLgzIpoKEnGbBFtB1IFTNSK+JQ8o
d/yfCKzTutRaq+mdGQaCXLHA9gs9sIFxKSeGEpUYlWlszOhPltrWCTePk3YHv3uR
t3p4BepzR0+273bEpGgosU0X4FJ8VoqiLJlknOa/WRsDh5+ZbKRByGPjtMsXtGQF
GUqgafosJigWCVrDvPtTSqTZTmqXIo/9mOIDE5bWtB4IzYL/rNHz2xllsRmW4+G+
57DcfgU1ggxhrFK+nZA0JXuOHaj/0/BEwBHYRQwkNYTStctJy6ES7RVSQxCnZY6k
2HSR+zZ3I3RuYUUA3EJQ0aihBGhq9PPnLhf81JORvbE4BaoLcbUvaRAVomwItztW
lAxJd+naNHSKA9cG6UbnZlmLpmMZz+GnvxJeH8YFVKOFzJmwQzUK51tYtODlxAht
6xKT4s+loufa7hI1ByRcnIwSXWK/++pz9FVT/fv2iSpQT9Wzap/dWEWvuJYZ61YO
oI0ICWmAnAqJO8XJRwAIbVNeHh8k2j93z6Ph/l5spNeBQTrmDhO1uWvuDBZOYZn0
FqxVd1N2XDvGevkd6SMacWppT0+tG6icCwYgCfrBggb9XfiLQ9F5jGS+VyUshkAB
6Je5HIytl1cVDoctUxNSiA6kLXnGqTvjy5ZIZ+JL5uPy9MqxWyiWB6usysepciGc
Qo3pR48pFg70UNTfNf2ir5Oate4qOS0p43QDLOLN0WfSb9tGiDuA0mfwDhCxU50M
32LApEOknTyXFHT44adDijwG+0Cu2Kh2hNt0oR9sBIFP8YFjbSt1VAjeoyc9RkPp
/N+ECyfLOgWJg+bATfQ+jLWND5eIxl9e9hXwGYQN6UvErRhjkwUh2X787TALLAOi
tzKif4Q7NuxhtBfyd/FteGk8p9QbCA+92p5G6clqlA8tV1H0j1/69aSoIX7GsnNf
PMWVmWstsj/T4GpNgzytrmDvUbf6QX13kZZuHMyWkZ5UXShcK5rY1jXk5mL4l+Yv
sEuJDzj631Y6e7JNYRfTlI3E/khny4/iwBdo9j2b4NacIBDinJCNa5WaQGFapE+q
tHhreapUBJjrbJ5QM0kGiw0lwFH9oPJ8KS/XCbPZp5FLWOF2jM5cEhINZWMrmHgw
7eg/1GiF7dnFykyhw8ApS1L6yvGH8THkkF4fHQoMr+ml6+ATBTx2QTg8cQLmNy/N
Pux21MuQmBAeRB9FXv/KRmwazikgUUnl6LHhcUeyCQNkbJcW5HLHHkkHBKO0kxTo
XU2MgS84FBdVGd35qcUiA1QcMqN+adkY/EciAJricMl2WRKhWYZJeCdqKokTWzTK
Qes16Pbgg8bkMooJLNXpm00GcRXDI+xd/YwpUufW/nZb5ztaZuaIBMsnkkmFRnxq
j9vv8yVikEKOohEeeYQjkAmQzlm/KLXRSKiOvV7NYm4FponN9ZP6hXZCsBwzj+Co
oywt4rbrJhoq7dCAM3pPQ9ph0+ILtYX3Z/9f1DCnD4zY0McudZg49/R1lt27sthR
whfa+2yHniwvMTmOhSsmN+HcpFv2rEfHy/fzDK3iuHvyItYTfq58SeQTpLT1yjnM
G57fXQXuYvBXlkhbjpmQok+oNvPh8/D605GWr5so9uUpTa1Ick2hZhS9tUPa3diP
LchM8n/h78Mt7aiwTO7VCXm4PzK/5LunwX9Bt2yXGQFLrT9HpzBVGz230dt5qfME
sApQZ4NUucyjM2571LDDKZ/znpqLCOv110AqSOQoCA63MREj1+0Ex46117m298U1
YBOPVvPj5iWIUsggN8YaRRZ9yrmHwymlTH/OMqWto3kJMJ72LCvSbW/HsQqcpxKS
UGabu/61ZYqYJLA6W9fz/cxwbGCRSvHY12phJIS8OzRs0Y8tSFfF0dXeJQONjUNE
V93Jewur6Ok4Mi7Mrt3PxSnV/+yW9FegebqMuZEcqbM2gVyzm8LBPtlSnk4iACxK
s1JaAxW1sYrOLntWHPLfgLj7YVdtXDOv4iCUJ6MGfaFrhLI2G8NJP2whFDeQ+rSL
pOMFzNtE6JCg8qXf8eKoIYcjhQbOBBmRa3kiydU+4a3YQIha/R2hXQZPXeQTz4sm
27SyxJiEGZdgRuQ+Kqwpa+qXI7bSFjbT+oBgKwF7HIwqxn9n5QYivbCaXR8fpMGp
ZS6cqq8c0vGR8ttZEogkAxfKObpdk1bwYHBNKhgv06Fn3Qe+5hAuFlT4N6iTDrR6
FExErF8UHTR3Uy8ZSwoZbNwDVGsKg8dS5UV6YtTWRNVNGMG34jkrfmTNvsA7iNBo
LlAMYZfYq71lb5MinkTm5FtdCDxbRMIJdhmNWspwYZ7USf+BRVpWuHPSIsHMK+J8
gLMjIqXO6LyvWnkqFL0syidM9irrppaTsea4EVONdPQZG/dB1f5yRt1HwqwAlHnE
QhBi0VxRXmSFlxyA9to6Pr8I56dd2w0RVnilPpWP2gzB+4pFAspo6DczK8T9YI0I
BetiaecIQhtQl62bQ1Tg+xtp5rHPz8hdRILUyKqf81z43sOkTu9pHo3GaNI1urDs
bKjdSO9g3YHa+fE3wAPoASdb/WV+S7hhv/O7TaBQzRFrw4txcV2Rt8jTQtbGmi1W
0GtA+M9byw7HV1ptiFOeL3lIFxivAx0yMQ6vpI4m7Gajs1AT2M9M8ltG3RUaN4XV
wIvT6UdkMb3JUuZOPqA/yZ7R5fHh8p3hRL/sU0oswpKrjBHZuRKW2DG1ZwD0rrdB
3a0jYks8SJcSKlXJdMlNOF3Z3yr797+qIGPkNIM50Allp8Yp45XEXbDLr1pjSEyd
tsQSl8pSX/QB5SUxJnz4Xp39uFjOQLf2gVLPMERTb5iInBiMChA39JlpnPH6ZeY8
HCHF41iFhhfWllJWam05VUUFwiFj7odvuLtqqJZ8RCgQGElsRmy8TmNyGXeg2Cob
t2wy5E/nlDOFrsH2Oik9WgHr9j0xZMDkYPv8UknSq4LtR0+BIB4ge0kzHmUY7/Aj
BIkCGx/j/1xHw4durn5oUR4UTlPy4l/vlMBvzbi3feGJCoTkWBfTaNBxOVJCnbA+
rQL4lpWZTG32IrfQqygo56n9NaLMRF4l1xe43yrxOZPZJCfB2PpQrJj2jBfhDhBN
7a4WJrupOcPCjoZPlhwluOdvULTQbw7Wae5oZwFoCCq5cQy2mVp0nf4OF5q7PHv6
m5I4UNrT2nbpJy3ZLcYfcl4SW3iQ3pXYxfyFu87r8HDAfcV0TQnrD3VD7MHL7QB0
4LF0Dyakb9GiNsawyHv3ILycogwARZy2z2o/w0ftd0z6nvpEH0Lg9qdtSm6Ujh6H
ZL7JyO5PGIU+jOcd38fTYK39HG76PD19DPCIdOOBYXdxIa7QuPcFS5THUOURhTB+
gPl4o/ukzkEoOwYe6NpWrjILZd8wpqPmTtZT7gTmraQJAhzKddPAxyxIbcipaJ4d
TzV1sFvOtnl3UVwt6AYOxV6SwIMaGwmGXPUCeYy/NRYFhbTuUY4bSrhWcaWOSguR
Y0eE9o+ESXBuMAZcNYwF27ZIfR76Mjw9+ao+GNwnfOiqFt1uszxdYmkZLWzZe/bS
rdLFuxJnb3mZoLutjrbW6o0yDlY3qRUyCIaoOPjujYA4QXrdLK1Q6v4/3Qj7dOBG
hQG4xQ8q1p/PLquOQ6TNrYa0HFAV/B+SmhaRjOoS0xzc1D610DqXolkpNHdPnfNN
8GWGvI1eOvnnGn8xSaHObOSXo2UDcL1hkghcw7PWa87gX+XbUTysHVlNrHDViwk1
k/hPU6meeh2FLlknvlkbEVsiOlE9p8DQvRZd9iCd03Mu3utRu8ByOsOjnSxbS28C
fysmtwjvo8jior84tjyimqwlE4uGu7I4NssFiQ1Dvd0NlQawpGdm1w+Qm31mhgvD
l9qQH17YR0pLvTRK8ciL5KUfOnMQzRqB6yXzjV6QClfh7UNcla80NhaBE2RNb82k
fAImQyL6xVku992q34JNU4Yjb1Do8o4cDEMAJ8JH1uKtjPWsA/AZ5MQ+A8JFzlX2
tcAwkZlDkeiTHDykxM5HutO6ZH1aT2tdt7VlTyDtnV6OEh99s5R8ImksTFkzmHeK
n6H+ZMiNXUBXPQ5UiqHq4BYYHprvf/53yek8JRPNFcgCFfPB55HHT3MBWN2NkTU9
oYl8E2kQ2IuXpq+i4Z+IJ69hdvM25713y+0s6XvhnS6rf6a+wSP03cM3xRwnlcQm
FQVIC6/lrHBRqDFjnECQDQcOR6bnFHx0Oewo4TJCF3ToNBQQqvDakl52ZrADY6DY
CM5wf5mAv5A5bZocG9VFQnDZ5fcCgtpcgbQUm3wNflkZ5DppNrHGnpouEqVxb53P
P7ITDxEewQWlyqYLSV7J9ntuJonhoKFAZhD0D2TiiUHWAl5Em3jHnYo7rZLo03FM
RJy/QAbvbSesrK2ekbaYadzdyn8238vePtBhN8OmErX80pkzMEi/RkyNikx2/EiO
tJWTyMin6zpgugcD9xBhXuO19TzSoexumRV3GrNIqxHevwIK69iMeREMURSngUac
yhO/qHWmLIiOSlmBg0CTqDM7hbzCoKB1UpCLQPGGPPCl5e2+7boXY1KjOyJMtSKN
dCV9EXWYtuiso0zqr07b6LARqXuPN7EK4VdLKxfF3IDsYJ5tNN4mUWz8S1gaJ8cZ
PHjEWhoy2j5TlrYZLv6LtWc7+/8NtsQyLsFgbvdVyEiCVP3ee0E6JfW2O8hRBVyr
1sTib04wsEZWScTaza8KsfwFCcFL0FOz2RmEkmj6a/z/bjLO2/xKv0yg+10Wv7VN
YSimThfzvwEHaLUnMNtC5pXcin780vSIQ85HO0phbtX0faRuMHAMKp47k7vDssZT
9HJ4h4aoz5qhjmiO9Vk6BJsW9d9W1zDbGjDpIpsak6I7CJjVVuAdh4+oM03Kpx++
AP+wvqiT+NVChwsuc1gSKl/pkCk3f+K0XPUaRKXJaiC2sB8b6695TweRVs60/Fsz
x5BGu1ZII/iJ4yEbyQw0AKngbay4rgQ1Xe10CUo6CFm0j9Zn2iIvSIBrskwAdY84
sCQ+qWVIbEYr/og/04NQVUWzrPR0ePFlfROKLqCdGVu45UbiLy3RnzHuBCAXUkY+
t83ym7s6jMMmBYDgCO0z41OXA5B/fk+dyuATa1UxBYrWxt72ofFb3aVvr2jm4yRd
gpBozkCVXmYeMdcX8l5xPib/lEjFeF8sN0jGy3HT1cULlcoq2mLZGapn8XWcmr1O
6VXR+tRgeAWJnXOoxvTj8UV0+Jb1sfxyvRI22GwtnOL69MwRaDUKNaQmdxXPzhkf
Q9Sdw2C85jf2vZMS1PCiBoRVJ+SSS3nF5i8zMMl34PmpgJIV2j7s6+NVF43d2dQ5
H9WzKQMQ5Dg9aNZV99syQ1MSFfefERIuyZ5CQGaZLzcGTgBvRrDIrP65FUB4pGoE
HunKj1itV1bVWlVgblidcJkv7shA7zAhVsgnzlDsYXUWSGK4P3OQ6Nh6OWhMRKrd
tCn6em3oPVkNZeU8L42lL4lfS+okAJPskQwuHawvrrxVS/VzkLkj2auQIy4YK9jV
KXME+6V5+sriaeJhgrMeIogQbL8sSqD4gXU8OmnWmijRZVdBZgHC4dmfrfU0yunv
FCs5SKjgZNdY/t5hVNTp+loqqmYbolVISwcMXitNfXyT8qKKfaYLQL3y/6zlBoKh
qhm+AJloLGVfFnSOKAh+9W8IDOmZyQMX6DjQIbt9bRdmYXSOQpzvt/Pv0A7GLw3d
BqRWHWtFHSc/W97tnXjuX0lA/QSmOeT87iokhjctGHfLYAMu1e2MJM+yelBscNNW
LAKamRSEgS4gCeuNt5F4FmmAwiZef74aCwWhyzD8++CYUDkfEsJoEMKiTrB9bev5
gbiAQHsKpwwYKPxvnquUJU5vsNB5xd3iveHzSLAcncuoXzyFHr9si+ix1Shed+Zw
DHMmPn3y9oz+kcc8XKoZZyOwdnlyBS/ScYyhKoSmcbNG9BwkZfNEQxujXsuyUktc
vRtz6Myo2I46sPsmXHrFnm5YFWwxcWRaZiGxsiQI6NxRPlXocq8KCMrO5q2hOKr3
jgU0oCGMM23Y2ddrMzzXMGetg+ihmxBkfKPEfiZeH9Ze8UZQZPjPN+EjiWOG0iUp
LmTlCPGYWM52M93Zsx3XyS5WMyGmi/qXaRjVHAvv6yT4StbyjT4jA/wxMJhbaFkI
6CrTJhnmb8jP+TnHMjPCG8qcWuuStKLoI/Zn0yugfIMhOWAar21ubaAygXoyPqnT
jFaHm/+OiXxvaOCTUyDO+Lm8+choiysKwqDxmzm4FUGUJz6x7hNsizDmN6LOwGqK
vFpLiZgNSWD0y5FcE0tn1rZy+u17twER12KauhOz4WVvTk/uCdpTyMX2atK6klKK
Z7PJC/nOGhvMh2J3s7623EZcTzTLBGXsgztwS1+fgDzdEQSxEAPIXiKc7N1dh21o
HDG0XMcTH0ybFgzKaRdmRsMNt+94LVPezmE7IQo7jm454BnOll6jx6sxG2sFtGEa
VTmMMHGdJDbU1p3dA/mgMthZfUSF3rKM7h16I2POnxNvOj+Nqq5iMXXKmQQBIckZ
dt3bfKypDQ0IfT109UwG7IWH+pLAJJutdlXHBkCbfjqNrUEl/xcNDX4MO0MkMCX0
FJb8c1+adQAjtojNsXrjvqdY57ZxqWK9o7H1H/g+Ir+zrHFWguNnfXbu4ewJBzZr
r/xMRk3b5hvNe5e8+0K1kOQpzrRMFccrojCjbQ7ysE3OfmTe85NkqzJOllzaHLes
NgNUlVNec8jHqPE7jwpFdduozWYumHnXpsSOZMxUS+lDtwcAZrLJzHR0udV1F+RQ
MJwcXiDE4HxZfuEqVosHvTTfsbp7QhuBUBXtXF1n6ZAw9WxGBH3LsqdlO6+Y+6wX
Nm52bBCPcPaxz0u6vB/xMHC1hB5q7aq6MfBHQh4oFiNf+6eK2zvHKRfNV2DZcNob
RI2DSL8k65ZGvKs0bEh30eVL/p96fmoe0d0Mmuo0akHKn/kvUXlxDf31a5hUAgU+
925RjInUE3WCgnuS/xZqWKqhYpFx76kxDoPSkDHOo8pEorcJnagqPU0KP1g3wL46
URp1w7as/iEepH+CExoM2eiM4O4QZupFMxQnPsGKDkiMhT8bJ1pyEeuXCxOPER9p
9yDKtkwFhFTPjqgjMBRuQ9m/dTO9sau55OalJWEEsliYwjgtgfJjNKr41AKXoizF
w1w7PWDHQ85erxZR6tfevOIZ5kYxAf+M6QI5ooQRUbsi2NOth6rM2Xa9gNtje2Ky
F3q3maPJJsTFiZyZrgdwXvEwO8qJ3NMW97WHpNmZAtsMjsFzMdFDtiUgiyE3s6aj
pLTrAaTDI7bwtk9brW17vNVakrWSEx6CMvbJVOXIiOh6k+r7bgoCvPh5srALdHKi
/CIW3MKP0xDVGvIMOJZnSZRmrJBxKbFX4n4IJ+mJpv9qhqG4hARmX4Z4CkahSV1W
atSCwXAZyCdN6i2azXb6WS6QqpnsGXRIT9DUxH8qdutweVAYc0FO8mqOaU9RRYQT
RKZskd6jZJdi+Tw1GH9o9EN868oWC+SXe9HKVPY1b1hFrPr/MDgX0wPkBeVi7769
t7bTgnlLtQMQbeQLDamxTvhMn3iTNV+qzwjMXNdvDjzO7UfcIq1u+wE0k0ADPAxm
p4ijr0Pi0UVfJN0eyFCWDMs2SPNrWiiP4Xi3k8Kdun17XIA+blxRaNPUpvm95AeG
wl9jfQ1WFb2QawDvOy1AMczn/dOfZO0dPvWULiBHIfJx8U4fK2tJiKXO8RW9Gs3o
f9DAi0zVIc/h9SQJ7o+kb3jpy4nBIV21z5dJ1qDjuZikEL5WsCbEZdgxCuKQfqGE
SUMJBaThbqRZM7qVLiDhPMkVQ2X1sUxxiudqimqtl2uot8m7Z0slaVYzV+DpcEoC
vJDPvhnBukBbFUSfDwV7Vkw/SmV/HifpqnspfEB+Pjiut7K23uCENao4BlFYL2Tl
Dt7IigQjDRa5KfaPUzmyiUSdyZPVKnaY4I03ESBzCXUMQRRqVYj8vyy9V4aA41YS
1JHwhFTPu5N0zf2RODv1M2wUJDmomOFMi/i+xoTH8ZH29McKXGZuOQZ7sIFTvqCx
aQ94/hzx/QWSaX+N/nWlNTJO/IV6LEonNXz2FLNji1sSTSr2fq1xqpyDCWfH6lYv
bgy7qhSgHrJ5NbGxtM8VrBBThznHLLBvfbMtlXjeptaU9nb2lkulZhiFn/OhMs/l
/Lxrhf6VGLxUta0a3btj+uYY4EU2SNtpqPUAZKY4ry2iCqWRfcJ8A7NtWgWr3Rzc
E7VOUKrPPgtHa311ZwzMPm6UnCMf+FZ4XE3ZbvwEbZeS8oV+2HJg+looF3b0UMLj
qBR1jQLvBvBVPUTkCPR8Q/68uIUtYP1LK9TsB0BL87QdnJudLhyKO+n287RSzhyv
7Q+KvAphhhDwFdvk3RdjOudcwTWCPGBxAFmDpQP9Xp+128WqGhg7fj+dhcZF4Xcr
`protect end_protected
