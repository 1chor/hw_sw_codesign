-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
cC4rDi6RRzHlI12Ap8RmnrN/yg7SNrQaaTOFxrzyO+XStlDIECYnkbPQRZqeKv18
qMPUr0f/272n/2GBqd8mAjLQh3xtZ+v6h/ztTlOoqiZB0vqAOPI2h+Ccssj4xBbB
0mETxwb2LPhTZk8GdEhJR15qvYhaKKgW0eOgN3n4JR1M1ewoPHxdng==
--pragma protect end_key_block
--pragma protect digest_block
hG2fAIgIwcCZbTXcNlWb0v+rJ+I=
--pragma protect end_digest_block
--pragma protect data_block
jC7IyJbBrP0T1LqEawGHrBzAr8tRH6y7YN5/qoDJQIxuj0EEGyupNwaJQXve0QPx
J3O4fAfuwUKF66HiJvfDTkL5DvMhrLn9lyRbz20ijaB809OC2OpptchASChS4jUO
ZpGfEF8AH3sPkYWCibK6SfQi2Ja9f1e6hEOr2Wbpv0um/Ac9DRHNKreUFcGBHmiG
uDfFFQtvp3mepjjHF0wEbg/jUAYv5cK6tQJ+sc6wBr5Obxe6FJ9lOY7sxE0jKFcr
sLq55S9oNK8YXFbUlPVOiQj4uobOdb/rzqZb2vmUiGEIVSrY+8LHL2b1oF/kKB1d
m3z9A6whnz9bHRuVMoE0CsteXqbW2bGEWC+tvq4YpP9PReMknR5QLQiF7eD6HNBS
5mwbf8JZwLNI33WICGhTN5jFzmXA1pojeoL87gESWz9QH0LSxBmooNJ3H6R1YJbG
jH/wq09pbPuWbnA356Kuq7cmPhDeJwzkSsGbDmm2IfxvMzRKwHpXnCzzVo6UB1UP
pFZW19ctpFXkt9AFxmJlU6R7noE3nN6YpEY+x25j5Az+ZSE+3r60NOjPGkqOos9p
0+lsw2ztDxIbHdjSR6YWU8+mA31im//uvJv0snk4YcMphjPcLoj/0S1QRBCl9tNI
3Zrd34IludqjsfXVuwWYh6Lz6hyNNIoRQtEY9cAcn1NjI6iZO/9jo9YbJIgOuTtH
u7pn39A0T1oDkfYXPDmBd8dHOKH/bgivbxMy0c6sOuCF8X4+94LJdJVWUCWzoJDS
P1Mtp2kejMW+skQqTKu7nFfnbtZfqstmxAWLf7S73liLJKlwJzGyRbMoIoKV3h6+
+nocy4rL7Jvz3Zth0i0VenqchtdDzFUo2A6eEkLCZ0IzOsCosmqNAU8tY9iwktme
sFTwNOTr/YtASch02Lr48IqSxdcEMQ8Mk4PInh6MwJgsQPE9k/SDwVpm/pQg2C3Y
K5g89Ran0G6PI7t7g3lUDypKEiwr6SIZrQg5pRmsJyfZHs4F5H81dWZ98a4pxUiO
a6Z9r9/p1V2NpZsPxOuAdfVxIHpIJ4Yq/QLpbo6osuCe41l2O3xw7L0wvPj+ApOO
YO3s6dn99leff/PtZy/hOHNwEd9leKhKX9qqqbROzqlRQwjNuF2CUduDWzUk01Or
zsghYiUCpFpFM4SpYH29xHVy4ZO4bgPQUIlmH98+pkwozSHF1EVdDgioCvH2vM7Z
fvrL0lKkY2WKwiHEOhzupshDk137rcJl2O1Ox9bKTFOJV+NgP3zw4det6axCzPa6
UA5GiZvbYwnuXP2Dn0fHw0Kmv0X44RN3zB8QwpG+bXOmDLESHVF3h+oO0Re65t3w
iwsVv5WCV02Ysd2GHTu9mOl5zWfGc1UWBnj1saTo1XWuUTCjCoYVK3swxLY5swQo
jOEeLqaCxG59YWalota7KSqRohJZF1asFzpMEk4cJGNAZwDkwz8LRUVTQjWNVdCi
eUTiDxHrbgDntbH9ZPwmlYJkgjwxnRawPfm1/FoQSno0W6X/Baq827Rubx9ZyuQf
NwI6ldKdzuIMlP53luOxeqmd3fHsjmeTUEWeQf1ujhD0hWTPCYyxOsR0nHmuit/q
OdOJgbBwNS047APS9Pu65Sq3e/qcDnZ/I0y3yKvmERBkoApaPiP2lGdGqz2LBXp/
VHk+KN6Ep+pI9dVx94amOz1wRdlakS0hNJ8kw7jPKIlq1Pj73Mq6y3g9zAr/QR4I
MZbZeeZxyWrh2VOBviutcSnd+h5mTHOrTn/EtVgj6tjsuTblvh/u9zSR/v/dbuS0
8CahYMqXe1LA9lVZD4A/a5zP0YjzCwo04muFJHxzmPVrvNkb3u2HLsE4SpqniXJI
iyTjzaKPWSj0tKBe+3cmlQg4W2g6djcasD34DSu6t6/rE/hfRIW+MqwYxhZAjHTN
ytLMxkXFDQDG4XDJYP3aMNr+KbBwcdk2kYfYlZbjd67CYDsBL+Fv3Va8ojLpnD35
neInc5C5jWe5q0JE6Lb6bh3kTqNj05g/CfSbLjx60l3Czs3HJ281NXG8dWaejP9X
whJJIjY9sAz1Lgo2XTx9pngRIxEfkTcogyMOrCEOwXEuMCpmpnzdj6gmMRQioxbF
PiBEg/J0ymh/bNv1zCawIbv7KZ2OXZ+z3eEYvVpGxYMHVAwCHq/eBZU8yp2nTmql
5YrMij5hZKWorIrxSSedyf+qSiOUI2I2WcJCZy7MszV4rAm8Tuo6xKVDBeSGY1KB
F8zAXy3bUikVpILsVXoylfBO0j6VBlyhoBetJsNoO8MELbs2xhTrFWz0nb2S2pKb
sX0xN2KxgxLLaUk+yBA5Zofunjgm3nm+9bPqQ4MCeHBPg+fz9wovQV/UlWmSPMkT
/+ZkY7aXeB6lrqWKztwg4zMwW1Q93ZB1Hc9IsHNdUivmgvk2V/cXr36Yw7p2oWm0
kSfz/AyUYrx4KgYF7RoiFlkbQ/I11t0cREmqjFGeplXtf0nkZbA/vAN5jsk2UbAb
S2v518fRzaqevtpFl4C0i6Vw4sQKkKHSUH0f+TO3HAZ9WwKgs5UY7rDwew19PVpm
onNT0lVVetNruosYBctH5K0V8PH+f2lKmwfK6PPQP1vvN4cKVCsSl8hptugsjqZl
1vNYRn3i3TzWCyhnMYnLRjMuFAeNXgK6g8QqFq/gqrucZw0qa90Q+px1t6pIddpf
3EKIs6LcUYxfAggGfNCOcaIu/fKR0w8XCdvngSwkelltkGWHP2ZQjkYxu72ma0/y
i7hTp74ObOD857jGSAV7JafYB6IH8P943qv/fDjy69sVqnh+60v4plt0GOMLo7T2
8jlmRL7JygzAfxw4GAs5O6/YFxTnGSmcmvbJQcxXZ3mdobUy3fyId5OzxSGy8Nl4
g76iRXepHdQJ10OQscO3nMc915jpOEZ32k3Ga9OEtLtfzcsAVCqH5YEucNeOtroh
GRwDq55J1TLzYn1ZzXbHipZIrBtxGN+8YFH0eGJOJW6SkibQ81DkBJmin/K418rT
QcomK5q/lJYcaefjM47LJ+sxQwkgRgZfCfynU9bVTDg//kgWlZ2tAyufaYx5gZ+1
60Bv7nuHDVQx/e29ZHJ4XgwOWdaVjER1LyuQYGeCOzj45xW35P+fpBW2psbSjHtp
rkJAZ8zmSCpyzn1wdgGLI8Af+o6/iksakuDu41NApR3QtbFauMpEYlmELtDX8/uZ
/0275e7k/b4sl/DZS7nXHIeuCArmWWsAuRfbZJGOyQhgRpD9BfdxFLa79/kpmmvl
qIi8VACQQZQjgbYGqsLRErgKfAsmc7P9pdcijgTnfyo9lBbXTFFFkKW1GSTIXna6
Zoa2ocnY5Ojy7DSg3AaiCu4kRy7C+695oyI2nnJtiVq6ZkWTIKj6hsyUPqKw/FhA
QKNQl8Yh/bdyFyNjDE40moVHPtNa9bj/Pgq53vMhkYPbBsmcJuHWO9pVKNMoD3uk
MhegA+PZlI4OZRBPpk4HtCZCno9rvLjpoWl4OxJ+IzQlTpwF/fCupETVyS7RzGjA
wJJanoGrpux57cyyHFg1GFqTDgUreqcj0K8v83+QF7p7MJupJ9EBNlwM/1UOPMIN
hUFw1ApFW/pmmD9BtLYD8QYJfuOpK66tFQJPHGrlTaCBcJbzbwF0LFprMXWLjdeg
lUnwKjQbuxShsO8IMXvu/vlqp9fKubRTZGDhYyjE2w7EqQEBTCK0Nvtw6UYD00Bi
J7sIHBKfzEGJvYpOdLD8c4/i6HyxQQvwatnh8EHrdasFic+V5pFXu5SbDHq6ZbMB
4lj1BfSPyR5ohgi6NZK218+GcombfD1DoYvS3UFrfpx5sxv4GfHviTa1c9rIjbzS
hKm+g7Fw4e+RXvFQNyngSNOSRbEOG5oo2Hinde5SRn0Zrxftb1MO7uzqbnSqvxbH
XHFb+P6rDZCLu9/dqdJfErZ/ShuZx3eA5ostVHRPmYkkMns5RYqfOjVh00zdiGiK
xSzuywbBOgAMLM+Ml3KtnipbfWa3+QuAiGozoJAJyjppdhfIrHzHm0F4mBPeVS2H
cqT7sOwsmeNCGo59F4Jd56PeCBfy0h84CrIU5LbLXCotRTXKo92MDlu9+3rnrhJA
aodsP+NEsTwQ9EwIFFMjT9S0HWpGWqkCi9G0LGcnOB7FMpMaG3uDaDzGdSa7DYn3
EN8vJYX1tneauGtza5IvmRu2wLhFmYUylVnQkSVKNn/ENfBeK747p+K/lmhNCQy1
mxREBHp80J8uOPZJ024tA2cp8w+bMo17Nh8k6GHAivjGtXwtaS0YXnPEMucirSqs
T9A9kJKcA/yXU8JOBPoVh1UfD3ZWti10oLCBcj7VzytnrnFVPbODH5T5PotveEtw
4kbNAsG6Ory/gCdg8HI8aygwyKB6RRTI+xpIRUhp0xNkPR/9KYXyxTSpxpgnr6ao
fS3qhJuh7UmroNpO4NZMDPkYyoilk5UTv/bTKjwtUFkuLJtoVC7gfNG6DF3/w0uF
OpAjnRHv+6G384VdBRREmQMqH0INVQX5nISSjNS0e35lsQ8y6v3bTdwTn2fe8TXt
Y+bgowViK7fbkVjS4Tr1ML3emGjVVynHuLIN6JYku9DgBm4XDymhTm2A7ThPBWgL
kXrTp0dxyOKCUKIpu/WZccFKjLTWFdgmYE8gR0yYVci1/BDCDWi2PP8qqc2qC+AK
JCnMhSuMfB3iyV/ZTbkq1S8XQX9g0a1JAtC6GmwujjZXy94bOKQPPnM5ueQlIoDB
6y6GARZEfTCWPY1aVwYF+e0/32zS75llddoPw1Y5oJNCqcnegH2oXVr5K4Lo1wsY
rMcDVPqQEyp0rBCVZEj2XIhxi+Bs1YgXbEw9JMAIe/Vld49Le0FXm8w3wzLmg7xJ
CdIueFsaZyexe/6VgQ0kO0X1DS/QsLC9f6/fh05nDkmQA34bT3QPAgAl7XyezaJE
0+FMNdm4tajzjmmRCI1JpdnFc3MBjqps7jJ+3JBdM732izoo+Ck337HVVrvdBqHO
eCZZuSeP8Y6gqvyymeFsc9ydWwXuStIe0QmmgHjX10nzH9G/GWAsYSi39SvuGgtE
Axx4aJd/9jctPSqWQISu4Rbzl4mMarhVvG7QEPG4ufsT3G/NePmSmgMvLQSGSgTs
uxn1HWVESqY+DanULVWd3LHdPDfUSdxFezXoS7v9AFuMuCD+o4NM0K3NkWU0Dg9H
3vmaKMoPWMfWAAK+HCotsV98eOJbG9KYdM6ozCVYKeK6+K+fSdPeayf3WjqKwhzW
TsMlYOUD9ACUgQpKvp6C7qlUBq76Jo5BOyp9ZVJz3GM8Ma3n1q98hRCFewGvrWct
GI6t/LahNr4VThRnUXS0V/6IlF0pYwku5kW7AXgw5U4EXuyPxYJMKqwER8eGQ5Zj
6HLK/4G2k4XS9RhWNgjzGuWvQCEXmXW4qIj7aUnKFbTiyY33Le6TzoFIwXmq4MtC
1mhvhQFLUhYz3fQkbQ0td0U5RyWf1P/et5gFrgclJEk9I1VKCnc6tChKLW6nOMaw
msxrtwMl9XxPuxU5O94NZhd5jnUXAo8YIkoPZ2EABZgN9lZ+TGBxhKjopaBlgmpu
WsDPydKTxMyElkkssdi0ZNpViu/YgrhRUCw9fUieOYmTeYJS5T5sS7FJapkTl9Qk
804Byd3L2rQ/zeLay3ehwSuObBFqJXr79nzmd6utUMY4arA+awitTGWnlmb1ZxLK
Of5X04yh/QPzSCDSWG8VW17SaomVfw+voq2jY+M6gMtbx3IzmaWSK7daiH06QCuO
Ep7fWndJeqoqJMdm1m89+EwCbvfJumRcU46Z9j4RVdkMFu07MN4xKbAeCz4pqI8O
MGQXi59HQbBgLjIcjkpDm/ow5WRJvYIt7v8SIR7va851Fzl/z7eKftIqciEMVFFL
LstKRe+PsAOlNea+K6iyqtj8yq8jleGLH2qMBfni+XXgiCSUlJO3bFmn7IQpYBYg
KwOil2xILRr4TI9LVCtWu+0eJitPQ515P1gGXuyMY6VlZhGpL2xt1ueSstAl3GY2
xw/Pjl+LYNkKacPfEA7ZKFVTHdndMnoU9Zflg4MriSI9puyaJOoiKtJsG1ra2r0o
P6dfSVIyYo1we5Et2dyeACZIjVFODU9VpCYONT7GwHRkuLmauSFvUQbehgDTvqUO
3BapA/o3uLObdjh9FbmmkhSmLRzAz+MlZzcoMH0l1FGvJ+e3sfpbE2N4BsKk3xwx
XR2b8Lca3H/rIfZRMa/6tH3LeWFUfOmxV5YR6FUwExWe7y+MPGZABzvaugKFPnI0
cnmFAJEDJJXyNjM4xruRmT+iTDAwTC09gQVlNYdOXvvxILNAgFwy95hjA9wi+AU1
vYBJKQ2K6ctvwnWIoHnwT/Ez4UoWO5irV4c029hFzESUUxdourkOCelPfffV9OHi
Fh4ah8MdZ6EA/yyuScM6vIhSYGv1jBcWI3QbzPrCgphNG7qjU1bjf6pU9klUJzmv
AJvVw7sNBKNHXu47aviY2LU0xZam0Qox1z5sTbjMIG7M4r2TDdEDJzLKjl7RmKCt
XJedQ49p8RfgSYrDataKSKbnj0PRYcpsbIqFHmp1E7lUR4fduh4awU8uscBs1kpy
4+JOrtyO7/ICcp8Px7jRDWlxKEYFYLh1Bj9vt1dYJhvKf+B27KN3uoCuNsb0aCmc
ONFMY2/MTqcvodSLjw6MQ6NGne+zdDb73hiQRe/V1yPY4fyGqtyepQZ8oZO4ZrK9
/Mp3dOvMNMPYPFHXwFhkOl+YSjSpOCpbf2uAcrR6ZMaZRfPPThgYO0H8KUF2qn2g
B8AV8kgR+WEylvYuH+Zr9VB/jsZukgv//jDrgX2sYPPWRhGHFNlK1o1VrqolEOWu
5tCANsMtHe9paCEvLY2YjE+qpijf0xLRIeD7AdeBhY/d1W5mzm++lO1WcAALCTJk
DpKOji3TFnnHEImZQUcLBQ2ho1JFZJKoNaCK2Ue09sl6VJ5cSZJ7VaDPMOKBVldd
Om2lcASmqGI+hvhZ7g99kM51BXrnVAbbdSztMTSq3Lq8Ovy/wNh0vJyvPctrYKOL
Jo0JWtEQllKwM/Ze+XeKyQlvjIxlL9vL86Ah3pbsmyxzfsTDXSzPq7v7IaTppMkA
pA+zy7CqCs3WDjNOwTYNtQ2SlACYFpvEqzb+ieV85K4oKNFzR6U4Xq+Tr+MH/B+s
DJxfev0P+lPc44lblYfBLxF9NMb+AMF61qDARJKJZEbpS4229OTpf9Wzc+CIAnHU
y6YgjKJhpVx6F/XaufT6eYJ39ctxQJrhCK1yWLBFtMm4bp/g2mfyhGsf+NqT43Dm
mvK5Bm+gYj4XTlTkQNAvOt0ReEhh27bVHE2JUZR8lxTkzwh3GGqh7Iv+cSlRApWQ
1b3ng8OFkx3BF3fSWF3zG4MoC2x+4HFiBXq/al28SXfExHe91AxG5w+0q3Q/Nln/
xLEcgUdB2ndOs5PNwNhjK8XMpCrmZiQfVv2PJWCHzipcpA/awgFf2BYzCaOxnIEc
yrQA+3j7wqUgaAAjOK+i0vz1HAATy5T3ieuNnsxDWUm2tCPsuZXzQuFlQovKTpG5
/2s3ziD+6yYn5ZltWNn9lTRSjot56wMLFDvxdT/JCJeOgsEU95JlZaXxcuOIBaMB
+RnYw+nEg34QG4RF4uZG23NPJyN8kE3DE9j3PZ5VYE+qXdsWN8duXP033YxYnwVv
G61hSfhwjXeruC0np3Ntt9sU5PQkb1VxfrblL4/iIEujTuJogMwGgE3/l7XCLbPi
0NjhkAm6LJrTP5a8uKtZbwh0rNhRM2MUTiQzccDFjZzurkA+dEK0/RxcAhtqcnD3

--pragma protect end_data_block
--pragma protect digest_block
QAGsGrMIcxQgfUcrRC+w6R6Ggsw=
--pragma protect end_digest_block
--pragma protect end_protected
