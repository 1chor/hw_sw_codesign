-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
h6EhJLCo7nlnKhyaP0/p0r6OAiAqL6zM+A6B0St567WsgcxA04JkBGk31vSSV1Jow8u6sAuTD15k
BjS59ZGsb4N/7wP4f7osa2Y26HIMJlQNTV2Qx1fqZEP6e/aipyagxqEgTOlhntb7k7cRAmQFeEZX
7RXVEKhxlmDbycCCH/Vey5gQbynZ6CmokFicmHixsmV9FQl/rhNwSu3+76A/5r9iPYYc43VAjuJK
b6JkVmquamzeaNY0Abgr+BEFrTc1lMplnT2rq3HHkVObxnA9uAezyA8K7I+j/V+jY3a/oIWsYAdX
zjdtii9bWiMyf85R8MSGfNUTdP2zl0n8E4vBJQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 39376)
`protect data_block
wfd1bm8frP+m4ZlgVzfRSQbKn9bE2ou0IHhRljKq9Ek2PVrgKYyYKz1cS7OjglkOiRywGqqV6aFy
wf/qmsvwp9f4QZC85OniLl23fZrriTZ1djrJTdh8JErSgEGJA5C14ZTr79NFWkNV1TrAmR6+bRPv
Q+N5JGazrMdw0N99m+BYUSw1pEVj+i+woug77NMN8ciZ5hzVB5SvtAlB/sgtjAO/LNBGszn/O8H5
T3OjXN7Y3XqfJrrB7A9333VZfhrZ8V4jwhOBXTKwNZXbp5w853wTiMr54FxbGk6AKfNVEZoqazwr
I8vZqUKEHWTvICj1stuw/uO6i1j9ZgDUlPkJ5Ak66NLt8W4p10AiWkrJWhlHF4ScwF+Ftootj1my
eUcwhbccRdEbbivAuvUV5h+T8xkQMF4vx4B/hGe33BokLaffo0qTh1yF1GBe1u5a6LJ1noJmU8Kh
29q49sg9qGDHifDB+UA1KtXw5RMMr0wDUVUzX5ZGaTiDKaGb+t2EVO2/sfdCVWdg6tlDX2czl3Bm
Qqs6DkLKfgW0VUcLM7UYkmMPsRqv+tA2Ub4TyVg6qtZ0ja3MiuhWhzGjS4R2cJNNnl7ZrKDOhB7W
cOkbbzNt8hWoHIAdidIfQslKIJqswYks/ZhvHZGm9clMqX05bP0bNcTJXlJWVTi/bMC7fOLqTmLR
758UgEsfNK5fwNigyr5pr2K2c3NVLR7XNyJAB0ZuyFiAW/CYZCyHdqqygmIczYSUttFtXMdmmJPs
g0FRw06Ib2xSbaAKm0hO3Xb2tLXrkoARFIFJFdZnJSntxizro8zJKJCoL2VRtaObe8aQUxFFaLBw
s2yzZZder+38wjSaEmxATxwsLosJAwFtfy7a6a6NLECUG90SWYhahmrWchZdUwlcXVW1ZMZn8voU
ZHDqCXwkWDbQodDgQB8kgJVLCIBsQnZWq78xCsV8W/AnZiqKgR4xSsoF/WMe/i94ZoT3nggM4SCF
76wmaU7/flFKN8wA9dB0xAAIbHR5FRysB5D2+hcwojOI9ye6XeORBaFP6IyrzT/mORyPfsYOsvtz
0yk6P2XkJqEGy4z4Z+To/AW18OXJQ+EFRCn/FegSgoEPcFi2aSP2xVhg2j3hFF/sDGqMV0xbsnqT
aif8sS1JNWQ30oBPr14KvhBtIPwP9KuY7UCgZP9deZXBOIKtfN0KKT+XwJCuu7QGLRpDUJfJVOBA
p2PWcXWB3PIWEOTsHIPQ4Ry7SI6UCXXYY8XPZ57jM2SHQQKeAxjvkpZYhPW0RSx/W3DV48DuirtB
F6gZaob7T8nUY3CPEmuNRFq/suJoQl9vGzMbMMuz8Snq+2EcLbUdNDZXXKo1TvH7++eBv1U57VdN
yisjrMYsv6BXt7RzYRN/U2R1NZbl5cXtdejGi9SnzHJWVx+LYG2FBlBrOAcCfYTH2HsmkOe67ECs
b6EAHLc8QljynvgsWkcPDuuQpEa+gmSrrybpbQiwB+WQEX4Zu2SSe6yK/sk15e/Tanf62vcicwi+
M4K/0NDErx0KrI1EL3muL56FumvQKk4EJyDIBffwDNN1YTSF2J9iyrPsVwz4ShRZDwZUjk/V1wCN
7JT3TWrQBJ9peDPLKBcx0lF7OLFfDnTJ64xu0BWhMeP9Yq/j6N+w9N4CccEXP8VymVm8yL5gYfVH
k5JHg+ZRNmxoWgZdK4v02qQvX/SKpONVxG7vlbZLpaxmhLsU96ayWPq5UORqUuTDbQbzl8iOaxrw
7HujRc/OmV5eqPGImu6zcFigvcgnQ1FSE/Ck2OGJHsE+FmbC9C+ljpBtWeipwZ4ZOhiOtGIU0zSb
5yA6tGLLCqvpKdTdLGgo4BYZDR+ZBNyf6jFGt98TgUE0Rzxy7Pka4j4EU2kNGgRK6LSGnc/K8vgl
0niaB7MBFaSUDVMKrtC5/azDGhLaiIRCmsiKBN1xf8fhS16yJm15FiXbHWS4srQVvBFO8UnxNdAI
0SVXZJSIza9pp3hIzcLOEq+w7ea6DmjVaayxJ2X+rCyzbEH+fbBGArqHyG2vZ3IRiowCo7linIBI
nGIGBN7n/gjUScqkhCd8tosjARYr39R1ciej2OWcoar0zZivXLcmst/YiF2shqFbCxOvqU3sudJC
kIgKFmtXcoPTUVtaCzw3TTkX+ZXwKWJui9nFledtG/PCIKt8/Al9sjUSLqMOAzjAkVoVwpNzKFqw
fW9GdM9Ck9htGPYsA1aeAq4NgbteVj7MNzE55t194FwC/t06sC4lVu5vVVWgsPEAgHWQX02bDg4Q
F9obYIWf1cl5XYx8duVoi1bkYFubrpvz12sqqxFtFhPyI6B2CrKZ1NM1JTiaN5tE0pnIt5ZBc8UY
4UUimbGstDBICcNZC1v7rx4UtjXsczalHscwfqc9/4efn3FR/UAiX92tOH4gcQrEWKEZ11DgFwYv
du2oWj8mKm6gl4CUzYhCpji8ZjZRPIH+jrhqYul0RTi+8c2FPm3i3c9qBrOTZdsqoH8jzfWPn7uc
4jgbaeiz3TczNYqo9RXQHGPegkX8OdoKPebmTG+z564AIp8WcVHPrpKnn6OhOFqBEoiYIheipc8o
9R1XqdpirXZy/969temU4ubbTKrFVvfA+YG/sRIoK3nuY9ZGJWFWxWz3Ri13aq0iKSrZVyOFdtBk
sMgdnBGMNS8bqho23jAz4Q/OVDQAGnzPZ+T6H/uFpCgv3qPW7iEl26lcZ4qIvOflf6UkhWGcfso/
0zdr9yYE6jHytgVj1GXZt7lFTXh2Z2Gik6kXo9NPDOoo62y6rnO3FJ4A1eNIqYx3oTMefmk0Wryl
zjp4lsmpWU2M0W+l0uhNVw54FssSv1+H72wEguZ5D/vvYyNiG4ZDpxALsi+vXZ3gZ01MxJo8kfSd
UEbZSbFw7Wr7i0zjlVGB1DLjvnAYeyU4Q5jUbEMsJeebGXzYNbcXr/prpDghB0x+qQSt9YRIrs+c
mUnnq3zqhWg2Po5ButXWJniy5qG6a330LlYtak3bdvUvElKp5tFseMfLwiESFmQue9oo2hiEVru0
r+FRjuROsrnreiEAO0tT3NhJHmy1F24Y1B6+PFi+xRS+tfi7DHuk/C4P2THoDi89pgPR9KVDak5M
9RvyxgL7nRb/I6Nt9Z9IDsNSUkja3X4GMTvUpehkFCR8ZpeRyqYfipyBNkpRUqxLV1iLHeZvvSRa
Vz8PqiHTOVE3fmmI/wD1L9f02au94HJuNel/sA6eXeB/VjAqauWYTiDev0iw/lEMWnyc8qV16n/4
HKKnAuVESh1zu748lgMWVCZE4Cu9WZLgKQ2rWA0EIhQ15Cze8wGZ6JXDUTdZa17rIWqSOGJ8H86s
t1/D66VqQDHVz6Lx3YMuvY0ZqeQe+nemz7jwXjdfKU8v6LBoMOJyzsqxc8yyAdGK1mzKYPm0+LRu
bPyUNrUVdFqwgpdEn4MEw/9tp7U5nNKA9/Ls9qh1sl3FqUpl+DWPnMQIoFd+Ofiw88il38IFM7mu
O7L9Hys6T7jKXivzvtZiKJEIuADTrU+3T9u3QpBBKlSVC6t6y5mYtcm3itxVfhTurQzgAwQ+6yIE
dXgyPHgr0UntNP4Efk6mvLDDRnEGSR37GVm8MfSkaag8tU30M2WyMpxEILNi94IaqZ9rxQAS7XhB
V7KzS98M6l7wSWBfYPVxj+3i7oX11oolweCg7WD6WybT45DmROF3bqT7A7GEBttVAAOqqWMJ9X+r
ALdMrwlRlYi6WPtbFjCO0xJM+qwS8k3PYwUUK+/kasxlwc/kE4GGxxXRn7ArKVm9bUYlA5Z4rc9J
xM1pWY2mx4HHoCdjcV10cBH/HspZZGSWrBRPy0reegheTireXujK82Wq3jwnOJRRrYJIlc4ZvFgx
264FHAICXdOQABfHuMOOAvpYDRTh7MYb2SPZllR1Jr4GfECbNmO8+ysthiaoWYRiJYa03STPdSrJ
6kB2c4xbe1KUtHeVd3irV5bpp1obBFyvIwahexDBgVj7wtYLGFC7YxwbvfGl4F+JIyN/FeEzPcSd
mExwBka3ovVYz0Qd5u7Haqx7u4oVy54VXKM5ItEkTWeGKxC0N/LtjVj0OKt71ut8pkRVkgvPTMUL
dWGBd9Wc0WWIziFAxkTavZJ5S36VYTz2G12yNdZ02jY8/2GrF0PyC31W4CiKVpyCHWfIhjK1qgex
dQM8Hnn1a6C1jPGPO1Bfh/yHJBuNVxdREu3u2f+pu0JU/xMrOFxK3M3w5EYKKMipBnAHNRRb6JlD
h3wkBq6/0U2ABukQdkcoySA2xuNARMHfEhnIJJvFvtnQkkYhYBkz5PboTlk3rqb7BCG1IEl+nbM9
AFgB+cS3I+Ru+2vG9doG7mv4ph5tnHZ3YnXWumcxvIkjkk6BTRI0zCZR7zOGxlxVnlqBz9PDxUDt
q+KGWKBQ6Lk9IXXNeocwsbktQSwVLaWQVgnUTNbl2urdT60GMDCitodq+jNCJYI6nBoKQMmZoQ1b
3+a+Rtgfpr72x0x9UljpD4lrSlfTBcHA9mxFPEoO9BwHwiLJipGcZsWgXX0LOg+cmFsWtT77S8w5
ZftBibc7VabXwiwqt1x8+9l5gpR6rGrIuwYw2DA88oEgavuOWFQRep+ey7kvEaOw0qIHghDqU0w1
mVjzQVMHYkIvGaAwk9kgFUNjGTgXRyXHCOKpXKiMWdOehJ0zyiOcQD53h6fdHNU8jWqzYxGAdxDB
KvsqHdDI49AUaHyiUjZbUOChD9c3jwwLZ3UucdBvkEqu2DytJFMtRFqIzCW0EuI/tcq4aItGmV9x
Lkk6Jxh2NgjGVOh+AhTVzdmv51xVzv+2Rm/swuVwnnm5/1VLPGvSmPieat0C6mng4KK/lzxolI16
8bh6FeHDwJKdlc6QjwDGPtgRQJ+iUDKLASLbmIjtZn91ibsiXUCPIPtkkns7mX4vA33TtzeTmDSB
MARnc8pbvKdTJaIMBJ0cY2NUoPgrl0hIDoXElKefJ6MA+v/+DvGLf/hf2UmFwpTA0qJvGbEO/LHX
1kH6eNlTFqmJnjSReWYklZUOLGWahyuOXiyDKnjtcoDwFGMnwNl0F+57Fgwy0oxpBaKlv1gaLxQI
2Wg3LpGPYg6OtnhyXjesC9zYDj0Lu7uBpnGsSG/otvVw+JK9/rBI9gxuH4wRxGheVku9dH0gaulP
3d90e21d1DYOLx8ICfWYt4WnAlF/lBOgFpYqhL3WXsLqgpehj6DII9H93Aw6PhZ6KbCtouTJYPMi
1SASuKII7FiCl1APNw6gSIhcsurwDQ+UHwVNmGxRhdQAOWyZXReaF7VK9LFvkFYbh0ZuRvYRsXA5
mYx7oTPHjl3VaQwi2hkt/7HeUtdiBGtASQXomehepOoKoj3Xws1z8qgqoubQI253KZvglX1cZ06g
jteH4tX60N/jceFz4Ry4mleisp+RSu9pRvyOUwLnVMPkH2H85BlLeNNOq9TOkPw00J4Ax94NhX7g
+vUY2M/p6+Y8+dbxQXhNKFuzvmI3jfj9KYeFktf0iMC36l3tN95zYsiC2ZtLN6tB80MCqbLOJ/ji
hy0gkr1xcF9/V+wY8M35JDkttMd/r3M7sYNOLhT3b+RV5Y2KlssIWYwCOcKV+as3xiYkmLWcH8dS
3c3H7zxBLuen9cTRI2M894ef0pWgT1Czi1Care2flRI/U+PQdV8BYb2OojJv7DP1JL+3FE+nNbML
grwc1t1tcVgsQcnLPEnSp+sLeZGZLSH+C0L+xjxEd3rEkh7rbzVGbZHlE+9wJPU0mlnFDKLBecJz
ba/PFM2ITU8etbV9qxRPOjQPk/0OeKruJL3uY+55swXDC1127ZYj3dpLofnlUeMCJutZgoUSYclz
fuRotqLKtC6cnOY2VRRUfZ/DpEPhw7Y4imv1GXVx2gqACvWuTUhj27NkwRBv7CsN1Urqo94VtSBd
NquUIGLRK4aPAhyORy3pwhXN8eTt4tJQ9rTCn6ASKZPUJhZDGjf0eAxIDATApkVHpRiaboLSF0/v
F97UlM9pgMJ7zh7s1mn07sP/hqvRCBWps8GcUzD4O0QMMBry2yCCBn36RByVjrVYAjVv0+WkPDWd
KFDtfAwDV/UpWFiuPKBPQSEyQaz9+M0iGWHpz5m1FDJUBS0jVYdhNwGFoNnfuP+y+CEygSwZ2d9f
CZlYvqqmHFQQKABrmz0rZjRVcblpworIuY0ZadPeM7aoM4MZ46ncy0lrCKNY3LEISu4tJeesa/nw
PSwSJD5RGIwSmLnESnyfgrMiAe7dznof7RaAq+qCXlHZFDmmBbc/B7zeapK3Z6nduAOLxbcT6iim
d/Y6Kp7zw1V5CG/33CUbNtp5ZlQHDPyRnFIYVazhOYqXlElsB6tkQmT5qwzIIOHDAc4DLWbbCTQZ
5/J+fpEqPSKgqVCVL+AoPE3G/w4299aUx4+rmBCm1f2sjFNfRZ+1EHhoaWUV+IfhANMfAOJaGvQv
qOQ7CeU679bbeyzmCBIDb55tbD05Gm+scWNMPyP+Rzs+yc4e56UsIWya1Y0XcbcP2BJHMlxfCIBD
S8OY3ErI8H3j4cA5JsviR/TkZQp/9MTgwf5ydEkKNGFpjAYBNA/tr87ve/0V6QEvv7LTdKMQmlgg
+S+fW71mvyjKLMeepl9UzC0lopCOvN+6NJfj4Fzm7ZCSnh4j3z0uGCONoKBZLFd4jb3MPs58DyqA
lnf8RZn1kBGnpEPO2YxLi4L4Yy71vq1tNppecf4kykRsPGVMFbxExLIDdRYYdvG8lP4PAvVLZxJI
yOst8L8YfaO2o4jqZ/frD8OqtFYqTQgBaVNu/VZi+aSbJTXPyRgYeb0i6qjDRr+0YCDbn6hVWuaO
es6q90xgK6GvFio6LDABRWDbttnqQ+/Di4Rhsvaq5BSBXNvuy4kixP+rd29dSNJ1ToIAr3TRJNi9
VAkZtZ7DRUjI8vLrNge2Ayz//6Tx6s20fhHldu0KyOrGygEiEFzPLfsMwr0NnpMrY0ltOydtgjNg
sv9muy/ZljZk+Y2rEJUNYlm3I2kLlNnR5RZSq+0M9PlTZ9g/WpdGiIE6YCBfkGxr8OW9f7BqM3k7
powexxz3kXdExHii/aWQRZzxO48TteuGac2suI/VREBMTdrF5do6LEPpvh3WZV/Fy09AXpFROsu7
cIWpJf6cVtqs5ZI8dKbp0AfyQiAu2BQOhlNCwvlD+pXYA5pMwFpmf3uzDmUXNM76xGrqHzquUhZt
QumoRc8JAw+NxN1tfNKhLINA3IyTJCMoilRykYCtAhKG4j+TFcOsGRq562l7ji/r5Ffd9jknJVOY
606GuQDUZGQUQ6j67WakMojqy8ZU6o5b+BFyel4NWTvp+pRSN3Tp5eFsxbm9o8Yp/FhrLAy/wVJ7
Z8gx8r8mU5AkOSvkB9EUV/UyEZLTauqIc2s9luc+QVpB61/Dzf416t4BH6doVFPfCHEdnDcw9+Si
r7IBKUpVbKNsXTOgJk8OhlJa2eSjxMx/fokunVhBfKJy+VsfTOBOkrap42uWMbalop5CiLUPJeO5
2PJjtiwYIq4NhHMbUoBnIOJfRU419xxdX2TniCoMttDHvOhBHfJeP9l5Bw+T0IIKARZEsQq+jRDC
LGTJrkY7AsaY+7a0CQgPzDOaqQUMzTxkOXx1pOFzQ07kU6QSdXTCOfDGSRiO0Y/zoAl9Kv9IFSc/
/+o1d793DP5vPVkscnLEXFl7v64TRegy4qQ8T20otEcvSprT0Cbm8+vxzBHP8BGLGXFIU2YZcUBG
te0b8JVo1YVxCRCLZWyzzZKgHsffgWM2CBBCEvIEcMHFDgGchI9EI4NL6cIwMTwufRgPimy+8aXA
qE8TOzSCYrOkQkeKYuPokHn3IfOQ9TMA8MbiA6lTPbdc6HVnFm0sD12LPGIP9YNHJSSc+59qgkaU
4IlMW4ulhP0edFK84s6nCYCeCoZzG+fkOagAyCPVbzFWi+38mmvBiW7+lQQwTU776BqAx/IewRx4
wg+PO9KBEqgb+kmlDG/2/lSWT8plwmAIGlpLBmK6weXl5Ob1lyWxfsP9+j1dT/MZ/CKIl7wa0WNL
mPcR6WiLrhN1k1dZe8N2FrMGY0hKf9lUfgSL6d9yAdosiIy99dQdtiK/o8GnzVuqPmVMn1pI1Rg4
0/fgVvOOpex+A6p9U888TIZdQb7QX1hyaBoaCqhfmIbT48gTbIOFMYBnKvwP44K935xBKrp1GvK1
lksGHwhJBOtkqixzeDyY1+8QfRE6S9YIGmNsH3RkOJeqBF0RJCU9Gw7A8mJbvrfu8IImbzjBuARD
j0zNSF8ZPPOljajXPu6lK1OseVy30T20CxytDpV8FzuD/nuELCYdakwWRWg85+8lBrHB14rnzTva
7FwAlsm0VhF2rDgsWwuEMvvPgpOc9fwogiyQtlN6FW5YLdQtGJfebmaAVUHADUC5tSdS+ZFEvnF+
mTq6ULKtruCXadyZPp4bNP1o5w3rezkuYVLqxqPaLuyh9ONCJHi7LCd3fCoKy884EoJcKI3lMJa8
c6QkF9PkGBWso7H7KvmID5ml4JWg9KdjzRLwmxFCzO9HwvfsLxzv/QHsS4Rve17/MdcNJLJXz49l
Z0v/u3wDSVYsK5aoyQT/oDmHkfksh4r+FtNhjzKtTesRNc4jFDfrEEpBShrxxZPYpOvFAAFmVe0+
A+YfHbOXVTCqQSO4HmfYcGrjT9s4lEpOEySYpsxvJdc/o9ECqG/IibMOl70+wBefZiQ7DUIv5/6T
PIPqT64omYkku6MzFwYUVUWKzW65stoAwpOSsx5of4e3nuzbAFvrrBLclwcy+WoPT0QBXvaFKRZk
Yw+aJMeLnRIq9SoGCluJRjhUFJ/asOIkBhN1wY/ag/i0em96WM6InWrQmdBfH5zjfQNhVNej9TDX
IB7qPQeeAt/Wzfnz0CupTncyVJeAy4EbzVbKCb/EXWq8ewpUVkZ3ArWHgiTyor1s33X1SvLNZf+6
Uym/G2h2tcb8bpq5Z0McuDKAfOhuTGYJv8DmbNCk358nAnCcGpCJtpQ2PQbbcTHxq8eU/3JjV6wV
elr9lOQeTGsuH5Inff8oINOO6Pc8HLhU+3m1O3WcK8efRIdTn/oMg9avIV5ehJBbN2ZHPZ4NAtcO
LDFGuU5y/rLbPPFuTYJkR6OGeAojGUhc6Iwh6rbUOCwyLBEST3IEYV/TMldD1JN/nItd9lB0j8PQ
1dNsyE4h+c0QOHox1vvY+EIQIO+5GpD/Q928iE+Rb2uAOhc6BBgFuwvtSdIW3MPhPIk79uskUqTU
Z2bfW4c2eqdomVf83Fl+/q38GySVpqkpL++7l+xU9zrXPRxgg7rtXMI0hkrwS5ak5F+LoXbQGuEe
faZYhY3Uw0qtA4HJxm001MD4KrbuTmw8feY1pP8eyStIiQA1IahDHnv9eGA4mkQRUyOVsJnu86gl
kE6GG6rxy2GmE1U4gAjZGyLriM4JyniXKKULwa6WKUZIQFWz+/IFiEEOA2RvBnMvqs9rnp93H48H
upWZVQtII6bngBeBWLWQxwh484X6PKjQFcpLBLEJEoHKIvybapoi4Eppf5eoNuevCItzMZFnNKTe
HayV36/d7yq0HEciu/SrL83XN5lXuWuoG1gRu6pcAVk/RmA2pTQ+YcR23hzDbqLsaTue4l61CF6D
cpA6V2mO+XK0GXsUXObyBKLMcZj1c1JAnfVt3XB38zsechFaXvYKJ5yaMF5Ekqj2OqP/HOsco0cy
/fGyXPQJGwPLdLrjHcl0/I687lyWuQVlCghlH+b0oy8Us9Up5DlCSV4JGQ5QVzhPX4SCUS1+FypE
JI4x5iQfdJ2SBOu67TMYeMfaZNIDGBtFyuJLkAI9o5nVTNFYKJYBhNzhcrzVAd1a3NK2OtuUn28W
1GGR/l0HCz8XJIwYWsj7q6O7py10DGlr4YB02edyp7oLlDTZwbhunkY7fJ+u+XhCG8sRhyfaYWV4
XGT+FfZlnME7QIkKrXTmvWE8kDzI6j4y93nFczXCwK3cRFCdF824+WZrtPiPZcyMDAPjGGOrQ/4i
ANc82KJhiniIBeK7hPkvik/VURwwgv20Nz/20Z3UpFQxUnIUSW+VejQL0Q8pH4xf4YDZ6e5Q9P0I
XtEcoUhAkNyiq+sx+jj8ugt90acsnPYLiWnzDJkbZGy61/gai6AdoPMVbEV+155ysXHLf+WkBugC
Yh/l+1eEVCE6msm5j7L0I3u1wBt2r33egVAlGvIdO0jH0cRI07O8LK0k5dNdD1M+EHFn8IHPvPRg
7EG+ciK/aDCZnWWB+Fr2oE/xUKeyr20tVaPcO7Y5waoeyruTuyasN4S/nDEFw6d4eIFl7nJ5u2wO
l1lpefAqlC5UkQPgynmqk7cPgSJHfxXIe1H0XRoBZKDXYNHJgw/y449TF4v/M9q3DR21qWSQkXja
1spn4VAhvzbNNNzRzD0Ll45AgzYSPHkkuNUAWwi8cIJ4qXBPjfZGWhxyGjHPmDXUgqS1VehhIlFs
6Ks6V2xPbEocMOVYhZL6gFM1SbXG1iKy5SXwIipOiw/kKapaMPH3GrUQvSU0aAwbiwEzAiwLX2MZ
1nhh3bRaizGAYGN0iLcQHV/FgdXIgDPd8SEwXcokn+kNrW0rQyi+44clg44PdVMYtvYBYUu+nIl1
iypzFtRW6YEvAaXcnjFJJIJWDw0HJcNPDNGWp5N9K4xkcAdUsNQBb+PKUIFqgdVX48Jstt7eQpk/
6FqJ/9OtjZDX641/yT3Bh9R6vcJv8KXb7QZfdK4kR6VX4W+Um0Ul7leyW1Ikdq4NVH42XLQHLnzS
QWkCKv8/o56eqxcOe7eFeg6ujKJwrw0b2xiJlJAC+qA9Su4MP2YOS8KbxYKpGSsxwkjMhGlHbTh5
lqsD5A8apqsBoyCq9jhpnl8sfIM/EnZBDSJX7/VSihkYTFDEY1tPRNlEeJytbQeJFBSTHyFwFLze
sOM9gc+pWjrhKE+wX2P8ovtHi/7AmaBIxis0yaIzXDv0G6hkfGD7HtHl1tKN7/gimT8hADM1fJOq
HdLmcafhJaqRigjkF0ki8fXxsiZrAtCV2iwXxu+dTtYj7uV/1xDeQLtt2YqiT3IME61Es7oaKu+t
iI7BwiIjO1fZ8KLZniN8TLCNAGpBA9Xg8D3brZBfoOLoEbmDZBNAgYewnKzaasLoEk79V8ZVyDC1
Mu/au8AgvTCsixRUGuP+3PNEgUzcR6TVKE9ZVje4lvTtvI2Yob7z5d+XZefIpVjFX/jc0j7Dxulp
CW7oZs/MSvbtpNXj/dK82lmBJaek/BM+aFOPr6IgnWvz03s8cWCVdqze6gSLZqqEuJOK8a0ZBCjS
kXCEqyGLMZf1t+cNxHsR5Wdnnuk+JNP3PeS/H67IgTJst3A/nqZAHa8mgktBCDBLdB3WXOX8Nlj5
peiFCRxK2oilEvdUttv/8zAiLNdhItMttocAdgesTSJPDJDC96rSEyay689/e9bAs0l+2M7lq7ZC
s0E8DTqxJ5SUxdOuo0HXESRWEtLU1J5nBuCza0FAeDIGsnB8G9tJqSM+L3phsYt0RNXVnDpxxcMh
calfI1+IuenujuRWH7+yrFOM1eF8VfwXyEssaoNU3W0TljY0e/J0vy3D5GgkbrMddeCGHxME1zcN
LrFexChQEkqerxsWxnihfbTDsVaR4hIpFZqUeNZmGrzfPwejt9lN63J5PTX3FCBMwF+nZ6vOkD3N
/Fl5j2CshJHvx2icOVMeYO02QDNXDyVWAMnvEhZaD7pI/DYviFb1dROlLT1B6dBW2QBn49iPRq7n
tSmZihtXoxMSo7ShWvRIZGsB+pofheoUJlfQJgTfnXIME462K/LmNVvML5I9GfPsiMuW0wDHt63N
cyckhWBUwLIWEcltc30cDNrNgUmxe/uQSvRr+xJZcUURDN6NSFtHNQ1zHzxdB6wf33GR1IqLYuyG
bQw/wQfhos4SRu71Z+FzgRbFctrJ3qAZF8Y/6VuMG0ZrWGADcb2y2Mrw5DMNYyBIMu3JLgZVThko
xqMsXjR4eFy+/0+9dRhXbVMWS9cLqlLCdQEFVKj2Mfn1/+CSbxNL3RI+wOpfxUpDsSdsCmKAgbZU
1E/+l3ve3N6SWrbCXV86H1Cev0s5B3AM2ccpLEXKXuAGz2k94FAYbRQo5/IkWuaGbfggVB68P9Cq
ZJxuZIDqYJw5JeTHeSxHbah/GZTCsOC2rEVPuZOr+1dA6WsSo3A+RAT6Sh1dYbknwp/WqUyHJSUH
YEUtUiB7HylfmkI36FEmpTAqhe70JeKJX/QI/zbBZXq1Frd8IPFXn6pPXsSBcW+cLnxRGDESgE7z
ELYyr+3xtOXu0D3pyro1HT7WtOhKvV0aAyvbKyhypIm/KSb1FpNEK58fhqIpDMMqGHFcqhLukt82
5sP41Fhmv8p8yZMZq97b7R5kd8FQGI/pRH6KawXEHmqu/W3Eht0cwUweidqE8py8JTEjRIoE4hA9
nZp0RwMBkifhS4bBEpB5kB+9mtUnoIOXHPPGoyefbW6QLFWGEcbwz18r8sKuaos5PAtodEz21tZ1
4t9mVJGglikwS3iBSrTGk3mV+O0xB0y3VaG7Pajz80nrh8vCBX1Au5s2dZS2IpLoScV+qihgbVJ/
Dvv/KwTaFgOwUICtr6kCyu+ulOPs6UAdFfoIbn2W+JqorelV/8O9ui0f8HBQzpIJrRKYRaroWADC
/Bgwe95qzAwRRv5X9b+kCRCCw2qQBNLlPeyHshLg2YtwDH84deTA3iVvu27ZAKRT2wDN3hIMa5cX
UrMTBgsf55+TvFXnXcR0wgsLLtDGNm76n9A2zH0uuoqSyQZNsjvq6uLOJo274iooiGsIxKu4655f
bKUULkdY8CXYpDlbFRmM8vA1lelO9IkMP16Wgeb/r1DCAEk0ylP3NDH/f3x0TNSgwCjMv9qF5kXp
JvJrE59aTIWDotlBzhGzo4YT9FNte6tAauFRHbyEuZDoRWeQGHe53Euak3jHWAs0NZrUxtwVkvCK
G+hNF8liMmXEGgzHsJIwhPRDzWkZMfGXbAZm1PsmBY+9qFZ9RWzmv3FkSaIck75F58H/XjukN70n
zrSTWjdC9LPZz6M5Qdwf49IZtqbdTyqxqpHgKICUhlgkdIkjZoJWgzWW9XbSuwI/fpK5udsJerij
iKpwQngtFDxffgO9Ah6rTAuwTfRGTBphFuqiVaBtdz8zlC5IoQBNOShrez++wyRFkICyHQFUo079
MivBpB8cp+EVnB9IPVQYuNzeCA84Hsmfn7GK8htc3FBgV1t1Q9AT1Wcw1bYjXMEw7sloBea/NVmU
nxHwWKXcB5nlwEkQoIjIOC11GwKHkBArlmkiLkHSp9breWVhBoE9T7yDeZOjPCUsFoIU/uRnC7LW
Z9de/o8tpp6HF4Z2Yj0TImS7s1u+mGGZylfFjHC0OwJj/yv8O3+88agL+0k+fPDJgRN7isM8XfmD
8QTqaUD0oowPA+p9UChmSz0R14ebuN8qnKQxXz2YQWyAMwxKL+8eVdTFy3sc9OQmO+1k6tbC8yoo
j2VcI7VwMnmmU/RbKMCTe+XDSo7/M220VdMb90GYCXTz8FejOR9/dq7i8YU52wHME9+G646drtDH
5LU8oepNZGmPPObfwXjVSWQmVyyHGxRuCzaYRLfsrdOmyJzgtSymHK6sD56+Pqy5sz16ME7MedVO
C7PFo9+bT0TFAMCMGx3sAUI0WGE4pcABxn31quMvxMkUxSRkcuEOQih3nDHVavJ7HPSf5Q3D5XIe
KET3e0bM5bdizEz85c/3RJOVqbiKpOsjhxIeDn8xnaHUnqia+83kqcxOgaIGDCux0Z+YQ3uIHqiS
FhRGw46AIZ8KztWCy5iW2L2pHxhYRj4RBcKh8NujRpUu9ZZOsEf+IykseXew3apLht+H1lYX0yrJ
zgCfpvctWzn8HWIE0QVA5SLmD8kmtGwbwDMa0isnCx1/jAf9Wlxm9FNLJu4ie25i8ZStFNqxWOyQ
dDSUffIIiLj9OPoo3ESI37D43YU9aXKtsQUfrA/NseiGSPy25cMgFGA+3dbgpRkFm5kWVexfdUKk
keA2dBE/IlpjHGywsh4RGZ9idcsnGCQ7HskkEnrr5mzQWD5cni5oexKlGtCHdHASTHhQeiJrsvB4
6P08pxYmegQfFs9kZRdx8oGq3lD/ew08aa3g+MDK4bWJ3raldxrbC+z6UMBlDSyar2VhZjBX7O8w
M/O9nw6JvnsfgIkTEPmJ6L9ejFuc90ci+FU9W0hWyArNuW184MZGnulrX1h7sfxGYbjSE4sm+sDf
e+l5X1BFO2cfJ6wwnlki/t2Kd5NWn650XJ0A4/SfzYrZHHDO+YNhGt1CY0bAlbuJOE1/9wo0WCEn
ZloSCA+GnO2ak1SAX5a70kRH9tEF896/A9xfmDSqIwI2817G10yLYj+iqeZW3bZcDfsLS1A0Yq1m
Yszi3cuD0HlJ1pm59f3EZpoqvpT0oTqKa11YMXZ43SJEq+ijqdR97EBgKUDOy6uzUKD8kV5Y+O4y
H8gH6cVCKXMOz7AkQ3UIh12ptpiLVZ++qzjau6MJoKlEpN1tJ6lgNDS3RGzaNuVtAt8C0noEhx05
AB70vWqUZQJLeHjW2qXetq2JfLc+NdVB+/r+Rturp0yiI4AlftPHQuLa5Q9PtrO5swFsNhYcFe2C
iXDv0kUIvUoB400JPJc6X7VhrJumV9FpGbGTZXTSgOQd4YQx2XBNHGIdCNSLyZfWSpAk5cF1hKic
SihIg/P8jLf0shhviA/6zWgBcZW9UCh+PSnaIzY0A3N/J73EeaUABwEUigrkofhjvkiT+eVs0jQM
TvBg5XacL8XDNCx2wk1UKCU/K1pIkAhdEg1wij0e8l+dK95Zg2YXwRCqGjDdQQTlrb105HelWG/d
pNxe/yRCGLTD8TgTUuxedoorE6kLnc/fADVI6+c4yagfDh4mJ8i864aMIUtvyraJYtYZlXmJFWzu
M1k7nDEFXVBQV0Wr1v1SiOzZLwnJkbgmlDF1N4WjkACfRfz7NigXCrvGd6vvKv7VYQMRgR4w2/Jb
NOy+GFsyQzoyxkgwfOlgOjm7fVGWzoFTRWqDsvQUXV72hTcyTtRESXsifERX6nyL9CGOfQWoEWNe
WbczagYdHD2tBmydhw17JasXxcYziA5TYCT44RIa9YEtOqJ53fImuCIC/FlHeHCrISCpQ4zw/w5V
pij/HeYBUt0Jid1Qe1Wm8bmrG6SjDf+4t+hAZ8OAXKawePGJdrOojySMGIo6kg2F31SMfcC549Q+
gtzbfZ3n/CCKykpLoaFnymHMXi9xWXMhC0EVtoJEk5HL+cuDZBHX8sbgfUTZ5chFlIEzIulJNkz5
NWIdI7zlzlWTKgtOeYSn3S4oQFZdHyPBb3ELMX83yws9Cm+uU2zVkOC0VZCvJJ+Cy2ntJvzbw1lu
SZLFJMqzdHtpSkaK2BKxdd8kFkzeUfremybvZxbLxhollwvg6THALhY82XR8gaz9rxSlB9RYAcYF
t8IIthTY67S8R9VGjBr7QdTMErYdALcG15HlRKMU2OtuLb76zIssxpAgdYk7+Y4plrw5orepYLpO
xHY4K+3WXtR4ndbQnmv5oP0jsoKUPQQ8quiTJt6TU0ZkTD+9Fhfot1fgoZ8X7spAczgwRU1f5MLy
HJw+uN2c2N2bjqTlT2rt2msEZgNhNFwnVCMVv7a3H8apyIKxwn5IIYulqqgEMyoKlC4P5rLwMark
nf3v8JvDUWbZSaZ0CDtQ09GJAAx+GNz4/8LLVcJPqIt68D+1P2soWJ0JmGPoGLRwH1VM7eakqtP7
0Sze7tWUoCGCZDsVFmGc9dM93ny3YJnQ47aeJpK4ju15Am+M4gLrugsm952PfYKenD3c4+7t3tRX
7qh36lR5kHIyPIGuEHfTHFBTy4e8TEUVsskF0n1/zmETCRYMog9SBs3Yulj0FWvg4pvWO7fys+qD
jze8iruA3oHyZFI4J622R23gLx87NXIkw0D+70uQxeT4deFDSt/c3m6WnaY081NvYNKDPiHivjB5
MxYQSaEAs88SMKvaRzUvt4ap0TBEydZ/P0HoolOOwSWliIh20MXC7tTDMF6Sk+Z9fwly277zXKxJ
xUF/I9bIJ9wrNEqmmWo2umAvQLurcw4wwgbl0TJIECI6jJmojDmxO6tfSKVth+g+xoyiYPN2xzZs
I+JXe9NkecdWBq0bOF9QZsA2HkjLlPSdSLhgtKr1gRVzvGR/Igdw6rZ2RM9Xiyo6tpwGa82NuwUg
wRXHMzJx48WaMCZX4OuXd7x2UR6UXsv5+92EpSaszRPf0GStNN6cPlRWWKdUwEICtYE0RQdRNFAA
zyyvObuidRM3JNf03+5lox00NeGKvbVF+cW+59i5r1aS80uXYYon5439LctfxY5aiiiYIQLjJztD
UnKZ8XsZEg0UhZiUNRArLcmaEj8cwyc/kg0z9vPbu+brrSkLxy50PkRC+aK8j5kSNA2xL1M5HDQN
m4lCzEdhG3P9SPzqz0+BQ305Z+XRFzvzt1wE10osOvp6GeSfm7mME7di2OswoU7cCXdz8LCKeMfC
uxJyrlST5hP5+xxSjOAbwMbGmaKxsZ5/iFu196zkE8KM2Um7w2bQIN02sU2KoH0zzN3HSjR2ckgZ
9fUE2sLmABbO5ps1VAsiV+X/ClXRjIGrTaCHZPc9yWPSEXWqQ2PnoX7rYzc8KlnMqvKfRsxu+xCm
qEHmUQEcwOW28T1EegRsaxVJzPJU//SUIOcV0+F97u+nWtZWqr2pljHxlUGIk0WMIh81sbHo3me9
6q6vbHsAMF7PNHHIelCsO7nwH9y7HRCk5y5zVDdwTvWWs+wGQiS6TpmOD+Te9sCnH/eDQOf7noSP
pUMcamt+0LLbiyGPBhJf/+UC/bjybT2R0VunWqjRRfNTuyjF9bvRXkT7AcYT/+JIyf9tCdjUHFyz
CSsInpK8S0FrOO3lnAkwCxuxtLir+hQ64VYFFPh0T3bi2Vreo+62oynHPr9EnLJR1Gw2Y3lveXiQ
7LGIl5tdzQE2AOXAxpK+r56WeHQHLd2abakHILHqa2f1yb5cCR87mkpbOhoDFkeROf318K7rpgqS
qPMykWskJEc9dZ+aCIPe8HIdOCmYf+OY6EfO1O+XTydErBE4eUAK0uTxTFOi7lgYr8XU22IwzG03
Xykyk7bHO41RiExQSMTeQKrt55AGBj2j/onjBOIvbf4CMztTF3DfNiJmdpgGcZD6S02Z7uMF9+D7
5+wF4ZvolDCRthI5ShcOanoB9gVazyc88aob0eI8VPBvGh1Jel5yblcJRHsauML54iEjUAlgLWxq
ZF/r8dTjMFmi9ZJ+oLRRJYcb/ag+bM0MzUIi6wvrqXYmNp8pUB9XFu/aS25Z7TZpB3xbfiu5uwbo
5JwTJkC8M+MjATEet2W4earTMzJIcW7cPGJpnQvmFEfFtTUT/VtRDr28mwfrsO/ZfvFzQuzFkafB
5P8HjrHnHqIcA3L04bFfQCv5qzw1VJDSScxCxjy1dcg3NaMWm8q8G4T9Lq14rWJ5z7ScfhVkikCT
O/fCWSXup2wEFTixQk34A8jgh1nnvLp9cbinatSx0BPFev3p/1LuyDHy3q1vkw6RBCpyHQP4eecO
Q2f2sxnPE3hia1utUpyesdMjnYJvWEF9+rI5I+eR9vX1nhPLBANO9lH0Kb0powkxhcmCotEYiSkx
qqlhrcBOvGPIzSZgyBY2PyVocwlQQ8AO9yNckCpFi2IU35uyulfJfZfem2yBfYsCVFbRlYjjy/We
KsHD4Nbfs0KuFCmWlNBLFutCBgd6r8SxC80gIQ6SChZTTXfJWhjFfzcx2BWIRxTWxc0R3MlzYh+R
MMm5q5OkmhsMWcQIo5N511jBd9fUXK6yXh4mtkYuP8n3E9pvvI66glsrFTjrPSETXWBSoDQlVLyi
eJ3Tn+/hdlMsxcfptWmYQML45OVf4slZePHdxZ6fqgmoJIj25dexeJjjqMFsJ71SACPchVrI1sFC
c4hUUhQ0YoDs8nMBBW3xAAElazX0VMdVhBmFS//2/ZDR3yEu6JReGPd41Uuh54pczqaMRlBINge6
Dy+/7cW+oXpVGXN4A0bKRNxYH7cXo1Iwtey60ofNvjHz3mrxzy4eHyYQvy5SJPvFhg6wGNGw+dz2
lLZuSWqjH5Qd3WrzuVWALg4VU1xK2WzaKCEYlfPS/r4Cwdy8/umO5wfqBAU0YoDRthyN3re38486
G1dqCRNkRUm2DAm/fs0s+d/xJL4SFarXyRP79ZOHXzzCw+71zrPLbJ2YNj5oHI4i9fb2DGUJZPSj
n7+mrwv9SBPNkyMAxPKQdXD2Eo7wae68lldBGl9aWwGWBSKPfyYxYkMSXHIecSJN+ViWT1CHHuyw
90tMMvopLw34sl56VoUeAa4HMZxocB8+LdUG7kbElbq1Xww1K3n+7jKmeKy26gwuWzVCxTWUwYSz
PyJcVrPU98n0kZHXTOWVVGFDUTTlCu2QKUa+L+I+MA/Cz4T4Z84bp1QP+QomigQuBkp46v+CeK0t
7x00VnFH2OC1Hgv/FFKUcQfceyU25N3DgMDiCkDDWXdnIzLwUgowHO9M/EkhGUHCTSlmHlTkKj9G
ttptNxBeprpkRYosalq8rItQrGi0uD0rtn0jAVscVbCVcGcVzOmxgtysS+VZ8jRc7qLTG1RMWEO7
rr9692gxLnMlCoS63EReuFX9h9GF/4I09MoIWmbAfNEOaNx6/iGIv4EcoD6kLI6Z4PKcYVKxJd1x
Pu3g4PbWHuY7IVOwb3TJq/tBLubQuQRwN4yaPDJ7ym/HlNF5rQAgtJ8Yz3Tbs/oP1tHe79yZWuU4
XWMVWYaKBy8nw2x4QzFAa2VjfvwHN/sRpNeHbfjriRvz6LOpB1q4lligrrUj+vNVMJUMEO3WfE5H
LzVH2LwGotAg6tUGtqRBok2G76nOh4cLTtQ/LeptCRt/4IGSLHoQ5El9nD5HdIrG/LASDKQI+TR9
vY/kIRHOK4hXLLRuT8Omur9lfA0BsffgqtpwAh1aiyIb90Dk3L/O74KT+l1LQlREMa3mmJ6W8cBv
4Q39Wa/0GqPMezHhawXwddBTtmaLrRQezMcy6zlmlxPxgraV8ScIcAIeD6x+Cdf5JOYMeERY/gul
+flPxr6GAMkurlxXzhlsK8evCHvz9NHULrGXXqhjINzWOF6Opv6nIu0Ntv1x2DXVxkgKvIz2EyD7
m/cG7/cL2gFSqARmKf9+2b2huzzDK4PdR1HDmHE9xBNUkI7MlLo22KPB38tFLZ/IloeAQGNHnoAE
2sD9EM7s5XMrL4Mn+iiY+c2NqlLTMDm1ppWzn3YiyprNlP11IGv71mJ+NDUd2n8WiZLFyeqh6A+Q
HCcLXkhN3ZspIdITHE12tBm2BYqzoP2ZG7PdnQVNVnJAMycJb7nMVVokuZxk6y/z/3lvIgZypP6F
ldTn3Nk5EfhIdPJ+Ea+jAR6HJjVIwlAvcwAwWOiz+DzvsVj+oMMQX2jDjXwIzIQT1Haj/XFKeF8b
2o2GaVMXENHU63EvM/eyDbjLm3QCbwTvoRoc93GpGqUclhLaP2YUGx+VbfYPAk5/UlajotTgTX+3
gzPG4vSfecC8g83BTdbGznnNYnHrwyAlw7sqEeZjs0b2lrVuO34rCKrFVIvkTnRRD6PJILB8CQ0f
ns8CVKGmHxRdfGMDxn4VQJ8a7VUxFJdkAkVMMtgNU72sKuM5kZcs8bLy5o3viP/p127Om6jxpQhB
LiPW0/3LjwyU41yW2aHvVivd5h2tume0Vg4QRzjh5TZN1+TtNHLJpm0jPLqjAxKyfpeTsCIBBJdh
rMnVMlV+k/kgG1gLKsa/2E0D9DoA9cKUXTsOOZ25Ajcy4auP7/xqH7iTGmZ8EeOmzeG83xZZKCTl
YrxLnT8Kcfb+/E0QEX4OEM0fg4StB3EJ8p4HqPBm3sACCwvuxdtJtmS8PGti55d1Nch0R8odsty8
tSzhIjxvOpFT6za/Cyz22qNRvm4ZaGDN+9iK4t8DETh0tdcgnV6XZyHnaIZ9SaJGodxBizQSJop6
CIfNcxN1/THYdm/7oQErJMOMdgNUzlIufwWGCh4JpRIQPpvnGoHgv0Zbdj0rh40FLaZ6FPrQcami
Ga9AZXZglJQ5bKcEb35L326N9Pi6VDGb9Jw0lwN+FyCbOaGvOUd8cGfHZwoft04Ph5vBUM62hE2e
W6KLjB0FpG+83Bskbr4lqClj+EiZ+gqWEWxkvQ+l8WEZ9ITEpcti+yR6bBsBrZriiykxslkExcXD
GwYwLJ3x3XsghLEF2s2vVf8ydxIlgqnrj6J4Aq2G+MX9RdQbc+w12sj6xQF3ECRR1urKHt0bdFzI
XmysN9vS2+LN80DRSrNHgXN54BVv3hxFIfhFXuGCGqyMZ9UamaEOVjLys4K+aJRTEHyPEyvNjfdc
xDfCzqTKZefOlpoFOstapikYmGSIwiw4Rx/ObhuQi1IfgUBKXnMcp6rmqFdUR+gOiL25QnOaHEKD
zt5wHbzfMjOEQETzsmVVg/T8RFF5UjjEzD2DC4ripZfrh3TlUG2/cX9DB+kl3ulQFvQppIop/j0J
/zeH0qhMW07hrNYgh5lq8uWfQ98nvt8xbhacvA4sBSCe6ZNeo2WWUnM/OFpLass7otTmZxSagMa2
VViOwVa1iWt870Hq6AEJqjH979nd2aKZ+VyHnfhipwkHY4GfVW5g8YjAI9UQrskF5nA6UYcgCGAr
MhNUavA/YHQDVT5rooS2HoDSjsAR24e6lu6gh1euzCH+MeAuC0iXr2jW9g8tiTBNsRewHXQRFhNN
sJpwaVRWpO+SW61H3dPSGPTeXN8rPW9BxnGZowLdljtr5MDfJ5Q7KdBN95jIxz4Qk88soq6xG8Wp
MiCScf4pJ8AuepQSThKFlHIb0SiDI4i7ASqwJUfPoloFIzhbcJn3N3wNZF0rMnGJtW/bg1iBg2Sd
Q6sbwNNKGgJfPJ0+urv6DxKh4PmQ2LbTlKNwNMBxN1wKOucLmEqQNJFY4acXJWBdcGF1AwzFFEg1
Eh1NFpPYZdvMPoXaTotOG4vXKC7RYA/7db9Rvs1/XrThSgFZ5fTOme/gXkzSMw5/O/y98u0AqW4S
2dLxbVzZVYjLyv1HcMC5GqdsY142FgiEhitBJ+wratlqF5YVK7tP9gxvYuMbtQSSg6x6vnjBdirc
9C6auQrsjol8r9ukaIagRsvUJIpQWRN1fy7B/JXilhGySUqrV0ePkLbgjL9igrApxM7k++YDnSEi
05MC+YMKp35ngGj2JVuMSAoPUXYka76UjtO9P35ZzFqhQ6Ib/cS+twlr5XoavLQGTQbucIxYpseO
Zqz0ulLEPeo2K0Woehz45qPW9FfAqqLjPjCaBRXJUcDR0T68yhg3mItdMwWADfp0xROOeQOMhTSj
B6xaGTBU1RWfwxVKot0QsbvoycQaq6WZ3Kw49wq7N4VGeHQ11Rpt77vwmfhUdj962P/o7SqEesua
f8E9I1SpdJdXL4esM6YqSTTmLPwr30d+/PKEEv1ln8GQqgNIdbLAjIBGBykHxhBnUr0Ds0bAoOPq
aRyUv+NI4KITDUU8WTZYJWDAQNP5AOd+cpGjCl7GYEe6cmNas3e8ku7+i9zjMg/u6R2gknpWqc7Y
I4oQAd20EH9DAwmXf5YJi2qG0Td7CRrMjV1cxAXla6Xa2c5XVJAg6FunDfzpAdtlLaHuZ9cTpEIN
eQtHwzgosO+9MZNB8AgNebG7Q68aSXWfvDsKSeGH9YjGF3hS5XysYB+uSBlXsym60IwDd0AotkYO
hfSWJFSHZ9MbRxDxE7+xPGj98OKRzsdVQZryJOqHmZaCq4/lL4tYPRYITpQBvmZBpu/BivEuOjLp
J8qZqHY6pXjHkUqRXQKw0Hm43tLmi31g2tjM+pEyGuskzRY4+TuOcMjS6Y1moUZ9PMaqpHzia5Ia
WZh4PrLJ09SyjejtEVjuyKcQixFcBSmQbDqbpo+0QeMy9ij723qyH5jxHrABIHrzWSdzpWKRw5a9
a+Hnu179pITjkOHDWmaRgADb6SQzLR16L8fLYpHBdXaQD12CH32ZSqOEyej5jkxF8QJShGFaaq0H
cG6kDBjU+VKZRql14iiraQ3iO53a7vEIcJr/lLk6jS9knHdw83pEfupiRhZmVQn6aVd9vXsNrg9t
LLao0QJTfJ7Dqp6uWT+h1xctQBF+LYXs41N8CWc0BRkLuxkQC6Td8iKN598y+6/BwR+plUxmmkDD
2Df2AwhNKod8vLOR1Y1XqVlM3wjAi6nOvuRaZ80OYoSHSZAXhuURFZd0GZOyaVsAPKczSGNlOBju
YElIFIkNJSt1jfueYlJ0Wpq3h5eLKkvYJXR+HU0ZRb5+SA4G577FI9CQjWkz1xVL6pVx8eag002I
7vOGCcuo7WzGpmKyUbGdWtjxTLNxFvos5xJ9DmueZaTf/CEbWh8iBfOVzvE4kDocJH+zYLhgInZd
PlZD1CalC+ftpzOt1nLxMrxu3PYb/w4A6X8KnVyMy9vJcPeSOeHKIsuJg5rq047bVwY9iezh7daF
axONxZpA2YRVilfHmpDJuHgNz0xLbyyQqP9WEF0QVBHXwGOSN0+Kv75v79YhG9v1FB/Xld+Jtz+c
imcE6xobz84Fyi8whldr9uLc321HaOAMtyxBiIWgBAjc8CXwLqlejbDP637mPnT9dv0lcZhdvxdB
DTPITinUtmCFaWrHIygfnNlszOc5ZsJ52k88s35cR5ZCLd6mx4z8UHZXs3xZhdBMrAuf2iPcjSA8
tJDRP2d0h6nbu0qIMNS7IE6/xc9QxaI/QPxha5h68cDzmeRMRccA6xGCehObVDGN03Zk77VSfXBb
vVVPzFSuJzHjOMncWq489sK/ZnscNG8lcFPnxLoenJhNvCPqL7Ex1h7HKApwS4YneJ18xhzMV5Zz
qNwKU7BkfFLvIMHsfp+QgjLSxEhBJEej/gw5T0mj/JyOywjBoSZWyocrss1T1PoAVlh2muwB8IhK
1W/4eRTuJWS1UYao7DWQ2I5JQrT2Tv69Po1zul8CxRXBc1089oV4yrThusqpt89zr98jfpnnOoSo
KH/Nh1T0DeTUIxPaMaw8qxg4D09En6XqM8dFoCvNlAzaC4yeKtXpQvZWP3OBPin29ubdEFRoEHEN
77IUxct0rhC4lL1RToaWj6IkjmqtUYmflLDa0w6STSIqxV4Qnny2RkuyWTzzO2HT9rUrbMXvDt0k
rTgXHImT/FSu1BtFATBdDnixdwtApqugNp09HWshUAcTTk5ffF/LvnjAOZkdW60M+kuNU6BZ0NIJ
2gOVU8zpGyLbGib5r05jRy5YY4sfESNDMZDima1a6BveQ5kxYosTkfU6HYdTweIE+KMDA5fiNWdp
xkYs855EVPVS0GKbqPTUYwv1RkKdZFTC0nIUu3Rw7OYpPQ0Y45oSkRAAt9AxMVbV9xG/ceaPJiej
Y8D2Jq609xpp5+S3qTDxm/KOmTQEuFiODLktHykp1H04/GddV27bcru/1cjyQGZ30p3EnoPHAQ7O
JGJEFLT75uyMJDnOlNcn5ErUILemPaZWVs40T7JvgJ4VHOYVQSy+tf+d17Fd/XW1G64tixmc4Ppe
ZcbiuyJnsmPxgSa8rXjZEOEhF7bA71EEiOTG6oC2XRaz0HtFPYpGnd55bdl/p8NPY/nTub3Y9S1l
QSvVRchl6/kkHojejURS7ROuOMw1FkuyaQXWX3s7hUSu0Nq/Q1Lk1vFYI508BOv8NI3Y5H2EQiR5
u9oQz6m1LKWNywCDSy0K6kPXS8o2gZNUs1eCflMxUJdlTGqFAcxLHOHs+9GdkDBPA4c2eP8OhPi7
QuEHd4f+bM8YfaZoCiwhoD9QW4f24SREhnrkLOKXtAlOc91FfygyQRReAQNPyKqnxL7OCJntFAga
Z7DlyfqBnjCNfCbwgZrL2RFCiGzaQsZ2jr/IaCZc/XTDroJP43SDgCTtv2zu81msKoTaic/6cwzf
byOx6WsIdqj3fS1lamk23h054puNIfg9odlsLJboLbnK5of6gDWfpT0Y4Dr9q82/36TjqLnYxRzr
5H2lyI63Ith2IALdi+LjjM/6rDEcLT21S7o6KSUBg0tx6W6HxFoN/vbDNTBWa+aLGm0QGRpnZM5d
Hz8EuclKdYVxWP/sbcgcjxUwqFEVSbdUzV3RLV36q3Tshgxc54UeU72xxMqmmQWTsFBfth5PWmM6
DsBUrKoLEq2xBafUVJwSAEfSGawMNePiE28HHtfQYQ+TIT8fmDbWcXW2Uj2UTaaBpCW3c6hpUgmA
7uaTwhfS5/Ki1DkqUWv6yMZtEGmseUtAFIw/aeHux3uFlbbrc8Jf3/pBkJD24wLoFiqH3/IC2Chc
8ReMlbxvscJddqqnyc+tzHIvQAlg6oUD8EI4uqiYaPHcFHVZLk0N0w0FMxoxXDgV9uTvY8o0K4PP
1BBd29vdZX82U+6F7Xz29eyTbjsi1B2wmP5s2WBG79D9GDl+Ym0Xa0JFnaDXa2OIfthtKabc+MW2
RmmHieKOlpB3GPyM7HkNOAfz19xN/q5qn+5r1jyhV53f90FWmhURjOiRNeTaYOsEK/VaLayuYfCX
tO/a3DhahzLr0JZftAk8ksEeaF8L4ISMzy2n2fk41npemLhAX++c+GiYmjbcsMPWlJ9KZywUxsgq
AgrpLgieEQrAFE4xp3rd3J6RVyFgpD6kYWd5mCucqkfH071s+c+jrYwoT8341Kofh/0Vn8njtaWB
Ygq8m7kybFN7u5nVjWydSNtSDKuQKIx1OJJEzzLSJu8YT0Hf5pRJ1OBB6cumFtFDUuA/0flnqFys
X3gP50deuJ92wkFqFu/tB2FwM2k4K9NDtRn764kn1SgNh7BDEt3+40+JBEMkh0ngXdpL5YQ2BoTs
6ZNmci8qmMoU67t7v7By7uYmW25+2HHXfR3aw2afnlWr64a0HU+LDjYEKFGB22yEv5Ot740vkBwS
23LB+Ri6h2ueMy8F4g35ml4WMdSK330n0eFf/FGXc9ZtvMNJS9L1Ksf6LAAR3W0PNaBA2QDBG+Lc
WiVkEZ8X+Tn86yXH0xyhQ0YztZZWf1/bZY3kndRTJ23GnRaQMhEd28Btytr3C1oTVDkMr4mUIk2R
abE/A6heZG2rBy4i9xtXzpdflkZe4aOYZnM17ybkFr41Jg//RX2gAhqXWte4rEVMngDHxdA1T9+o
X6QboDv7ybc4JFyoQQ841vq7E8tE6jfPEbngLzcBOO1ksSWVTJu9Dv025WCEUkV0lol1vsnC2ODU
ZBcMZd4vEpdVdjFe0otlFZAMCeaeYaMi9aPrVt2Stjlr1hRXCxsiga/IsT9Q7vc0Gtoq/TM+8CWN
D6x8IPgK5d9XcIs1EhM/tIg1OTCwhqWKETaSZV+6YWZZI7MaoqftxFq5UP0F4TSi6SPeEd+BqExH
WcFA1hkwfdlnE8FqFfaaj2nOR9FWGHayFBrWvTZZU1nSPDBpQr49R+BJOz88THX5N2IvfiQX0K20
xAvZlmEJtcVs/xpV1kVpFT5KL1mDALyaRdbHuAwoKzGohA3xDf8xj0rSDW2Dj6OLOQyQPrLEpvdP
ExqOrDoxt5voHuyFYe9R56cWyCNvvEU+zBHqJXSAF2pjhyNTk5gWJBc7NvJIwdjcxAUOoMJOJXPt
atUt4ULo37IPH0moHfLFY28mmO0Jphu+GXnolVkIl4kLQjlROolcWmLvcqsq0AMeC6IWgCWdO88G
hZAC9TZfHpJATNQqHPgHkivsci7tHzahV9yhcAizravqT/MUvYYmvt9tTZkOycYV+jjRYJv/5w7F
/0h6gMmWhz9lLLhi59CBTZ/hf0BfqmJwvpbLFN1LDNufCmrPLvdehw1/q138LjmipL+Lf1bnph9q
94EcnA5E3Qo5askaqkMsdJLdBxkPWTkLWFtLgDLrIyaP6JixlvFWK7NTeinSBBOsmeLoYzgd42yC
vT8oaPFNwEwI8rdkmJibfICYCR8/hjJEsJXClJrHhDllpQU/XBS5x4rfHrpt56VMbUJxOiEYG/Np
Fe0TBQtIkUbUW+iFPDj3bZWktroZdH+U9nxuda3rxiEJbom5ocnAekwbrvEbfHHDbDP4W9OWKCF3
gj31mDENR8dWmo83f0QGbRTjclXn0y2vXQpjtovh8svHZKdAON4PqkCKbJZHtiBJ1TqAu4XpHjlP
7X2xSpKCO26XrOUm5ENof9tcXVBRXFgHYO7jUWaxyPEb250i1VPLe+uyGEJOq51U6rUlpVvnIT8Q
hbpAwu5QorIoAD0/DMcx6v/NsOZ77aU1SL/vFHsvo0xHDEsQfW+JhEMa4ZbRY54YBhheHc8VxX6K
ucKgZ7AUUaQz5ztWU91FDyXIWYaz88ABq+TykfLmDfYqk8NUhkedfY3aEmW/7DQvmd5FhZD3jsLG
Mn99Wo44bSpqAbvhStDXfwAi6iIeL8U7+GHwEuRytBs7j9qNkPRhw2IrkophMKdeFwPq4yKxvpam
XDtHKJXUQK6+MNkkvbFKS3y0UvL3Xz6qlTnJen1Ila24POY2vDbiMkoGPrv5in2vjam/vnah1d7o
/I3uVBVoWZykKXuFcQtPFQyrRZxq5YJE+NHWYwZnNQXi3aBR81T8seVMtyPG5vBS8SCiBrcgEedn
/ziGC7Ue81Xzbo5mYFPyvkOh7dgCBblZZFU0yFYQ0u0zR9cj+KhsQy4rvKFiuqUyKC+T+Brn/4fG
0OX1l0huxySUxhPCCs/tKSYvmNbrJuAdVWBAYHeUuJ8m1k1f2FlrE0VTXyjITKAZ7qEzsjspocou
tMgl2WCQYlpA2zXt+ZG80q5v9W1SbUHZYRmBF16xsJ6HV+2q3IOOo79YTC9hUgdkkXuGYUUSr0MN
30WoVTXnv2YmfSagf1zERRpjCkYXxkuH4iAKdVPzkWv5T/NevEj20DokcTLulgJIPy9qLIOGl0RE
59623uSzFVRkwIXg0rKzeuxCcENAKk+bpqeNzGJmvqEECw8QQd2mjdj7zGjUOlD+Cn3SKIQP0XZ+
K3OgnxGIVq8qiC187ZfMsUQghCdp44PJ2TSJPb0Szrsh+EeuItdIiOH5sepyKQwAhXxalYhBOCB3
OQOW24v58oR21MnDHSNTo/pq8qTLqmtt1hYqwH6RKG4H7KDmZkL0+wx96A9DjmU9h9cQt8oKzE6p
aevgvY+7wrqEkSCHyH4cfiAhPcn+/IQ4mzUMvz7LioyDje5veGjBj5CePEKlaTcXnvOw5N5/5pLx
tpj5UkpAYnxfEAIXrxWVBMntgZGBEL2+y8UwU9SjdOZ81fhS2zb6Y595zQwKvbP4cChr6bEFWRpH
hmvbAJ243GT7kcq++IHe+XzUaFQUZc2CttjV/D/dSy2loWmoAiEmv9VGWoI7CwgHEx7flve9Rnt+
NEQBapaJ+64X+AUVf2I1vHFGlMUb98m0XAX+c59NvdX/rkjpXvWzILyvUd0ikPnc7GkJrn5G6s60
oaTKHGVvox2dfz+c3if84cb38124K3ccvIxG65UhXDaVSZluKW+BAT/BbUYvHmEiDHZh9f31lCi1
gLOe17rkEtEggDfDks+1wNTL7QrOzHQzdDmiINUcmUMUSRfjWj9F7So0ZRCSS8L5TvCUgtKIueGn
skGwG5PSQ6sR64pgKH2fh491ZNpjQs/L8eNzA7pxGNITw6yUsFgTL4yGoa0APp9KO0aHi3iUK/1Q
XARbHI2AOIzFIi/2Nut3gubXcxjfIyQtzyuhROn221wPD7gRDolY/Ls4HbYkjHFPLK+SK1ocTgVC
AbXJe9juYxnjcbbQOeHxtugrVpcz77C1XOHVgPtflb1HURpVYLkBN7QzDSzkD1CN1RJRzWY0nnQY
+0Uq+Gvp1X+VGJ7HGRsughXVQLKdSOL1uMRlPmE8nNOcXnQdB2tAl2CSmX2QBzz8OTgPMnyU8K0/
ygmllbzQ99CiNGQ3bL5vPu2XklBjdLBAalCMiYxjZq/bXivRg46mlS7FkB39L99Gann9lu5EsMVc
OyGugHgOdcZx6oqHdrC7toVnPBHtjHbVvg8jTohXETyHK9S8uHlAVZrzPWi4JPVZ6znFD+imho3z
Dqg+3V7pnDsDNG9tkTFfxqia1Ncf4EmI/R1BIfeu3yErL/MM9dukNRvOYESXpfz6MuOeLkOUQseA
lVtZNLZWTXJWtxA6EWrvwn4p9IMs4RsorjI+MsQsWvlVmC9zPr9EmSe/2VYf+O8kZLjBRdEXolSa
j/xAaW6EkT+66MQ/t1MIsO1iinBIY2sEU0HNW4ne/NfADb+i1KNySADs7S1VParDivlICvWvpV11
BskeT/qtfsqBt0Y1+Jk3fhB9MCANaOmy/2QJWb9Vc9VxH6PJRPhhweR1A5ezwW3kBbKmjVJsDaal
IvTuiEdtbEtSJXssw0I0m55gK6I6mpELPYFXZbb9HjHWz2pPYSboq3smIZMR/bDBuH/f9VyP8Fcb
p6E4mLxFYNQptgyPemrxfWKzSN4VBNJrswxWBRAxIHlDa1gx59X/lDWwRqGL5pxq0a7UkJokcvP9
3s5chmAyoLEzeCb7poG8cDEGRcz7W6lMHZTLRQQgPCZ3DBwiNXAR0tPOtFUSTk3SRBYB7GWXZutJ
+3tQQKg7VR/NGIVttiE38nhQJjb7FycWeZ0THVTPIV26lAYdjKhvpoFmYHbRDX9thtA8xBgFCEX1
6IKq8kNwLgCrAy7njHyAyBlCxJ7yUUS539FyTk0RW+ZKNZMk9EcNNti6a9HxrpW5rFqe+1vX6gy1
/mhHl2i11whqh6pOmtXC0WwTzgV8Wy/Mok538S0pkNVn1meF1soqwhWKUs1Bcwi2UlAzU53KkPCD
iSp2MsEuSouAcAPHgWXZV5tArT2dh/vFYwLjCoMv5VK7BVo2M9vQPLVbyIOQjR9DKLD00y6xz/rV
r0BdxQJjlPfK+HjukJiddhCXi1RTZ+bnw198O9nsDBJ5Rc5jXAxBJ7ddy0tJmY7XVinB1Tl9m3vb
zUU0G2FcV4Fd/3v4xhBzmlYK17YmqGjvonDUmdsZmiJW4dXTp+O4o5SimxSdku5Ryc/pZPNfVhnT
kK+ucSJUNKB/w/SD4sceUHdua7qm8bYJ/RCa3ooPXn/6bjELhS5jYgxEHKzZ8ujVSR6/HjmC94E8
LI7JZs6SPUX9yyUmmPJvpzXz9APLYmFkwQ0GGdpxzXwQFSwB9fYsJ+3Gt6e9pgtdH8NusS8pjFju
h2bTLatxycx6q1W0IBWC/e6hQNci5j26xw6RBPPmDekFn/NCOW5nSQrOu4EyjBNy53VYLnkX+AJX
8lvt08vzq5gEvgAcLCpDBwtT5F2bI+ixGN/LUe7GYE6J/pvWnIZ9DAdRosgccEDiM2AuTmuv3B1S
PnNozBocV3BlLBVa49xsR2/JNxXGhkf/dhgndr4CQUvLBcUGc21IM3HyXj7c433EsyA2ByxqVgKH
ggZ1CVHe0rP4icRqWr4zrNlL2ItKcFeCSsXCGI6dZOCnLcGv3RvPomlal7Y8oD8XorfSgdujl8Es
kf1bz+nGvCKdLm3rQxkAtE2meLGUNeQPjTxkL4m+SzY5xEmrCJqeG1iH4fEjzRDqTTX2qjVwxSnT
0z4DJCjlJs8fEJZMyFs/9C0Pva1r1222cU5OuNrJfYz+M0ddKs8XE62l8IyQinPCqpVpWVouRC/h
CQjsbOcEIS0SkKnzyJvaevpOkBSOappdn6rNYipl+Vxy20NhMIwvXgCfvluqWo/AdQzQkjDvpuHb
+0cfYV5w2dleN9htZmD5c8ISLPLjm4mz8tA8v3w3fPm2PvMl/DaDaQnK/u0kn8vikhATswf9n0pc
bd9nre1BrmnulqOGSiW7rKFKAgw+8BnmrHt1iuBDMccRz+eUxFT9yFRTIv+t9od4dDzWNz3Mafyc
geAc5RnSWwZp/MjoocaoCZAmtNfdeOxHy82d8awQd0F68pDlB+HxRkZKCe4oB/NbVB9A9f1qhv7M
W5gqvi/0IB7bMVx4k6pOA5Gm4fZ7IgUPpHTPoc2iLHfz3QDxXeeWY0XWwP5wSFxvAyndEVi4bRai
tbwq4PmpgzGCwX7x0zxka7x/cuI+jbmQvHtuj+Wy+oaNL4W4aixR7iCo89a55EW+hRRfCCvv7IYR
O4YiFEwZ9jOXw+jVezYtvl4mC7fmx5nNiFU+DVIOh/ZrF3Qob3VsTaTkd6aHyoXnE0AHAiSsdjpf
es5DST+Eo7P0d0vOked8YCdwAxLedFPqLaOw6tQWPkdESbO/e0PjX/rme4J9gWsK4EuJaIWF4PJm
+9Ld+svNaKTrEl9cgpf9zcIZ+eDEklP64J7ps0laWuQB75FbeGHkx1mmkRz5e1hhddAfq67BAK8O
G+2/brMlzfbAySuaqctQ36BAsAQw6a7achn7Ox6Ew7IZXyyStvpOCfDgStPo45WWASXsOJzRM8u5
iXe7KnzjCzrWFiJuW5WuRlQ60+QY6dnxeAW2gpULmTA9iWy7ABArDwHgu9+kLsdeV8SWHZsWdit6
bdI9zXE3D/DDXmFsFJ/9soBSQlP4EXhOeRdMQA67bEV2zHKfnTEEf278fQrV8bj9ANX99V7cQMGD
eto7kZhv6JYawSiMLRMGsbCFwIpXaBs3QXLVkQI7yHTOVfx/Xa1SKtvOzwbjgyFE0NQuOvv4S9Hx
lBQ71YhqOqOcKXRjOlKGti3b/wBFi4/KyblFy8Wn4u+zuyk0J84eI9pZ89Gxon4t+cfPfY79EbAB
qTyTUe6Dfoy0RxpcT+LKp4RdPOP2trn/19zVV4hWn7q20QyhZ9YBl0JeAd+rsniSIBOpPgu7uDxd
1QxnH+dPqAgA7r1EXSDvg/pG6fuOWT+4xKkLOc1lV9LCVu93Ig06SwD2uhHBuTm9ead+OuTrf5OZ
+oYH/cxWhbWyfbE7+1tmpHt4xTwQcpLA/sn43BoUEu9+VcUejX0VEVtZs/9CRm9sD2ey7VB6M+9m
4pL6XwVFlAgEz5w6GX4Mo59IXCBl1rtK2gDJMy6Of+7nyHVvhGUSNGpLD3TD+LBPRApCK25huWp3
CignyisxSsoGcdFf7NaHQVL4qL/AMIoSK+bElU/Wi59sKygkcUMFqUf120dCo9at01LGKGzXUWw4
LhJ0vrxKSdlJqTGj0eigkG+S1z+LChGLS0seNQfnLFX5AajlEnWKQi21HArOCZHUs9SA+A36Sl6u
OoJURugVEd2Xe3lbRm8lqZN7yBe5dU9V4XYsCyRwW2RSpTPkxFGYX3VvLsDSh9MSHBtffTCxgrnx
4kgFmYmL8YaEKuOxZf/bBl5MQTTx1fkEHtj98/ujqU5eoL1L3ejk0IxMK6Vyfe0dxhOSBWHe5DU/
ERAZxvX8LgepOeqryjedtklBsM0zSi+DtA6Zn0WsgqSY93tM3J0dAt2l9aGMlZd0/vdFrFYHtcVI
2/D3bIoDGw5toIQ7DzzLokHcoulRMN2WvywjQTHXYj/pcA/VB2AfYoLnMpImRM6ulSNijCM5HmGj
HJNyjFglgLKmsQS5oxIB8eo4uHjxFlh8hBrEiB3SRBDh/mAs8xS1noknBef4H7/jCcj6QzxuNJdf
NMt2EdS7nQnYBkqaLvKTrZdDdYNBvS/4VtDNDLDzOG+zJ+3lojlmfakF1ybU28TIYG5orPpdOP2Z
idX5UH/8p/Pl4WAycKbqLfVnDAwm3omUf4Z0ie8aKlyr+nUHzrGtxdD8m7vgmzFnbuFQ5WbDIF++
EOwJ4DgdhWk4PsqXOr2o1JaN3zQ+sGfCh0Uz5IdWatsKLEt9NQx/7pV2iyWMPsX1kPWxy5BCNu3G
sgv0lAcD9gvefPCo8mIECUTz2P6tOtJKdqTf+VH9jXw3K8pXfuF+zNDhxk55l2vZos0FEdlUBPlB
OoOOP/m2tWc4XIHDVwobqcQXWM55B8TlyjMJ+VO2M8elShAS0Wr9MKLKWgCu3xtRJ/qz0dJjwv8e
HtCvQL8794LTw1IxuGpd9eCOibgCdg5MAHgw7QDtqLtXbs/xBmZJmlK58Vg4WwasS2hj6LZzijTg
JSca37LBwaf4YqF+yrzfHmhpXtLVM8OHTrndMpZKvI+K9K2tBxZmONCFLd8tJT665op+L7dCxo8d
zAPNSm8U75UEUOmKpSK6WpTjGok3vt3MRG8I4o4e9MhYRA8zHd8mJM/yeDwbgVS0EhH8XOaiXT29
L6PBM9x/fwjViGzVv6c8iC63FamQCjzWTFNlxWJmQxzetO+T9gL9WTzaS5aef9AD6soB+svkcqyT
Hl2GZPu8Fc00biasafDRSZTbmh8YnW26q3axYjqP/tXV0cuO17ZY+9rRn50UTlgcZtjMJGx5/OCA
Gx65u4opGbQ3XQ06h4x3qDnNbQSVsQF/sxbuV7jpHAAv3wsB2jzh1COHAfAaJHSGQAKYzCY0aJiT
hAn9WovoUUP2nOvYZ1C66La+4uJFFslOMdECZIAZxv/t11jpxNaYKK5vG3Bj4KrYWXwSJjRP7w3q
hI4hVYhkO5IK9NKw8UvdosPh6trgqeUAW4JfK+9Bx0Fd4t1MRpVJrOlmN/YSsU7QNGsSHQt1F/oB
Hk/aCk15ie0Br3q6mTA7eQUg34nyWKUjcYyWY7xaEQ+3rMylNHHQZrUb8k//HYPHvKYtfH9nLiAD
hofnBlmeTrVaUo26TtvL3jw8tG57PjSWZ4rq2WFu5UYulNNzTb/tOnSUx295L38BpqinP//Tv9E/
lNfJCa19BO3XcRPvUBpLjLVcKZ8RZm35Simb3B9NGiCr5kxjBxlSfv6T+GlPVAuKIb3rpaWwuBUf
FctNKuHjKiOrz6HeSxTiGKkg75++K7bXvBjv0BC9z8YvKUSMr1j8K2cIiC0PKtkSLRNDuUzIb10T
e0i9qzXqGJGPbqqhUkA+7sNCee0XjpHZuhmjfaICohRSfg3okGNagK0R7pseK0B+VoFNyXWB151/
qFeu4VYrMN9srfKuwcrOVCi9V7xkIUUY3gNHgxma3WdtQqoDERrjAy3OPqjcGXMHMnoltZPTMi1k
q5V1hVq7glkMLp0KzfXHeKbhpUaW4knEDtGgk8Y+st56OrF+oTwj7adlR1qPGcWwuH1LzvN3j18m
RTgMoPHP9o9s5mOGNEgQcCT4FQbLEjZBiAP5jYbQhUh4TBDopI/eVYIX6omkHLNuNEvvfvs/SfKp
yPX338D53pByHRtqsNMKQz5Wwb19mlLjzkoaX4M+ESUlgNjmQ1+F201tvjiiijvOtrj9y37Qp9TV
XvPGqVU0+0qiQ1fhC1yyXjhmQJHVeF5TsMJICS+6HzcOQy0IA6mmcZbq1TBP5iQ4TAF930uTO5EQ
mU93K8GyZN4X9/IqZ5MdLbUEpB/uubZdnH9f29zxjtWb1pVIem7X1vVLl20rriJN6d+KpspI7xGT
b7M9x+lSRKTMEHxWBcND6mLRCMiWPUqWcynztEG+50fJzQZFVBMbfEb5PFLKoWbIPjG6XGIxniRB
RPWMNcXFYf8aRQeUG5XXuqkuD5TpzIyK3nbZ/oLVufio8FYaT3xvLBUD84wx0NI5BMcMmV2jzBoR
bay0OUwIHPUxKxhfHkKk3zUii2oqv+9SaMD98Tp7F4Oxr3xkWE01tLtO+aFNVRaTyGy7w0spWknw
OOfbuOqpr4YlqyfZX6L7/KKlZdcukd9u/nkAXVYp4+i0JxR2W8f4wBcJceY1QpRcG2uxLXUC6DME
Ya0TOZNAIojquN4bCRt8PPSNHo/fSCVkiDICimNM28Jp2NUy2uhi2stBe3kh4miMeueEXlf7l9YT
5sNGZnnufPqTzkt2okmTqyDxX1nvFiAkx07ZFhuxVhAsmAC5r36FULjA6oHA5y8toAmUcIL6FyeE
CfbsoM4nuz1/hiCU2tYIZRxf2bsCLaYNYbkgnXxLyPcpO7QaGt+bjVoQO5bRF3OXkBGLtbTJ6X6Q
s7yQAtXifNd8TrijZ5r+6bf22RfrkB9rULpH+b0qDyBlff6YpEWGNOSu5hxijCh5H35umrVrWC28
rGAFFZIAMrRIhYUvFiOsm3Q4T7NlD6htUB2ztMgkNG4zVtrVyZYLjOGMQjdnI8avS01wf/DXje6q
ejgIN5WxfizWICwwHjjLPdmRtOrN5gaiEu57ByzePSese7mL0L4n7bMNFg8tMSqTDLVWlTrqRcFM
dua3wj4kBA1H4srjYO/7c9FstKhjjk1dhymVdWg7YQM+eKsmx7TJw30q3WXGRhY6govDjJ75wBvr
/2pw+yvADlmup7XEWNefQOss61leutZoGbSetH9f12QhgunJXhkAwYGbEASyxpFqtB++zVnBlLeW
rC5CHCfI4D4UG4fbKzbRbqpuK3jL0CuNXq4UaOyKZkY7VpKTUkEPFTdyGyeR3ujMxqrEJu+/WH7w
y9aNljjidLBgf9oIC4CEYq2Ni607Nq/25O32Xk9TbIMeF0VpnvXh9qX+T9IbM7vXWSP/jGjhvAqe
BQ9KzS44roSnaRNmsfKCa6QgkCwxwwNmIqxlJJGvLO/AX5wyj5N4LfcOLENHf9D8ohBVmNc02aAw
VAyEsg/ITsSUT+0UK4ZPYLlg3nao9g5dtNYwNjvXF2vPAGPeuZyR1E1Xs7U21B8URaOQaiUB7OFy
ocDN4T4d8WHwe6pexqF3mRoyXIsONGNpnpHRB+GTONDIcio2WsYRhLG0Xpa5H/UXoiGRkVGwlzFn
xTbCbYXZOPtcyl8SpLx4aL3rieZGtIUYvtJKaW/xSszoFhxTgjB+H3UJXjgJC/8uProFUIWsuvlg
hIs5+vi3izDqNj8rr/wjNIGq9V8nmWgxUuE5wbbQpVSBTArT15WTpceqwbKlaobxPo4Xx17mJSqL
0jxIYfIgij72DXQubb9eYr1s2x+P50sJNHTEA9fs6LJDq4zCFRWqJ3Vu0+5TV8/61ZF1Evx/hg0e
HEVDBj9OsFuoKJLLuIrtvgEkPnlZk1Wr/C/WpHU9jAC4ePHablCBI59jNOEUOQTP/Jw2ddHYyb4p
U0XMzyUXo+vMyVaswl+4PimBVROrZhEc/6ryhWXZUaHmljyiKzqmZEKRjpXs5dRcIg9BooFzSSoI
++u8rrays0FXS5vJ3grQYL1HaUKTy0bzr3JH9evQYprX3ouMPafoYX9B+uZ6ArjqqJxg93dMwFen
Cnh3UjdJi6jKNTF/wqiF9PgElTtcDV2v/XYm1BZOt9VMII49XSEybX1ftz3fyb2CUH3CueW+ahIR
1C1NxIhAGFiYohr5LJzZiPveS/aopdp5y93F70s9uyJe6TPoRswwbu1bnS32RprHQoS3ZR3HkO3v
fJTC79SBBErVyYTj7IU+kz46r9Vd1ebM53JnD9nIwv51QZrLaetIy95lGchRVQ0zTAflLnYDmV5b
NneXOfCqJOmft3EmkhBo36gWfujXlyf4J5B1Ki5mzIC8LlhSHAXN47eyEH2PKp73dGxik9ALPjts
1x+rzEuvhVfcLIxKmgD0SpsiL4mqc/GsrCMmX5Pb2hRDhui7O1aRaEKzdgyhtwkQlRuZEgesExQk
FBz/GANIgIvew6hGvnvjxRCuf8Z1AlN70Au/Xxf2BMG4Ii6cAQ8lBxf4eXl9uRg1UkKz223IWD/j
gE2+DjHXUKblVLCJicuaFu8MrW1rdr3ofZDy6w64Ys6EMB1JCrN46P64DmhHvFQGgsp8hGJwnIIN
2eOv1qxsoyPffycal0pBXf2n/2j685fgB5KuadvnFnwN7fsVkV+BN57VbMM0zYRX59bPPStBUm3Q
Pm8eAw4VqzSjoHkDUJCEfmSxI1OAeuXnjmy7KcG9cQunzZynTeXJJW3n6gVof5vMxGHUaxUAmima
Wl7F5ME3AhfQhVJnrn7iGphLRrq3MHzH8pbWTECFEaRfZJN30016J0A6Oc5H/0LrK8gfaEUAQsqt
WO87S+Src5ykOSH9Y1x18X3QX36zrqCrqOsKbBlwUlSqUT9NfimbrnPN3MuEG+0NhkZ+pulLAgzC
9qFcOTJ4degDIakktWUn8jX+rVjAv5CG9G0Ur3QUKXSWIjudVgOsPzkAW6+g/3MB59SNuAO+wL72
uVzeYP2LeZumFsl8/wueY+g8ILQXNNlxojXTTu845f0K0pD7qw87enkWf2vfjmiD+9A6u/Xdr5O7
4A+aP2gH9k2ZPpsW8Lv5M+MtVc4oqrI4++M0w3ik/SWJ/WGDCPyd0lfGzuduLpDTyFAT+wWlRoKG
UQDfTbzw5cUMR1tqeqUCz1TW+yqk5nAx9vCZNNpxCgYZvkfrUZaXYEw13BR8WF+JIHxQmxD3UXmN
c1z+LOVX3Z78XtIo0hLJIlIwrIbJ84vaiGjiIPxPUuHFl5gwdYtzF/OWjVZuRBjOzTxW7WY2tyI8
hKI2YkHTNRQFKF+fam1eF9fni2vQNYGaQUCEX/ew/O1tjOJalNBRI7jTahScrhg1iom9bd8Dogri
v7xHZKusUmEKZoCnRyr1M77qidsAbQT7jnAM+kMGHGMaHLz3zY4U9C0+M1lTktDny5c7b2jzv79v
KS53yyVBQd7bbjwTJMQ9oWsQXwOqLbggYIdTpQrTKoGBsBaH1dCybaZPacDzW01wiEcSum2EYjtM
94F0MNj/xwwK/zSB1MNTXTTsxF83qJ1gtEFcykF95PrXr1xJLsnK8HM+V1+D514VLKTlf7AKnpYo
AzBBWr4u/fDM3LTaLVTxRr+5Vp3oqfnG0ipIoWJ2vyMd/HtMg6d3fEpm1U3C+s09oKG8xY3Fdp7V
dhz16XqSz3qd1lIHs/+18ApUFx553Y2XVjbI55mgmPowexCrh0Wra6xihCefPAtenFvqouoshHj3
XZdYw9ZcDANsHDF1pBcUcwwfz84dqAK33qtKQvRvmXdpk6Rfb4TEry3QHZ4HEiWsQ2KElpKGniLQ
tKCboNgwTI5klYb+r5SOmvr+VCI5pgFGW9hcnBYgJicSHPcsE4YT/GIvzOsV8VorVEacUhpLDwbI
PByzcqjiBdghDTqsXsynbL84Julk1VcopKL8XA7LMktKOFRKqv2qzq5FaLuv4SvqT8GhslsMB3NI
Fgv49vWbAVCnsK6RU3XaqBxbLg0GYkzPfYEr/gprIhh5qZDm6uRn3qgeTxmM80l4OFgS3hxsakmt
osVy+lwk+b6ZpWTN6YLt7zRQlOk6CublTU9U5YWZytVIDl0fk4ZhohNlkFUr/DES2e2gUJrlhMvH
uZLvFi4ydjZ2Rx1ahMwpDFb0U2NXmvHUVSWkcNr9Js3d1zMPjBf3Oxyg6LR8QShovgV7sFTtJ1Vz
YwGdJuGYf/tSbhbQi65owYTo7F1dyP0ELlBsCWq4wjRRgzwJ9ua0Ufs/uLU60CcLMyCn/BNt6NyU
IJLUssloeLraMh8ajVl9clz0x7snM48GUg1dZMnuB7jjMruB9IcgR3JxSeXZcpUMXPWkZjJMqzS2
LBZfwpHUycw+Q5eDMi/+WniSn7YaCHyAGXin+IPI7FMM2LfHsz/bCxdZYkqUPuyMEzEnZZRekZAE
NoMQ4QnhDdDZcPDdqeUT9U13Yb65sPGzFI1KH8LTvzQcFjqFCthHSEA13lj3GRZxUFSBT6gzcxzo
3V9tcD5XmbqAcFAZIpRZ1Pd4kAu5W2LNYOgxjCvzlpnvsE0EZqNPfXOLo/kiuhbWrMNJNW3hN4rx
7MSOE1ToYs4Tm2vt6D1Ug6fHQ5j27zQ41ahqrZmv0gx7twED032Zx9Oryv0ZmqTDDR+yY2tGnXRN
3+E5Yie88TQgmt71aEb9xGEpEIYZa6SVUOxBtprUZ9g6rr7Q7jEcZ9DcrIn7EWk85gyH6qP3q3fo
7kCs/av1n2NORk/e02iZ7ZJWZ/HCoGFDeczDrJDAcC0MOOjMyZ2azwKEnHX3oxBaVHdQI/7lTXS0
V5hZGnzNF5Rqw5tA8FxqBR0BdhgVKnTCwa76PRO2wfS6OOAOHfeklkATK0vM7e/NvnCth7VhyDER
l0QpxpB8IHU/RXjw+/ttZ+YNxhTwfw1eDGHbzRhk3NUF3f1F3SGp2HHWljdAst1t9b7MZnqndBgr
Rco0DKDbi3Jwby9lK2QMAMSSso7GafuvW6YjpkhTidHKbmaXO6DO60D49aQzHjn//GbxvbcFga0b
MJL61cPOe4v4j6gCGF8QCaCrLdiVY4yOJvGJB4pp9cRpHvAi0e6cyWQuQRGRMNNItzpPNbdnF1Yx
p87Fn/NG77aXYogNOLJL7/gsMNAhquBWtXXJVzZHZUv4zNkck8iJp2T+HB3VT2uiam7kf6i60v8l
UWbw3H/X/qZC8Zmw0LqInRYYX4V8Q6kZz2lygaolakNvxf5lusfir1bPaLjEhBbmZe0VP3uWpk2k
g4h2cO1vMQV+JPg9rDeyqtTjRw9kkmM/YRCk4joeJlbggZUPcXfLyc/PtcKC9sb4hU60uW6WMkpj
iWbt2xWGqmWLeD4shLUSeDoYMmpXH0rnREWkywsALQylB2cMUGBwilsEfvd1vYIrMZgd55qGwrmV
PwbYQeRQUmIpwO7aiPK2Zv2Qn0FImDRHQb4cvXkvWkWT/ziVbv03jJIZo8k0AOqfxd4j80Vca4ye
kLi3StAL7tjZ/+ntvIHDNkOBKXAG3YXh8D5nxZvCSVeFwwwkWZaFksOPQhHUVvR+00tcfqxbjFF9
TN+TlMDakpbfkWXNNUq+wRpaXOCNhHDJvAS2p6Hcnh7iQOvdaQ4BVUQBEoRSGGNgDkI/t0IG2QtC
oFVjAhrd9ObuxQRx+wTuiUavBSq/N8+4+N52/G5FSLzQYc/Ny6+FtpJiYgENcRCT/t9XgnnC2bYi
oBrb39ERLxavlcDEUc56AYYvMjds7hvjwNUoeY3tk093u+0EWBRTUssweLuE2t7U0vPjA6yJrTdc
v+cO2q3YvH7+NsVR5Tue8QlQfGGT9eJnj5Jd0/9/xnglH54GyJsaXd4Ke3kH4z+/LCyevk8axOaN
fMbkH3gCM9KTG6GiX1rVGMPvQJ7Rn/q7c17NqT+mHyMSVYxX/mQa1bEnopREricpnrjqCirHbc28
qfJ4oHJ5IWH/HFi97Z9ML2s9ir7fE3dehqbgkDuju9E3lHOh0M6dq3/pfsuEdGkufflPJUnzbcyi
XUEXZe2WUTBjoJRmastp0XlyAkn4ab6uO1q1bqLnC7o7ahA5anNRdqt5tQHJetiSc67f3Fh9nZ5q
V4m0wnJuD6IGuCtML5/h2ceXGbjUVOF1bTqf9mJEou2qKLhqQnJ5DzLYrofev2ARfJQ0KQXcELIH
UBXgEPlyROPs7NNbRPuss7iIa3gfWKVuFs90brtoDcySjbFYIRzkxv31uFtenvpwk5eLhB3AZbST
eWs29WtP0CgJDZzeo4jKBP2q8/O9toHvbyYlPEZmyURAPUkrej2pCvTpepQaC0L6Bv82CWFuvelX
IubE9kInEo1OZjRAm46u8G1wF2eaGX0zfM2i+ZK7mHthFTRhG/By67MkNr9A6BfBa+FLjGhCRQs2
BbR8Ww3wdwgHDgztauSJhxkcc5BkgWIfvF4LwDIS1uqSQTik4ki7a4sJ2J3d4QeD0C8KW5fP8H2E
svblIDhUVOqMTQ9ID0pIcmI228YsstXWPZhczAqCUVxBSINgYiMo6nMAYOUVHWRuseUmmnpTSVTd
twqoMkQ+hWMHd7JmRe6YeDu2bn8EBGwylbna5GT0PTSn4LSNjh9qVmtf4Lr9Zvzb5QH0LMF+X6AW
+wyyoJZ4MCO5A1jtlBaKsKKwyogVoffczffHbaRlDdk6mWWO/5R0sRRtDYTHfiiYpP5M1H1vCkTn
Vd0/CrQfckkD28r0PDkcdHCPYrvQbpvpA89lH0DY1qR3kh9l+L3PNdymETDBG9wn5+xnikaan5lX
tJKnfA+yf/2Tx5UJN+LE9gzn+xiU0ybAezX8F7dnzv0HyM73yNgxRO8tAwI+4neA8SsyfDsJHQpT
lhE7yNaF4//drgsQckwdSeDkylDuJkcW9ZFtrEHRzj8PsDj7gUjX2D5jEbNLrh2/Onw1MXmFdDys
pHO4/CIdusmb9M/Vn2lYPMBmIE0XvTHnp3HvuVpnYqeshcXMzz8AYE1FGb6zVAm4kgvt62hlOBbm
wgZDf3CF8SMwDk63NphPyEDEJcoJftENnJyRJRWwdcmKMIgTQvChsVP5wEvw4e1tAOQmGHVrahcG
7M58oGEI3Isv4D6d0rU5zXlJ7utQ4N8Y7q1iFMZWS41OxW3it5lojGPszgjoq11SSvrZ5vfhHvXk
WFoNxOrOxd+2hb+mc4TG39RWc0IpOXgIqp2xaou6cL1pO52Z/1ouJw86GkZ7NskBay8OfTlMunbE
w+2mQyZbWm+m66cqnMW1ScgEXKPDZNlfyQpDrxaxDjls0daiWywHgdhQn1KlzxxVg8lAbTGKICP0
RNueXAFKGM6YaASD9ISjtg9O//T+jxrZjDZ0UE3AWHOjJWN6xWPNphaYpIzzea4aEeB2H82LDaa3
h60vapv8ACqO2A6lh4w7whVVGgDFtgenqH4xNlMn0mIHwKKN2rardmueGpP074vyxfQX5Y7iT/Gk
McUm+2vpvUr79fz19yubzfy+WPEGcazFcLWTzge98SQWhauHfmmTs4Io5BoczgZu3/7Jm0YYWTO8
M5YkwsII0gPb0s2c8eGAMVqsXM5hatlwI89h8gFNzlMfRHTtlReM9yu20+5O5UHoIY7KidKmEBsG
4vS+UPZ29jmZlVYD441OFurH8BwKPGxdFghpGnRUCfB7xWJFpyt0BY+3PjcxYA3C/alNz3PuDeXw
x+RGnwYuqS1GaKJJAlT3KNwHTNpLgSouV2GwI45VNafpyIWngbR6cZB/pEBGW4w64vEQAE89yHST
QOMdEmOhZR1JIn1cx+HmPYt8LlqmVLHss0C9AEh7GJYfH/2CnKCqaf4zf3+VKhwigJi2RrVPNbI+
5EBi3MHvWbGUzkFBg0vvuXcNpcWi2Sr4s//0GA+yWZlw4/M8Mwyt1e8t8mysMbwhlICBuUt6vdsF
8G48kclPyN6azW4TGTT/ZkWtViJ5Zjz3wwd8P4x5V1jOZP5onh+egEBqcz3gTDcj7DccvmyDdjno
dmixNY+KP4Yqz7g9V+eR04YunlKQ/f2ZIPW5OX5JB66LhTzQleFCqgCgQ1Y3NjcvJttQJW4sb2sx
WHEB1lEmo+FPQwU235gWiML0VWNhVc2AEqRZlg7t14J+BlJlxSRe+WIhuvHRFponszAZp1JnH6Gs
jpxAVPxorNA8eoTgQysKt7KfOxsDqjppJnykMywFOzrNsM+AyhTKGQVLKp4KZH8k3RNylJCI1kKh
ba2ZOfUej654g7G9P0IcIb8IodOVlrda1rZJ6dmpZ9wAdgZqO7OE1p1rv26shJKWg4syzG/V/bmU
ZWZi5jvTeNdAliffVQkdX9rg7Ie0rzXjoPHQbv3TxJ6t0BpiiaU/l+mwHxs+ClMPubbGkXVx/Ay4
n09GySmjJllQfTuJLHxNOBU3tolzA1z4xVk6OGPhXg0J0wAxhYojUuSV5IkfhKD/xieJxDsh21qy
9w5ZXtUxXmEcIYGbus6Y8D5QO7eBe9aKaceeHqFL1tFE/bJQOVvmbBQ5oT5uKGi9UujdoKF8Ph7s
SAsBz93pvvHMHL+AgVlYz4L9GdSS49wPJOa2hZO39EIy395U14Da0lGXJCclcssqm+jBIhN9bS+P
0fBKExC0Y2+KKHitrAUlW/YxMdtbi15swMvuMAaFMo1LQaFP8cXwNBR6W1dgzEQTF1Pzw2CMSF9h
mjFr5AgU4bDAJHlTb27mAnhsXO39AushYtUR2wKoam6pUC61f96YTfKkIlR2ivSC4bVs6Zp/Ngyz
N6ypt74/3ga/WG9nXsspu0GT3THT6dSuJa4HGGPAWOECqTs2HEFMQBUtAFy8q7sLVh4WQaSIRezP
mDE8mcQ8fgtCz7Hvfo1goeOVlEe7k0DN3S2wA3b5Do1t8itP5OkMLgsmTavhnnROWPxPAXX/Lydy
XcJsONJcA6rYi0xCYjE0uJkZRnu/wqPse9hNdMXlvkwj4VaL5B8vJD2gSnASZVXHNzULBI2RYT8u
4gmbeZvU8g/7pr8p9BGA4X447gCCiCezCVh2zr5HEN2PcLym+RUgpQNPoDgZQ3lV+yzwJR5IB8EI
EpHJlmZd5gDTptXiXarkQGm05ixIIgRNTmbTU9zVxE+jJA2c4TCViAP4xueGLiBg5FLfvnY53N8j
Q7TW0mitCYJbqUWpkE4/Nq3nhMPtgczzkEqGI9eQYY1ySG0MdmeaaQwVNDNox+Yr3Mz2xd/upMTa
38jYILB7XCju/gmWFNx+rvA+RLe0sr2WI+tNOFfeVwCZALMGtLpAPVtBmxmvyTmzqLws1oEjccDL
pP2uWm3uf9T/iYtMhC+CJVWSXpMpPKvsdqOYN4CbzJdYv35VDw8Je475FbzZcQkNvJryW4fboREh
Xj3qGE0f9WoXgZWDpKQrk9YOp5AFifeZ0/tTg0CLVM0jGUnm2/u/piWb0vLxWzuzn6ZvR0OiF1FV
Yf/jK5JAT4CUz6VA9gApvFmt5OHP07D3ZmU550vn6BMpbApBWNyh+stYsNmReNWDhrKI84l50ceT
9WaWjwmunhG/hRDuUbTWUeFosuqS1IxXr32nh/SPvqQaS8vYBdch1qH6EazcyQLjE7U9Tj61R4OE
QW+Bwf6PhjU9+myepDNLdeoLgzq9sJ+CN70mefdYUVm+4Y88NeSQBfjogRkcp2WEW09gWqkNR5Qg
Vv5smUI9aMKrpYJWhUsJH1nZSi2rQ9cMV555rxqTgVaMZcrDOh5KoEIsdtssLYFjUps32WWwV8Za
KTQDRV8T4xhCB+7rEwzVvRU/xfhfDOHueF5YRMbi85bAi8dH8aYV+kIvClYDRXxJK5OnmAwpUl8c
4v3qpJsjHvDmmyhgN2bAjxuQ3IT9xHoRIQFeNekLeDtH111+mpv9yKWGZOytTh3YF8q0eO7p8aIO
k7mlchTA9sVkJxAfMZN3hGYnEVyZkpeLOnHyVb71BQvKSoKp8FWfy8Fp79TTbAxv6TWtbsnIRno/
3qWNyGZOTGCnsT+u+oUCn0JW4E7Aph+Hg6vFT73drmPCo9s/Czx/tI6KI3VFeMu0UeFwVDogLFm2
flmVUEnjWMVU8hacivZ5nctQ3MI5yOBjoisv1MOjHvPOgTeZIs894Iv1hpJr08N1K0WnHrxJWDMt
PpBKICAew6CsajcMc5bQw9qngD5xcNoXrMWYx1S804VVAPzqSIn8yJqm+lxWTztNI+0UDS/o7yFU
KXl19UYaS0G0XTRY4Ztn7LANd7t3rCldN2ijyW2dD6871AGOGlxPoJnHwWU8LZYXxI0dJDGATgHD
0McOi/pyJANWfPS/ReWIBv/TSyVDwmpPP7MQY/WBpydxvebtYVMq/c8Lx2NgbpmX8lcFO5cE4ZbL
wZsC5wizd+jdvVHX1VNLQ0k838OpdW+MjRMfweySqoSHFMo18vY7uc0+0H1fzaubvxA/7eG6zqzn
d9UsvSGe5YgZGd/3aGLxDYhuvLBIA7CA1xCmFY7Luw6JlolYjRt6nhiDPkdtBVO6w5QnAmoAg0rd
yUMSlMMXxx2CFXv3F+uvt9wV7eXmnDaeZ53ef52kRQCqAOHaJxUa8k39w63O29UeVYqfyD/g28k0
Z8gdsoT9cIryC42jfAvCwdCl3Hn//0GROP+6HlduO8vpzeETL4wXkhhPgKXDvdWvnyepjjrS161o
1ear/gXw3a4a3dAEY07rWIskvHDq3wC/FLFWfQO8qZWjjnNXWEwVavkEtXauDBXmkPckzCErSDq1
5bl59u/Sb+904wkJF/cccXF2ukJzolhmBCfi078yxjopRaufyaRwLTL+PYEN3PqVtelZ3TQJj31V
Z2k5ouMHYDL0IYEHXEmAAAxCYMv/vFzLMf1pJ6Yl04rZXntO2ABZFFtl/IN7kBP0cuqpWFPjOZnG
LPutrxnYKk4smLIjseN9VWxj9zTZupFtxkqTZV/OwG2ndoa41lb98g7sgOrNmeB6xYwRYNsAWW4c
aHHrli04RHiqjV3P33xEBwVLhXTqDEcA1CADOMBZH43XdczqV1WwL/MZZJZAR6kQSZyDq46YA2eq
9xqfXoKVhsgwZHAh9icXmCJykSiAdrC6fma6QvT2xU9ALlVc7BnHcWCFg/8HKNVJgwkXjXRZJyGF
l1d8/OkER9SJLbqMIYWcXIwyQSB3bXbci+1hspS6gEpI6gwKTIoejoNuFX9GIj3XUiBWWiKbFsp3
DPQUvvqUOoIe8vouPVBlqIofVwOANyuLE7N9aTFJpnWh9L3+MVQiCCMveRo6skogrNTXiPm3d1uF
D7rQ0dI6G+o4TUZCZNefsuVmT71V1PPZvAk7z6yV8UdFKUu+PVlmBdo6pg1EI2ga0m4zTb6YQOzD
AGBcS72Qy1PQhA0n23UaLbAwdGXV1a2kH2ebkiH27cyWS5uiEhti63Kb3S/Pj+C415Csny0ymi85
nIWkeavB3aKp+8dPd7VjEnpiGf+WWO3jzijjeF3XkOTkxz+K60MYfFuldnw0i1Td3cMXvnGJq7Xu
smQeTtTb5QLVn35B3YjnBtCFSH3uUPgngf4vYcMQ5j3bfOWexmdrDpWAg6GrE1wujqc4hyCkN4bY
3mhyik1x6wfqWLEsGRtVx7CZgLH40ro6xcyaPVLBU70IbkG/nNuryFgdrI0Q8f1dLS4kgNPNr5ay
G8LEuOkRYxx2O66Qlz6WNzr0ZvBv9dZgxF1wzwlRUIJOYtoNHNbrdjY0rxVCTiCkJQCPFHvIBuOn
iMqCGebTnEWtIyHU0uSTW6zEZD6gsut3Oh8f6OCDaJnLa8SyuC2ieycYiqkX0Mm0P3DGvLHdyYiV
T5/bOufGnYK0pZabcqABEIBRiVDlOR5mTUGdVV4ZnSjlTvYSKVCb3gTW9trWBtxHmmlo8COOfasx
SAAspJSZp+p6M1TsWemJ5A+yE/Reog9bqrwk/7icxggjG6dUtw6ngNQKd4zy6mwglFc41PN9AQbA
FU/HE/nf4vmm+X18dh9bDALK09OPalZCH6wF0HZ5/ntd6YsSJANrbC+Bg5m6PutFFdrRhFqDe2RI
Rkl86qljHw4iuRPvyKVqdBsAlYhrqPa9T2HTsqNafvZYTV/MBISNbrzC/kjszfBU4/fFefqH7/6o
ly9YZ3zs8ArVEjey0tN3jTjllLTbcgWkvwfdk9y2TT7zD+9M/WLMEBgG3KZOUhZaILaVU8RJIb2e
/NAPCD9AEY8BPlCfuCQbCcWh9+w0m95b5qaFnSj+BOQnjj8caPUBlBTsKdiYB4xX6ufF7pNJCFOE
HKNNVuncFJHSD5GQFUIi+/yjKOM8/Y8uX062xf/gF8K5efu9UNpG6bXMra5tsTUEUcoBJAQpKo2W
A39AlYjYed2jMUwGwKIfGgkNk4lYXViUjgjpVDZLhRZ101Zk2k8qT+0YFoNUSIf3PSwK8jSgnw28
DDjWWsBLZa58EMravVlWYBk5p4NUsUwLErNNsIsYjjcFxlBJJ+IGy5cOLQsAZNKdk85VPZugCe7H
Vik/4hbCbUK9u5SBblxLlKHdyGtg500DM3Eb6e+0vCpmhu5tLafIsba+fUkJUyORfDXkVzUkTPkk
AqzrJlFyAgcfZ9IS3xY9ipxLku8EOgCHKSgwQldZMOGo0bJ8+N+A41UgcY13MW4jSUbo15n4sRVz
V7yVBw59hpLkNAVNgYcmNnySBbJqkBjZuE8BePCaN4P+61DopIkhpdr39bnuB1pwxj9r7hD6hYc5
LB4RsIJaVA0lsxsnKIm1VyzDyWWSeL2rz0EjgOwecjZ5mvH+BKCAl+3lJ+Jy9YCQ7vI5BrZISamR
bCaE2w2MQeCoKzuRmBebSrRgFGgg9tL2ZvoO02Jv5ap0gTx31YzogQhGuwuHk56rNijjN52l7C0y
O5JxxpuqmBemqUaGT5Y+AFF54SyIfB6AfhpvNUnB8SzxR9KgxV1zY1qfww/Ter3S74VOvUcivUvv
oM0yjqJ2qy57aIj7NNK1+Yk/9ueq1NIGEyTT4E4yw4SA94co6e2OtrbAAFRo4AedakN3iFU/LgTT
EdbsXiaJ/LuWbtYp5N8PsF1ctAHFGuuxZlZCj636FkZQ0YesWBM/IOhXW+Nb2qXd1TKcWdqN8ynW
a3AamAzZWNSHwOlSRuSF4S0nNg5XP+RfI/YUkTBxDoSazl62tpp+MeasJ3OyJfEdjtjkvlRvP1WZ
I3RQjj+EupgX0LDPEgBZF2KDLQlXMho4AAyNfnWBTR+M+IIwzCvouHTjrhIn10gEcDGQ3D1uYVRn
CJBBc9JAcB8Ka4Bgn8oZGFbPIP2nK8k6A84IRrfiyOmHHz1pV8fScrlCwnNbUeYurNx3RF0R5mE3
M8lvRsbzQ04/2mwwjSXQsc+IWR9k3CgvKnYTciSXiDzZkqX0uMWA2GYjZzVjBhPIRU3PQ+q5ya6z
SH7OIEPEuzT9Bb2lwMc8kZ0l6Pd3+twWedVy5ePu8blORPDYemob/zrpJZpJKmiF3hXDdpy6nuei
9sejF00STz5nMKDYFcYNgN4L0dhthnDtk7523VPmQTvBtUTr4BQt1+PNGMmaeg8YDzj/Nu33oJQK
XxkSPuYLt3cwToC/VvKt20tkPzbhZFOZ/+hXdyT+SGmCM5NjMfA3EY8qHgiURGNXD5+yXG72/BWd
TDKkqCPMVkJ4j1Xi1187pSIl/gaBnbDxuHJbL20ng6darBFNiOiF1r4CQbJU+gAw9Zts3qjDPbkN
CcZmpa5DQMkOLv3+5uX36Lonj9oyiVEgOkXhA/e9xqLO04nE0RSvRtCQrGAQ3CEDFMXFDmOsiWTG
qVCZn52hXWhJ2KuachXXhQmXmHVPQmwmFQX8NiicREw+TeSeMXVEVnTCLXhIlB0uPatr0zK+K9xj
lfqyAqoiJDs5zxjIQF7GJKW6BkkVwoPMeB/07+li/vqfXUahxnXAzulKmWGMwqVbcVx14rM0nS28
oVVUOaJ38UNbdCOt9IY1gL0/o4oC1hZyAXm8HPIARzLvHeFLvMHwDIL4usGdB/za1JPE6c+Gjzp2
ekYHYfmnMRsiJ0UoiZ9l4M4zwrfEPVETfjAu6qa0XjqypsOwcZqa2Q/WEcFpftrs7Bhg0I1voVWj
iu0ugf7zFEtpnlYBIPYI2hDY7nK+YRt0dDBXXNwHKuXGwoPb3q/ylJkKLQzh3CZtlZh1jS6zS/lz
AK0RKo2A9GUMH4pd8foJnsbohOEvNUyUpIzFd7QvDGANQuBa4fl+NhvM3GNQxEZKmj0ykxmasmSf
GrO+TE5oXy2VltLKqL/SIbSJ0WP6DSWfpD9ZpYMuUgUJoc5UyAE3exW/tro6oYGZLn5gSdMjdZdm
U5ax9M9z4fuiCUU4gVNSVvmLrlPJtqIQXhOwPv71aCyZ3EvnxieNBjzlztr7NEFHS8HkOfK4CcqT
UIj0uT55MToF7lPHP4HIoDJBC9Os3OxfnGVUc5ECPG5qrTujJI2ARp2hLJnAp+43fzvgFRPdKHmG
V6mmJOjeC17Qxtu9aEJOUlANJGjZPquDn8UKBlXQsYi6qIXmuUA38v2CKRBkq98wKw0jFoObnTMD
eKsKyB/C5wUAo8jgnCCLeAKLike/xrln06BYPXhBre8xl3FLijFguzo/x2S4QUKQUPyFIuzJ3RRh
PmO+NTCrdJgnh+L/JSV+jqxPvhQfXNDDxQakAGWDXKG3iNx8F2NB3GDLikAxb2auqHm8hbUSrkgn
NhTOMQOPFYO8c5K03HbOU+J/cbjzZY7zjCpF7CUMfsUD1ghCGikF2cRW5lqDRdej9zn0AdXwZzbB
T3elKCdpgFX/TKbP0XRGtYCKWxIf5tyQmPtFH78lcjFsqKYFS4md7Rh0nMb9Uvcx0O6ZoS6zo/uA
uhYk3bazrRYGr1GEdj21j0jnRnZ2pXZbQuR9PKteK7oT/3kvTfjfTqvgggjLQN2wOs+jPIQt5k04
5/Wzn0RgEmrVZ50lzxcZs/wuwxz0kC4SCmt8l9qjtWJ6WygBy7yQsDD2IkVaeeZCdsX+OTDwWSfq
tWp0j6nftcMruB1r4usUzD2peELbEV4dAjCrQJVnxZ3WWLIJBujBf8VYuauYIKjKAfL6D82jvf72
uE/Xs4IWRz/27VKSXuxBw7Ni/QTWVWThdhW1mpZ+Swx4MbzGRSBFZyhlMWTAWSzDFzNxoU6xWhBS
RV5LJGSv029WOC2Tqb6cnv2k4FX5uyGkyZxKDlmkEIryUN4BxrwWs2Tw8gs1W38e2Z9wqfvmlFgp
swHgf5LOdLQz4bV5jvoq/oEV+h/qz6ygHIsxSccGShY5e9dsj7qarkzh4OcWHS09DCqEE4Dfs5Zh
h6aVFbVxAbmE/nBPKeCS8bX3sUmTkvRqbLgxeXXJFd53TBW/sIoZcy4mto85KZR3RnI5EXFvI5M1
vMhP1jWTnSCH9FwDicDR7afVPPe8SeD1enVafE0GC3/FEqMmoSRbgK+mQzCfcyrYz1tr66j0LTi9
RhOepl4/N2EAPMhlaLDmF1Y6DKWMjO81gpfuBor63FpnWvAyOsqNxSoPLTX5SwkhVaY3pMQXpPuE
5TUTp8HqwTWe/dtb4Xa6HjA5UkO1mZkO3XHLqwpldGvK+VBPuoD1BCCZckxpGSwLjOP0TjSdpQih
zGrSxjMNZGC0mKNHL/MS9qLcUpbRdHW/v3unMEhzsq21g5ZqdNIwui0//qG5NWcPh/p3i7FXCyap
G2N5hIAo9u7bxPc0rdALTOw2znMox3qTf2KfpGzRnGRgJgL/LqGf5L7ZTaq/zsa6hTmtCM0BGAlR
TOD/04Gcq5P3/kypJ876MsWnu74gbBM6RsaQN523ZVtqje/HCCFv7/Q/A/fTjf1QZ2pT7+R3JjAx
qQHEmISd8JTbvWnr1p0J1cBFryjdfqVIerHy0nPsNBCeHwhETYfuKKyPoHpNW3yYyuATshRk6sOH
gzhJMiqjIanCr2k3niwwcibu/96XXsrXYqhHIHOVsfMAh78VmVSqHJY7SctzIpNb+IzF8qWjastq
5zBlaGoyKTCPzb4/OfQTck8j632Kotcd3DrDwFwXQjm3HRd/q9nznXlZyNCU/lJ2bt1lotshgQSA
tz1ozxohko00WsGhDMcCm6cbp1FVGin+vDsUlhNOxxkXMG6aGSCG4zd5PzU7rPrtf6QtBIPCzqd6
EdaYNQ5KHjzm1CACYYMt/nl4FztL/UXuYLOnDemHOGdEnmvVsQFJJstxFinA3NVKXaux75mRVW1Y
aaiAZPrZc3dSuwCVF5lf9hO2vhYRY0Jd0CtpWzByTKS0p0XTXuIWSC1wCuvzFAuGV0Yk8vA7OKuZ
TeT2pK682wKdXzwa9c/39+irsxrFnfGPQvKcuJcQNuQfjxG0EA7YB34Z8VJg+lvdRtMo6P98RYbV
y1+Q11cSMj51+7N2WroQqXJU8P9HfXwMq8FC1R9kqJxzy9O71fqP1UiR7vi5RHIysx8B5QUdzalk
4Gjg+lnmNOvqf5Giqqog+ZV0xxbwnxpkhMjVdEXs0yJnJujQDuLDb1BYfdK6QHblR3W/pI7KGPTw
dmxyHBU/GHg7KvYjT1jB2svR1avM/e9S3PDSsvG4YExGMnQYtIss/cN9lAPATBfZPn12WdU3R+tk
I/60M+wEdx86cQYqEj0GUXRpitqZoXRRPd9YcdeAcxUVTg8tGcz4uiHUlpfi9q/CvzbEZN9CvYOO
WGJcHmeV4AGV4inAx5YRhm2ve/Rs/jZSMat91vkpI4I8ED6wH8DmuaQ6KzX/B+cgiizBHG+UhoPl
cFsKnQ2Og6dBWIkk2OBce1tAfJtiL9CJMFY8myUBX03pULkCgSRTNOH2yFF4Iywyq68yEUd+M0g2
ESWHfiCVx711zixaZAY1WfyX0ZRXYU6zU/lFNz1vLjJ0NDgCWRvSIpcCQiHhGqN2QE92CtP6AAb9
jrcuO5P08WUNgO+4uQOZcNHmV5lNxeaW3zPxmGcU/Mi5Irh3529LNdoDtHt+IHFg2Hm/WC8n2pK5
VvovtnqeHkff4HV1GLu+FIO0fQPS3+4xQ1YpX/qSOVfQFtqNpcpFIGcgMMCSMhxS+RqXxbSNR3bk
8LPAu8vXPLNLC9ET8f+ob4q+3V+KltMUnOGIDVip0fyI5vZNrPdn9AtVYOsXj2aL9D5xaFjlJocX
2E4CTpdrsd6iWkyMzL7Gndg58/YMEG+PAm3sBNXYqhm+WvkqnZCmzIo6+M72Q6812FTfwuiYr3YA
xkinCeeEN9qZydwM1uqWCnRhhMf0H28YiJzM9AigZ/kCiIR43GY+JRoEmbOmDJV3B/06NzsjXwfc
hds2+heZlBLrgbfI2krfeLuvBZdDWH5/e8vkKTAVSIRfN/matfjoZbx1gvUmoxwsORplVpoFECPt
SHCpdTUqmSXG8St+3j79T8Ez9adcxDtc7oWK5Dv5TrcsfUkCWrMRsSjOYkgrhuG+hwdzZdH+LfNP
Fbvh85AXOU3MylkfL8TttxxbJ0sPn97hrmh5ie4DCDBBSDzTeX8W/Qg7OWsbu1YV4YA2sDVNWeOC
ihxKpwl87ATCLe4ukKhwKiMeJ7ZAYyBZTEMhSmLBFK9lrgNhFglEIsNLV4EkiPzipwXuVVO6axiT
knPGFrstGkYQ/ZeBUgS37TwINv6ZolfwTQGesLKYTWdtDtS4N/hfn7v4fwClG00tfIMrA4Gq9lky
2vJmsSycn0kN5qjvfK+xrDfEgUUliYhBTqxAcaXVRYIHp3PTPIrs5a0fySSq0aNWiKo1OaPc4UG8
D4LEP64KLtqnbRX0sb+b2+m0vZmDXKSkxdYL+tF0cg1OBtsjV4nG8xVtNYkX2F9eYanFJEuDaluI
td99GGD+D4Tq8O/vOh+StK0bA2wKuFTVRF+cl0ySV+6OYYbo7Lo9BZHHvakeTTdNGjO+vWpMwfdp
pThylzuy8agi9QxO4cNAgm8UONYsR+oSjVbEC+7m7FTkQRF0CiWEDSu5LZe2SqxcsJQn5tln5n0U
fQzm14//Zhj1sNFytAQKprmmcGDNTsV6EX/u9GTP1I/n+xNzpqUQsLdL1DhItnLuUnnBbTL8TRCt
VXy3GLTb/0CDMCpfhDqhp2AqOL180rUJSMhUor/i1HKA7eutyQywsWpuRjD0N6IccYLN8FTNZnoo
CfDDK2VXGJ3LEL+LKYp/y2gDMD52dM8z8yGBY2dMo8c0x9hyKfHYoAKx7x5WYSAK/IRVZT8FgE8K
LfVBrNixFtoRCSIl5iSwIyJC8XS5qXIwdQ1XsSCraNvQJmn6hY/JvIDHrGmV8x1GRHccMXgb2eZz
2jNc3BX18gYLpCM4X1Czjn1wOXA17IaJxGesTuLJUEvOVMM41fNEM7C423xMme0Q1JyfDI1bdmS/
gVDn3D4stEhQ2yaE0UJibv1Lhp7Nge9aFvLnmWOcflczuVHA6wEagwpYbw1YcVbhMEDS8uUjH/KY
I3YzrbpWfwlLJdI/so+EeRk+NQPtzJXCtgJm9SB+qCtGmGYtwC7wEoaTYAcW8ZCoYw3WSmzHvTCg
cTZMcPKIpZ38hCTv0iJBsvdpQCUktdhdEYpDmoCnPpWEEzbs63VaMSCDlzlmUYsL5dLBag1MIdD4
Ky3CgHJ2Vg0W/cqyePwr+kAi7agI5PVReXHgRNxF+YNSAq0cpRYqGHmrZIQCASf/xAYmX4NVy5+Y
C2iLdma1RlPobBBBA3qnrNI+kz6gCpqPEV2/w98BO8PKcSHV71liOTvtXeIQxRUnEOzT4EhL4qSM
RuG+c4csJCfy0r6oNl2tpvJmBUF//70s2jGAk+eX2iVnGnJdOG7pJUn7r5rW3dJxJs912kiFzdtY
gTwb+fCSD2/EdvbfHecKNwVwUElMaF8dv3aQN/Fut0jrjuwOf4i7b7iV8ZtH+Mqz41pMw4pmrRcF
FgJ1uccPa2LLeXAv5Ncn1BAn4KEXDePtOJ5X5HN7VUbgDppe1GhDnj13jSjh+tz3fWLHQ7uRMrSN
e1WzcX6JDMabuWmx2JBhQSt2hCom4A2VZUvmRSN9R6PMu2RRoGdk8DtYghsLdCFbuWZji5wSZ4QF
07Ic5L6JCyH51ksslFBzE/ejwFrzJ4vI3ba/r2sfS0lb2lCAl/3isKp9qs5G3rkpem/V4YymTSoL
Pl1Ckgp93D3ezGIhGaQ+okd9lgt1R2SAwB13wnnDtar9+uFowJrU9gXplg3L10oHR2ZF8je+laGM
fQ8phAw2N0EDhQh2/JSklmX+QpHMR/ds8cQY6Q07oIf8FsGBk+G6jCOC0wsEL2/EjtImPGEb343l
zIBmp82DMbp3D/rdPZ6s+a5ElMxTBIS4O/clAsqgth3xlaDWrzx/5kxdMeqWgQixHBVi8pf4tsxn
02cwUzbUHa0J0gn6qsABxN3Zu9G+Z2mY9wFRd8Pbzj5o1Fv5U/+q+/wkerLhyQ==
`protect end_protected
