-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
jYrBVZTTka/eH2F0Rql2CiQiQRG87r/jDt5hGSV+PBxNzhjdV5rIaeCHYTx4XgS/GYaPwhv9oC7R
ttsSHaiQJ6T4sipkZflwG55AQ7PB6NtSAmI3krLjOD9pkX7hFr8wqxSOes/d/J471ws9ibS/aj0M
0IRRNwJPmSg8oG9VM/yL76nq/Ye9HmdMnV7YFgU+9qIfh3gEA3bu6AUpxcUS9cYNZl9c74BPxzF2
Vj62bH0/Y2O8RhBi5tLU37TS/2umYcMQvIrM+hS4mXv5zyOEZtWPD7JKavmp9VGzxM5CLvpmf5sl
pwsVtG02qAd6F59GBlFmRW+nhleaHoDpBoyGag==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 70960)
`protect data_block
c+RHRvs5R4tLj0V3kVSl9+62b1xxq8/fyMK1qS01DfgXgnwF5kUweK+hUoqRewISgF0gf6UAnK2Q
MRzaKnAv4jlFa3N5qNtTY2cupMtC9uGKnmdeWvbDHxNCMalfuKRNTvdYts27TRnRVBEOKuAKlgRW
wz+vlcIhzFlbTsYKO9X0gC4w782M1JNZ2i8LjHf71D1a3UG1yHwd06qMq//6de7JaYA/k/N79Job
n3OIEn5km0QFi/SF1gUBIb17L+lXoJsp31PQA+VuDwN66B5AOd14th8IwHagdjMxWWLA09wqhoZo
J++la4uHsBccvauJQ8GAJTAa48u/NnEvr57PWiLympLLXBVER+o3r6UMZd+d2bHOLlmKaXDjJbgb
/n0d7CwdjY4bxztvBJr/CB6WrAXSvRHraSQ32t6ZxbDzZtvVB7buSEXA/sIUNDYC4YK4EWO51yOG
keCWwLhkYNFmTQ+NuCUzPh8YsHSu9Fs9ll4pAGwIFiVBSbPEUcaEziMbWzlx554O6kC4w+g0QscP
1GTfkOSudBfmkaQiSMC97Gqs5Djuxg3v7hVup7Jdv5+mEdp8jHq7KWDUJYptOg2IctEn+1Nxylyr
SReg8Y40oFH6uGWUFfy80sObBniK8GGfIpBHfTZOSMqusqQWMZo6awmo7dtcG4rJFQzVQ5GgLPen
iDCrckRwZk2EhLfyjnIIEi0s+lfAZw7BoBUSLuCeQM4C8vnMlkTv5qZEWrQhNTO5BLT1IYQ8H5jC
K+jcGAAgZCl5E3b1P9cgQXbHvRL4blv5NDP9sPmvRF3o6OBkqmvfXC5JJFqiwZRV0EIB6OKEWBjQ
vj2AdmHqVfLQudH0B5EafO/Nyg22utnjki5XXKew6IjFwTmDWu+zM4IXxJl+8azAMHKgHYYdFZPj
Jkg4wGR+OF2isJ5BvH6QhGb1E3Km70CcOPEP6YzjabILnUlS3Hc+zl/CJDhSY1X5g4kxI63V3OjJ
hVl8VyNA6yRwDn7Np3jCFZ6AWuqQyc6S4L0QJ/BJcDItsnXOkwp7Qj5Fok8o3tNySjnvr9OdZCvs
oh630ETY/UXen1a0D6d2w/c5IzxQJjB6ZYcaqKRJahEFVW9nioaFknPhdfVolgFOzccaMI4kFXPK
PxyToW2ist9NO3GEUMTYw0JMQvcQYbN/5h35OaUJVIbnHC6VrnNrj7xk9tg9Z2qdtAYzAxySacAx
nROZWlcdcaCVj2qE0FWmGcjHTMPTqeoOnteEwWOdZK7BGZ7IhbgX/c2mSQbxcSdVb+wLgAHJfdsb
rXLKM5Mew8Dzsscqy7liDAe5BGhuwxgNLtnXThsGS+MV1Ad8T3ZNK+kwCw8tErRaYIXVyRC0dElV
tDLTB+S/mrxYdKZ0wfGIF4NTrJwL6nhdibCi+RfStMgfRfCbSf2+EfRx8QVtDUqIACamLBYwIwdm
RdgxKUj1FJmMxal8o9rfhBxZs6Hk1oPanvCm6sFT/4Daj1OLnLyV296zbOE53XIb+stRbJwk6zbA
vxdaBEhGpnqGz0NBtDpZoKnWQ46EJazagTh3rAEZyoiC70VV/GN1F5KOlENCOzqmefBEybSoY8hc
rJN1KrCMDwzl/4QEYinkjYfYN9mQSr8cjTXme6NAYaHJI+smoa7EchWg6eBjuewJJcCgNJt1lDr4
vzsfFFnh/LOOZmmZuel5o5rLANZTnt31DrbGU4jcz3FOnUm85f3WI1vmKGKJNBDDHysUP0TDKqGx
Y4qsUaDErIu/0So/sVJZoO5fDmuofthFB/LMS/7cmNRWxGfH6XBUXjc/Bc4dXCKZgXsPr4K8/R85
B5iecSzNCwsWaGmrE0p6QQZ48FzQwn3Gq6LerxmsBXb6pAyxhKWyuarm2IphwqWcP+pxmBet8gci
HAiIWC5kX2ZVcUkHiGPpLJSQpGfwwo4qWZ1O7zpA/F8AmYTb31o7dRyCwGfQup6SDw2shRe5vwN6
oxwvtxEMs1vcrc/vfh+tiB+hynFwAdJUUGxJFrU3iGwxZYCZV85PE6AhT0RCw9QdpiA4AVEgoL2d
460Vm8awWTD59bxxYrOBjiBVfix6s+oAGIY2McFIYP8omU5KtCI112KA8vZDxAqaL+gANjqWIXRE
8ZcvwAk3h7UZDDiK9br6b9pXA4C4ES1v965eYQZvHHN+sEYNZqIljQkUPXS60+aKpD91sTYohjhs
HmT4VBcbFRzGGC7B4A+gCzyPnCdSayNcfKxWFIt7m2Nh9Rx+cdho6M6vFgvB0ntpcUAlRYWF8XHa
j/OSTrZMNwUUyFg733H8xt2GNsHKfnNPR7JbtmrKYkOR2KGaA4KnfOtiiOD5C8AzmCSMPUTXQoqd
Le4sSGhA3ckz6uRWOPlnXY/Bduy5uxxfv8cMrzocqax7avdrYhXkqbX/tFwW60IQ7221ArJLy9Gp
9E8ztT5f0fUWdLwNdxTwsmahDNQ5NgetGqqb+BzOqnfxzwMcBmjbtWiiXKX6wRACMSoy31d7xS7M
REgqAqYZTakBTSpjWJke/WU13P8EiQs3QrS2vmCpIbLVkr9VbmQkPGDStcxLNmqA91t/X5ePPc10
ZqCsdf900Xo13V/UJaGp7ZFxbCkr4+UoOnhICJiVtmQglg77rPDE5WBqHnWzidW4KbzYdbc90AF6
8RBBdQJudKhsPuHz9BWugI5ZxOVCEbY9P9kMS8VojBwpxJlHVagOn1yXmun5GtMhu7r50llhcAx4
JC5i1IUBSbHbqA8OQ676U+XZEBy5+I1BKxcA7jbDRPX/upwGAAPQqJArUBrZT2lB6M615V8Q1+lR
EXh0F8nXu3U1b5IswuyFvb+skKmmjeqCOzTHArM+u3Z/LwXR29GrDVGlCmBxPOSuX14MH4GlTrQd
//U2AQAmQbj8Pp7kehcT7i32rvJmz14mF3dra7lneAnIFjqrXhhQ8A26TfwadchlHIWOq0lhUueU
KVCdJxhF6KGX9MdWiqgZAxWHbF/C+KdXPMZcH5UgIVxAJCipj5y0dpdUTktv8y52lTchnO4VOQZg
QRNn8vVYDip+TNfraDys4DhC+OvX4yr6b9XW85p2QXF1wxdMIBWMHQYvBK4unEl2cluHj7CZmqHF
456zhV2XIHsQ55F/RXKJioXmt+DRMw9e63NNZZ4gBIkle2DBM363EBAUQdRuRD996hwccknqNF5x
vlPTm/4tLDE8jadnaxgHQhbBX797gzAyABWcq27fuS/OHhlp3ApDPBDGaopkRG+TgxCPVBvDb/FL
ftVCgdkoEq3EARlspxmRTQZjYqNnO2vHTMmQaU4nOfDQAH2N1fLCGtTR5JfiRw2iDvkngKge3JGW
sgZU8baVdvgCrH95q5ASUry+BFBC70oDHY7Y008V73NwzseJxn9yhL0GWKi9IOUT+YHy6Rg88CA1
Fx2aYjfa5rv92MeGhfGnljC/sENTm7tUYUXU9awZEqJV72wOy5mk5vlCd1Tk3K7dOuI1NkO82/uQ
VDUxRld2Psh/VfklY8Iaq5J/YUfkLGp+tBHDUCiDyhhbAZfZpUSa3PECLXjIU/RnRxAgAnGwONNR
KCs1+U6RDlTEBnBCtaZ1qSXfD4IyFMhmM43fD0ZLyXVtN8+RIL0BqBm5qmjD3mLkT6OLRghGy0Yr
OtNkkkK2HtA98eGxN/dHQfJDdNUsFzpLaDq+Uw0LkzZrluAuBzjf8sJeLIlMuNdOIYT+duc248Xq
GM0MiQjcA9ES2nI/qM3eBseFLp/sYfkD4zVQbAVeknSG2+Xxp6gD8+OlPrRs/QWSWTBJeZCAPX5h
ryDDm+CzqlMaymO1wc1y3qt/LG3GsDeyxod+j50Mwl1g1nTjggoPNAjt5gRKk7p8akAPdhYxirFr
J539zy1oSPGvmEd4IW+jHX3lQZjdz0VIfF7ft568iHCcUcAmsBpf8TYWtlP1sSMy+OE4LOVfWbbg
Ps3QmZXGnAe5nY2LXLx8iw5Aq5QJg8X5h3qIeH6RRT1QqfrjTWLxqBHHQzNjw59Er52XUH4+hg62
NLFhwukb6Qa6jT3u9WngpeBQnzrKQOJjcgJtUirYmCj5FhkraIVL8tuIEsNvXltyJz3I7rxczRO9
NKhh/nr31x+vfsoSb7cDmLLynRJG3QbC7/UdIFHri792hhY99r9FHK9LNBbTOkQun+Es0Q3PemE1
HzoqsMaZsWnrHPpgMt7roC7DY/Mpyo0qVK82bKUReWurNpEXuDSMI/yuqy0pTrTFvxpnnb+INFv6
H97jLHnUMiKfRCGVhoGWC9jsKBROsKrNNN1S/KOZ4u/w/GfgSfc/cOZXK2WyH9BHVAj4rSGggWEw
W+whwLwrj9jgWcCAJTNZGHMhI7CCSeVUvgkejV0NHHNGWS9s/vyYlUZ8U8ErGhY8onGsyp7EoPL5
g02kY582c59lAgREZcFdRntCraY2+uKw6d+EZCprp8QSOBkpbgqRWhPKsJmXMsiN7p7VTk/DHiLP
f2EMoNljxz3k1CveywzY8/rFDvxFtwZzzvRaFewgwfvRzCSNvuzJVa5rMFRVUDijonD6zWvrqj6/
qmJPH06BqGf39A5dyUeTuuvsncmBQouxjoeSnePnKGVTeQ1hJZ0HVu5C1UAdmZ8kiUzwRSYg0v2p
h1qYBJ0bXh4H9mH9iJlQlVMdIX2OJfEAU0CmN8xgYSAA1At1nwAHfMUIcf4chdGJtSZb3um7xPeH
RYIW8HeNTph7tkq0ZdQisoV7yuNVuvsz5Ys3IZhQ3WNdy4i/Vah/LMntMA2qY8bpDp55IGmJG2XR
T3r5tAQMzHGsV5M9SNXZdu0ebP4nJQepzVRYygyKV9OL1/+dxiEMB4Lm75121vShYZyL7UMBqIuO
TNUGo1KSP0xWFhd5DXKUj9A5Si2ITQqc01CIVtTmEyio1dq+iJZzZvmDO1M0v57SHEG0cu1K+I0w
0qI8UljvHyw+ffns+r0Mbbg21fIpqbUrphuy/7x8RaIh5dc+AwuP03MvuA/CH8omXj+iqKean9OX
NOwdrZavCmojPqkPhBMjnU/UNlVzqQzhsgnp44Ie40hABpfinr1Y85h2lCPFdbGXbf4dvAQgdiKG
x3ZXWe0XNTKN00I9U9mEK68j8RbbNF7tZDgy1CTgRj0IorgSIXS0mxvtxPGFGMt7mVsnnBrG3WA/
3BQqF3d2mbXectWwS+W/pUK7PaYTcM/E52DQIzLhMORiRQrbV9TpdNR0r1urmnoJVxA0kD/zaFt8
qJbBHeB6aRo7/nbCw9RgDRsHIWGrDOkY9l5ISRfPHbS5D1Oi8r+2lpEpQgdDmg7L7zyr67FI7UN2
StCxDmcqa3+9nwZMD4MHA+H4VnIe8Cg31bYebgWAiIL6qW4yU/Yt30e6BfVJZx6CdzPix5KhA1Th
/vo88iB1BsH4LAFzd36B1ioJGqy+DmOK3pu+hnRKe3IpVEMJjg3NAe2DEq49GjU4r2fzeL52soHn
aW8RfI6D4GbD7Qf3sfv9pb4xzHtK7ta8FBmwFnsZZv3NagJUO8HWdIXTTyAPeDED0KGwll/Wzd//
w1S7P3OMIS4LUdlFUOFNGadqIQ7duQN6MxK3o2jJalekmvlDoIjJ5N71SfVdzKfZhCXoWaMC2h1Y
lKup7kD3637jCOLoCkOWSB+yz9BknrhcoO5QX6ZX281rHndeAT6OQcu7ie/jb8TFs0sO/4mGwuZ/
qdhO2QigOqJJjPI7S54W+nNL3V3b0gIpyvTmZGOvyc1AAHlxcrga441VA8Nep7JN8ZL2SkrkiVzS
0Rmp9UwVaHqQmg/Sjj/EJw6EBejwdpqy+10oN7i4c86z33ImglxV0ziRLI6Gvs6Rwv0ExeqIH8uY
a3G/2DQUTGBjf4UGflLlROLVtMPUC/BLFVomw5jsIzBPJTr/Gy2FGC2WqOyhrW3vghVLEvDJ6ATG
aYhIyZENIm/7rXqbglw0CuT4dOfkeod/TmbS1w1bDF2gRN1wJB9EtfdIS1uONe9p4+VbD7ckkXJV
qKiy75LCs+GWuEg24BUTP25+BVNaAvpfw/e4S1MC+J/UjAHraHugxjVkoD9F/1tdcUK6ZAxhjWBz
eF+h7A9XOUF2XPHGclg3UeNhT20jlP8IStZdu0RpywngRuvf/BN42wxJb0yjY5qcVmB9UZYmXS4f
Il2AY0F9o1UFGzrde5Rsam1jc2uogAwvOLE46FqomZkOdyn6V2kx5lW/SYquDBUQDstg0c5jvtRz
ORT1/kzrTdWatGN5WgVzpRHncCsNzI5E8DRRop4L0jVypks2F4NA29qOTYYf/UYnBSgOQeR4ZIn1
mV1f2rmAnaYb5e9Av3Q3up8gbPFtq0E9cb+OGUaTZp+o4Zc/obMn677rWgp8e1wGeDqmk9IYDBWa
eZ9BEnoeejkPlwFjWfjqdkHBW2iPL0jkvevU7FZKCIUAP5zKu7zTa7zweTm6pFGb+6HZ2q5QD4wg
ZNuLQWENs2x+tICBMgueHN7jVJT0mYTh2Q0TTxNxYJsWsxzjz04qFUpkyOi9F1boalhdXU0cncSZ
xHvyD7xPJyiot8iCn6Siv2pdVxMzDy3jO/QKr7Bm2x4KfdmgVe6DvucPELJmN3zop1kwJ577esZ4
u7bJoBkqaoXNIMjx+M2eD0G0RH53nSqBRrELPkUBgGlb4YCH5rLfcRCR5Whf3Yl8Acvolqks8ROf
r9LXrr85VTc1+6uNgAG6v1HQIRZ9XGQZOS3DdKOyRe6hQi6gZg6pyk0vG1836cEPp4DkA4/sxd7A
JZ0+e2Y/X0CLNqyPN5QKaiRYSjhiT+yxf7BcRDqMA8GCmEse9BzlsJl78k0L0O9kdi2VYd39Y3IY
zUo7SLUe39vhc+9ktUxNFkA0TYl6wFkg9hfHL7GUQnGXUA0dU4xZ+S24TUbnJDlTz6herusagY9e
goUcBK4iGDykm04VTau20XBbvhYItmpS0tg8e7koIypHyLSaV5XqdLv5nTr457/3W2E0CNcYtmpT
0PoYPtJ/+Cm9ZfGFS1j8e+zyKtLHzqidEnBu8OVt2kflKK2If2JaGm+MIceIEBKvrGia+KX8ZwTj
cpp+B5opmMA1RF6tfHXNCXdJHLWJFNEo8Bbn/1W5jP8d3vf8sA4LhXD0yL0GYIFGfx73AEEfVyZR
5N1eP0ARE/h1TvUDjH8IXTQ6qW66fco+wQoZmih8M/uwnvSxb4wp9G1J3xzisjOBNolskKAJEMqq
N0xVCfDPZUeRbgDo2zYs7vcnQeChh4goWPs5hH0AAl0ftl4UtlVswXXkWkidN26hp3qYypeHqOAC
HSo45n2wf0fBZMgSauRnOd8KVMk42EzkvcukgI/HCiBHUnlCFOVT10ChTNQ9x3DVgzNFPXoihqX4
gixXGqs99qTnTOBO0Y5D54mY9mwNKiKudHZE2czASGEGQR7CUYq2mvszPlsztTiXnge6qnojmiSa
haprhkPL6mDQjpA49C5NTBYcG7q0SwcU2EyIPa/52i1B6jr8jRKGGnBO7pIbmNJLb/JLEPEhxNjh
8dWhDFiZUSACEIxV8mTKf/a5xrl78r9BB9gXddz71gDso5RoCmdhzEl3DsBx/+wTsxUpYcs95kZq
kDeGm73vJtJwmtnzT5THsopsMMi8O+hjXpJxNlKYh4CWf+E4LmoZVKzrFb0zN2z+CPiy86vzmn6b
sx7S6QcaTX6R4w0HjSmxzNoQFsENmlt/021Ohb4Jd4GFI4UUKgqV0tmd9lmgyXJiqf95upE6GqCG
HsxFzpvMw+3ZlsgTfi7VISVoqB1VD6GtPX11MAXrDPzsrIWZAGZ1H8mErpQ0AO+K9mDulSaENbot
dL/TLpcI3I0ggyTXB8EF1Da9h0MStjg6SCVGdC7teK1t4LGZhmnriEjgfJ6gaOyim9+QZgpDz2KO
xb1tD9t8aKqWAGUA1WF+LB5uSQEQ2GVaRPnpjDSblSAAuxRdkvvO72SGp9Y1uP1qG95UKiQOcd3A
lea9YLgcD1KjVVXLfNOAzpEZ624kZpFKWpD8T/s2+Ydg3sxXvPuqxxGM6WgeXq24YnygOyV9s7RS
tbSpXEBe6h8hvnTeim3BJpXegQqzPd+ybMNqs75kxAenZ9d76ax6YDtholg4dPDym/aFdHGWqtdM
qmt7AwtxZzHeEy4FmG0581ntnSoDKNU/V9kv41IG6VziCiJhYFN+BZdWCPaCfuA3XAiiq/Z8lOEd
Tz2c3lhEtqwI2UQWJ39391ZpDrrzTDVaI052dnyJr7yCVvM1E+OwsgcXLlrzwRFfyu+zLnaIBdrg
CVGil8Kg27WGxX8EeyhQnXfBRgnypwTag0orLX12hHI8yJMnfa+aQMOHbidiQZIl/kl15F3qjRpe
9DQ+nffnE3BFzMPAjS8n/cUAf0CLWsDMNtsl5YTEb/H54z87RjjFAvmTS5hcy98GsRXw0wBhRJh9
+ywYuwFogIYuNwOT8DA65yC7IVo4EajSgxIz75CGdbnm4bSWcIk9vv1tlPX5lFzfVW1ixLrjGrqb
DDWXesWcp6RN3Da8l2KbTZqMV6Wjnya65HOQTmynGIs/3Rcfa5nM/R7QDht7f8g85KJng/0e6Rcy
0PqHb7Cwi/unLB5L8tlBkmOpW3a3PGPhxTFSK2W3xfRluxoVRTt2wlo2jst0Zb7Xrcr3nyPY6ZcC
suFOpNOR0AeH30kRxUN4dng/HlmD1MlC2K0lSAqARWxuu8gErliA91zbeaUMtdC2iAx/JX2yT1U4
AgqonPgS5Godka/JfCHZpeHUB61ATsQFu3RZ4kwmjj766aXDRoRj18mObeGQ2EppDCFmJdUeFPmd
kMvDfXYwTR4aFpDronmCOPt44v8/MeY2xfFSk6iXt+PyRy4wyVqg5OmZWfT+vsTjt8EcvwJUc7nZ
Vz/xGX1c/cFvw7O0TUDSY75XvAe8RCDEwQzTwNO9fR/cW2pWJRFzGoywRhMo5r49Wb3HZ8152FV6
+6b6kBIzMzBsbaLJf8fxghIacQTtd1tOlGajA4WQALHMtfbMYCw3qZaDE6oSPrj678fs5vS6viwL
vV4AltkXJ4jLpU7zTaUesf6tW4fke/iOqMJCBpPIV92ZupnAhxGZwHbG+UP1mHt2urE/NKo42zRt
Kvx7YJbhwerDXIIeZkxoyYQOmi77FmBnobvJlhyzECuCIpA+SAbYq3UE7G8NQQreEf+tY1l7zsG5
RWLv5QfCPwhPTyv703M52TzShSuJfoixenv5iSSZXaHCg7nMX28GMYIncJexyrvav7bX8dv/Y7VO
BiihSr7706fzLG2ailKacpZL/yKr9TRfzW+5rQN/lu922WTa6fs0hUYWvnpsMKdXgRyWg91SqcWW
nRMYWLwH+7g5SngqieucJi62Gn9Y1PDLlzUf+8HL5sMwM+yeCCvxQX4m/EFbmcl+nQQDxx5/AM4g
o2EWroyBomxVkbQbL09I49NgQmic5FUv0vi2G+rWjurz/wrZKIHk8JmeZOnPrudtVeszKGX7Hpbd
7epMLkl96OkVa51pgChJG0z5Fed3P9KvhkBBC2sbnKQgh2wXXx54oXctu+LHDCbaPx+PF0iU0EE7
90vU59KVGv/oiM/+/gSPsKoiAA2UKlnYhJsCMA0UMzMsED6o8q6cq/7nrGwQSvC6eJTQXa9KQvv9
vssokW8ZZn0hB4/ENM6qlOnovArGJhc0/AkbQWr0uVZB3oTsHlUtcEiVq24ppTOaAjTyqFuWMmBd
dvKfBkau4CTTCs4UJwf+yoC/o73W0gSTJmJfteJ7GKzxEwGW7JHD8H36FoBqDi34AO0sPxUuUo8L
Tow8KCi1P8LbWf6uwb5TZXwsDHzYgniKaZ8d+ouR4B8Xdb9a1y/E+wc84mFCNymJsAPbDBb2mNpG
gh2KmEVco2ofeOQfbhlXgCNTkUilkFD/lD/qp0I7ejhqbOxxEo38cgcrFgKVPUtWlJS8bpeI6G9C
vKhAFUc47XGKqL7j+8ekmyKQH4gD0gxhpAQTntYc2Ybp+ogwJV6Q2t6YCBxIPVt4NJevHFGdWOh3
GgpwNhSQfxzAa/ZHH8OKBc3hyWnhWJLt+bbapdTHf51U6SMsynITSVU/LuP/jHvZS/QzhsbycoEa
5I++PvVWlu0Xg3Hnz15LI808EWn1chzN6JReSIMp7P6gNVFcKs45z3+RGG068FO0krjL8K0HSBUd
YezqKqS1YIb+dbFkTzzg7PoFtvxJmqyC3LJHFrhw5b+Gp7GsagbHO8GUy1927CRWc7nBVwpnaNkx
9StfGVc+Oex/E1MDHGNMWQ0bP12AHJM6gppGLZzsqyS51GUqeC1Ty5sbFRIoui0SWqFCEvUQZg8J
6MyWgcDLjEuPEe1F918YOtOQfoAYlwMpptQkDKU5QX8cmtGd35Mi/MDm7PBMcovZPrDBuVvV+MC7
Lvaqu5vQ0KFtDPtReezUvJdoW7x+BNL8wKrNtq/xwj+gPXf7VzprYHrjzZAvHHeGh7Zj2Iu+uIMZ
HPOYTaamU0fKnVWJkR8Lwteg59QRXioTctizASCKkdGW1GVc19X6TKS14JpcIUmoDjy2bJUNBJju
3MZYCTc1hSrJj6H6HqgR6EsqeTHq1udZ9bHquHu50SEVCoOdda2EvfzoYFKWi0GyZyiitzH/EQH4
e4x64nkufg/bWSTccZ8di0pr75cHRTw76HPnn9+LwoGmg48mFaPh0Myrn6wXaOlCVF9Ep/DZv6b5
JTfyeEhLaS4o6L/q7J04QlT/tts3ameavsycpVqHB7fGbacAuxRE132GYCq7esdTrFfZYpZ71t5c
Lp06chInd6rFhNmV9PacCMaYcFvsjIQbVxVDdCwpm+ueYt/MXHiJRZVwN52Hq+Ng4v86rqE+jMNB
j1eEnbPDFFqne8Jz0VxRwknXXqBFkQuxLHoQGFyGjW4VR04IrcWWGNNGRnzCyAdfG319AiSCQx5o
d9Nqo/3o/u5uZrLJvuDWEMYuimy6IVOJh+9E2GdUBO8N8BXOhgKKI7xyUmisAWSUI7Aprqnc+aAk
9ETj5Nie8r7cnabEGJCAZPmDwMNQLghodQ3eUUi7gfkLiXKVJ0VEfgmIq3y1l7/MejWnQHN7APuv
TKLex5A7ae//17HiWRAsre9NMBY5CjvtuJUgGc4LlQBjZNTXEpTUkzviqedOlPrxXkomZ5D1V4Ek
au/xM9jNDuHH4ZBOcaPpnEctyNwgMqT0OxbYyyzIF0s3YZ887GRh13aiI6aQAROpJrYLK+igFCLi
HG2ge5bVc/soegY5pVFjRjA8HFTjDDdAUfwHLRp7QQR/OFVAluctAFtk4072saE6myoRjAQO82s1
oCRgMNwmywClnKA3lgVQmotbguE3HL0SDl94GVmwsQuH+g3nD2mLtCzFfFjIzFS17HSDioRNB8AQ
cTgsgfESROL5Vg8DXUfLT9coO/mjqj4YiVSQCPoQ5vG+T5Of8LiNIhgRF+N6c47FuTpxIn0do7dg
L5ohdCj/mE2TfCiqHYNGYhVVv0TgpmHm+MdlvcnnMUNRFcssmGhdNY0Ffnl1a7+ram1CysGosF4r
IUmcoqkpBpDzlnMDn2ubXB5ANxLeXbRmSut+z6CC+0W/WJpgvwMe+fzq8xX0FqOMjAqMVJutCfEk
0m0xU9gVWO5SglKzMd1UDSYN2jQF2tOh4Xw8wafMJ+AlMfueoLZWYc7OJsWw6udODtNcKrkyWNG0
DGygdC8XQhHsonVSYnirYjv68z5dKZje1Ex1JBXFR2w/3clx4ntl8tdOkCHKIrRWHfQeWImaUi00
LUIqYJ2VVL98fGAbAg61PKZWMOLoQ2j4w1aIQeUCQr0zl71HQiGG9f66FaLA+qz7QECOiu4d9xFv
QSBQuYD2J+lu9erUHLDKfy5zJlQ8KmJdgV7jvf5WA5Vh/CIfUhs6rIMoB4/XzmglXJi591QWWC3Z
HbQzbK1z2P0QfzaRxO5zibjcBdnCl11u6hUMJM8wRc5TZc6bDcMziZH0qH2GwuRgIUF6GWrXQDeh
Up6v4wzJ+YoxVvJL/0NBWAIykZEdDmVlYNFIXKkBWjv5fjZPoAHFQTqR0MB9xOP5NVjmhVI+Jqyw
cravJalxgcTbxvS//0uADpk6C6FJbTWyIhg7KFIiJ2OzPIgTigdgr/t6bluapd+c+8sPuiQYfSqI
CynHky1AfADzyBmjGq16pDKo87h1lQ/araLheIr2FtjNPAMtXRTcrO+X7GiRO6/GCieIxGoxssm0
H1zOwNrl254bMIp2BDOiDgyeiTdL4SQPfDDMyDBzK2L/4vv+2ZeuCP01hTR5MWAHCJWotffjpJ+O
QW5tmDbq7gsOsPvkFZfO3J8zIvfy8Z36Nd2RLX5dzJouqGWgouD9V6WNdMCJVjk7LD7OJ7Gku2XG
w4CC6+SXCcHplyuL4jG16kHCFIJY80yqQSNuvdtkpoZ3ShwoBNxMw3XhuoOWU3a4YZo1juLg9mS2
PyCdgHK9UsTnO/pDoPji5nwg0gga1rvJfDtVIs5syYiRRFV91KY80j3iF7JK+5+8X0Kn5KYOR6QN
7wVxqu+ts+jJ6+Wb2QMM4/qrBD3FMXk8wWBnC9d0ZeQBv0++3l4VkNurnGA8yBjFl2YiYkBLOZKa
qs0ppNoZwvcaWi/GvbdOWsPzYKb2/0s4QJGiuOIZaUcxn0OPfmYfGOlqYSb1n/JdjzymI6fJZDnD
Jf2NNUx40P5kZZZRMR5MDWkWhqtPJU+VbYfXwub09r5+dOkUjmQYYHcZa1k/RYsnshf2Sx0VhBSY
2t6go2zBLPZTBQj8jcM7IohUyMOFHU8Nz2ngDGlTox3//CcC4lqmlRj8e1RsDbLfrM1FP31vWVvr
diw0ohRbOB7JXXUPSINqPnmEF/SXRMxMEU/NWdvO+LoA/4sOehEwfao445IbyuLDEpOBwvzHZEHX
UUKL12JWW0iTH9OZjDou5N3G6S1/Os1pW4YKrL4tMa7PSpGOzh63odn+b1E69HRZ6cb/41+qWnCi
23b0MGJSkMWDjRbL5DavROCoOB1VmlOsPUadnEUyArBQz0vR80USv5pPltip5qWJaKa0lMKsREWe
5bS3HvYuDGwa+Y1nXzyUVci/z9vgct54NbMH+NWfylWP++W+YWy5ZnX6QDR/AWsKhJ4p3q9ygPMk
dFAJiST+Pndm4kj6wghpZdxDx/x/WxLw8YpL4c90CObfnkSS3ahH/nB3jtPSXDGWzS1+TTed/ODJ
p7uLFUpjCKMzsh4IaPsx0WaclFRDiW/EpJWjyPC0pNzweFJQLSCJC6rdWDOJ//iwXI7M+M3BlVHw
SrvPP5f69OsZz1Mcpa2N0rNOtx4Qoi0CilNMfeu6nzna4k6FZscFO/CdiewER6KpSRtXkxqMgKrM
TT8fprmlDMyYiuGe8DiGT+lvr7ANz9sOO3R1neaApiZ1yyAvYoJfX1UU+hh5XlSZqVJUX5AViKhM
S/xJVqpuVZ2qnj442dROr7DiyUNwmtrVTUs9By5KJciQlqs2RCYjU2IYk6uMTiiht5quw9l7OVMH
W1Sbsd9mtHkGOGwfkxSFZhgYDkytoyh0bLtJf4sFskGI8pH9zsycuDw7VtxAhke1LZz5POk5DP4Z
nqbysHZJ7YujspTxE+3lXo2gycyw0sgMWoauFtP4RLSuPZONTrptge+i+CNpQetv7pQ1yYhJnihI
UNw4K4pMve8KBQNJ2mdOgdKQxS+PjfwyFKVV/Umyto8gh0w7h3mj4luhIDY4GwCxuAJpdoAJRkbt
eyKdijVc/vENr0bfpT38h6CYBYcAVqTKr+BUGOnEi3AU/nUADm0oNtqvw7O2XkdgYxi2bgv/GE2z
+UPidKndrRV5tbfrH1jFwQNqt/xMZ4Is3vehPpNQhYhj7dN7ReGhtrpMq4X3NctfBX4SxArMfKFZ
P7bRLNtBYTVn0APpCWND1GPoAyBcjTBm9MHyIOhZLCl1opyTyu4QxcsXK1YMDaErtemYybpolyEp
fgbbLQ62oRpFGwHVSXvxCVyfFYYZJJQOnhKfsN8vlhTrblyyUF6VQWlNxZ9jn5JWdr+Hjw85I93E
CYyUUhHly28goGrJ0CrHylRKD4qtsmA3kS8/u9pdOoUuLIZFdITHNDRvUULhS/UO+LjBxlg72gQF
x7IuRhDlSDyMSYZHA4NVqnwaA7yy+wlG2XMgL6qR4QTTVmRkPte9kXKyPtMuvwnNAJTrA81qVwez
knqpQcY0UeGo48J3WRpSv3BAKPKv+3ltfLdGElOOM2A2K0iIIHL5hCatL5fGg26Lw55FnTzatFBP
3+60yf8FU68z1A8LUjTc15E1AtjTfWrsDOBFgj1PoYEpMys0UJ8sqBSmocgI8dTPxxlbdFzGy8wM
K0/m6cqjuFtmbPV8uRZ7JtxDKXM5UN5lJ/i6rcDFMyY/3y54oqqiNupXZoaGKsjnJQTLzGLpvcR9
fi1VbR4gg8NeyFYpd0aGCJmEJicIWuI0H+S+sPBqbDKTw5Ok3bobd3Mp/McNUYq7v46vrbg8qxuL
QbbPfmZkvNtr1pkh+qFLnFjIsMmHtPf+nydP3Oc+g+jTGpwfEvEquo0IJmFvNnEwIT86Ln+wfFWK
gfQg1asoAQcoBCANd4CDSv2cfdlsDlnntOonmQuv41TpisoXCVt6jsq5lsHNXnnCKIrpn8vyQE6S
+/Uu963KAD7ccxg8tiAHiw8yW841bhQIaThTbJt+4wbWUaoWZvQzBVicrHzmIAIbvG20AMWe5VcD
kImndrUngj3+6CgtRRmtpYXRLTsSs3O5DvTocrFLcW+l8BsGIKbFAGuH8f6pj9W/j2Vl8cXVivPD
eXdjEeZOzxOI0zcH4PxO7DwT0/1aCKP63acYIiEvhfwWd48kUhJ8Q4ERGslHbcJpqc0ymcZvwxUF
To8CAbYIDwaiQ+5wmJY5NmPp+1TyMpTj+apnzbNnBQ1LieBEFMsmxrOXpromnr+LyKUr6UDh+s+e
q5w3Ky0L9jJSDu35h0Kxr02T0ooq/RmIIluAt5KmavXsEAxzLkoZDk3oEVHEM0KDNhmhf0X1TpO1
jYf87fZKIn0sQCcUHIvbneAH/z0DVGdMOq0v5e20yJLdic9dhzhTRCAMnxwUplygkcAsd5todt7I
HHTh03Q8bW2EnN50nk6gAJ935R/Sqbmqsf/SVLWxSPbjZqwvVHz1XIA/lWqvF8AkLolpM7Ld1GKQ
9a5m2ERirPw2KVNuPCHJS6gd1Jf+X8A44p8aqt5iIbiv7vNNUGhjFiXUgN6QV+EpmGNbgFnzRnj0
KsuUZWBOe0chSvdoU2BQFR9TT4gNENf3C4ENHPzA+7XWX7RaKCbkxhJ5FQ5EmGOy9OVMmhOIxe2Q
Li8/Mi0nsfup4sbYzAluAEb8V+yeqmwZ10HVIsC28DjepwH49DWuD+tRMWkvoPBpcip38lsyV+Ui
V4kqHgCidaAWlRGTo2IVtH3w+QenqmLJwIdIMI4ljzVnXb1XnWFpHcCydLzbsM2VXA1DyY38tIZa
8RG9ZoI9YuKO+Z4nCO360apDS6BgZyLdHz5fJIzVFGiOZx+hrbA4RgAARW6Nv6kLNxbsd7piDgdp
KmD0V7HTZtVSg1jVkh8L3FeOsx9Pogrq5rY1xxTVl4Cf0MOZer/ZVAcsA5wSaV4HYogqNk3u3yF0
FyrcwCDkpZRcfYpnWEGZ1SjQql+fiXv33w6qIWBAKr59adFZqSSYtklW9OyGINQQfIshAqBjWOUg
UxQATDLE0PksdC2Z0+PQMtaBIP7GOy4X5CPwyX9GKXK55NKCC2hkU56POEjWlk1U4qZtrdVWcirl
A93r0gv0TI5toHTyr2rKcA8QsTL7K/33dWnbI4pN9ydMwabJuvEZuKA8UVuFed2Ym3SMeiNCJqzS
rwiaExLmjBNtxrws2WifGqgV46yxL8dHPEWjJW1uAQMKM1wh8KUZ80YL2ECAg+08Gngu+qKRtAmO
l2UabkSVozqRUrUVANyTiaLfGH7CW3E+sOhCq/7laPnHOMAwUF4ODFJQd0Q+8XL9PBjUq5kVSxxD
zkj6Qwc4iXJNkBhTrvIQ3z+gkcZR11iZHimo5ltHSc58H9yVjNVcHPwjRdkgdBk/SS1MAny+LiW7
oEOHVbuYQHa2MymHjP4tyPxiIHca5/wpztKfLbgpL8MKj+VMFHBycV9uT6qE6txlIIpBhvjC6CV4
vkoUHD7CPf0u4NvsAi8lN2mc9QGd7lr4uwSwya9D+7fXzZ5WOugETOMC4BA18S2VDg9ggIGvBhJX
sqd3+BKcqHl7A3ZIpE47/Pc1I/6902KSj9eZ5g1hqQohs0KkmgWSf4O2euZ2CD07ALCIMYGSeter
oePXVhL26jc0/rUSALoFWVXMkvAwYNGefukBSJr2JXMHd8Fqx5SSltoRPC+jbkyUiqKFbOxpA5y2
TycrLVTo/Uqa4fFIo6NIdxFAVs2lAp9NCPLesz7SsreCrMKHyQ82SJ5OqUeBQ3RkgUIp1Ddd5auo
6aiRU5xvpjOIKDF6lidaKNQaN+e+uhaUcoesmTaUEdKVQCxshMG1TDmsLRSDib6fmgo6rpqRpmKR
mWi3/KNtt0WPeoC/caRQd6RVZNo9XVrxvCkiN59aRO1w3rAjGpynaz+PfMVQLMt+wF1+Oocb+pnh
3vw50IdvJ48SpftX/KL936SB32fPQ5s4webDOReS9PccqWlKStU7cVt+Y0hpK1DLhhZPmRBD5RQI
mfy4cBhIgMqgnEbgXUfJRGbTiKWt9Y44gpsy3LcICDcV173aC6x5qZ+0oPgO8oULEIl2hsIs5EJT
rt5Cfwai8OwpdTZTzZ83OLjffUTyehTUYpQOa5ldHnm4mufQhzUKqUKOpHHyIOkZM7NmuNHM1EJA
dplWFv4Vzw4+/Hp4jHJemF3Irbkw+d84P9VzSkLnZHyc+Nb6US7irO8fDb0huKFserJrRDSq2SjB
VCAllE0vLDZ/kU4kvkt8gyLjvBA+p8EQIo7fA7Ar6SXI4bSzZbL8vkrlMuUTVKwKPjfqGKQ8sTg3
avmZ/F5HmULbM86s2Rlkmkc1ereLIoN1pxSHqxyTDg6jvVsa5TfvLoOAlMkL91fB+T4zw12LyBcG
8Fa9oRsfrrpomPo0Y+yhsivx208wJwHixyX+BNHOz4yaeGQCAGhPKxM0D0CqtMmUNnicGgZHYhOV
t8QOTIBYieI/xRJzvlgSuJOW/i4ZDKBI42G3UYWBwz9Q0QUXHaKafYB3dNY2MvJ1cczjSxHhGXo3
hPxhdAWCjCfI3zRzbSMNYNgkT4U4iGuXaaZevqvx8/Yw4TpbyzbkEy252WaN7q42YjjTXVY04/Pw
sijJbR5i/BgooqNknxzktdSsZdnW2kU8ZCDBHPCAOReDmwOBiX2wfQGsgfvZBPyH9PeOJ9olQMvO
0xfyBdb0i4ko6bOfM5JbJ3+NJYH2gjhosbqNHN6MDbHSpvQRl9APpbBYXskZNard8JQKx8MsXZ8e
9/tKkEg0cnejNnaP5K/4cIAIt3kmJHhUKfQMO0GQYs0C68uEb0KAqYGmmRRji335sP56VXC2mluG
DYy2fLlUvfjkFlLZdYqBC+HWd/eb1YqVeVMONeiOP8WekzYlj6y46JlU4N3Ftcc5xWKqkod0ehqj
uSRetpfzz51MXC7R1dwd3dR9gguV7ZSli7cqqc/PJVJIRYPk3SztPwoUozmeNFK9XIDIpSdrsBlP
2uL8f56VDxweu9fEbl2MXfvPNDKOwj/fcD2g7OX+vD7hI3QVhleOE4lfEab1HB9nl4D3ynlCKNPS
E4SqcUpGp7Z2QwSUvCfI0EV+AnJ+VlBDK7VDJU6t8FOjjipPvYN2jVv5rx0ZpNV6wyYhOGc4guK1
T5ioil862Up21h+l9yJrgnp/HcDTGR9ZUEAvRB0j0qsv4OFw0/5pwS34AqnDWv/GpJ1dvX6uxl/J
CINEdPGdINbSE7R9KfHil8fSGpZF1h9XWN8oSD2LjLt5fy68tXm+ZmOswQ9XqPUFThdE5o/pFZjC
MpFjptd4uxmIcHrVhlb8xI1nXGTHgPTgVHLZoX4KtG9bdLNkuaWBDu46JS0rr6sOtKRAO0Ijmqm6
F2xpglDnIUbCoTuP8zZsfdAVxfBvpN0PwKuUE8rUDa19OsO7TlBRzX/+4pmuCD85qMSG7b4v8ZD8
+blEUAuH+1zoEVSHS6r3FvfeDX9dOVSBlauxf6nwq9i2lqQzRKsaArunNnb3ArgrOUL4Juz6UW1y
ZdxchccCy7U7TYqJgz2J+pUn3GMCo1Qt2xIAKc54npfWBsESdJTOe565kUQg+FNJFGQlRjHZUze6
CmVZfJ32IZb9mRRJNzf80giC/xrE4CatBlhKpfZ39mf3iDAszbdrUUcmOML3cjfUoCl77C3FZs2z
k8uB7Sjmq8eBN7+nPXZi7gAxXeoG7ApwBRm7cjQFRD5s9a8avfvigcV+H37+oQhSa/hkna1eRA+6
dDO1KXR96kQ62vdwNHzNHh3jlkTGrAFX96bRvveefFHkv8MDfjnAgmoEau/uWg9CYS9qhqgJbtvL
ojI1ni9o5tuLAKiD1c2Zm3FOiMDpNE2yKIClYp92mMS8Wet/bx/OsULJpg0LwjH/MxJK/ckfb6b4
oEEChGCpb/4rnN215onuGtdsylnpmSaGPcJ8M+WJ2Pet7bDSkLZWWyeUBsUbbW4c19uW7q5j4CAY
/KJjEd8596TeeLGGa49OSm+v1rS439owkrskPB+YH8hrnz1Wa3aibrT12VrbJ0upWFoy/hCu2a3x
YIxVRHbOr0JKMWy/zRt0HubZHG5abnBxvr45N4Iap2QOlRSlBdLpcLfkba5AfSay6jQliTWj5N6s
SU/0i3skfT1y77sCSrHSoxQQ1uxyOs7/+ab1rcuOHBcrEtnRYLys/u4FkNMXXs1obL9tNhl6K3fq
6pgf6z7TuTfl5gZ+ZTRlonBBbcX+jmxur1qALMUDNG1XgRZ5KUhOd1Vcl/g8hzPeKNCWiVm5Faj1
43wTu6SA0FeB3mfYc7P96Jy5BpT9uD0nssLgXOAidGZn9NVXaMLm3Bh6qu7guYsR/SQxxJ3rA4Mn
wGRTqeMMHoc9dj2IRcqdNmPn83VvPfypnn9IKQ+5AbTt5UbibFHt3XXd7Zo/t4pn/LCctPjFzCGF
PWJdqV83xZn4mKWcmUqpo/EmzotNdrDtexLPLbYjnd1tYtIsENirhURKTfrdTjyIys4iv1WldBWF
HBuEWVSIQrFY9t9CASyHQKPejSc22rDN+HaXdmqo7zpWdRtXGLqzaaqzxBQ51tvXqCA7Ztuj8h3E
DCkemtPHGqpBzH4wmS/Y5xWFg64z1iPWyW9uCU9WcBMvfz3bXx5BJvcLtYwraUjR2E7lHxTgy6aR
m2A+ZdxC6xhp6dcnwTepic0ABVavPumWoz9V3hgcApwFp70U93m9aa/Jjgoz03Vla+QUas8mHIHT
4DhVGKk8jyQ31w/lk/bppyL8heLIQP6cGk269+Rc28p9AJa4+fFpaW8PkkhT1BN1RhrmnkhB/FFh
1vx2qUgYvcoGRtKS7wL4BAsJexuV8N3q27SyX4o0YIP0vCLVuRoaSLZGYQZUkW0jMjuf57f23aoG
7ITUfldmEMjqSuFEMtYbk+VRbCFrIHEJQ3A5MscdX1UqzVuNKpe94tdIDBKgu04r7KErSllDcZxK
e6CQjiMfj3nXcxw+CSrwCJt1TwPXl6bYUk+D4lHgpbn6H9VFmFe2d6JDKjQlLczWDwAZ2PzoN2BC
G+o701HQtlkekK5qLOsI6tS7pPiHWWkdCO4mCptFq4ALta4VTO94vmEAoS28fLh0p4O7YMdhvR0J
zS7yoC+3/jMPeZ6fOG/8ON87fKs5FOIPjT6KJugEan8MrmP0nWnf6jskqbbL6XakFLLT3tSsdjaB
1gzDu4o1/APwyvaenVCKdfjrwLZ+fVy22pc1sLMtI0Iid7+QcRUGXMySugRHndi8rrFJFfWlEZpZ
my6Q39+MYd+Dy+XVwEEf7So7832wpfKcHsEZYEH71+k/Ldr93imxNqgZIZMOQT+wi3dDVnth693m
C1cGb0NLfkkbP2HIfIoGT9ATfPv8Ly3LqooCBWPnJ0XglhqxIZ6IgHae/XDi7jXQ/3g+wCYWBxJA
zKdRlxMogeFOb1I0xg2D57UDf0/8fU6suXT83L//ZFepMQEH6WLFEerjaldhP3AJyCUdOIhNP7Kr
47HR2LH6YEURnMioUF1wWXEozYqQk/v4t74OejM90H4V5ms+DfKook79EvmUUdcKYi2Np5Oybt/c
aoYL0S/7+RaBh0ukPNP+LvIf0cXVBqu3qUDlXgs22CffaIVLHpvHnjhSPFroIdj3bEnL3R3dm51h
nKKXfgV4ab8bQkZ40lDJbOJ1WdikDNG+3eMFDMhyior8mProP3SaWIO6pL8W7qepITd5Di4mbCi+
xfFWS/SuDrDsTq7DqN6Ey+GAfnm75ZS4LBw6D1NwTV/ql3XgQtD5i7cQtlNW2dZwTNJbbiEljTgV
TxOffYc5K3jCykwmF6U5u3NljlxwwWS7aRQfee4KvCDarU0p28AsgiHeyLLBKIw5nMaPISIXRhmF
Dc3D3unqN9N9QZ0bL+bQYIbMLtW5KXaE3+u67/2c+GzEtaoE32nZiOqDicXkySJwBOigbKf/SJxx
QqqVF8i/pSCBaQEhJCPq24YrMySCplST5lAq8c0V7pvrTs7tOZqXCORc1bIY2Ucpqml80W54aoJv
v7DJiAqRSPCdm+GJQrniYNGASxI1Li5ZjkqQttMUHDCBgnBCosQFbyGdnylO1T8jfxlZ+izBxm7U
gYF8Mn4mmSACgWJ8KWEW/6GhG5w3eh3LtwfhTfJ3a3S67gPAhnxTYxY4x6fyMvLXy25rmKXig1r0
yk+/QTSMqJL0fe95yXzg/oWkRdZq8ap+MWpOSzYRPtU3i64LGBtbmzkuLM/RR1NqAs/yYAA/KMPC
5db7bKu+MhwkILO3DUT1N3WRzwHT2eu2piHdCWfKd8HN/X87b8mPiObw+odgelazGcKCilq/nfUk
WWrEnVAx2Yva+DfHUu5a8Ykt6Ao4mjosANIdKPE20ySkinjuLo3ZXTBeFFli9fM7dVA9iF/t2BlQ
UU/fL0PF95QhC4MQsgmfcA+NuYC8qIrDA8g2fLcoAUp9ieFhRIoZWWaIM2nWmPcA72X+xXWWu1qy
aUYBGjz8ePpNWYCS20ORvHk7SVerydI1fli8k18T4X6sg+MJdfsvvn3PTBnY15GNJ797gc5yeYjH
Z1DzV09wrbK89grY0hiHXfHPceYJF6f+ddXvfsvnqMR3Kw4WeFf20THGP8nXOnFbgrETIBxyvzDV
1W78iqME5lJJR2yLFM1P/uKcfEknbe04++JhvPhW+zCUA2RRJvSsEWkOqeshd5c+axDimJnZTOdj
dAlfijztWKRv7kWPhAZpu/fBohxy/Zr0Dv3bmZ+1mAW5ElA8Xc0SgT5HxY7tCqNgWgIwgcZ9it+w
2d7eFiVZkmtFTj6LABGd1LYIhT19BroijvDjHhWePSRvMSwFwgCwgpmuoY2PA5kbT5E9vL2nElNr
K3aG0f5M6Qp8fnnXwghEHoSKC4u7ZZoKvmu0PvOY1woEj9Y5X8HvV8orKJlBAJiIDIWHMxaEDvOv
jbrnqv3HSPwp3+8StrBIVTq/gOm6TJCrlrANLVCYH9MlviHZwF2WUhQ7vPiHwr7LgE/7YGjdavb2
d/E5Wkicu4RJgiZpgfcrw9RWoIgUCMx2fObmqzXYkbv4SysAM3ARSU61tLOddOOnc1ehbpohM5MC
/Lga4ozMofkrmZYOaHeeWy8bf5a4nSpiqsLYJ8i0SR0p/q3B8nBLpDz512SYlZSf4FE0Loos+cuN
+hXnT+wouHcCvS9o3vRSCylSHoomOBRO6RBk/wq10Kqt8kjn/1c0RyUs9OQrUaFUuClDYHllr9/N
xzYLMyD4J7j9pIbNIazgPKqzun1ZQ7l4xQA2ELGvVLIniJDaXgYLYSiJ+N1nUZivyzkq0s0/NVVI
Nq9/f1RUlMe6lO/7XC8InKemXqM/+GAUzB57oPvce+W3kPD3omC4pSpaDDXf8TSmLFKq26USqeUl
l2fKhUTfLr7TAHAth92DHEtlL21dJUornhZc8DmnkOyzfpNeHyY4eZugBFp0fjQNZIs0IBqZtngC
68rQ3ihJmqIS7FLtRnB+TFgOB4kFQbwhcqytB29E5lqtg6MnQNyZCwhnIeldjULLrLw5WgLpNDvR
bZoOOvzIMA5EHj3YHX/jK4pw2GonRiutnxszbzZaNVIqgT8Q6JSpSTBRI/0vP67pvN9xC4iWM5l3
AJAxpz/oobzB9UnWBjbUOxKwnYg3N2Fe0+jGfg/ZED5gcHDkoeinpKyREXEg3fJHAYqUR8fvJU8d
8WyF4mLCgy/lzw7H7xj1N9pgYGkvfBe4nzohpBYJOmDJZO4+Y/Io7q5nfyK+AARd9fEw0+a+uGHD
cjgNh/+nS1vqQfrEMwVVQDbDLAO6mBdRvx7vMpGsAaehJAAjPEcbGClIi0D443KfmoCMVP32l4uH
eqjTHn8u7Sc6bmtj7M9nl1Df+CQS/AdNOG4iAaNEPSGlordYDAlrnQyz4d3MZSeOgUfLuoDb8+nN
aQ/pIljBWrx+5C4n7YPRE24FWODfSIn8Fx5/DV6NEhEzp8cyM6IJttMmBWA5IsegksjSP58FCH/k
d8hU4Xe3L25eCHE0GToGUxKtLYgHDkn59HuuON+YZyThr9yzRWoRlLGXu34Zw84QzYcoLhY82VXu
wMp3kTRyVmcPkUgalFRfTeQhMh/Xqx5Yzq91bPAaSSx2CosoNliXyCH6IeFNdn7SVsatAXaxWkeZ
Y36LH+qzYbL4/TbQuBsdo9wsgGKS8locFpQBm2hpDoUf8wpz0GFa6x6zuJtp4CXXIv7v5PWFQXSg
t5FCTJ/l+OUkyQvUvAMZX7FjBpFO9lUS8PWWrIh2wnSM34TFKagKSpACM2c0TZx4ATpoKtqgvcvs
6kaTOmlEK+RsuHqvnv936aLj+GFBGGAPP76V999DJqGhbVFLZxTUfmgvX9QJy5rhG/Y/S9xWUCzo
3bpR5h+tSx2xeM0eEdtBWdC/X2UbLG0du/aTAkE50LqztOnyvQh0WkldqjpCYBsDj2F1j4aUbvLm
NL43XxvuVZqWBYRrRpvW1DwxN8/zqS7dIL89WyRGtGpUovkqAWP7CeI/cyf4VnpnhGdSnGiGimOL
cI4pM7PabPlIpz1NBD4gaK01ZV/ZPrZJH9m4EsbV3szJ7OoA4fEcm7clWBR8i5GhpOPL5re+Qxev
5Pp/k5NzKZdWkw/WVDFm1X3uohjHhM/xCRfVw+UnL7Mi5SIwo2AidKCdzvad97ZG9+sejk+d0o/s
WPMQJ7plgBas+fLv5egFXy5GQTfvdn8qeuNWjfGQ5B4ObAiINA/octvPOiaDp3cVvy9d9tlzHIcI
KwGQhwiRZZyI+8zGX3Q+UNu6NqqlkFyamRQiGBp0c5J7x9WDILMA/SWjhuqS5DgrulnagHkIKrew
4x2qZLTm3gj2D/e/nnJE5fHCbCRPdFVnFn4Kw6Hq7nLaCtKkwH7BGjORt87+s+Wa4hV/pu7I5Fn2
vSvSnm6CedjPOderaPA+ReUHqgvu4d5M4wmyasmUdu0LiDQ1w7R8tmrqsUDSWsCzRjBQP9Wo3kGs
y5qY3KmG9zP6f9GA3zFK2YarnQ1kLkmiV6z+M7xi0Vn+y7KKPvpIS8BqYTGp4XjuUSo+WLgqB7Gq
HJRF1ew7nBPB3QOla/L1aHxlpzxI3vXMgT556bfCKOUNmbGAkI1tAyYi1SdXV8Oyxm9r1IDox9tN
i82uiEqA3IKfNQkN1KWdlXzCcV3O/bkdVnG7WIVGM87b7Gueq8aceGHAh6Zswr/EAsraRd/qAvqQ
W5CwXMfjYK4YUiKVe0/Mi2OvABS6UdYMs9MY9POlXV274B/sRJrSpa1zz9da7imQkdoPWI1QDzlM
Kr51WtEx6X0I4L2TQm7mLzFpJDtpPBg5WbTdf8IK6KB2D48xIPo+F0OvCKYxHut0oBSFzOig6GTd
ByoWzXRGqxK5O6NNDMy7MJDLwXmjcHv9Sr5ArLuThYzVXZJ2JCyh5NEKLxtFTDnQ7K6eNBTU4XMJ
MAIOzjWmad2qKbQO23nDflUSTcoKQLPIROalFVf2L1zNvkuqRwstUcltAfKsn3i0J6DswyX/pWW3
tAW/rxL57CDebU/0mPo/oGow7XFxDX8ntahewISLYiR5+Fx8V/0Rlj7KCdMYbE+zopr1+nqnvSGX
UrsMuYmvfzZT7pmSt2DSf6vJBv03YlUYRRONETWQCbfPIYp9uwK/16Tb9itkrfHgm3oQ+Yn1H7Ei
p1tUNoQ2OaW95zpGvy1LdLk+rLTa+w0TEqnWKDNaoPpTk5C2lILJgcvNhTt847tSzL6oxUMoUvgi
Y8DzFi5Gd8KtI7A908L9mYdpxpB7Bg8+/P1MCCOwbLPF2yVeSqNyGieUCAYnKwMtuvBdLUBUzBBo
85smbHZRcEeMPAXugLRiJPJi4DLvUB/0oTRJRDzT6GgtW0D+7Yl6sH4om/EjUe1fJUOzB1Cb+F0H
Oxtkv4jFOATV+bPDYLztG1OXne74yVDgldxFtwhErbFyVuaP/pARWR5nSEbb5wT/+YFt7JXO+mbu
7QzZSAjdvvNuF8KStTMyqvVMLAbQ+z8cUvAMq4S5h75mRLHh/2eyUSonxl9TLgygFl/q8eUkGGng
MuysJ0n9KRb2s26k9bxGOSGnZO0chb8KUQRy2IA5AEAAqF87Ez92JLmu/YBzrzkswb/NqbO9UVYt
9iam4KCWz+n9l0hWdD1zaHf6CPgVdh8lNdklPE18Zo0en2ko4111R3YKgavQzerTk+A0yHr6L/KV
stBYZsXSTbrNaoajBp+1ZxBKBqz9jsF+xXJjJ2S8SwWr3T2bFI5zBy2dQc5pPtd36pz1hNjlHU0g
TrRkr7Us57lbDyQ2XOa7KYduFOcUYxZhg2dO2eLFp8ZGzXyeNnE3NDQhp3MHysCy4ZNbGuJRAJW6
V41DzPx9xIB+bnnpGaCig7G+U4AHio7PqZ/KOXbWNx0ljnuvxVRS274fmeWIMKCxhGaPpf86hczG
Rm+kO1dt7NcY6Bdm/caci5kfWlW21UjdLoWfzDQl1lJZt4j8aLnJXAj3pvpAeuwi03idtrr6MqQv
mw4v2nzTBveuK4/T10BNVpm4+W3QUyg6aGEjvnLcuNusicJhII6a81cfl2g4Dr6IxqxEdQrNTrPi
hrSa0NLbImNp0NJCMF2JVz76UfpCl7rqs5MUaAiUUOMxkSfeVmvYh6u6bi8aMZjMlssff5DmLG8h
nEW80ors4M/NnXGqsLSMMkdyd+kYEKnn8LF3dthY5CBzosScf6SWyJB7WGzagqosHkYsxg4VXj1Z
uQ/fdPC2OxKqEeRPrnvd2VcQuAndROx6Dj9E0iSQVVOAjA5S9wGznOjOnnKUZEvdJUN+hl4dlIaf
ETann/L4FdclW0COlEHWDPWGZf0eXou0Gymkdbq5WyusKdZ0QdQFbfD4B4aebNh2CV3L6Bi/d3xL
Cd//FNlHzDohz4QfynD3lX0W0XGju8gnk+tJzZahtoDyOIfFj21AVS8ya7S8oR5UoQLxx+6P4OwU
Ba65MMCm5j4/I3FwMteIRj7cB3a77LO/ZxYVQr7EGxGNtgCNkt0SOrC3jghjxjUGUCYrgEynxCyU
BJpDsxzTG1xTBIUW0wlKXM04OlbNWAAWD4THaeAuWR5cvgb0KnV6pKDz9eemc60B2am7fXusHczT
dq9gxANNnrWGwo7DXObKz1W+rFj1lBgIPP2Fw+gkiYU8W5UL9yraUjUnVc3Krk+f9VmaoC8Fj0bx
ZwBfRJgv1ne0Kaj9Z7ROOnI/RWil+eqz4/F0fgRSbc8bMgb8P/Z+iigskmplb/zcTXy+1crSKpNz
esazx74vr9HN4Lx6z4+I5FTQ7UwON9M848wzW7iByyVaj4WmEcvxFOxOtqO3KNcnm3bvJyM2qIM2
3wmJ5hTIOU4SlTJ4yEXUjI0uG/kyGNh6dfB5WBcFGGPiNqJ+hubtFmzjcAIM/YWs6ZGmFgY4euNT
lenFNL0yzfUDpNEiyZm4vK3B0PyWA0S3h+jMGfd/GMYpJk+25PC0K/kj/6Hk3MugRB0KQSiAifA1
hQHq2wGV/+hbw/cVoe3tC+hIzjqmQvpX1YqpsGKK5Aebguatq7TXV3x1bBvwJDevWqmBsDNGlCkT
h4RbfRvpbOMSIK979Et1LQBoORWvLnI6g4ouIW5YVm74QB1PWaF/QdYKQtFsvz5Bc4WQ2XHGH0G0
J4SOdyr13FKZ9RHMSTSVXlRBxJbu9+QDdW8v8vWWCj3kC4C6UnjSagIE49cxqqMbm8Tu/hIUTNV7
q5I292NhaPMd+7HHhDwTlZ1k3duFHdk8tZ1TwO/30xFtCnVKslH4F5sQwagqx8L+enFBw22iMeVL
eiDlehM/OR6+bdwXvWbKYWhnkSaGLJSIpGYRrzpa2LDLGwrxFvkkgUDKg8Xt2Ia4AlIJiPa8l45Z
ZiAEL2x1gy9Apz6Tu1ftZaqPXfVgp1T5NDrxeXvmnUT1UcOGGY+NQYe0Auj6oyJqrzy5JlP1iY/e
wYySewcIBIdYOOL0nXjG8D/3bHi1WmyrSjBE+7YpZdEjVck6MjNf7gfNxKr39fTjU3hvh0CoYFBg
/kDiW6wQPGCpD9bzAvsz7EqG7fNlkz/FuENFnkGjIhyT7IoK2HWKTDe9rM75wCpoE4tsmg/SHGqs
DaZ8ov94nyHzanNiATQnYxJqrunlAuYfVbGD9zf/S4zVPpJBDu8zrGF8UgbpotQar7SzC/05+jAj
EEwI1zyAzCwcjC1CztcsAnF4X1XYAUv8PCrXCEXaPyc8+lsxuzy3QLs81h+TSiPqVWrByjmtPW64
POAMq9qdTkv+u0D2Unph6M22n4UrabEdSXxMGLnmXVu4QAUyTeyFDzKkGcO6AhzCpMBSqIOKGpt1
NeMGHe6q2VYDiXs178GOrKh4tB4K6pV/o+MDwbB35cwuwiM6JaZFyrr9uz2rC4OMQci4882cP4zo
YT1m0dPObaVQdX99G81ES6uwMZ7jx/LaBBow694y0cFavjTi30UH0TgomaueIzpBcBzFZL9YaDPw
+RNwZEfHgm7aF0MYOkTVCzPi0zyCLdC9ikhUcANTyAe+3cwP1fHylAmsBdyYnnP5oVUcmrXN5GFz
2KAdhNP/2Qm14UhVY+WZ8iyWGkYfn9h3aA2m/mSeNnl4R0nFq8fke/8hBgL4YKDktZr/MJv/AeR6
2iaxdj9Sil1LrP2hI5Ycgn6nSY8XCR0O1u3IxcvEzFXfiLFle0Ls5Ao1j+N4sylHJREkKqXXqtga
Tbgeq3roinmRUtLyBXuw1EHDSMeEuJdzjjYapTXae7O1u0VTHD5u6hciWEqEaREfQVOokWbK2GKV
qf4LxKVHqnLc33ro8AQaC5RzTDReihXbvCOZEmiWSHUzDMV0emrniSRV1Pvgm9AdMP2oZfNQLdY3
wOJGzea9WHkinKjbamQpCKxFKTZvVdslZ2ji8zZKxQzkJxUjkUI7YPxuj/iXL0bD460UVd08ilqW
ibZyyyUirEajr+PqEzQShoIQEDZvDJzRoa3xRkrjWE+tD7oT5XIgL1wg7fXOBa/QyA8J4yhM5+Cb
ykTfHErl3zV4xLmE+u9/0VkGuX/Awa3WK4Uq7aejKjxEFpScn6MxOEggbiJk1RMyw1Y9lecnb9cw
T0hlHVbNYZivVY0Tn1OgUNLbL6biA4+sNx1Yu6q88aJxb4uPa2omKbgRPSk7pkHarapSVKktPmzK
BIPHyM25gVD0+XsiK9WHP7XkG9MMikTdw1TtHIn9QaHCIxBQFRRGhDH6Ixa4dh99MOsapR9CNCv4
80lJLVdTuP3x7yrK7Dxw/6jOFd6LDA4GGzSdhP3iMDcdrYdh/36EcZBaKCL2Qg7k7MX3y0ptoozg
dzyKM+ESbxdRTIbCvXeSx8GDUrHAOtyx0PqZzDWJDFvOYZmcj2UtQtz9vWVJMP//NQMUo1B/zrD8
cHwki3/sehSkari+5Y+BrLP11eJj2sJcRyfr4F5vEv9qT4ZAq/+V/7lzZAWWN0TzGVA5aDmDq1Tu
9ESGf9B5q2WK5Hri3n3CEcmxtWeHfkP/9THo6PxsgmodLDcVtjlYCj0AhIcBkdFVB4idfe853uoV
sUpz11sBlYwOP4NXq1qUyY5BqNhEzLVmSKqwlDxtwqNAZoK2abYbDfOcYNC4Pd8Zc5wexasi0cP9
4ICF8cpHRbEGdG9tmMSWGz5DP0uBA0h/jcynwjNgBVgmiFbRgpb/zx0LSjZWrhtfOafgRdldSLN7
lDWZC7ffFiauBU++uQ4WVJjfPvaWp99jg7rMNv+GVzXtIZSQa2/V+EYGyikj68/vU7y10Nmvl2jN
F0p/GRONsgMduDZTXw3hMLA5sZhTOHnuHUiFUc1nd8x0Q+OqBRc0wmxSGWQ6k/nETpEyhbHJK75t
z6KudARvcnQ0x2zHh/oZR9Meh2s5bQLzUwQwxFhagKIeEY1clTPiIvQdOeTc8gfNu/XdRRI4D4wv
9vKiq44zCYPcKqEKx5dvvxdA3UTIIZGH90jpfPZXttIqA86DVfIHh4gCYU2Cjawjce5GUpaaMRP4
Is4q23Y5Hne9urH5WH3f+L00ZN1NWR9JVQ5lckD2PWEjiq1KKnkOPpAwQBF51qIEpEgk84z69S2N
BL73h4E9vdrghdzsMCS1xXbxXy19EOCkdMym6pSTS4TeKXWT/U+6pgqZx2ivbyzbljNxappsXJDI
P8/U4dKU/i5pupRmUguIXqLUdo9hzf0AQ2es5tlpn3lZ8DMYGEUvzm8fnfUPnFJEb6/unh/ek9GW
AU/UDbJL6YucBkfml/FthX8T4vMvw2JGdKreHqlPWKyPe0lyDUn6JGms3zOSTER1WmWc69b/qmeS
TxyzIf711+GraduxacAjBKppnfbrtknoUBZ4bG2Ja3LLFbpA3GwVN1laRKe9Lt03NV8EGGfagxk/
c1z//jn1vcGtcIf5Eg85nFlpL2BSqkrSElssohhkLLOjGuI9Ypvlo5Pcd2yItQnEsytjGuHlfbUr
Mp1bJnrJCGX/g0femB+s5cMwbmiWuHm5bFpmbtUuDmdFm4/+ZgbSgK+18OZDUEPXT2SL16PNJjz2
BRN759mguhCtkRl5BCwLaLt826NUU93chB+NHpY6/mCMeUr2SG4T826DqLaY6ukvSlreGch9DzP2
8ErVfBoFw83Ei38Y6O7IBILpKHmzo5FprDDV1w/rplpluCESrkCKsNrr6IoN6Y/39D/L38/AKeVf
ujDS3CHfqBbVs+84DaBL+0r/KYzTXYxArD12O88CJQUlXsPsr3mY/ELwV/E/YazyEs9MWn0moo+Y
emDrAvR2r5RsHl6yC8AC8VJdX701w1FDDOlLxbw1NAdkMFN5v/yMtX5NmLTVnIqKpDdmt7HeLOBv
zafgTmjxn2fZym3Bx6kdwKVBRPvS+ofh62qN7WsE8Euh8eg5ndxgOaZMkAkjEykJD5FOVNCtx8Uj
cxgD0FOdUKN+LMFiSw3q91GecYSpS/FKh/+uA3JLp9FMcDUsmsSTGtvO814XLNPOQCK7a34JZ3a3
v3rxUEt3dNNFsZrH5a1R3mbixTDRCfqfunEy2vUqkLdjC9tEimdnS8or3o39QgKAdbMszGeSVA5F
85cqB1vDivDSRRNZBufhSboPckRsNTtFg/XRdzEejY0zkTIEtq5NP9+rCZ1/dzntbCVmeIvW5NPT
KBgaP/m2ZQM9ItkYagTqfmuSTKTJbJV7A3AovFt+I8ekQcWdBIFi1K5cwrYg3NTRnLFM+gPs+1m6
DcUfPcllQK8ftARmBgjjKBNdkd42TRvi9kxWHG3aY9lTDM/L7w2tIe2FuIPE/oQxLCBTH2MYOG2h
GD/e16SgYxnZoMUlon67m9XvuI8KWu70mzKc552h2WrlKk95yukZbf+gw4XnYYudkIApxRYSb0ge
9vGfMST0BVlxusFSDtfZe0WstmSclpVCINqnJNSxHZdfh95+Msu0Y2erlvvSOP0MmrpLzWW8A5rD
is1lZ5254hJM/yRy/TzEujCfAiolITdqSpF1rybhgtTeywCmu72dEkhBujitwjszFvvaTQXQkni9
bSkOhbh/PChV0H7AyV2/lN3QlKw7Px7yqYXUfhX187KO8/DkCMtw16Mx7oXqRcjyOYWh8KnuFoU+
fd/V8sM10w5H0D6cgapM6oZY0uYe7VajVzUJhen/tHyjvba8fuqNqVdqOF4DUFJ8RRj0GAf561ES
g1EJlNF7aXKiiBFyhan37EkxE4PDe3pFVKOitT/0K4snwsF16jSjvTkxubRUehGcCbgWgoD1xz6D
I0PYBjryF4EETwJ2IaE37B0qW8C5g1ToE1ibv1dzDewX8kN3nWbMIi9gQy/1Td2qVVH5rsqeTS0t
BtubOLrFUcgh+jRhGY7Q8Tu9jRXDWoSMYqcXdbhR6D419DD99PVrHJxf48SLEPrecRNyCBV1Q2VD
uIW1M37x2CTsy+R+9jfSpNWNiwgh3OcwxH+H+DJ85bH9LkFaf2PPEoH5HkHLI4pWaHZ2Dg2FSRKj
megkaeZpKE6GPBk/MxXsijehl0vVdLfjGhpXQ/Ugg6uYRTn6YS856yoMA9CdnkvikyEEm8XywIXl
s+fR+8uDNPyQn2bV/C5sRS+k64O5jIo94xTul3qOFO5sdGgqZu6aejlKnkHqmLKhJIuBd0R1LVgp
w6l4B+H9TCO8jX5Pankstnkvf8Pn/n7h+2xBM5Hjs9sbrc8x2msAjQOYW6Ao24XUEmJV+F2OOuWh
RTJlOBsCtKeojJ9rlXDVo2YnD411JreagvaBNazFcqz0OuEsS7z3P2UgmFsiX+eZXCs7kgM3FQW+
Jlgj4ljeUDThTvWq9gIMs1lqBaHoenJIosyH9APtMLyTD7cakd0paULY7E7nobA5WY6mItsB3yrH
23WU7jxq74VJbmUvX14kjS1p6OEW58ovoU1RYAati2eUl+hSiDscSVJzjLBowY/0ozODJMPTj8Js
n/2eHtvk6/TeEAr85Og4fbddS6iECwQZsyubPn1GxdGkT7SrkZpnFR/HMNYV4wKie2uw1uwvBgFQ
gNFocv4Fc2ssI6JfikvsYq51k1JFo995IF6obYBwwmiBBviFt65AReFVyXEtITYn/L9DPEBUx8QQ
Tpfk7exvRCwGcJ9/T0/0nGSp6abGmn95eXB35NDAeUqxEDJlbBZ8tceOmcRmOIa3wbn5bu8OdUxe
4gTR2oAsZysmYI8D3jurynoO6/Uto9PD8KqMmVd73RKd3WXp/5k9ZuVE9tt6lc8hDjzSjem4MlAz
vPQRqJff8Et5wHFwuBgvKi67yJZ8Vozl9QhQ7oWgVIsNSCqQTfsLfUg1n6K/0gI8hxUKlexuYY3z
/rzsAJBAvi91D6V7+SSkpy7q96oMDW+FBwVM9Y2may+HUGbX9cBW9FJnlNUepj+Dh575zvC3VXBG
udDLH4xjzEjwkha0T0GspsB2YTYbAYgRQDaoYY6NggVbMdoINLlfsgBVQB+iAxFbt14MRGbGwpgu
mY0VIStdrpnIqKeABHsuOI9SnkhFLetXutjha48LKCt0bxZfSH2MORX8DCw8YOT+BYuOsTRvvSWe
EVsehkRxpEqp8xzfz1/iCBBRvUcWOwfUuoFTPU9Eny+IjeecaHMOauR7GCvVwf5cYTEnXkIsWUu1
LYUG6L+OijoKpArn5KPNtsEnxU6Ch5J/7yY637BcUgCsbwKb9L34BuRiKaBo7su8bHDEP95TnjRf
SNASgUmL8jSHX6lFO+lPJpus+WBBJ+TB6h6kPxMm+eg6y5eaEthQSL1iuTJLDqCmzM3XmE/4rZlV
D0JqEUyNyaa+1wa7+uv6+O+0/mM6G7Y9AbJ+6bxHCmF5qX3kbnLR4iyAD923ZYy5I8HUCd4n+7xr
yXfuAuKviAg6HUtfagTLK3hpcr3gQ+ZpO6f82lVtZLMIl6HX+FfWc9WUOFSrSQH0rSC0xdEQy10d
OPtgxCmCq0eKQwgSgeD+l9t+WBS4P4oM2A9UoX8MagQojK8Gbdjw8pDGsOPLrbBodJvya+5LS0CP
pWl6+g4o+fqqq5TVu5D39PtA3HSDlZrhPK7YVOK2BOUJhLcxrmV7gLjRQGnOzHfhuKHYdqBdxM6t
eP8vebgvo49NSLTWwGjqq8+AgNiHAdQOumCL7aqbN5KlCyZ9xcVWU+/fF4L9Xi2zp5HTALt/bPzD
AMJsF9ytEvdO1A5QYV3NCN5VNIsfO20qhPXmYSHcOm3LQkqt0ZOKoTueOKumHG7UOHalNlCJSOIp
Bi36FdyqxW2ULZ/BFphODFKrhB2EeSrLI/cxWnNrujvswfGSmI31OR/9nrzxS8KVmbTIiRb5kSHk
lWfvD011PVNzTGMvSBnQKYF2MBJBfi20SjZCSCgH/Lk3oWK3RujIc9tRB02RZ/3FOyIdm1FSnnTD
WELOBKcVvwFIJoMV+HfwCQfW6+2BEUSASh+Pwf9opjJEp/a3hkLUlL+aJTEg4kCMnJKl4IOtPICO
bRTbu+wUdzvj004h3zDtGNsmRtHoAwk3BryaGyqFOICqLymR8UJW9coa7E0Dtk9TeA59t2jmfChW
53B3PAz/NvChMm3KhouRUrEqV0rUFj5wDvCqxWJbhBx+oCJP6mddbhEdAU0KeZFx3bbD11KDu2vK
7sv09yUYczfxkRdh9TpuHahqLKduRJv/5EWpIzxAd3WRh9cM1BUgHUQTYVTDk/843Uq4gXb0SeBM
7O1em6w8X1/i0MtSIPzBSLcolpg0PynpiLFDJ424YnPICr0MwLIqcjxHu5Qbzpj/ebtraZB8Xgyq
kGBBMx0N6ywLCs+kw0KeK1YUGoP3BJomWO5eZXZ0634NQQy+vphVu3SoayPHGDpnbMdxfSAUPInG
Vguw+69hxNFdDMh5TSV+1MGapeMwXuQT1R/WcsyFcPYE3ibaqhse9QRoFEGKj4ueOCI0y0rDj8KG
8slh29B7obvZ3Kkignk5Doq2sxrvz4h2qtBeDP4syQfrejNCBjeMp8eLPHhTVaoSLufvPwllSUth
PGialm7zl2RIjwXsyZMHNcH8WBtCV5b5EqTp8CgAoRfAiorNlp9ew9rb3XW3evPkEMN+CGM1mPPN
lwLVaM2rwqVe0UQTmqiTZTc5BpI/2L6wZ1gkI/DpT6KkOpg+P86mY5TG24J4ofHzzbD43EjDTQ8E
lMSzTJJLNElDmBAPJpG8JOnBg8g3tMQBHkJcaa0t/j24P7ElyOnqtTm4EbYmzeIczGrH5YdgRxEv
sQCfjhOuMO+fKBE602Z+Dghq7sl5CmssiR8sKRF9AuZPC3ZHhrFKBlkrprqZRoSc6Vh4g1hfKuzU
RpSEPgMn8SpW7SkmhFpU5ZhKqRuvpmbTngs0z3N+0gqI7/AtRn4DojIs6+GERrPCikEXRFBOeKOR
C86jlO+z90MJHtY22sfMDBgygV0qmyvfooZALC3EHMH45jV4q/gPXMABqM1TTjOjKCVGMNYjMp1Y
V03UBFPzq4GzlZHDNXj5G79F3VEMvwlMBBNAAYkv/CAIH+haOaxwH8ntFAzffMC285JGXxXCLG6G
Ohr5UJXV9LR/qluIKYsGK8IFM2EWbQ8MSeHHBhmt0IeWPK24+9/EuH9JxSuwPMDqrRGTba+wPOup
RM9TdVi6IneIAg7dH8WFPEFybGgtOrr/TvKmcRtyLMNrgaXykGgED6+wqQjROpc3RT/xO2qPM4YM
/CnA+suZ7gg+3rjiCpWqDvxeEG2sGp9Q/vzOmf51QZktM4mDehlFc1ZqEjywRs8l4RA9UrKbzv1s
fLPC4a7IwqYYOhg21nBZ0SkttV1oDunSaxzrL/EKa4WQr7bN1xlaOXK55ACKLQu5yfiRq14SoUXa
HUkifNs1W3teyKV6poXbBbcA76Cwryjsd522pWT7mey1xHz9YtdEXizYEPK1k91Fd4QP8myDBUJM
WQ134wnHxnT3htnORv0hog69RzGkhSWGHxbPIvIW6Ezy0tKSdicyNcWlZSg+jsJvBr/DNn5veNEL
UiAXiGbphKExSd6D2nvRDzSFUkBkdyWNcEfnGppCgucjtLbPTLuKaD6BoMpHVZ1EtO/Z9YfQtEk0
dzSzqPvub/BwbT7Rzzr5AHSFsyRNWoj/E9wrkWiEqRX6AerdIcEryTeu9IN8KRK22p4ShjcT9Kz7
esMp9KP2V6T7WRa0a4IZ2zR5YJYMmU3MOtXyrJR1VC00BIrH1MaGTGcskNP82Zp6BwVk8dfy6/GT
jG7VyRzlZ5Tz+CI1jIXswymBKPiXWLHlK0qAyMGFWVofYzNp9i06ZAmgPaxrifX1QZPdNi0gi65v
tOYkMubFMq4lrkKd6PQzGSgYGSKDLGIGulbuV6nNsJllvEeZ/9O2L92cRVpdfKzxJ/UJVQNXBC07
pejQu2lrvnb15mtcIzDtUg62/RWaRjVsgGTr3becbi5rC68Q8QauEJDVXg45/vG/U+HItDh//h5e
O3Vn+1zDgvupUUiUha4Rb6IOQeqygNP0y/Fg0OkOVw3O372Z6o2Cwa0+HIzWKI12qFlhb4d9Nn1e
FUD+Uh4DAaX8B6dQW3H3YngIX43TctbpgvIYmCznwP5PhXt4gCa4TrbUrnjisg9Y/YQ16A6HYcPp
jUXIpd69x2jKy+l9UZBFehP67Q1LcK+603YuiqDT4F9nG+QFZ/SAzoAXlWk97f0GBlgKQkvJ/ddI
uxNEOmQZyoQz3dHD1i424Hpo1RdWjRmeQrIVLEhJMD3efs1pEswBDokLevf+rZLpiOR9g8V5VQFo
MllrvnbAfE9x2kBJAV4aFY3SsjSNSBXtnBt+H2zUyWxLXhrum84TLUJNpCAoYRlKRvG+Yoy9Llmo
lZ8lUZ9ZLFC06xBk6001JzFGCRUXV6W5iWNv7TRlOerzgaTVmmMU6Dt2bbOjNcvbS5GxNhJCujOF
RNOB7Mad8CLdnPUgBZdlnWB/yu/1qIZecDHmo7N+uuTebBHpz7qT9AM6vyFicY1oHBDmW6PIPe/A
plXRL4CA4sGx8IDUDPgYaeTjAm7AbgPDPnxeIdTm9VP8eQwA+i77vsV0KkXFP+R0CR9WCS8Ac2vg
qnV4HD6UKAM/F5TQnWMzdX/o5NQ0bJB9qFiijxz5mmcjjgVohUX4BC8xQn/U12XOCS9CzWt9Ljsh
e7OUDinUPbDy90oDIe+611/Fxy1Lu0QIhxO6z/eelnpXUlqw0Esa0AQjI4XaeOw8F5SAihoWiIQZ
5LhoXhVq8zZy2Yii3Xjwl7sW8LnsyVtWwJGG0EgpCwVqE1qF4UPAL4ffgenUf/BclYyAKptV9+xA
lfbQb8hszE7O+pexLrfvMwpPgv4vAFyNxlzBAVnlxbioaXsTFFjWKuVoDrZCxTMHUzbFxqeX6qdU
+IwFzT+XVYX/wRrb3jwH4RvMQ8lMY9pb7k4dP5zbrUyjNLu7MSE258LDIi9Ip3lpsMoa2QNeEB1M
f5mAhGZT4hHdSJAkEboxz/7+5rAmxCtGtfhC6QuJX2ZhRQwpOyt081D+bI3sXI4DZuWzf7WMClv0
kSjct6ZGosJb+cQ1Y/brw9ZOfwo8ed5s87d6jMptgpthdb+Cr5gAdzIg+L1CByXvoL0QRQd6vAVo
qj0GxDiijoQnSztpf6/O7uJEtbdT4AblhESbwfToO6S7gmuscNXmEsme5NAcoN3GCOOWtb7dUlOM
5fqRZGD1gjxLeFy/DqDP1x/fIN8cyL6PjRyrU/CRJS4rT6UfkpNlEosxQHgW7OHdb8SE/1vSBISN
rMtJSQJZ1rR2Nybb0Xt650iHqYFNUfBLA1LpgOaWiQp3udSXly8UqSFIr4W9D/Dym33XUPRzzK+6
OLcQxmaD9AmyMxnwx45XQVBcm+uxeXmREIDqDqA3tuG/c6ZXyIZv57pVA6J6LGQAa2c5GuGHZpMo
XTslefUP/wKox8MO24YY7P/C031RPJaMCMeQU+87uoD8J5/USUw0e4QQwS9bAeowJltY0OpoyEcu
WjztORUzErFOgfwh1YP0EQ0YjUGbzIcH5EJZ83XyIOPgcgahRa7h0MTTd3bDRygX1saL7NEHnZBT
8aAINdTTi3cJbokqCqB+ofUS9wmnarg16kwthuieO/apBriuJA7AuYW2xybQ89SO0IYB4yXCMaYs
B82NQiDzR8VoLgYKBARD9oN+5o/vaJa8OEz6fV1vjHptl0pSiRV/3T/NYSiKocMxcYMVHBAj5NR2
1Y0lB66oeCyAjV12VqKaspLn+54ij1bTV0gFiToFH2nqfhdvBDx36vCjEeIuBZcmiaU49O0eNdgl
BFWtBTwSIDlr4YUmk08tIdiBkH1hhH4SuIPbS3hUAYekTAn6EH3WDzuBbqYLVrZcUJS8gahEpn9r
73SHfcsWUEJWkuF6r1MeSDPma0N3BPn6UhjblE0lZ3189ZfJLvH/rSZSXgYhJ/DNassFk/tOhmiG
fPiv4z5MKvhrt4o6Pme8/c4E46GYIs6BE1bFE1pzycJfB7njHkwfVkQ/parlpLQ39aZsoqGg0XIr
AcetjO0867rYdUgGSVM3hQdku04y/NjPwjUaimm9MY4zUtC4npYeVsnoxAGrwsXJEwLYZR6KIVrN
K2hmBlVTmyJe9pHUACHIuJdVPueyXkgDekG+6zqnGNqf/a6BGg1gl1tRKpslyIzdzaG9Bnncpax3
y23V8LYXD8ZU2e+P2+YEyQhqMRkTYPoRYJVAkV948utkLlP+0/1zXkwvOscYbVW2mCxnt2ansHq7
g8/Ll3zF3n8BTn+FShLjeOiIbMVfcnVvWHwWTc4zJ+rl8GS9XhQWIAhaZCrmVMH8w9fZSUfoD+ho
9ZIRINYrbOHAj62/VyYGnXlJuH5Wc0sSj9L1Lo8CObdbuIBQz0BFtGK94/I/djKoWSUCpBfaBZS/
ZqFuBGbUTjakiJ5h6RbD9tULxGEL15+/RnnIoGlCFlwl4kjIQKi5bvc6hpbHv7XWsuTtt6rswBrU
wFcHw/PwXNsCfEx6ObpBW9sCnMoeXS9aQs9sF1/Q/i87h7N5VTmLQpdF2b45M7jy0oP2TiZI7uCC
9bqRPlD99IJ2wgvT/BR5RWgNg+h93ug9CwQ+zsaWkmB8w/Tdk1Qmb1pxreuesmxCVjoNRybJuLhA
XmnMT8KNVudXPo1rXigp+14u8xbBAslmAfLx7vYNZuOO7hcgDcna/o5eXjlbn2Zg5Z3026HmX9P/
SIa3gXf1FXStgu+o8flhM0wC6F7QUSexQkXXvER+WFN9U3yrJ/IuIvoN+13qsvnZkDoQ7TV5euSu
P9a2pUHTVbSnJJwhRIMQ64+ejMFga3G3htu+jS2ReyzqAFqiFJJH9L2cb4ttZVpkWQ7oXcadQJuC
jQdfUUWuuAMM2YZqeASYi6zZh0BWZcqwQf9W0y2FF7msCsnMz8kl7w8hXIyu4FShXBGsM0woHXMp
O3lC+7jA5fqqvZ8hkH/nj/QJnkSqECoyTZChtiF2IYaaap7/x1TXeeEvwNPZM/SUi3RHupkMopp2
ccH6qDR38u2NWzJesty6iyN3xo3yanQdAzpT/lrAnzHQtjEXF4AS0HR0msEm03Brfe8tiWnpzQHh
bUPyR4Z1vJFcOjDV3p+vjWZrbMH51HMKYfla3s/klXlUFoNxpKB54MvJiFa+mxueq9gWRp1+1L/Q
GvTGki7Gs2/tNxpfDuE5lQZtqYERrnRa3ytBCZFGULGr/5H3WBGq1cUuWeJFIqrYQtKobvMcqiDm
yHn2vrJiCFT6TZQeL38wMKiX7EnaKYE/bdRCjlNfjSBQ0uyvFJuFjQBevb2UZ1WgAjN4fY9zo2n4
h1Q33XMAQSebgqktxm5OhgXdrPVcFMgPNBzYme1KLZWVR/ITQ4cszdDQO5adExiphuPmfoGt6Ds0
TwyqOYYHEBdp5I/2epHwHRBqix7f5lZgTQ0ZApdnYHo4LSU6aNswEZPnJV/BwqoD20g95CT3YQM/
QWbxV3+tmzajgqg0Bdd7FXKLrV5TZii7Cu3+c7JUKzpp90Asy8a6zb+j06CcRYzWvb2o8G3t18mU
KCpKa5Jcv0pgmby6RT1R0i6PFoZRqJNlvwCJijwZvHb2WPBSGCFH9n/6x+r+ouyt5kSJjyWbQiCM
p+/b7Z+liYJy0hQpKykRTfOWfQse5RR4TCAbtlRSsKXnMshayoX8Ahz46ISwv2mHvtPvxIlvrKl8
fOCW369ebOt1vAv81aIw8FQcIASefgpgqQ0kdd487NgtdVpWN2j+u8NHqEireJfDVmIgBw0TTEZm
pgkkegCGvo+ddD9t/ksjT2vjKt1TxUQBO1wGWSKtEQ5ZKxw19+Tm+/2TW9YFlfynY9xyQtBhQxKj
ZpWYxs+IOI5Kv3+C2exlk1guYAmrxh4vyh3lVylU60Yr9YCn4UAB1TdeBsPB0F5RqvtcV00ZY4ci
rYB2OOqx84yIiDJogYLurv5vejxviZA36egOF6ZirYqIIir9/ef7kDrZvNr9CnnHdxKxqBT1OS3v
ERZgbsQgix3N/nI5V3S2p2C+1/rAQOfUL2A79GDcSor7ueVUo/GYt/NMwHvpPOXFEgNTcMaatZM/
Bx7tcyubWypnLOOonkWnC0i7IBNoqcb+wCxp+maYjqdykIIp9UqhtvkaspeJZSjp2+vbz47Em91N
ft5PBH1By/y/9H7HDuJz+gpIWy4XThBUgFreZAonIyUExtG5hMqIHvAsDRnGiH0XYbO0RtS4Xdql
FtJG2Z7zF5CvP15ZypGuGIp137WCUcbWDD1/pj94n812wXZv7UMYz++g/1CqKaDwiBrTe+wSsx9+
m/F/8K8fSYOFQpJr10QTHNM1XPZjFG8hIc8kPUubVsO+wdVDTmBODcUi0pAlPiAiKpzCc5pMg63t
vAwhilYW/qvIf/oG2Ddde93AOtFkKVxAycMOzRING3ZW7831917d/QO3VHEgrOuTeIXcOhSOULkc
7DjNkX5V0pmrUmSsbaUrCCKz7m6kG3bIilzjzk+46LUUo20mTIBfiq9Cp0i3vn5MjuPrX9TpWHY+
UgKYZn67rnHNFBqZh+rjNfryAXPMkw4gkWF90s5/FMMEfFquBKD360dM//sb5ibzwLTYCDzI0Y2A
VKLC7NcvRSVEAYzmCp/ItcGHWPM08+L0QA2758kAtzpMkrvkI+D3tFAkqkZXdaaKZK2+MOxsJiME
N4Lf9UzkI1TDAoVfR8mqLl7BXepm239YSFFsPsNVG1MjtgDLLUV/5Od9JCIqpSbi0DdLziKQNhAh
+baRws0UCOYyQw36SP1T3wEu7TzzUJO/Uo92giXAUPIsBom2Uxh36/WRoQUCf3LvhVVZMbgd+DHf
ZXMlx8GeJ2dy/pQnb3l4WMF9uw2dV75zAo03mwrJEIo3YiCSEtQMiE4qj9JJI0K3/KTVMB6O33ws
0pmb/YfSVCmkKDnurwOK4zpBPgYMRl8W4pyXiEgy05UuLiazeBtDBqlOGZuiqS8g6rDwVZPrhLqX
KQKrKBSRHbU3WhG8s0aB8HSFesg09yRL0kNHCKFYKmakcnhx2wWCFxQ2Schk0eQGNwvO+z/SpnxR
0L0Wj3UeFOYUNhYcEMM4ivTjGUVSwIoM3mM1sgMoOG4OIdG/umRvrPVq5XObMnjdUesas4Dob/82
6keHUfe2bnu7nkF7NZA0fLlAlUm0Vi4epf4sLvH2pNwmju+7I+k3AMXRDYNiVhZKQa88EI3BVm2H
RGJThP0fRkorqvrbNn23bvxAjZhIA9LcSYjIx8mZg35mAan3kAK/uVJUDjE8Cnu7ccDWnZniMhml
LhSYDYCDLkSdEdIYoxe0+zjyQsO7kTbNP43FqIJAHR5+veycRKspglsdO8n6v/a/nLyk31c/ARpt
aavC918wEoRX03XsDmjit6TnJUzKNo0vw51LuVQwOJA7rZhMHkTq98LzGxGajTvYzOrsEd6Ol/UX
7HXx+CyLqKeK13UEB93wfKx3eLN9taH4/16acDfukP7r+gg7Oboj7fHoP3Wf3SEoQK2Ex5T4flFf
oi7ex/TLfEreePOZ6R/te/LClV7i5uL5LLMKUa2JpfOEtDaeqBzzy5U+qJDJHtJCS+BLMUcNZrY6
oZnKLKzMCE+kGibUMYScaVqS6F3mCnQuluh7PKTaNyTx97wR8xDLzpbyv4kmWqnTsE+1s1vmBm+9
PXVqY6kOHTrUu1aQbfW2rpVwYPqugBpCW9befm93Sfrq5GSwQVNXIdOnUnTaOfgHrf5c/tn2vJ6v
y2zA8DS2o//Daxk2F3zZLo7nLL/qksDa+OGGX3809ZysGQKKeo6xqRKdK9RChHq93yEGK/XTzpPl
QoZf7ZbG74L0jc9QYCcNCwfOKmvTOetw+3S5ebkEIkLSVB+PZC642bonN/MaWpw3xboZRHpZ7tzI
3VEDmRaTmkQ3fFEC+mdP+9rwDaK7VscTznLoWzA6C6fq3vIViCTB7iV1YNkzH67bHXRkojknl0Ax
3464rAcP5s1M4rxZruEThl/3LCychPhpv2octJ73AeAju/2W7LvJ3pkSZRsrek1MV+kHJlnsdDSg
Tvm42GbdTjSpIOdxxMoR613BZsC3+Atvvzi4AJuMvdGv15UAonBytsmGcnM+/xOv9aZKjcxOFOAt
z0viraITk+DU+YfNxTDs9q7hmAmtGqhlTzVO3dGkLVd7pcUS1NhHSpYo5cxqDjzse7r+6qalUtY0
za/cKouAnUqInhZfTucm2wsi7hr/OdmfGoG0tpTzPW/041smKVMhJ+x5+Mw2mWdP6UKX15j/NoHu
QaeAj5H7TSQy5OXG/k2LqjD8cXEXznaxMRUD7wUJ8cDG+pU5M6M0MPdJfE0DwkX4RRbT57SwuRN3
oc/4K/pWbnVqp2xr/X31ZhRptlQDs2mOfmYaUnZVj3ZcUpvo+tM9vkoTgVQRLU4K0372cESRskCp
Hjyulbg1sVdCsHHt3j0p7ytWgUZWO5LwdPfgbcz43oWcDSNKlSgS/HyQmY0IM0OnPtTjUEiGZ7+v
bvvrOgRQLrTW8gDXu+pTD7nDeTpC0LKyixDffG21HApsVlzf8z8NeH3jCCzofgNubLKcWayMnHyl
VMuK56bh0FPmEimyD62TecXNUjEwO5wRMxOCVdtyiHRm2BnasC+kt+cDE/jsEjxu2fH6P90aQxIO
7s2x0uAIXgazdkrUJprt0WNlHy6Qv/oVjO9lGJJa8wJ4t/IlO/dQpsIt69L5qaiGJ6avBSKpNsZ/
22EMKr3kB3o+HV78Funa8fQ+WsQi/otlDsKieMLCTYlGN6rqmgz/Agk5K4cavBWqkML+s3RTsOPZ
qPSGQzY+svyqe75cTjXZXsn84/Of5xc4agDdymynKRLD8v1RZc/8UXj5Dq2l2/DQbdLqTfc0E2CI
PxhQzFC8wHlbZeFwDF5G1tLC07qiv8ijBSPGNRUCiX5WoitqddPDyNn/PqVLBi3+l5wY7j5Ct6Hd
VX6NqSSS1BseLyl+zSyFjEcqaVRjv4iHNTq0rERRQ5qfhKC+N0CnI92dJrLSGnHg6n6yCgIcLNCe
ugO4xywi79SpmIJbafozjoQVCAbEf4bMu3PnrdEZaNI6SjEK4AiXiEQJyFEArYtXURvabHge0gfy
f2fVVB/JeujNDKTqW5HZZ50ejhU717b7VlDV6hHH6GQ8tf1ek6UXDza8pBaA/TEM4PoqSlcZz1NJ
APyl0GCnNiwDh2EcX0+5PNRRNU6246mFQRo59jMChvO9OGILD1FSL63Msd82Xjkr+k6Io28ALhwK
pLtuiCOfrfKDrk0pasKaauRYA7hlgjzH5OF4nhuOomKNl1yGslOMslR0Hkl5YwywGjkZb+JB1ZNq
P3U6FdM7S+EN/xi3L6BUzliAeETwGLkcLxDsr4zDlnWtoDIndf6kd9RNOBrMI4AwWwHF4V/Y2c1F
YToPxMXSqeG43ipJbCDKrznPfndCjz5ajr2YFEs+7igqIzbkzMy32iWVq6m5QNCh4CkGBT0g9v7d
OazoNu0/LwvPtWTvnPHvx6oaNtCY0v/v5uEHFr03hvSSCviN9NpUzYtBADi2kBKCkV7eWVE2iotW
b/yRLl3I+Si2o5x+eXQ1JabxEn8R1bsMnYxO4aiMbsPD3HkGLQtK3zu+tltE3fLGrWyBYWjzsZhr
ia3sL+Ajs8NppignCni9gGmOzbZ+X0DDNXfyPC01lEcx0WB5utsbLs/j5Y6CEV9qMOF0TJ3d1GAx
PO59BMgmr3VfMIBkUcHGF0MWpfrA9DShF7leKXVSM1FQiGcSdoF19MbTUHhGaEicYMjfUkeQURJt
PY0GA9GW2umIX1IUPjKnA3yvMpYdgxHGtDgFdEJbTqSShT+PAQNPTJzaw6ch9PPy1R/cBXNuCl3o
hP39RPU+womLvt17+VFO9REFmlnrcVt/TEhR8pfyESrHwOEAmmoLJvjOzw/I8VJefJzoE5HHNkye
HxV8DN9Kaq+aZbBxjp8vqYGQhvGly0sl4CQc3mey0ezDbp92A1FjAom7Kjl4NK0Sbk2VXIEE4KNR
cGkfPfjKWgr4EHTaIgXNqwRH/WXqNNyJpzukS/M4fb3Jx+/XItH8OKHiIMuroHzfl6j/KFXOKNBH
I4puN8pl7geVk1fkfliBBtEHj8nuH/fnR5X3h2TTUo06j0R5gZCTZNjrYp/su0DMeP6gc1z5rqbF
rntfVp9HrPipqacnSQJVMiNg3mQ+xTRS0OnqnYJ4TfkmzklW+a0PfP07oATvNDOjmd1hzLpLnJi8
B9R3+vcBitcsEOkckt3NYXjhA/QbAlLo6T4jO2ZtNC4L7LoxXyiEh4nhUDBZVUvjlNIvnjMRrGuI
SUXkwPA2NcotlCm70Oa6BrYvA3k2sV9eAw/s6hw33nUXchinRN12XsxVp5ea3uVTmqc25VuPupmM
zTFamCMVhQoZtOHhAImb5MK/LaomRHDFvVtUbG0bXPrWAaFzHKwJNWdyIMxsBdQnN4ZxRznxW7KB
vSBbkoYFUMHUF3jbXQCZSdB49uEl2DhTcc8rteLgJXrgP/MXr5rz1PsWbKl87V2fNA7D8JLR16g2
uW6k0Aw4jXq1wE0/iH7iwY1vwGzTrCgl6N8qkD/MmHBSp/ImMMxUaRtwBLrmo3GHJqfBo+6pozDM
OKqG8r+u+Whsaazj7mWWqJMbB+sOicjLOwIWxlT+uVfvGoTmeKIBIZ9jnKVZC9H13O6fCVEa0N4E
DvBQerF42ne5TCLMGacqVAtHBK8TiOf4TYets4XkF/WqmfHS5K69NkSSEiN5VeHwplyF9XpDxY9C
BDK6WsYccVd0E/sLN0XcWP5Uhft47XF8JEL0WXAhuyZJ0ATQ61afRzV30os8TYdtiYhSjCj0d/B7
jZ92dwi/RtpyL9sngTX9dQRfuHsjj/fOKzYx13ihRf7fXFXSfFuzZDwJr6Gc0toAmfrNSSkkmSoz
/Ft/RW/OfAVoK61cpMuDykN+q8KXipzElq7xlv3M/ObAVNNzOPxfeEnlfoZzZTCYgm5kFFV7lTFi
Kaek22hl/lB3sFoMAagIu3V1MvxBVG9Ag08n4q1HeBU/fg/Q6B91Ubt58AnauchaLg++wp4g/nN/
5EX+3akUGF/IPnYr1aWS9zg5JMOdNiS5HjiV574U5gtNX1wg1B+Dhk5IJ6wzi5HPX13fiHNvgOce
j9HbyWOX561y639w26HS4pZk23YEYC9dojw5UnmDhfq0GviCfzTZuxgveetRqjvFjaGUUQTAt+yc
izMSkCkAtoV2HtmSJZOmHQwNnL/9ZQlTkS3qyUp22cKOJeCfjvxV3Esk/Fd9KbnnJjaYUd896PMR
NC0UyyxxotXUA1NGA5za026cKXK6pnetSTiJbn0BKlic75PXrT+uOLftLHBwe/CEGpF+H8g8+KIw
GSz1PTPv0r1GgdgWbC1mgh1xQjcvQ3CoNJMOEExcZ1aR1VL2S5aoNBX2GIoI4lp5BKCoSfVvwYxg
RJbpSamLojIoXggB2b4vE4kPupdDkeuYQPIxfmHpxRx13Q3z7oINt8r1zSLQPnDZY0GgFIzHiwBB
F3/s4aUXaR2TKzsPu8oHVZZlmSLWcm8F2ObO2gEWWDfU9xDg59K5+ZEW2s4cVAP9ugYXB4P6Pubb
zbEjtn6Srg4lnb8+8Ikd3SK0pFPpQQzNhgYtk5c85Xib3VGDG7BBKs6AAMmqK9eUeF4MS5r0HYZY
dcDX+yNYEOEuL9JuH3H8kqoAGARW4cL0BkVYlQe2JvqRxdcVAXTp2EgSoBH6uzpX+d4JvdP45IG2
C+aY98jwi6vGkxWvm0Z/8fpGrxGzsuXVyMJQzZ3bTnxYYCLIkd+TpdPCr39Vy3DY2liYLmI063PQ
2js/F6IzBJ3rHY8+t6xJtvYzvwHlMYRXJNjDYeLnncn+ublroNy3VxJLRUpfs4DbiEBcGpn0VINu
aP77IXi8tXAv4qrZYBj2FoP7neUkjrDMhdwx4b+Oi0xxeXDDlm0cJRNYD/F/hYhCx43uCfRjHq+m
JHZDsJNIjo7He14mVT1AdY2d4tj+XmROvP3WCgscy4LT7ERvVB0pq+BYv/7N8R0nk4/TzY3BR2ZI
VADWCRFVylBCmD4ks/5T465gMEZ9dFzFZoW/JuMp+uE2Iivw3LfiCni/PuD8HveLFBNEiWOMGF+h
oGaK/YfM4QDRXVjsriiBL0vjgr3dpheMCIyKcpXJCBvKc3Z4aAZy1aZ0HiTQ5pOtUwR489gsfZbo
/V4BV21B2E5vOP4QtJb/zLxviHNZ8m1Hlo4b8rvAJuwudV0fhM9XQnsxD61jV3G9Oi2gW+fNLgsM
KGfQQ+q2zzqFaOvBJ8WS1ixNVM3uafEhBIoU7weG2imFa/Vp223myDwapqmQOT6/ZV9N4pUD1hEX
6Kf6kK1GRFgiT48n0MutAKKh/HyqFLeswdNohvA7vwisL+qea4PuFNp0Wlrp3dzY4qax1lXHYTAO
DpwnKyzpNtta0nUW5GRkIIAf8WlX/Ql1/MK93xTUy7j1KaMLzyMb4FYIT5h0SnOu74qILu2vHIps
oA2NKX0poeQOfrnHzXkfSnIi2N7soCCCXX+Ros2iK4rKOfD2ydu7/gy9Gge7MZvpEsRa1Nr2O7HT
wOWleGkuLT6Y+6Guw8VUeiUO1DxYJAoDK+o8o8OVOIxCB+kJeLaZ0gTjDxgYsP0kzYfMFVnZcUam
BnlwoeLIoiZWRbDvVQFPz76CfBGsFAzf/Yk61msHNILj7I12ZStL+n8McD1OUmUxDKoVl2kcEyBl
Qciz5utGuoh9nMWzXQ9s3aaNAEbVfD/Ofto3M2UCP3dmYz4B16w0PYpjieyhhqEagfXCtNZsO01f
uSYG9T9F05RqkRxoeBaUFgo5lyrtPp9cRFsZa0qXRgRxlGVSuZWFU/1dbxVyAw8r5lIAhZ1rhHFM
OrP7zlTWeuQQOqF/6WyWt/CoUgxlUYOPqKCgzEJBXY9X18n94ShoU6ajFZAO2IpjovCtCNMqU0M/
/ZBypJSTQ3uVpT8I/WRIM6+0ifaP/vDBDsuaU+T+VATsVu3nmS3+g2cPYh2psUlEg1KbaXvg4Dmi
ifatvUKF1MJv+FIwTsmp2H8CxzpUT0sT7toSTJ5B0Zx3EbHTJrGUhP4h7xJnjQctf91gCa/+qsX0
bgtEfC1JtqWPFNBbJXQSMW8Le1yGgAk7NRiqj7BjNMenAQ848gwHK373tHB+qtKYnHIyexDJIbY7
Xpy0ug6ce3lBxK8Znx6TFc6B7YtuWIPAniXbU78ErRPSBib7oodiX6du2tT79vOThtKhlIjiIUZA
80xc+6z0ZqaYQ64svdlBRt6gWtRqh9ToU51uDWvET9x5UyBzjxs3W42g73u13oTEniTrxdsy9cIG
gAalrPo7HBs9A6Ogo+Lsg6abGSpL//1tGcv74iShVAogqLiZhN6ACvYKsF9GXZEuvcgARElgsBPO
8mc7Pq0lLbJHQOSnftqgpa9nJKjRv/adHd5IifbNzY/B1g5EgfiibDHaYTBBk4tDIZu8N1YVhaTs
m/IDbikBNDF0omLqRwN+s714xWXmSk1qHdZ8txiyhErTMLP6/2yJ0MaxFHZOPY1V+3CFcpq6Wkob
PciVg6kX4GZnvIA7A/f+dDRZdho1T+jB9VaJpcpQdFv5iVAQXwUSEKXjNgLFQe8pj/mf9Du7YWTg
3NsPqtV14OCLvJplCIx8llhrrFuRGP7WqbJrwoOxaPCyPr/DCzsvZPmUqjI2a/086GJ05e1nN6I0
P+o10836iIVLfpjhQwZw4PhIHh/2McmM+cwkodWNwzgm4RBMx2W3QCLT+0IvGbHqgxdWWWPrJW0E
Gp2ND02gdklPEd3GhcmImssRIsKKs3Eyj/YJdqcK1RhEiJhk8TEXfhkRBxLdqsei9A+nt5Gi/Nu+
0ffJ/CG/omr3cF5NoZXdeqHvXHgKB44RGbDVVsXI4UXYpzgcLYxWId2vKDDwJhX5kMt3thzNPPxf
03+PWw2mz4bZ8Y0jsnv0uIoL4v9VxJSrRDxct4ZsR46OvtE1rQKC/wjUVh/bB+5SaNH+NTjNIZzf
jPqxHIkGj/98lXzACRWBnieZNn6xGw+/iRzKpWBqsQVNLM8oNaOJ+8tag4uBCtz3qB5Z78g4B8kB
eHFK8wW5QMS8lH3EnwFBcjULYoc0PK6IudUz109i69oXoPSuNodT8rKOmUaJdoImt3taTK0tgkR9
CmONKh8D3EiFjIByad7aJ/e5xc0HG60G5ttyejItEmokWZG/50jx0Ra60zShQCoNKBcut+MZpUCJ
LlrjWGILS137jV1eEuuvOleAz1wDfOfUV2/9DPoDSS7GPqI3v0t/bEowKG8ajebCpxicKx9avEzS
8DF8ns3Afu/1AMGX6HkmuDS5kT/TlE16RstZJ2uHI/5qRZwAkGxjQz67URUnxiTTGIlcrXMqHBI6
tPmCFFmHoa4NWuwQUlA2HxShJ3m0EBI1v+CjAkSM+zH0qmUy9XJGIsJdaZcA+W524suHrcAosxpO
5gOgq33/qt49Y3KVmfPA++1N5mplOe7AvHSUrlvTsGS2/lP95vWB+RdVnwPhRSMxfD+p1bSKnCcC
ovxh0jlAreHab0A2THziwpchr8h77MWhTu/V1sAygFVVs5DniAfmByp5g4eS8YJqmm2XycqZr+Em
+uXVZzWkGn0G/P2+xdAiA4NaXq+JyFrcXsSB1OnbYph8FmotVr5KLg+dZqbsKM79NF6opjxtkq2B
+135jB9toihd41ubtbXEyhSrJzmYQ7klkxTfpwhXm52udeabhslSgtaldrQBGTI6izpPcf/AyC/4
PYJeD9ismPhQqjFHZpSEVd6wAnRnZWPT+O5W4SXCCbpU3Oh1/148NBbIFLGI+cYHFCIj123cwqPL
Z4BmRQ+S/iWKMhUUfzHla3ah2TsDFpT8xiuvOKtikETaC2/4NSZ/vHYzE3uuSdVuyfulmmpbgMKB
bBTn3cN6EmRCJHvbLxBAPE81boXqHd7LdEKVSCpDj9niW7mwHBGwGapewjlry+DUZkwKvQzfULhW
ZFY6LnExkVElp5mI4rjOQg33Kg/CxbT/tkgQGI4B0lsFHlLc6VBnm3xd+OVvWFJab6tsSPNvxa1A
oRr4j+EdvKaJK7/9qC10dpzDTjCw9wpJSwCQsqvXP58V1S+7y9k01q/A7X+uRLWWkyoGwuovWIPc
XMXeUxJ6JaupeIUz+agLP/X0YETAk61LZDljcQbksbKje2TBwXyAbvAZ7erFep1ojVx59lrukceA
vtXMexW4SaNTBoqAR2IEf56OUyRRSt1JxdnYQvbbowr2l6B5D1qUvHrcRu/xrh57Mzn8uIZyiVfy
c91SWev24mc6MV7znt4t5w05PxYQmCkmJuWAU0UxPq7TbBQdi2bqPqFnweMJVDoVZADl9QjNJVYG
E1/CU8pqMh4emfvOFCMg1jq9+pp0SZTP/GknKtvRE3nCdWFWybQOKklYf5OfAiuTtyhF+S87dZWq
3GKApVIRTIaux40EFGdiuhPZxtSoQxlVtblFjtnmMB8VSoW+pyVgPbMkkQug27QztpYH68CcEbWy
HIbWdF240N3q6YwnKv8jWBzUtexUFPlICwjaX+wY7oOgmnRR6Mf8qx+HH63Eh/2QC3xaPmZs03J0
Na18DvbepmQ4qzwlKkvyRd29oIzAHJcW7xuRXBxfaRIiGoZVrDeEMgnYnCw5/agfNvo6byR5GmpQ
y30vqrNKfNHoxsdA8Cl4QnZThXpGM6mDtxAAuWQ5gZxIbFJJbcMw8mXMfclpHdMdzrvLK1a9sitX
VJwcY/+vg+LGcuOCKKP72K1KJ5ZLc5e5xULlv0dBd8n8YI+9xCUsyfZqhWe5pXMIOReM/skLmaPX
UoE8lmIw+ngJfzlDXvlZ3iB9GOXQupgrguwx4xyLUY4EMJLOH6FijVFfkbcaQI0MV3QJl707D3cx
FgzDhX+nojZR24TQ4fajrkP3t+vrt8cjUinh2eyQvBEMDWUA6KSL/Tlf0oFtZgkdJ3wtUxNSPqqS
hBiTFW7JYuYekgXaAvYbhIu7emXoGi8efsjBlxIBqdnS8NuClAK5ei+UBsSs2/68JYjJDuPmz2Nb
JB7b2pxGmn/lA0olC+cFbTLXnkY40K5UIirxtLqDSGlBjUaK6XclTyq1tq1NTs7wQEijQP5qHLfn
pga9B/Qtt0mzLzia+oI0cX0OiIVocsAVA692hWgq463UL4KTsFVFowA/2BtLFT14S3MjdbFvKEx0
ZxNwD28llqAiktk2QV15TBSCWcVEz+z+uICEwzl2V6pmqJjXzPcAHi8rl56fvdt1FJnf1OV5+RfE
X05gC6JrAG7JFZixC6BefGg3c9vuzKanCA967+Dkk3cOi2sxCazmwsYe5USfEKKdi6l/mClLnmgd
5/SANLu4erAN66NbR1VpHUvMak4t6YM5DqQYydF/EM4xZqEk+iawQC0mx+zvnPexA7M06eIjEHG9
svvgrjjH/nO/JjDuMInKrzOsH9RWyfQ77WQIRovVE84RdMS0wEmyJemy6AFz8EWFOC72PsE1QITI
q+qv/ye3gTgaZXloquBx7WjsnKEXSF+yt6cloQEFWQyRP5LNh6uS8T7bDIIuX8LL+4m3sWdJrrrF
cga/3ynPRAL4MXHAnH2K25fRvdWQGU2ZIWpIq/FgBr0XIbE2/yy9f7j+zPxuz6e84IkPCtLkiOzH
Z28sHkgZEEJ3rrT/w9wiqhlEc5Qfou2ltNiUagS4dcVD2VHEiuSn9PlGPPZZmOAp/H0RrmosjsjA
JogHGu8zXNoyiLibWlKCio9mDut/7rnFeBLxEQwu52IfUZ4YpkwuTKisSRgFDPziwubZKbpSCdqo
lJAkLoJiDkoE6UkCpXMhgEq+J7BCXEyh/cdSAVjQN58v2noufZSffj/ZLITBHfivJYh70KsEjv0g
Uoj2BWFd/xcIX8INQ8XFwHfKpLhaivVG4sakAD580s6sQn3h8OUKyJdtw/3VcAEnqMn7pgfMyhyY
5NlapttJ87oeoQ/9H3RqLq8arQ1k16vepDHHHndKCwiiOxS0GCwLQIBKNst+7SXkydZ0SbJk2lIx
hxl+crsbRoOsT+A7LhHUwoAyBybUWkwrQEj3BoAcfigyW6kyCAgtOe/OwhkuOr8lkOK8WBOQdCGH
ms5zn8oGXBqN9s1NcZ9HMCo+J9+DPRshf/NhJXfZn7wEoOj8j/HDtLDZZefe5vo8aDLLiFIxnfu0
CqpDLqFsQFQFfkPPUk1bDDDQEkOW1mGV2DlEb56k6ephJROqU7WWzDz5+t5qMFZIA+zSFzvD8r7J
DONMhPV+4nIZE32TsaliuOOiE33+uo5fB6oUw+YItPXWWAF9smj7hNhsCfGkcEP1uxgwgYLlSFO9
Xr/y8mk0dLu1ad1g8830FleW2aHgsG9NWh50fekrvOad3CSYMRtBOqTpP+1cOMIfoiDMfFLSzzWK
SVSrIKQKexhiOFpnOO0SSTndykSmSRfCv+X6g4OtxpId0QQmedNEjCGX6bfw8aO/niEuTpUU3Gfd
9rljNWGMxnYiyxGbaB71zb2ZQDAAPfzTenPrhTqa5zy1d1HpkGS9zlDs5D57nbRNvJvpzkShWGfd
8SwrOcRpsphYLmroYJSc4J3+C88nSvEPm9Ex3jAxSN7moKHl0x+AAvRbD/k9piUYjQqsoEbpJkPV
3qbiC7zA/zq/ioUbdRxfIS6REO6jl2Uod8x0EPo8XaK/iOBjBmV2eRivGe8Q+ygCdbPZuzoey4nH
KwcW5y1NDR1GEkzNvUUuj0SzsO00FdWx8tmp3Iq1YO0z5QrqNJ6kkIJTMgE/nbcPJliwijL1lVDc
d1eHfDgmRXAII2bYPhXvSkp2DjBNn9DoOvXXXn1uPmGLiVO1vrNxbMqplK8dgaWpu82ZBx7ANtuS
ncwH+eBsTjy40+NXVgFk9ZbOWdpBi3wCXhjM91f0RKEWQXGB5vdlGNw5lxsZWxT0zqe0noddobLg
1mf62eW2+GyksovGOrYCRTaQb7dHNKiQnyEjjgYqhcqBjdvKsT2N5BQF5QXDYNeOVOjLrNOm/L5T
4h3eN4yrx5q2Mheb/2dQ03QIPgo8Cqv9BD9A5skYdSKoJpCNaDr/PgSlHdhVgjcJeuUaO52Qjwii
oXJTECdBOC6yIg6LVoN8tX+68OILGgAL3P7c/kQnFMjNRvMyTzXCqn6c6s7FofF+4RnICWhedgSQ
jJyLLOLaw2t0ws55XQPBLpBzu/LVtyVKE5rGvgTCbs6guKD5Ld2OuzoI1Pi34CzwhsuFZUjIrlVw
7CEFzMACVzBOW/Ij/bL8UtrpmpgXl92O3i4JtXNgJwDcjuF7RXpYrB6HM7aoXJqGxhTXfXBr+zqb
dumxIAOom/eazTVfjxJhpo/BW0M6FFqR82uHjU6uLDq6fVrtQyM57PQsOk9tqM/rKjUdZO//LPn5
jZwmtO+hQ97PR8qAaLgE1QX4cTERnXOuE5Jzr/VTCv3dLaBfmGT4z4xPEkuQNl/fx7ZXnlNwD2nC
2fRly1p1C8vjTwVwuZs65i3at2b5SIWMPUAobowd/lQe00R4oIY2a2Ha1gsruP7OB6lyDiwl1G4J
HM0SfFkZw94PFR1mIS6Mv5Pys0U8wxvfgwGCl0PS3Q8QC5alntBBtR2dNoberOIE6rEkpXGKINe7
xvm3fR3ldO4UkqWFNZYa7q3eql6/KvslEdjBBgThFOPFctOV50uA44pVgT4U29teWA+lCjUNkNVh
2r3QExYy/q58iusy/+jjCp6xI0DIute1d6tQv9U5ss2PCjYAZrVE9vCP6Ua8oovQwxlpbfdFkzon
1ZYPsuW43UJXev/Hd6Butu8HdKgQ09uNVi0iqaw85P/RT+XiKBbKl/+ms0oO8NqpY+3Nk6NG6wT5
tZo22L7ZuQFmMpeREAneOhfe5NGST4SOaujcJLzm1Yob24sBww+0/M+IP+Zqdz4YpUx7ysPd7GYi
n+Slm6tLnxa8XilwWYvWyR6eBOozD7/sUbXYc+2Bv/3PexKDU7sXUZUdYTozoNomT6t+krzyNP19
hcHKd7t8Rv6IVkZhuNXyp7QGi6KlyqLqMXNUA1ALiy2fiDhN69juytR65jC7qksA+bVLJZHX2qut
j9uuuPn7l2+3nxNnh/kTjJdozp9HInq9H4mWbD7meHn+QGEJ29rSX+q7d/fQPOWjZA3y9JRydYkc
Hj+ZiQFfy6w1jJz3s+zZccsiwsjTiGdKBNAMSG/lIZmLLzNeWJUftckY7OX/WafRaFfS5rkcl4mg
cr43lqOJyf7mDcSYzQndWltEnJWhxmtOJB0zt+DJVHXICG2whYPCBCZxbsW6olNmciusP7lJtckI
L35ak2c8JI6ckV6oQcENdg9ugC5FUfmPm01BQ2YLFvkMyQxS57tclC3qBtRxjCr3uAm1dcA2IXZ2
TglVuAzAg0JnlGaBpTUBwcx5LWFC1OLi7RhDzewLfuz4t4mnVMehOS2hkYufFNSDaL+B7klRsJda
J2ry7V2yTWc1VkLKYWLHM67f6qpbzzKfXsFaxn4SSQ65H22ow9NB9eeEeIsLvqt5H1czOXB8DI9e
a5JQTsr1q28rlwrTsynX5lKPeCgQZ3JPAeAyqfXO571LEgXPpipLxymHRofne6SNzOw8Y2qzQl7P
8CP3fktCgOiIPvJsF0V9YiNvk3nrpYT0XehxhkkoFnBiDq/tRj5VZbS+YVDkjap1MKL2Ov64j0Pp
ZONFiN7kGMafAyw1li7wMqLYsazmqrpDOmodkNT8OqXYmICAHvxVcGx9IinP6QS0ri3N1x+qjdE/
t0XzLcbJ8pO6YA41qcLs3r41PsoEEwM2EKREWdokdTHx3DNFiM/OoWO07RVT8PNjhoRB9VqB8doO
8ZqDzmyo9vOn7NZLUoWK8+vnko7E8Zxv5atUxncJ3pE4YV0vkKlIFDtJDb5qbu0Pzz8h7Tj0TKbh
HO7c5K107ZhI2gZb8abk6Z2BaD3YjXkC8h+NQa2g24kYvCjpk1A3SJApFbujCmwhTKTRAKlUXLMv
mDlzYgIcMmOL9OYmFQQtlnje5e/DOsdCvgrlrIobA8LsWA0rmP51gAhiXZNELcheJc+alxzDim5Z
4rtArrF0OXch16OaE12DbRcBDCZj/09J6bFEc85NUQjpn7w+4T3OJM0GgTK1ihkQe9tY2RAcuMED
+QeOtr/gEOK72wQS74jp2MGZ7faniTO5Wr7/qVYS5CBbB2KT+rwYV/Uq3jvLERiyw7fJ48WkFnGk
9y2G0cWtdr6SxDRUsmEWXOwXlBRexxoXauzY5gWZQjogmK5qRXspabdA0IKDezAQiGv73gfKcWGm
qURRsGXsjh4mQj/7qB9mzG4ZyXXCj6KccJg48qVYhmswEH6vLb1LLCSMIsEbYWxtr7aDq+MBDXwF
OVcWj7ik36nMWAn2JUQ3oFPVFNYRUGvpEZOy5gzD0i+6FVbTTEIau6TN2PFicaX/cGIkFWkqVBua
RaP7Vjm/0YkkeVwUUgtBj1O3QDiEZM5Dw9Ae85kuGVPFHkcK1304t+si1AQ+fiWRr432hkjL8yMh
EVQraxVqYrG3niBsP0Jz/zd+LvvBcXLFCyYlHm6dhBPSYwtbOpkotfoPmohnFcv/9xgrPqAlE1wL
bqoKt7yLncPAMuUrgGgh7O96S74aIVtbT3eGoKcJLuoFqkN4+Tjt39Ss4I047wNs0sJbyjamhqdP
zx+hGNNvev4MDqAcdt6Wyyjb/31qhL800/OB/I+NW6vML8urGzCInf9yH5tHExaHwYvMHUR73hRH
eeE3D+bRz5IwIgHX+KyeUgxaD7gCk37celDsKLkagZ3SjKR4zqCd/NgvM4SEBpo3Vcog9fQwd6Tu
s3smZ57RCYdQcPh7YGSwExw7aQIpDiKuyaH4ORyIjFUNyuwU6koSAUr45VeGDG9tGClh//U/Feg+
mxqlw4uslzcLcoSX4ssRSoVeNKQwCad0jRpBMLlFFmL9BUrVCQGISRfcsYBh6RuoK81kpuVrozak
bYPTwDAultjRV4nr0IRbn3RyR0s5AkZAOjemvbMqgpLOa1jmwqXh1gJSE3MfrzhB1HQAyMZ19Tt2
a3WEcHippIm8T4q86ogzBp/NwbxmV35fZCr0Jio9/NUMiAnn47eeioXAWCmAks+NOGBLyk/Aqlyt
coO0xyaUu0qPM3uKNCpNZvmMeeaNEc/WMlnRyYLoMFzihQjeYfWyWbkpmSybCFAHSJiiEIAgU2wU
DdT1/Mq9UlIbuzRdyvUThDVm9KV/4qOrFDBStmBknHdfSVGAoPh2hudX6F8kZ4d04/49MPVLlACD
rcnAxPc/AZsuoulFQW0EcBeObTHK2B30Zyrwju4+2EDxAKc0quSbBeiE2gZEfyyfdUrIrPfeSqnW
U7mYEre5lkbjtlEE1bP+GYSrCI9ytc1zSNU910r3IonElbB7bmmR4QAhvTu/ST9dUsQD1BQhqB6r
dRsMhZKU+yzANEaecKD9LpGMKgAzWBZTDIwMpdOAEIP2HckT68ICmsNmhTGtUyDGPuCgyEuGdbdK
B1QZGjtiqvj0wKmcOc3tTKLijyw7C+phoAu3bpGJr0CNWgn9jTXNPM5Q+ogo/D9oQBhSSsgQ6GBc
ehEn8GCkiNeMGfpnYc0L3YZghJW5ZN8uimHAHFL7bqDWJ2eueBhQ6VE+nsgZD8rOjoVLosIF/psW
N2TWWcrmIExWsR1mBGyRIkDEzIZWqiTngKJQBrUSXWwXCIz8f+AvGemZRLk2XBJ1Xi22oS8D09wf
UAmGMNVJYJzh/W9NmRjhKpwOxvWxECAbzRminp4b0g/70Avpa2tQThM+wYyXy3zjISuxfy3Cvs+I
Ia2cr4dJb0bbJ0eA/TkfA7Uwh1KbchT1VgI/RaR1wxwgI0ruWE4Qb+U+dpv9s30YSeTikubstVJw
7XGxZYVO3sU8ngNbH1NUeJ2ootj0g56cn3z9E1NFy4eg0zyEkymntfQpHprMVcHVhKQy9AQEDHNb
QYRERLsWWN0ZlHIM8zVO4ditdFKxZqGTNd0pT3Uq+6XoYDZC1Nuvt1yrPwaZNWF8GwxguAdtKO0X
yjCsprT4HvplyIPdq5ijokity22jUTcgBjscNs9OIajBOz/0ntYpj6VCAdqMin9yEa5fILwugMvD
LMOgyuruJWQ2P7WDzusHqqp/rYr+dV9OpgKcqppCyWDvfH3s8P9Rm7P2XSVCPkKy2MwPWCqBbqbZ
obPa7wLNCu2GaDwOVGjpFv8LLqWSr8Lkr4VEdLI8TbFD51Cpjs445zQL/zOpq9NPj2niVK+u1bQm
vHyZUcOLaliRopuS/vf3E/LBz7GZ5HUFSwVto2JXY5zpPztnk0eawPqymda6xem6VPZx9Y9Gveih
sedc24QUhr4LH0lAjzJT35mu+966qRsJ350I20Ifry4VeDf7rb5QMjah6a6VYRRZTxjXxAXnoACH
xR7bigvouYYfJh9huoLmvXnzuc//S5l/ZEHDJduirQVGJlOHXtDYAaPffNw29W8i7M3pywk9fSzE
Ep2B0w+8wfNKriQMmXuugMPQRsahNL9eK/eO7I3J2bEdzA2bkTNqI2A8Oew1nCe/CvyvOR61vOdE
LR5gkMULh/1RK8EJZz5NzA/SAPqt+wepacwu/DMPk5QOS4sLlm0XSwlzHTfdpLHuWygZ1vtg892V
PdFaFpD6aYx589NBY4eImMD/CkOHE2qnBgfgmVORgg8QflMGgWhP0k/rbniFgfyLj+9aAsF3dQNX
EzEvvsBiIvQveHD2u3ko1H+ef7jwCD+kXQWRGfVLUA2+b+fVjgb5AmfNTiiBtoUH0SY+YRybTzKt
awj/ruIyh/FA2Q64mH0MaxYDevf/x1lSdg74BKaPjDcT9Q5QUOXVe0cXlMHpAmgZctE+aIWnha4R
PBVNBQsK1hS1qtvz3TcJK9NkkXqZHbj7wRVolm4mzPpp6ulIat4UJJuZqgkfq5hDEmQSSipv9cfN
/n1GwB7u0n+OMMFXXp9YUNp3XRE2+i0SHICp/PT8t1kr4jpEnm3LFSzGLlVcBreR8df9Qq5TGiAT
rQPSMxL9v24V9UJv2mRHtdWgZwIwjflpU89ZvwiiQJga5xlsVNS5g7FXBPtZz6NQ0mexCUsduUuX
FvX3I51MZ+HzXr5d+qQfOi5NFXDl1LCZgkiE7C/kuIdUlDJ56DujLZvj6CP1L6jwGD0VEo2XrSO9
62TXivArrwdsPR+ka71tAXxqdWEkbgp+jCnOf3F3nwSgUKN2bSOdd5y80tXmTOUdIUAnk3swLcmG
vA2Tf74uPJNzsOFkP+CIhVutg85bIJ68XPvZ4sNadftCRSnMzyRXnhfDZc6daJZihHrRvqOK6TTj
q+Ho4RNImbHGPkfG0ApEj+eA87aX0uSnbKAC985nBPooGt6Z09s9A4EUB+t9yupcr1LWwX4xpky8
jHu8HoKJJZfYks+TmmYJfeckf9ydiyePn/9P3Qg9BY9Kyl3LJ7rHgCGufR4Nu/W+ANv19n7/n5qj
2udJUJPG2SHSNpH3EsZ7Cbl9F8jmJ5KJ9WkOyBHp2ZxYbqWUEgBYae559/8CMZrkl6QdIkgn8nZ2
fsBo9uWKTTJsT2RliLmB8iW3UXAJ4CJgX+5TpJUhhq3dMcECo1ZNuBDN1RR051QRlPi9TokVCDDq
9LSXiKoWm5fE2EKodFMde4MwmKrYIFKTylU6ls/VIc0G+6NXqwYN98MLm5421O1dxuPM3DjCJuET
CwOVz1ntXtR6lJfDvjKy2Sebrk4EtOvs+PekQ2kYB6lVvBKFTRxVa8iv99bpwSuIqqk+1BFhZUlW
QL2mKo0rBFpYMHtZVPiEkzR+E9H/ctBSRfFey8GhqT0RI1uu0clKBxmCY9tvyONq+1c8z/jsTyRf
8uPNr3P9gW+RNFHTikJC2N7vi1ay1JoLeZ3bUr4xH4g0IIXXxrtU1OurkXgJYGcz+mOXWHil1TO+
b+9paSxk3sbaHjL4JCi4v5hAK1u3c/s2geSQhvkf2W/Jq+J0VgAg5k0URrPDvovNyvFU/phKJjhj
v0OJTumkG+a/WIwldHO6bHBAKP6cpJp7eA3Vp3a1E5V4XII8YQGKUGHzYu7KGTJCNFkuKZCAkPkL
/c2jVrMR3PTJNNlyEt+K15jGmPi1RUikMkXYMFGaOYMoLgSa9gH+EUzU+dWrA2YTdcVtssEyzABm
OZXVASLgjYzhROazD7Ym6sPxo07vXPqhjWWGXNkVDcD8PAXSM5hOOxae2IBPmMO/xHY6vWURjT6s
Pv02gRmNNJQ++VBvGIQUDnt1Ob7EsziatXeTlvRm8XWzESq0XCI1X72AcbVtnFTtpmTPcHsXFBOO
wNBPiKJQjWGo9Bx0bHNJaFMf1nrcdG7kU+Dtk9swSBqAHJx8ukPvqVhhsYuJxGeWJnf+RfXxEuYg
fdW6MKgih6KO861w9RdsuoXuzIqeNZh4pbWRvhUNimq/zXsmKup1ADWrh8Mgu5KIZW/ZuQaLnDW0
UfX40gwK3irTq6IfiEafyYplUTTXPpJzHvw4HrNa8NqD+lfPdWFux1/k+AjIkxgVOCFHFGfP2iJj
DEdOmMmxH671kdKWnu6SXVRqQOhk8bH/Q2+dNJNdNZcaO1VrCNNalL5bVp8EL4ZQlckhKVq+okj/
Z82Q7FLuS95+/qSBGjF5B7bz60Eo4+Xy/qxUd5+y3t6WgyP6n0PHAwOjYLMQ97rMqQzDwy1mBiU1
5lLRnr+XZPdoth6wUDTFrZraw7bdnwjDCUHWtZTSGBdNI3PJwYOXF5shK4Gyn1Q9Dikc33kqym5D
6Q++DuoQw88dOyLE3A/OKpQPZ86lKa+AERWElvLmfcs4wvNnPW9lYGzuo1vwB90GF4euZFBuQrCv
zJz+HQEAPjzW0mmVGpYkKR+tfXHog+dzmWYZcAYmklUKuxQ9EFlNVvmIKuWLA7UpnLDgHe/HogAu
IOol0mtTT/AJDnO9BBuUIkRaQqVsbDvvQyf5p4gGgEhEHJB5SPRnOZoHRqfs7bNHgVtszd93bQhC
QXYyeoGZ/tmoTB7X5oCxJ0XN8T/QV8/Uq5drhk1hegQlb1aIXHJBhn/Ezzm7A+j4HRV7jZqxd0MO
X4448XWN6elGDQomvUKMHfIGj1DxmD+v8/2F4EAem8rTYGF/vBb4e7WWJi2o0Cj4RtscGesgzmv7
T5DTpq8Hi8ky6OVjdbD3+IP+hQ+RpOA9nwirUn3P8E6F4+5T4dejnMvZV/s50EQqUjmuKB8jBdmK
yKqMOi6w3z5N53z+FVJthQ5sMRNas7PD/m0bzPaCxiZUQXe8liWMVMfsneLxOaNG8jsvIe5gWyuu
Fc5TRtJKt2icorIohRNbcA//dStrhK6TRq3EUpIGiD3GJkkRAysdT8k8bY6IbL4X47nr0YsVwFXz
z0xken7J6jQ1Rv3JCBro7saBAueN0P1tTPqmHDXnt8dB/huObWCSUmpVWOltnTLBGTHbPs04W1FK
G0XgY1hahATNTRmWWmL68SPu9cLUPKIAOBEAqL8yptwOjaAKvExHYI/mg+nRsj26cE79NctcEDDO
aKfq/e/PFsGcCJLWL1ml7JoWCBtOXXfPLPykOVaBgdJB9Rfyc6NnrWXe+BFN4eaDaLvEWN2jCv/a
ubpRP+2Z/4RyzWCPTIUow2+JaddGmNKz9mNFObfjq9ErfLMsU0VzOypcHdEw9DSKijKtZ7YLKgvb
bdXWZGgiiKI+9YkN0EpNM6MYtHyL9Tw0Jw7WG9vVmRiO6sBOVc4aqp34BgFYJbesTPY0AqiQxGrv
u3U7FXBYG7CB+IMg67ZSpwq4KqTWSxLOz2NcNgICucILyDAvP5Y0DAChLUSrOJ0Is1zdY2XYilCO
iP/hYJexzSqIxQS28ELBfD8cCk7LiB1tnqGdYhk4R1cn6jdFSBOW7FuQMRITvapGh5bgFjsyeHvs
g+fVA/VK0kIgWNYtz0aGr3fnhVV+CLn74lB36to8K5PvQZHTXpMAY22/n3faeYMlTGNbsne9avzP
aE9gCOWiyUUnUBCNHxnLkn2JFQJ87NInX42IEVRdcbi0Tz/+L/sCAnxBoRVaIdGcXH1RzM6RQQ/i
yY80HKTEosscj59uUvuLr4aE0EHf7GVZGpx1GhO+TgeLUAWVa8OKREp6072UTk0kzfF2A1j9LvRf
QGv7VGYdblSXF1ekrTJ4PNcGhzKpriXUecgfoOOdITE4dNZnl2SxVXbG3aHluj2xStN8bvJcs881
FYIkZzB3wvNAbt9r2UZNt3UCDJa72z3U3hqY9DB5nIhc0a36Cpl4WmCNbaJlMM31Qd+4eECEiQNo
k8xFtUZ5z5dq9reDWkHyQ243dqSpndWWDvJzrYDRPLF3FwawZlheWpAJOPWmU8EYPOiY4ALKiGnE
VAjdG6wny/u76Fb3HveFhZgnQizji1x2NVwkKNS5AqwGFh3B/aTkr6RuAxJKCvI9AwUw7AQfxTbJ
5drpmtcaalASZaS1zu7jzWAfMB3RQvG5xopN/Vj4/qc77VAypvgAa/Z9eYgKiAeVGk4N28uRnKpK
chg/c9T3ii/uObzdfg2GxzwHkBEVRFFhAlXeJj8IVW47THMSo/yImg/OL1bi+NimTHXZpQwFy2vW
1yqr7Odg2BdnRmfUtSO1xoVM0eTwKJ5m4TivoM0WpWT126rgcZPdzdRCjIAGdZqfsO5fAlRT30gz
QZHD15i8IRKV3mBpMaQ861uLY5KNCKicqoyKyIEx68GlCRf4b/lkmtNxa4aXWvCIJMC/lOv6ms+A
JWrMyFl4WGhg6WCVMzBJfafGvI0UZSxRDQ7vRa6A58deu8Wp4YJn4whk6iCRa4F46h7XnHfCsLx6
V6OAs3BhglhpEmFWzS5pJ5M6DHcivkn4zZi5LexvJs2elLKOyT51TcOKxWN4NsqsYMxTC+BKjJqM
S6vID8Qd3VjBCTkJqgMv9uIJ3CyClEUR5k8mwA+2+KfYl2xEMKqNlz6qkNk6O3qbic9zkQZU5C/Y
SgUV19SReEJ0AYZkaOZ5Gi2/yAZW6ZtucqM1kC14JJyO1X7bemaWangZe2TomIfcVqs35KgCYspk
Ecz8snlNkx3NL2UkN5Iqq4cSk8aESGnBZ9kkkO4AhJ9txLvJ+sArXpMvuczp9jx4o7Pi/vEk0ijp
tEDMw06PBlEuUK9eXrScqtIOMnZMWPuS8cVrvlUydfe7MckR+dIEmGNoTfofT9sA4jL2CbbmiWuO
4inkb9uANdNUwlpfnhlZwOfIP6Nxw4b6oIKpYxFhdQc56igtKCscaCnpOMOWPciq37yT/YfbNZL7
PaR+CQtPU6c/Gc8Coqz1v4n2GEK3sSX3iHmZ7TFOVWGFl6giV2D/CNKQJFkkRu5V3mBtfPexqR6c
Wl5yhokLuxndDlw9Q/NqVt1xbw7LIEbgCwOcdoZZ9qbCosx5DkMG1BJqxiCtkshgyL+G4Z+sfejN
aBfK+WWVzfYOUz+jqC7pWnvXAijbk5EJrkz79RgWr6VqNrtFg0y2+CkxcmDahKgf/qNal98msyKn
T49+2k4hH3ZItpIbjzrQ7+4hEISu+lvsctyXn+gzjYMWhrXXzbLcvbMZAbJOCWvZB/opI0sXzRGB
t2YDqTVb6JUJMOcgILEOA333NbS9bkjs2A/Ogyzppa+FYKwJMHxgbBtulDtmhofRLh1ld1WkfSul
ECDODYvn4wjzHlrdKSJc8BOq16lfJnsNDr0wrbQbLYnbvM6U4BtA39QN4W0zRFv1fYIik+A+WNCA
lpuy+bnxLOg5v2ru/LFju7dq9uUbVImTPsvWoM/9EW4BokVYUJxikaAg62PmgWQEA87z825ybbVy
3WthcffEEBf3QMOF2TeLdgJ3umYeOe+ildKpC1hlqJr00yEGsgIsjvS0i4OMG+yoC9yOzzdWHSBV
XdUDrq/6ZRnfR+8F9hb/pzWEVR0+2K5L4MqmbZrAPP3im0iE4MrakfpuqmtBQLtHdf9HPaRjHwvq
XTSMUOFZArhS6mg6XpPFWq/YM8vTxvrblbzMHhJg2mUEGL1tKY3sQoM7oGtfja7zCq9OEIPmHnkd
ngUiy/djDa6TIAVliNi59LOulX9jkJDbK96T4OdLweTtSIwOTQ3BBoT2CjbhCva+eO/18z3ROtAM
cuWlOO/RGcUmQYnItu+Nhw8iiPMBDZx0Bc25p2XbzNn+ujO5tkgYCST5138L8HqI9zur62K+17A3
lTDeHprA65rAaquqMUu4BW4E+9ALzDk7VKc4GPgtrsZMTzhmPESdv9sWrxbih5fEEAE8IYeiNjmJ
maTPGXmpubOBuYODf1MoVMA1xGg7zA28iq8xXvGXzmzK91ySwGGDRownjlGfxWz0eobTnl9wpAmM
ucinAe62UscCmpMmNHcKxK0eZQi6guRSL/W1noHXLyNnJJqko6iu4ChmI4m2y2auuyfs+wbDlmWp
Ol542KeUOe3Rg/UGx2jIQk6YLY72eAlmvTXsInrmTjnwzT1uPB4sjkIx0TtOXWIoWzsWUS9OsJrZ
/aq9HHiXm8x9vwUhMUrtAjnPHaZDcvhJ3iYDCNy0O/AjggtuPCI+Ws8u5pE6aV+tX50eaYtSscR1
oxmotxDKgj26GVFA1KvS3t3TajgrHOUHueIIX72DDOo2+eq8/MsVkZ0tL4/9USmaNEgYuSaft0cV
AxLtzv/mOdXW1AQmi6VHTVZcoBboegZtWXnTuYZJO7BgcVWUjXrFrka8aHJ7E6j7zT9lExrbPfPW
ZLSTFTaEodM/5IVVVw+MdGal01D41r94hSW9hG/PdBXbV4iHQ/Q7wVA18dcDi+bJRS/Wwz2CvGah
QTKuzSIGkj7fr14Ly8wqHEEP5fcxTTMLXTJSkh/YYD1VuwPhUsY6aDjkgk2up6Hh6Fn2eGGPlhPE
JRdbIrLBnZVxZeHlfvyom10En8O2secKLjSPFJ7kH5bpBc+n5e+Y+pBnW8RCcIHo5+Gnfh8CePge
PGYvfyMhXCJHIkCdQ3RroINkf+wbGrZSgiX9ie+ue+5BTikNLecR179CA1zZVirfx+sTQC/G6edA
8sLssQUaOcBIqn/AEoeHJC/QsQo9lJx4l3cwOWJDcaYFXgtEWbsJLd29cyzZGFn4HSzqVU58X4s3
Pl9zIFFtMK/5i0QsYjQUAlvDmn7QTToj9qW66qEba/eq7Ags0Dhd5/j8oIB5gyyDJTG5yd1qyJAG
OGVDIOkBUXV3+5X2KIAI6x7r5atnQJjqp6FDvilqC8kRyPeDZj2+XOA28WIG9995TM+rQmNbe79f
1uEX0qIsviZFeZ3xNlFhA7jzMHxdJZyceMfB4Y6Zt9nYZMm/xaL7uBDPuFl6wjeHWSN9HhSOeumG
zCKPbS3R8PpUK1LjSYv+NVxKMdDHt8PyLJCkh9XLYGS1RyVdXIM8g+9emw6Ychx/jc21A/Pv69wK
M3bKYXV2hh7v+KfHFp3bmtM6XVcCGEBaU1+0G3fxTNrduOdKna9NVCsoQ5R+fDK7v7yh0eUhc1Fl
/XQvI+2+xbXtb1RY4fY2yS3cF4TVfC4A7r4FqciaGFWOp1QLoC4o7Z8TlyMAKLFT1cx/7pYKVQKg
Lo9fjgVyqHJO0yCwhGWabP0zjpEtvejtgsR/n1RauhKEpXCLMrPigfbfJkVgYxv3WVYnH1lmZzHp
HQ9A9Re1lYy1ewKgMlzw1ukI/cdrUpEMAAI5w+FL301YDlVW1c+pPcYApVF1Gbp4828/XVxUajRe
+2VF2j1vokQVRa09sUuwsYixUo48dnvzaslgu5nq5XiW4pnqp+OL1AGYIoOPr9lzGpYxhydt8G7+
5qfmz7sWBfdYoMfiXeeEzPE9uEMMaR15rQSq/FHVcRpPkKODfTGTCBr7lLC1xXsZm1a4tDs3BKPL
Ljyf1201k02RUyAp5pg+7xr6AEIOb5yXUj+4qN8BJ39hDnFInBzvFcVKlGZiWmEYdHKkq4nAKic3
C/5oSRKQ48IxWFVoyd38cPrfQNghzyYRSMzNYtSTuLSorVHw0KB2liU4G5o7zkFjA+xkzJC67tZO
kEx0Y3kJUExP4nlJjWo6IeT0MvFE/HGarZN4IM4Ho+M3KOu4ZSNaRAUyvYYvEj8MK667bK6bRq23
/W/1I5puuSwpHyPvUlrx4I5kU1RXkLYqcQ1fhyvnLpEZdfu8JFtm4aBS2Zv3ETdbW8Kf7Ji7trRm
p41X2psaPaoQdXlWoekeqzZ+ZYU7m2pxjaGczGglczScuKCrjKy6bVkdQY38ehrbDrGxNYY1wgM6
sgbFY7s9Qv/gfp6+PTpumfQkKzoMeRYPfw+8o2xXHSRsHLHYUuBT9P2AFdw9/zQhcb3GZOhdDYU1
7x6b9e/q4bkUX3M+5i76oUzPBOHEWvQSwMe2hLYl4dxiA/WKAsln66+XCaEfYsrGRs914veHl5Qm
Zjkgw+RaEJTU9BpAo8n7jxMQ1DF9A/SQg0+TqxOmqNKJrZAlGeiL3b1PyNH0HejQa0bNLxoRE9sQ
+51KvVGfTBVbzNj9YMUQ2NMYZYTOQOkraevDQILN1pYJSs9ywU8Q4wGbhwePHITmrH05z/MUBeV5
jOGsyof9GCC4y/ft3pR6or0mYiXPcSw/pbX4eoW62kgU8YvPl9Zs+Wom0Wpem4xZbG1+1YphKSiN
+3qJAwQTp1aqQgdEii3miCfjWsCx6ljEchEwfXgRroEeaSvt0cjcPoX8FE9r0DUOp1/KmH7ExTND
2bA3W7L+xJZFl1F5U8lkYD0lExEFHjxnj8cx3gExWmaWKntwwDV2ZR/c9pwNTCYJjoF25l3rYH5Y
myL8QsKNxkGl9QEtVBca4GQoESGBqSypcRhinDYwQGbWxiyB6QUBjThSA9VLsftH54eNnyDY4zL2
6NZE8IbJv8FvMn5gjjcb1/I67AKfyc8ZVcPlHX1nomLmstYFF39ETwbpIE3Y0ovZlLWR5vKZIWM3
5Bc62/sxdEIcs7eBtcd3NAPePbZpsdtAgEc8nhWEwd/et5rEWgdrt5el29vGUWtIKNq1V6bRZgZD
xa1u3IQ6rXWT+IPayDOogYHeI3FTBeOVn0CX7NABk9XMOTwK6XPp8B7+ygWPbkA8RGcEoexS+1KH
ICe/yae/HHyutISlhf03lrPDzB5Zy3jGyUdWxiXZaJaYYmv6ZaiaSMRvpRj3CrtoI6nYvGubG2GK
l+DhDCIKXlnhv9v4v9KtjB2kxzPtIyUaqKLaPbzQX24OZXBzbytNHOUtIp9w7dNanxap646Iknbi
ZSj9XrLSqdBNn7R36lpIwo6lJb33+mmt8UdYl4zh/n/r23yWeCdbKe209FhTdc2oRuWh7jp55SrC
s8F6LR2boLtppSoOohnIlFLEU7TirZevn/jWRdu99KcVgXDEVcsw3uLxuZRK2xAHeHXmafHY8Kp/
pEYTanv+muZnCa5qTqLHqMbhBXdy8mWjYoeAnk9IWO09rHRzsJ/CQubwWDdnBUCnhZsJsZOjtiyP
7TLwtC37AKO00lkDTftnqwB+VDpQEPKSXuyTe77bHI8Xkq11umonCumoEnX/jlSNga6Yzy/8GScD
enJ6eWtiw99UlAvLYfjSPF3yn2Fq5uicVOVaIsv+H2F0Wg8k0CqUxvhP+2WZaNpCMXywn93XeUNR
x1nIuXqiMcT0UJBh5xUimJgKIPw8jiiFIvqtp+WjQPJNkmVBv68UMGfy3qbnx58Py/8NSw5ngKTS
uI6c87ft+I/rp9bfgGtEt3FK8igTJNrg6bu+vK7QJW0uhnE+6W5Kei4d2hUR+0JrLABkGCLg2XZD
fZ3hBt0pSsknkE4eoqo0iiaUxjLqlyXVM9eJLKYjn1iEdY7OKCnGr9HSh4biVogrjX1BSkX4mC6l
AzbjZyF3aAHSZ9oToAliWpG0RRQeczFADW8UD3jTGTppj8MVxpAOWYFDILFa5oA51xCn/jUP7CKQ
+/U8LY9Owx6PbOPm+y+pB9MDEZ8QiZfFo+vV1qcn3KWDDXLgNVhcwI495EgSqyyNWYFk8ukUr55Z
uwxTbTygOsEBM/qEZ1VPhvMBOO8oSw9oLQSFsKYpeLE4rLlTya0CcPmBWSOu4C/66Oo9jIstgimK
9t6eOYXylDW0JULyuXn9ptuJXIoOTpZlxbvYQcmnGKO/6sey2Jsi5scpLFx04E7kmSphOHEaorid
gQ7NQUWJI58XDYhKVe6khd7K+z0wzSC7uy4Nu6Q6TClOaSRSi2s1kB38aGXVhlP8AsNW+jRGLTDW
fcIr5SbIMj3heou6KvSVLabh3SzbDcN4NlX9FFsxU2Jg1Jz7ijblNJf7DFij+DV1skTzfCf1tuls
2kaUgWq89CD0QTwA6scPM3W/s8F9fJ5a1q89HzSvPK81eYe8w+v3j0lIV6Fa7DY9d73GrOHMBshP
fhWHbnz7+xMFn5gpBns4ueiHaNReXnN3vRQYhoOJEhWGxZ2EKvk4Ncv3ZsKexDWy/RsGUKfYsjTE
vo77FYRyuS74yZdBYAP1JaVSSetAa1COCnAbgJMCkGlU0/sQKhob3HSWILV6o0y7+29kEK2lEf8W
mpC98gTqKH0cnYQaz7z6Id2kdMarE4w9WYj7x/7XdaHAKx8GbzGSgNyn79QAjU196omSC30p1LWH
wVe5icH7pk9i+cxw+ztL1aYOCZoEBkKmKpLqJ2ykZWBrgnImfg7kjpZLF5Ec4htiyAIyN6mV08at
lLaKW3N9V6wYZJv5olWBmhyjDCO5153CPsdpQqvevseZhsa9BFA+GF5XqunQnT+Cah4gAmWbAvZ5
qZfSLTlPFrE9XZRT6r87i6Im7pfSdGO7Enn/jrAGFndHY/FhDDiQBzPaJkHs0/9+qzN0a+nV/ADw
xbdusKmAyQR1r/Ei1lzW2EHImrRUG3ffGEQp97jF4MjtR6oT1piUWh9ZCA76oQwwqcYdhEd8ADHr
pbE0z99G51lp4rUVklGVJH9QZ4LBDGsbueBEOskvOdKVh3OzwQtn7IkRSkkN5RJtfTKi0R8QoIDC
qf9yC1e5k6plZj3nqTU5t9mJsDR8lhQVl1QSf9YH/718K6ot3P164UGQ8O8jyGqbUB3VTbtTqm9q
2G1lQAMFAoRKHz2Ga51jj7pMLenxVJODl7L+ETvHuokQgYP5ZN5sIjS8LVq9vv26aeDFhjUKx8I8
cEp4+9jjlyhl1U42U9TIf+SdfIjLjiTSZPJF1X/MtxMLBFxhYsMoUzziv8n38zI1SJvTfGPYTmXq
bgYj3GOB3U9OQfm9F8+Tup97njYFGw/P+whBdPipNUX4BO0Ind0ThT5SP+chH5kf6BVAS9klfNuj
TtECp72y7qZ/hWhN5J2DU+D4oFyiNlGfhmd87RwwLrAYr7DY6sS4sPZLxq8YmLQg3TNsMgY0JBz8
Z/JDGJq6dWU66wRuT5ykdT4VDADkldnDanw7CqcM5dEDgb5+H7yIBnAi2uuMlofvje3uBUMJ+V88
ykt86NB6sSwjACESKeuiub70psw/3+Z1PXteSkq+iwgvJXL2/IG+3wpuoJCgqn1lOBbr8P85lF+K
LCpAamYKSDGAgE+Fi3DP9j2jZsiNgx0gRPhlOGYDrbkCJaxmC5j36/ClTTtVdR/7QpafJnBCgLb8
tUXJogBVd7NpAQ8xpZyw2WwAZih3rrC5J4+WcV6rDeETCe9rSZJMe1/1RYWr4JQ2RkXmoY4lHTVZ
MKeRkRTFHMtrPCdNEaPPQh/USiECbQitTjOJ/zLgPAv4/KO4OsGDhm5rFRQRJKSrmD5gkbvgU/zw
3cfOmU1TynRKkMLccct2f2a3OYXpIFKnBT8tkgFnHB8eH1htDwmwFWe1HOSrwjDehW67YzqcDsc2
u8RRxpM5z34X4be1Sab992LFe9ZNpKOa6kevbOuqKoQMBanU4RLC1AOK9e4WNj7TGpQpZp8r1Ucf
s01w0hDVIkDi9J/CACpctY7BU0tYb22oqim7x0MMGtgtfZ8qlFxJgGSAhOWRCPv1GlCnUZrNb8z9
cwAY1nytmhG9NKodqRPR4/B4cZh+3VZeQNBk/aaTzHBkLTYRcYcF+x0pi2WeNjfnWv7lhTwrAbF+
0rBuBxXLj36mpdP2827kPYVjKfMXNrZYLTXZOlthR6e1EHQoc/pRdgAmTqy7k4rCZyHt4z7v3Q94
M2fIWmkOPd3ITmMkAs2mIflrsqsvzBxWFa6hYuQfig6A8bzi/yP/2UET60U7Nu1q/tXWhApJawTD
Eg1IGnVy0OnEpCZELeeciMTxBQXVYD0FjLNJkHNNVfYp7wDI08SAwEycxBHj8sS2jEbqnSxdXkvs
lDGKJm8mQllfRddkX9mseVkiQd6kHJzG+ZvrhBN7RpfLFQJ0265FAon2gA1nY5uhjLyCuzR+ara4
+Ey/YXSMBbM+M180f0SgIMdzrjK3+lYceUEGYrhQ328Nc2W8z1wfD7nAKaB5js83KMcKyOFPDAN+
ChwfYi6RJhOb2Sp6nwzRDmIA+U8Y2dhdCPOHA+gxVJXU44UxnmWXLS1i7ZhzUXEY1IrlBz3DR0n1
H+6+CM/96+dRkqPybSvNhJYacHsvMrMKeJXR4uaPL2OD937f4isU5ZvMnDleOJekhVPdetIC7Deq
EZ+TgoxBXcBPSZMcEeHMv7RnY38UQ7cAOdT8jzvPKZXaoxoMVmw46iDWPzRnio1r8/PQMHtg2gfG
dCrxbLUqakkFh0frn5/l4uv33n7X3dT+/+xyJ9ubdWGhx2xlfsw0yHzRYjI2JGlQmEcNjQQDnlG8
gm9a0vHBXRbL8AQxXrs4OAzwPg39tNK9wLmal6P017Pe8+i/xgmbN6ft9PBLSn4blBXdM0x+d6vw
m5SKXBv7Kqj0yFC/MYYl0DQtJQq0t2Wl/Hjaq3yrFEh4ft1ea/8uOPh1PocatysQTV5Dogq1xjaO
tOaDx89coq83v2YMni1TQ5eZcPujDl6HFq/XBwHJenGgZIAHlmFFXHyaNHnYilx18/p6JimpPHd0
hcXEiEh1hevDU0rc9pdl4n7EwCGHbzK1ssI8tICZW0v7X/5xSeln8aNDxYRVGBijBXzzNMVJZzaV
Q7XfboLpf2FbrfQKfcSP/oQP93m+gBDFkAvXdIvdHOkLiCthkjfwgOLH73jSo1AeM3CPoVRMK/Tk
mrnM4BMCHwjidTA8pzNeXkz/nqLR4Iu9DPP2VSDg5mQfrkxSm1Fv1P57tF1uNnr8ezZQRh1B0dhY
mOKyMkRv0I2xeZUebGB5B6l3USrOdpJNXMjyAjbq4VA/vm0gI81c7WKP8iWIGjQncvmjzUGanlrF
ss6klki5msAs/tiGtTE/zHyAPdb7wi0NWva7eNmnCrSgx6aO7RPzlce0EcwtXdvqozgwd6hQfi0d
7zM8Z9aVnMEjkE8OqSCRVB8xCNH5tzxAA2Pm0L2hODkY59McsQRzSkW95HB4jhdN89Q58Dxh9+Sr
93Z4eHvBfD7bPhyBJ4HpH6jGtOo3BMlUp9/Ywcgp/pLPVHsGBGIyStBjzUNohhxsdL3J0A9Ff8TT
jKK2A8/4vlKrHJUudmRH3sZNkq1f8E53HUbyEsKsgDKbIfsdzgbTIoHQm9xlVftIUuuupS5J2GW3
oJQQJzX6Xrv/jII9vNrrIHriLRUUySdg3gtWOz0wdZL0QPwi/RBDuz9aDcuXdPQG5Dme7enPpYsO
lm3I2OSNGpmpWJqC89fQZLeMa+Npg9XoqO0MecD9UPlWKS7Cjq42dRHhj3nwYzvhP3dNjIfp9Wq8
laLj7+29e5JT2GYjDp6T5SVvyp11Dtn94bM1jgxosJq9rsMDZyhw9n6YnUzO4SC2gI5UPT1+GZjh
lJKtThGEvMx1KKmjMKaORiNBiVX5pkc4Om6iIjNpCMddpZ/dbYFF6h9cn0N5Kd0IIohHc49DM+QL
rgzJ8qAYQwJJrtKGqau2nCyD+Ry705oL8Kin6ijU1dAMEe9lAWd/FjdfOR5BIxMQ0DZF8++Sg4E6
HKJKLBGdTPIQkZX4+Ymkx/89gm1YXxzhNU9RJMuSfw4BxKuwlaeGQ4zkWQJ57lzBsX2amYlKYWdg
cRA9avmuoNFWfR1qeFjgkaCFqIaXgNciGEn/LSP01ynzmCGGgsjeITUhLnz9PuAN4/7cqy58mb4m
LldVfkEtQ14GVXS7rwBYoRDrLVCTi5YJ629R8/kOSgFZdHyMKShT+9MyueB6Z6C03rLk5aJz1WrG
aaEr/9aYz7IIU61I2EdxpeGNKH9kp1w4gOnni1MIqGfuuIpqJHX4bwnJYWQToxtEqkQuhTv6ZEGE
dFzhh3ZSbXLnFTt966Gmj9gCiJXQCHJE15o5QStjkog4vMfVAUf34enc4proBiUxB8cS9NN8gun+
AmV4KVpu3pPKjSvqpE7Acmwm1Pxj2J6rIqujk/tI6nko4TF7wcpPI3JAlBCSVy3t0IVybzpcvmSb
wwqScEjsjWQim5Fk7yi7DHht5cBwqiUvsSptu2fobXrKUpJ7pGNO+zq9wli84rDQHj56ZAVlrciQ
OFhi6QcBuxiYiGYCnZzjsoO9aw4hVUqO6OWz4mvldg4zToEc6B/mOlY6Qqw0UPkYhtJrZ9eesqCs
RHgwR/9FqWPc5fBf2HOR8mBcHBhtfTmKRDsXbnixrYCnhsWO6Gk+DfOpxOMJnzyFducXoIwh+dbm
aO+WmRRdRPw954F2DOwIosZ1DU8xiZs0Y9we+AQcFQMXNQtIrRk/xElQCw2Da3nIUZiet/K1UBEr
EspmlpgVAIWAR2FF2gtnsIP91JCtLrIzfvRZRHMjHet0DT21X+c0RgKF6VVUMx2O9HYXf79B6a+7
VY3IiPvVFb55/fG0ulk9MEGcZtLjRY5PI3RZcY21G1n2OX+va/Uh7TAbWypXmhpdsE+Z4Qtev2oR
yITR5sV09RuyfGlGYqPKK2yFlmiqdG6BnYyfV7mXVpGn3fdiIptg77r186xQHDig0reTzDbPm+bc
YWf8RjLola6/1SUQHrkujsQaSRBCXHzJDjZGy55z7qxLyZjMxyYZ/asCyc9H+q7MLcWXhyMvvORk
IWci4EsXUn/iokhVA9FIERdBBQbIAr2zGFvDPtxWUt7AYNoXFgg+SpSdr/Whhp6qPPEXQ/2b0572
L3E1jLSS/lt1gPWT0FjNmC5C0Bb9q3i1ULuwHmh9OYwD7tpxjxww6WPGBmKTRyMfbBu/j9U4KAWD
ZcdcqENq3kvEL+fP5yCUMEn+RGeCTVtcZXMyrZhIxLdG4Dl7STwBA8iUe2JW48UNVExzrzSzUjsV
IJVmGalhF5hbOCttSPBh7kL7iicDIx5kof+6Oxv7H3HDp+hMPiRX++FbnYj/FUO3ItDvRQkMWRls
CotGEvCjYcs5U99u+ryqQeyT5c5Jb9Z95KaBiHsyWWaAvKOrLbD9QkDy+Kt2dsVTydr/5xCqPXpB
1S0X0cRlNJAx/ku0CQqaI74oZv21/T2XHB/HffgYzj00VS7y3mkZi6aPTS4kaayGXEVbcRsTrQtX
WQQ5edoIsVelDK2zsAoUzvbGxZ4pVykzyFZsm8MA7MZ8urBWUfE79OaV6hkGNQMYszn9riWH/lcj
NIOj2qffKUP1/4XSuTkKUgHW+gUGxkWrNmJT9HTe3jcB0BBjjq1aQfTLM2FG5Zos6UQzHQiGmc9R
Bl53/0FZq+fLhjcZ+DDJ8/TnHBe44QUaLLMtlCvVGZI2L5FEpDkDbxyGmzRnth3lLdSkrDt7Xv3D
AhHNX8DVuG+fALbxoOFSQ2ASbptSYkIFXrygUUpS25kk7cU2wP6Oy1Uw41eX250Womfz2RCXq34m
EZVYfjVeazCRPowt70pQVgLOkCcLo53K77LpRL6pDwZYlyGAflgC1o0Ac63MshPKAVnVV3HFvewM
ORWXnMkVrADYJHHH1jYEh1UvL/RLd4lrp8QRywfOaohGlNO3vyfvoHG5Tj9XGoiet2BCX91Wl85I
w9TYYeEGQ2EWvspPoIIAHElnp+BUSQdmo+ZZv3XPzirSvRWTl+PM0iIRXq9HoQscABBY6l5a3/jG
qidZUrbRhsJ4fjM5dOF3e6Sdum+O/fizDvbAJKU5gwmlaWHTX/AE3Tgj08qUQdueYs7Cg5s7Vsy4
Rf2xlnauIIHSDyao/VKwzOLwv4QOe3nAZpLPQhfNEz8V6Pt63cu5WlPsP5kzBGpf4823xRkUBrcc
TwfdVTb6I+3wbYBS/zVtERofQUdtuyo5V/eceIU0zYWWokjPhoHb1HBdD0S342rQ4z/ypgbw8Fg4
rAzuQAnmj6UkPxMcnuMadNHOAX6mYVeNtkAEz5fCQbPhiW5VKUGu84lgIy7eoh4C9BH/RMvR5WZC
BSpd4Kro9jzAOTw+gAC7rwTHnLmKriYOv4SJMrVjMI1P9oaqk1dCdVBLvAZmUf9oFQnVz72pM0GB
22xQmgEr80mTL4qL+YYVJ2dNkk+0221gTfHa//H8lgW+yuYvhgjepd59yvQ+pOHVvOdDD2A9PMKd
RdZ+sZWNO4ReqyfyMTwp47V9ebixKmI9tpdye1RAIM3PAqFek4NH1HnIPV0mq5+YckHnmPlBc8Q1
JPKWh+t9wIkIQARYbMBWA+YvYabH4NvP/pf1ZTtblYj2PPhxqFmxb3BIs9IY8j56YmcmEyQN5pKt
qPgnJn0RdHm+2NC/qLzfshiiyKf2YsnUTDBseyy3auxiD412D2LPlh3Fyj/K2WyPh0PpIIaaRH/v
238RxoYsX4AJZKw6EKw+Sr1VZyEbq+2joQ+OFubEPuC7u7GbJgclDH2KtP1fZNIVi/+QYzgONGfp
9txw+6UonCZQ09h8U8LnpNRnPTkUflbNWa/xxVLBFj5KZuUVsfM410M1joE91SR/45HkkLCRHk3t
DPSG+b7g8+I/Lwwp2i35lqI7j+gjpV4OMm+NJu4JZThtrfSHbbkFxbHY2DeWB7tu8RzvMiVaFOaV
r29RWjJ5zz9jSOQng6ueKHPnQm6Y79XJcKTfztHreX9iC7Q069IxZOXvvRFoHjoHO54xfhzja7xj
XEGcJGMjDxmp0kDaZy1BSyKIk+GAqLzq81rsqHsf9oYH/MfUn60q4BHWX5v9PxkDv/uCrdFRqXoz
8VpKxGj7aeo25ZA611d4/KpuP7evCmO+Oz/iZV3U1aA6N38w13gSRaUWlzaqlks6t8yPhOEO34Cy
xkiRgERe4AZtC1m+cSXEDDmPC4tAiohAQlR/VlQkvD35JZX1lj/Tc8b94DpGOiISa6Wz2Qg0IqWT
XflAVcgtrhrn6aaJPVx4Udhu+fJtNl/GWd5N84MQcnO1u3KPGVicnZMgFuYA6HTAt12fGXKiKCCy
0N13j13aichQrB6EkwNJFGSverhHs2KpkmY4WBdiTB9ZbQXC0KpAHGKxTRf+aKgdlE60Ngom2tNR
+sr7EavqXwGPNiV0A7lFc71m3svux4D7I+HHHnVg7EPMUBz9Vcu+PYZ8C7zFAWbsICEZ6/WKiQ/+
SnBpVpXhMficNNKnguyaZqsDfjPWI0JO1iFj/k+hHfJyLTnzixNhufLDcW2x5Zfbn5Epg3dq9Qh0
C5hweRy2jCm025M/XlIovfcnd8hArDjWIfOczOF5e1xWlR6BHQLU4vZnsB1tHFqJmCTqw8s1q1U5
cH81AOtf4RfJm8/9c/5pVvxeyFfPh/uSlwrIlBODEHF0DyXKn2cV4qFT3eWajFo9uPO9xiHF4/eq
EOhCUzcxr9afaI/HZIbx+ZbypI5KuKfBOzalOwSco0q+Irl/mcEwakqdHI2oA3fMd89sP2Q6Gxdo
TjaQQgw77unrkkdSCZVWOmOe7r135ZLVPvvQTSAeXtKWyoyWQPAaemY/q/tKzbg54FW0T4Y2+XRj
8bTYXbJNt5v46EpI8kHTSn8SNDaGprtVpnTm7YWWlsYLi2Bf9DzhOs6J5GC7dkvQ4szqegbLPMpe
jOeLT6flbAgDlhTnOvh8oRzQnn5J1m3glQejpsbG+Qz4RkYNhVJadVa3CYHbkpe0/pywbDYplle3
NsfmnVzgWML3Wdbw7Q/Yrpmy0k6v34gFUB85J+NZ6ctlikmeGDegK25t/CyzJMBA3OOxTSbGeYng
n6H+d/RvpKewekO3MSDOy7wXKD/ix4cCKOHnFED4yy8OOrlvc+9WfvHbODHJdujzTN44Ks4UqxNo
SSS4JuKPW2oLOy6008xDtpczrhW1XsM7cI9MfNjhYuryN3jXl33GmSzQhNR6PNHRqDC4ySXSw+xR
TvGafeT7CPzEfO0fyVD87D2SkfCIHi/WQpeRCdgVZmCi6Vhta/jZq3qeglVKBA3bKxRMHfr8ialH
Fkf6MFmXAPOMN7if/BZsAZ2soGuVOKMv9DCqZ5easgfGPqwnDD4FyGf1OJINywqw8puV3PP/A0JA
+Vbv6Xyzmz5olRxKAce3KMbkQ8x5MbyY1kvOW+THSsQTCe7+krKp86u7fwI25XciHohjO785ysEi
jU/Qhq4ASG/1lgeRuIDV3z0iot8GJ+d+doFhDBxgwhqAEssNzT60xBfZhRlOk3eYxsTt0lT2bF4n
YsgHiYKBufKdpYvDxRWcZ9YgmcvoF5KPiBVMpFup0Nfrev1Q7NkvN4vZ+nEyWI/zXFlr7HnkLzEf
Bj7k/159cba6mPtnkC7x3QONG0rm6HKwLmv+12qeQX2KaXxpvTCv5+u7ledb7di+UPFf8BCta/FR
Q7DPcfrI95pxgW0hMmupENymuBHie8vr1NrA3GusIw1lq15mndUO/01AWGJ7hg9SKbwpfKxoLkA7
yBjsvjYHj8bfnK6OIblp5i03hlLKngc9IM03wNn8ooyiaNsUr3a5GJvPyEBbUu6dBIdsyesXSu0W
8hTZVf9bUut1+hATVNq+F5XF1n0/BdTpEeTakb7NtZTuZZL/A6QaWjd6xzaJHJp7ZXyIa5FFTBSA
lDWNKM5ozk5BwRIFbjKptrxyQFAisKmuPluOS/VweabS+N7zoZm9rsYS+L9OE4kcMSsRUMbt5G7V
A7mxRQy2y3s3qA7KGk6rupk3ma/l6rwbf/eeEUsx/h/ENbZI7N8ygFO0y2sR2mZbg/6OO4+x/74v
veKHS4c7Qfl5N8QlR2oQf76OuNJf8tJNfPHWRsGZOt9TR97BCIQIoIqtIKf6OsIEKOPUjmdaVZRN
WTb1Vn3HjpcoK2A/M5mQRa4EzTolVGPLFImO647RKCk7L/IF86rTj0DmboIO7OFs7GXW5zQK6Y5E
dNd3HZhBMXvnOSQKgwyneuaxdtuqNhTrnKrFUT1lpuax5NHB2kyvEUWgiQ+2w62HJ7CoIjv6QaMY
RBf7W+NtXOQXWF+nHaMEK6sn+D6GnF8mlU7zLwk8xWaGP66+l+GoS4R0l9HB2vb4HR716za6icMU
5+JYlbYFhCARQh3pZF+IyC0OA0U3rDjfEW59FCLoqvtVkS3J0RbegQ7WUwS+6d4MLlPd+KtO8Vpa
tj/1jtbPLLXA7U7BllbtQS/F9T8EH8ZId3XrwAk9zPY1gMf4Qa6LpRFHF5zEOwu39ALLDO7GeoDH
htCUPyaG8Jj1AE9GwhEuMRdFfm7CCiCWnDGoN6VruGgPrSuCIFBFIbytSIb3/ZXsWhoSEr+SR4xw
LdlT2BO7dyNFWNdQl7OGlfR8VRolsR63biw76qKHQykuwaZYkvVgXAOzkGZK0bi5oStYbJlb3uwt
8V6xuezOCWPYRRPePdaI2S0kdfjRBpJ0FZrkihZgE4UwSOM6WMT6/xbVdMkIVv9t+XfAZmc0KIDR
j34/R2DdTz8ni1DVfmv2LxM+z3qZqu6POiWmt22UMJBAxPErPtw51cdKF8oM3svX/uFL0+yf7yfW
kY5UgP8UKdJYYdO78S09DiaRAM6rodybXEA799jvJ7SGkuY6txhPn8wRDBdb/wp4++Yl27dkRVDt
y+t7Ivv/RkRXDhJ2mhTHm7ng95MiE5b7fZjhJMwt5pSofDFgtTAO1eU+3nR+2fKw6+MkCYBCZSee
f0LGZKOBkQYXnOCP2uqIydy0+PaKXw3VDP3IxI5cit4/LL7XT6QHosXP7NmP/r0F40atPUdAQa8r
hfXuOLuXZyQ8F7799bg6vSngzx3HaFFLt28VP0qTOx4YQo1C/RrIwJlfFfqyWp6QR5AFGWuSDnZ/
DEvttcfEgXQ7zGpGyPvcmEqOtGKUctc2drAEJAFkOB5luLJ7r6IJOlqlWQKBt/3luvHTUSR9Topz
tE2RfoQrA839XEmYUZpjM6VwGvEAEUkSSPJuiwR0toYm4cWfgnGEB2wsQU/W2bKwTX6CMJGWu9Vn
7P4nrzOjGoQXA9d6wSLBmEALh+yeGe1p84hgBUafqoVOQFH54hRvKRpcwV4Agb9yyzWG788Ru6B2
a1crCjdKLqtOmYhKrqU6Dkpa7V6Js3vRx+fsm2MeHoX4bcM/jimNuNtv4PkwBEXqCeDqVt1FplWL
c/N5UhwJOeEFBRvmahutEpA5gQxJQJYb9RSA5whRc1ZpXMkxGDf2GSpN3Vr7kdynUS5LmEjvVe2+
ZWWt95XSZrCT+WiYDA+wc6E9yrLlWGU1IbKz1F162ULyjwwcWynvCsCt1sh4sUzzIGTZCh9khAHr
oTOiIhOaLFDvjvVK+Dfgy1VlmENYp7heVAd7dEj8DbmVLIZoTuNQ0W4rxGWAupQKIUIRmhV5+nwi
eoLO8bA3zg7diFldfHHHBNfG+7RGvDXUfd+cuFapq7IaNtXkisn4T0SITJBeWOI5cvFDQ0n5GgTe
LGxyZjhiSr28qUOYk8AGsOZoLWW6Af1LU2F98eRtZxLv2tdQjJtppTKp31fe5/6rkugP/7wOKXPJ
mz26DkRQeoVnqLcKlGpcMt2xA+FBvPEBcBnx0e+lRUI3Wnn2jJTX1YTU9NtG0ijQtajsLntNC3iq
vfyhuvO/5O3jEm60dR6LUBytMk7UacMofZ4jwL2gq3DZLXi7vnl4eyeUja2zYf07D6pcCi9xpl44
G6KushDCFVbkkyDKa/+hJKAFYBjygQedK7qYELdTjred5KCCyNiSh7A9rc9OphczFCEvcona1PYX
aQ41Z2h/p64fGBZ+ktY1P0YFsVUg+d4HH38BZSVWiN7W71mkqJ1GGXjwk9y7hSI+TX1OvhO//+8h
KLczODnKB3ZzU6cRR5C3+QgEnRAKOtEYR8onnFGoZK8UjjHC8xY/wlGWEzYSxJ7K0XYT5T582frj
sbRAyI+s1uTQ9tfbrK1wsPpf4C4WUt9ua8qQjvJlBUkmLHqdOIG/of+taHY62bFsvSVU7UitpShy
mqHEFyP+l98piuDZ3VP+JR2psttqku3996FFgfwKm0vFJHWpNwFnxT9Ca4y8TXCRt2iGjhJO2gYB
XwXMuOKpytMimsi+YrZCDlMIsQ3JyMjYkRr5h+r2ozYT0ICBmskm3egVx/pk3WgWc5rcbirMw4Cy
ojKoPM9rQ4YMNesnGOFJqvJFfrIPXBOug7Oh2CJJRAnbm4p5nXbz9c7kQW7uw7A3KabJXVPGkWA9
yK8om/Vkof4m09O+L9BmYA0uksjmrVRkP+k0xQnw8xvVs0iZAh8Ff+DHp9m/YjEh8P9sff0yRLTx
LjMUJx3mku8nLiC+SJ6n2gxMDi51UhX/BEPBnPe8kk2KsNZ3nb+UulhsAC6dLAELr084qM36ArQp
gfmYBFVAnnik/jMGnK4eQcJhKha/N0ili/2mO573CItQsZiOrs+aPEPoq6EYiUTRZG/8x8HeHpl2
jyRSlQMPxpxe/KWe4GqNaoTuD/DvAgvlT+LpedbeiNUGidpsyRkTTgpGnSd8RHf7PulpYrN+y0bE
jnSytHIeLRZpmXF5PloSz7W/IN+UPVfxEkDRyV46du4xi92tOPZltW2g3V7j7axfPrh6Cl5aaUCo
FZ8JOS9rsJEtbD8zaGLgimUP1lRpDM7NeAhD5m98cwhH0oUhjqMsRoQK6K84vlpp+EObSFMqJ/9c
nWHh4hSkJBOlcSEgbQ+cAyb4ibFdg5/bLK28HhZp0/AKnWxQvQaVxT+twFzCx3SKRTJaZXdgUxXp
p9emYaq6VkWWk5n6RKyWB/fWfqPJwx1HEC7d5XqnrsRjdBmS+f7FSDzmiSlvJRnoQ792KOrg0ZMf
yw1qxx1nnqgGA5X1k888Ps7prKY1cqKfCGZlChZbedLgoBTfuGWgNpC7NCUCBYhnnK10jwA31Beo
m+/LaEeACCt3PazLth21lfQ3c7iEdIXDMyznKC0X7mZCK8xqwHnJYcuHIPloGoXdQgFbiHCsEUOU
W6VoBCDGPQwH3CZbOjDNSeXGNMjQ3YxN2kAQRNpj/KbZeu+tNCCntriIYpcK+wa29WOAYXaqKNQG
RRf8Nnag9BFP4HA9Ja0N9WPcGhnsbbmfy39ukCj0t5wiWJBgsjLIVZgAFCjw8/FLy8Wj6nlmHdKM
F3hz2Clul0FYxA8ZNEniywTYKE85FJUK2au3VIbhP7OlezDBW+gfxYwEThWGCAUuGmviH6yjtJnK
8PqPij6TQbnTgA3YoxyawIuwtdSfvEZi0ZFxOxT1rQA3AR2cA3EZ99NiBmxYHJ6dLywgJmJjY3h0
71GZplE1cX+6T9ceV2rGWEC/+z7LVjBYcCiiN5CXX04ZpWz2ztXbl4OrhKvrpytuAFWAYdFYF1/i
6DOb8D5qvQJXaTzkJhFSvH/o0j4F65tiR446hDyB73IJ2mN00NbbMgWOj+qMCghrWfhtDvNdPs/m
aXlaPCIyWUkz4MGVNy8ecUSGsVlKj0sfdM2PHFMVMGXFpsPk1bYk1hOiLZbz/64XjkjUQpujDvi8
rQczvtLbu/9hu8p3R3fUrlmGxZMG+9LLD5xNhgjQt3UwXUCMansAE2En2FbUXBNAGJhH2/TfmQR9
jQutLsuvxcESj9tBztIFes+2fa92PztVrqCukwe99kBYbvW3BeTBIw2USwVMTimdJLAnuQf4/TCX
NnIFvslXooLT6QrUPp1G6JvdUX8LtbE+kcsuaO18VCyx2H+NSYdyyRzkFggq/18/4SlIVLKT6o6j
0Z4PbUAdeKqkN8+oH1XO+DMzyd7J1h5q0TiircDF7+wF4oFv0Hq8wbu59rK1OiVOtAKSdyEbPjh9
9fusEIGhC6iNZ7/JomfspXD4xQ9AxQQQHoCM1VnQta2vwhPO3tlsLIiTe8zLDqW0l9YydkeW8zoe
duzy1S7o/1Kyu7Firrzdp/BrYumcWUcIRT+CAhi/Czhe6nkxshIc9STt8QypxR3NthU16lOBcHJe
ycgBWvJ4hr54IU6AIIO7UFGo4DJuV7MhJoy2mmmVdlQ8+Qe6258p0r7tFkLqApixJ9AMzrrSe6yJ
oOqIRoJf/W00nY1X+6Uw0PzZeo/FrRv5Upq43yu8DJKajRdyFgi5ORp6SPRE688PY2JAR6L/U1Pf
kmZTuwgaUNak7o6oQc8bqle54s1QSSyfAEPlWKOOOKm8gUFhgXDPE2VXHs6c8xh1Oh1IApZnj6fO
Y5giiQrzivkMM+gl0IEnIIQpB1nn7chZctZSKaFEjRKkXSQO7KhKExb015BpHl8sI2r3SyHwNtP9
95u2YblValXlyV4ilxVGo4l/mD1/9mZ86++W5mHK1+w18mmT+OQZwgekfKU1GE33SwYR6cPhBArG
kg98Jn5NsiBH1meIkWZndXOTyZ02JgY3V7mEMkE6Fc64UlDjHlJMJ/O+LTKSLGi1B69sLdJXioc6
hhLh2lrFMV88dD8Oz1qdHYQDvbpU2HdfmZoPWZ4iK/Gffp1R2j6Vy2xWfxYI2rvC5KREQQSRJ0xM
9fw/rh7pxEf8aHLi8psMKN/KQG4cqEETRk5w6MIuTVFU9/9bg2hAfjOZZSfyiFZuJtWEA1ICq/ao
bRvqvEWSwehjd72jH73d4wIsq8BAJqNj2yB43nWlS6X6RVAT3io6oZkQ29hJNmWuUnN1z8FMxT6D
6fo9PClhPbgvGjnwyXaYaKODyCAr7BjybBLlaOfvkHTWb26wbAPFtb6EOyp4XNzmkMTVeBPN6VlK
Ld3Uep++5msKkNNZA/vxuJWyKwRrjsC8ITRQR+K5ggMT7ZEviZ3QNSEPWJ+MBpXU2z++6cXhkjrr
dmuJGrXbTtjOyQ2cQ7mMKDZmQaJZj0X7xx9rQ5umY18t7ZGKv3NJDxaj10DM/od3CDAvMJvbHio7
VArce9eXd25ivF99De1Xn29MBEpTLqlNnLtRKVsAyuxgn88SALcUmHA4j3EoEOKTLCZj67LZckDK
QYTKGiA0urnWQ2ZfMqlvLR7XAZRgf/JT0XiTgDU7w5DSUn9jTvdzzwScN31xzqO26lsAYeoyeYKb
xpQQcojgatiVXNWUoQ6KZcMDZrBPnqMBCEZJPF79lc13NothhEZLwy55Wn9hb5lL6w6NHGFbhbvr
DY8UO/Bp+woS1Fy54Fouezsn+k2L5tVsL6R0kRdJ4nfdlL5Hbb6/w3tVXTxn92Heitz0NbV6TRyN
4w07VzZORrwEO2q89nyjtPnrpFtjWcLgUj4Jn+PopkkO4hIpdnYL28DpOdzte4H9/eWQ9gNcLLFB
SD/w0X+VRJKA10R8NbHfiJ9g3cmjbeAATWgxmoOQRwM6r2VCcyQrAz1hR2HwPmEdUXavnUEJR3ik
xdP+NbBVHSI822EkxQER7xxDBzVsTFN9+T/mmFNjt5AA0OtTLKyCYG8FMdXArr2ymCVMkbYL+9as
ATGdbLl0bEtEG/7DZ1NaDcp9/c2zQAQ0rRZv8rnURmfzFtJyjXRwYcyGPjrHpjhrzD2cSrwzdLLt
tIv/2gtFip5NwzQdqfli8ZqZqC2MClG/z7tc8XjyzSJ5bM/BhL2QziC1SH6Eda47cEZLflDm9eMr
IuhyletR5R1hN5um5ncVpOA+zFmeTjabYwPRlFNKlLrm21E9x9p4xcwqFItUwn4mIYVVhLc/d9lU
ng89YLMVJf66Qe5QtdPVkFMv0B+Yr6HcpNwPM5xpza4d7ltGO9vZKhrW4jAGDwIF+VGrVCXi6Kb0
0/w7ldmEXg9NiYaR2XW0Dy9zCuEIV+ejELJJ4Ed1aPfB/8csPo50PfnTC+6EU5lZ5ps+0VDWOTbE
plvL7Afw6UXRfu16LsF6l/+L63E0/578c3EQ5wK9Mb8lH+4FKAOMq9fR7LzyNhgEcA06ZD+wfDVE
pMzTKYaykyVB3ewFnzBqUHp2ThyMMqRgVFQv08NzCAGV65i9TL6/JIVtRNf6EhJ5HHu3OphaQxY4
NxMu3yxfiOkkWuD9/5+LlMBDxBOgbGrdvM0stTe5Mnmhm5CQZq6rp69zQJCSO+KowxqpRCuXtI+Z
SuYoaik4nGji6MCl/vCeUT6SoDsRneHNsVGtSp4zzLXYAZNNNlxZGfXc7BdSfIQWqmp5wJTStK2U
8oaqLAHLUj8xCvqGFRDLotj1iYce4PIR3Ze9JzlYd8kwEuVptqKQstqqQ70NPVu0cUKRecgp19Ta
04fAM1WSG+4eDHkCOEgr/o2kB96DJjQ717NL0qiQeSuMPEPyCa80LJ6XYQeai7qXkVMXcnmi4hzj
siUpirCV0FeGsAz8kJURFBT9PCe3AUqkzC5e0Y0UR7TauGCNrAaijOprqCLLjwhcGS0/niGiWnsN
UaNTfX/swFInnhmgdt7BnrzAtju+LmfZ4WDsTVw6pw0RoVoYnDSl7tC+X6BuD5lHhnQpjU+Fj9kT
ok4kuIlsCCq4FvlNmkNJqpkNAI+mvtE6dSocyGcNMXhNUNHjwKuj1+ulYzl72EvZ/+hR4giI33EZ
CHOSQRLnLjrYvRNpIyhti61/ALnmFzGGQl6OghzIESDUBz+ZFc8SPalqBxLJOpcyo0C3zxfE3J0D
6Qw7cpA0edjGe6fihKZSjq/Myda12r2LLHthd22wLAQkzeyYcw2Yu0HUl6YvYUSdTDfrfKMiq4mu
SWnMMh073hTLjQTDehMAz8BCcgsae3QC0qK3VmcTtrvn4fFMXXBNq36ldmnI+HuiJ5PDvmRvGtC2
GcrHS8DR/GU+OfW/iNZbYpAd46u4SlwRQR10EyV/iaUn/COZQoqX4iePtYnGAfJ0LxNTfPqhSfF7
x6qyaiIfBR+UoRT71XOrZDN2h2R5T1tlJyi2zT8DhciFAD35g+oVRKk7PyEDFQi8BLuXFR6rVnvN
6LYUQ2k7BQlnJ9C3xtftJ2wqWa5mWYzG5s6WeqBTaUZq8UrbzaSJ0KPD7I3jjO4XI+mdGHc7njCG
RtU7oC4ZyNZZe+OS43ij3E7FBt0MvbDyXINeBo6lpMmyIrNwGrISFCtQtlYzGAM9pWI9bt2yw1Mr
BA/KlVukeVxgvjyywFMluBAFDvFrU3WSMGCcQbt2uSwX/MGmi60CngfeZi6nq7ve0z26Yji5nhEw
wpUaiCLuzRrcow3sEPoFHzkkfsoOhZtLCes2zNXoWG4YEvR9aMmcMZdPgCkg7b8H3D8/k7xMWx3m
P/HPQ0B6BYLxkbmEKV9xLSnw2Mf0RhkuuY5BMCWdiuTchP3LikXSo10K2V/r3KVQ3imgjNXElfEp
L7OTkzpS/JP6RF6zsJARCvKw23RTPjOZzo56Eew5+jD4ks2gxUHVa4thuZ5g297m693fqOsWl7n/
gHseAh1qvveyISB/eJRTvdbWPc74Qf00k2fEvDRTTOxLkQODWxqiIC99j7nwe+b6fAZoO9aa9DqF
2/NpQd+pghnvqcsUXVDRs9E0si6wgUxp7iQXXK7MJ/noMJaIp1mNlGkbVjVHmAGXokWDR1uHycTK
OpQfpip8MgDcNe4CrOJwLg9RkuhL4yvsaeOfztryNPkMpjw8Ur5PF20uSOPYqYNmU2+mMMzJhrNh
9vunCccJaAWLw5ZBSmUqWBCvog5du5BQdXgFSsllyCW1iAJEIFlOy1s8F87S0wsl7UxCbugEYUlZ
5GVSPbY1JFdtYxq6GwJTwzqGdeit3JZFVxaeA6nXzpnQV7M18HSgI8KO8FKfwSLH83xsOWkSUXuw
dVwkQyC6/hwDwg+nUKEXc6sMv0aU7sTJD1ul7gNkn/Pp9g7pn9hrajhY+3t+9iYYQkpo3C0j41yN
Piufb8hEq5yHi/kscNncgMyRMpyXUi7SQFkpOIWVzXyisEjozrAK6GsSkUykYB7gNcbqbzFqNoxS
4pIO9xYVsCJp6WnZAo23vwXsutz76uUAGo55SBSL2U8RGMANIu8J0HDD3qqwB4vI0NS5oM/I4z8f
XFoNm+P7Pj6o+h9nV9vJqld2KeCNzojN4LZyscKQ0tSpZeCO/z6ayMhnia5SrD5hrkJQBa6AB964
t1QztfPqaX1pkucRU2/kFjQufRqVyYZo0WoK2QEvtq1pLzCoEw7vdc/vwoHYaKANMz4SL+jBEbrG
DWtbuiSrSVlJzpN73NEv+3me32ynMLsU+O0irwXiq8WbY8JsRdj3v2k4VCEuGpe04x8he0yy7AZ1
Rwy7LxZx2MZrYBXvHCsegdyr+RKB3tyFYlMwohZns204zFHliauDqm6UGd4FP+V6yjC8mn+Z+p3H
LkPGGq1ixSuTLj5HXGMHAtrqGrnQLRUV5aoC7tm5S/Z2rf0fOvMAfvdARBbXtBA6bmxhZEnOWMFy
7Ig0d6hzkiF9bDLM5tGbO0ZaMeKQ1IxQ4UVyW/NQ3RDdb+aVG/LmqmC/pbmjBiKpKLzHC4xCZlmo
cLmpBqWBkf8TdmYQMuh9ip3jWQTgjWrPoX70mxA3D4EIQT8ngX8CzBkwd1uVOszjKBj8nnEI3W2o
RyI9fg/UgNKp1HOjZ4hvFLivc8b5ekyuIl4ulXioaoide+VbRkYWbTwe2t4FM5GS1SmjENc8b7ol
W42kHrvIWXfo7nCttJaeTdkiFLYb74IHRycLi/qhqwi2R20pUHqp4meVw5LEyBYU+qHLrDHMZv0d
jmLfwdgAtzh5ior0sbTgAkYAcmzxGfHw7UlVcaK0RGtjXyuGv997ArweWsX3XSq2B8rEm6O2wRwD
82qwqYXhjc/b1/QJpc3QJIx/L5v/N/4OaLwdc1r8lefjiGnnlpnA0gkSNRb0TQADTgTMciXadBFq
5dkXmCjQmd3WBYyLRj3QVLjlA8stx6a/dXd4TS7ZvKMCPDRB9gZN2seEogx98biv+oklGa0JHv18
GmwOaLIE/McLV7bKfxxoSD1dOhKStQZk+rl+wKdyFJyeFV0vB5oYDVmTgEINrjbvWrwSeuHE+r2w
rdfcK2v+mS31M2F+n6F0wVnrXQ99JDirIG69OkVDTHejd3O14ny6yDZyjZYxXDZum7YlL95FFh/p
bGP10KvfWweETYUnKoqOZ82AaZ6Kh8oYmAlXLBRZxOO5x20qRK+bTuZ0YGQPYIVB3oIyqeMyq90t
iSTqSRF1tjVKacOFHmxyuIKDj2va6xTUhoSfoHmT54JU5A8v4ppk+3gXepXcmljQHNipp7JKHYYN
tf8xhn0psC9MnocvR/jfgUnKLLh/JcW3n6uBR+GyosoeVzp6ZiirZCe0PXx+C88hdLyTHhCDi2O6
QUBS8N7WO74KyoTfK1nb62kUum05IZCEDD+UmA3pS9g1at8/IVAKt9TzuYbeQjT6a821CSzUbx7l
z6bpNm/MpS3E+fySM4hF4MlBtXLqG3SZeTGCYtRrndYyeJo8wk+wYnHVKQezOnER/+DLL+WZZq5K
+NqyLMPpxX8iN11xckLw9vu6rA4o0b0UcMJ9h493aeZgso0KtZ+YEXAGovO6BIcgH2vCHwvIsAjq
PwNx8FLyu6GEeRmP8AwCrFolIe0CKObP2GPXS38uWWW3q/If/r4UnDYxz+Ti6qcv1rixNHIhnXfq
cpW9VLZ+zj6Eq9UV49AI6AhQzpSExx1Xmy8QgrJE72oQwVK94Yuk80FCbpq0lJ3MhT6fnek+owIf
3OkyZeH4eCG/c269gQiHgyapbw11+G8kZPeqHqntNA00PqMNkhHfotXDXWFJ7arY8PvHd2hetsvf
JIFJikFx/8LT9FLZu2yJ7P2+kDWFrYg7eTmkWgCs/1iuSNf+HEL/reURtt4qkcnun52s4RJBmagM
RBLW/p/u3dvqU4Zi1c1zZWIYlEz+nfG+S6qnHXGjF8jzlqlltOmyUulPYVGwnHoaQlCLPoKZx6lk
wjA4BLeU0Ws28a3TnnT/EHA04jAdAHNI1HUzKbkaoJuxW2+OpUkz90kemNPAXzO+AKXERs3UV7RH
/V7aleWbOiLGHjMk1AfXFCg8icpUDRE/rivcDkZ9iJCUYY/h3wOfR6BTsLD2r940af/qCldbBnqY
akTSlwXpPLcKYe69w3tkVrprB3rl/uHJLL85Qjjn6GluD8tsMrzxSbrjsy+wlFPUtuDqiYb1jH6t
GKm116ysgLyILFFNYdO842zxBd/weoGLs6fFAPC5ChgBMpKayCPOSiqAuFEnspDELTxDCsXHnIes
9G4SckI4lFBnmpNgG6GOqGNbtD6ss3OfoPBfmRkxxliy94eUs/L8gh/r+P1cN9KOuAjLra9OFzZw
ct8OHOy2KHpB/VHP1x/geZjpymBq/joM8OOG7YofWOcADtpTbXg9bUcsnDcM45XrcxJ4Pq57xfRt
8z4ZmsFrtdfFRqO3gEUp/77PkJOUKEocTJn5w6RbSD4hVflYqn60McQl519hjqzdhHJAhdT5awKg
4cPTNNtEHE6dYDqynrrtlDFXzjZedYAepOiOLaReO0Gboric7rChz4wGwmuAKoass1R5d7+0oUmX
mb0x3cit8Aa2pML5H6VvgpikgbhaakL5LQ4OeWlYxugLD2ngHM9yp3pTPbKPWDP1owQPkbKpNuzM
0e/DrlgBQQtFE/X/z858iwIbofbo4hj1DtBf3I7WSl45HddCWcnKt3qTuZZC8rOnhy8nuogZFVCa
eUZ6WybKBAx8D2H+h+YqOS/63UlNo51/bpv9z33KjBPQVfmBMJzuXdzYeaWXQzvaTtxrV0WyO1B+
y4LfDq9YWsyAfUggjnKOQlynssjdxrLj0aVIUCB3iMRvfIBFPdUt0k2en0DDaw02BfB1kqL/qs7o
fcj9kitgqFFvxyKs97a+dNEk7HZUK7u10icuxrttHdt+ODkrWzqsjF5dYcm1GPG3KYyRCqwtEWYA
LkovpzpiR0QePM/5+ZfQt9a1oBCfORUpNd2CqyhNLas3iV6sEpYgyQyfk3ZNKw2VoWhBLIev/dxV
4+E60gwv+1v2dG8BgmGa1RbY1RS+LPUgxBwBVnpoB/+ZzljbLGKQOmcdV0HEMRpdB+Y52MBiwEn6
4dW6Z7A+4J7TioA/v56z+LCjEAr3jiM7HhevsHO1VUHxLHpZNEFGJf70cJsHT3wCkHc3pEdQLyim
Sl+smAxoghecrqLGiShyVpo44ybOhuHtcqg+Hf4JgEB/7aJp5Bi6/JMX3EynD6uHzOpvKpt4X3Z9
sJoGQQJHjq5GcCDdx3xAc5Utz9fZO7njDtnQJcgLQV5PmrqYBccJyW+KcMdNrqbpmMOPsy8tld/P
J8LPkJb0mkjfXPBssFn/LO0J4n6Tz1ecP3SVSFMTDT6uJ2JIzVgPgKieZsSDeIeIINfNhd44QO9c
UAUefG+xii6W5MADeSCBha6m3vBM1qTA/QWaFlB20HpdlXVKbvmzTPicFsVt9Po7K+YoHqGgtaQ0
w73IM10jjdbZ4ywasr4cv7TK5C5wy1avnbvPXC4LRcWQ14eFIdexrVYhct9WlPB7bQR27CGcG99d
8cAQZLMvPKFvzXAbSIDMcv/WC54XVUiAYy1uxkLGfRLkRsshuVA8QWcCkPXDP4IRiUtRa+flbS8K
VtwLpk+8+n9KbyhKX51q5ZOpISk+1gTa/j2xKM/gM9CYCboQEitPzv9VnpZ7EoQka1+FP184MLq6
3rzl4tVdzIAWS26n4+obsAQ7oFdjmH2Zthc78ud+KqkLErHpalMHYXzMH202Ge+Uccg2KJjJb75V
j2dfqhqqZ7CHtSRn3u9jaznw0hQUUC14+kpQDb00186AUTiyG9qUWAfvh7aACfEFQZTKwsjXn5s5
Ie7u8QY0uPMEbinXWfWM2OCtKRUufNTkfq452eLV/ebelZXTZGpBj0qPPj4w8TYYsPwyu26VcRHx
pgOR4hQAFRBKaElbmIGCvyHvWK8hR2shgkHloUqWNdZ6Vh5VdVDEZWDcoDTS6qQz1NWUTv2CGVc8
w1Dl3u/e9jCkgXP6Yl19z6HwKTEvLhDRtwjwOz75CBxeye7D54xnfGNweZso5utCfN6FJWiXLqUi
CAczqEegKZD1OZ3JxMoO6EfvXY4Tp31bO1+P3B+dx21yqqgUOSMarZG4zKk4M3LJV6e3AokksJNM
XjXQQD/n00wvG2Pr9H2+32GfpPFbtMPUrQ4vcS0Xr2tpKcuAway2ELt+bfrSwp5Vpw8lI4hox33/
6CIfgqZzoxkSCAy3bO8kaQIxyue7YWF9AJsOT3gf3fItLq8aBXoAvVXoLWH0CnWGP+m27tawZicv
Zvdq1gpEwNtNiMTrsTRICH33AkT5OAw5nq7kjASFfDCQ5xabOnzCmILNo+UnYMJVJA4bg5yUBfql
zr9ffmGyVBb5g6TtlVXPnumFsL/ecnn0N8G/KkhEv9QUPWVMoFVqXTcdszKFqVkdokZkGoLrSNWt
QaxBKX6szRAB6xIzoZzroqBYTsPRD4U9gPwPc/oaiEVlzzF/gv4GhUZPzA0mex+Xbb/16AcEDMKc
Xb0ZowcxIvjrflQPnVJh9x7XP0cKlC3pVWftoAG/uEZ2Lhch084pfHSQ6SJ++tWHhXyr+ceR5yeu
jgx2q9MEPydYdkibiexdiScEYaBfSf34CoGvNvz3pBrR0iOfJOgdf9IAo4Qo8fJn5MqpZff+emf4
FzOO4Iy/Ow3l3+R+vx+57szTObLcyxPxCSTRaeLw5SAj+pmA6xm/jc6Y959Xdp7/IyeXRdpDfUxg
63xQsbZlOobOMloXp1zP6E/y6CohSxy5xOWtP9LzYbNT9woz5/LjzO6ASC2oqwvCLJ3gi9kp5HlC
olmFUPkWNOnQgvb4A+xDwsBHoQ8GhuFsfIKPUer8jjumPaEf1ATvYgtUg6PDXKn/7JO81ciZOlhu
QG7UIZQMONTW2JXj2u0T3FsxlBQ0X4KC//noqwYrnC795E/QIs3sEIFbQYIDS90tNEneY5i4SL2q
6a6Jiu1wqDQUhxdrn+b5R6TiCTzJEJqITaDdfahYcHgpvzs8J+Mw8/8rn6KgW/LaWza8yi8WaH8H
TS/M3kxXchJJhW+1JMWXzlfpywM7Qc0Ph5SW9cSVZpvuYZu2ysCIoxFqq94Qbap45Oim5uT6VXII
O0BGBaVX+jrFbRO6y7x/quk5Bz2UDZ+TfSP4o/whdJ9u1aGc44ZRso5poE2OtCM3Ydjpm5tOL78C
rgsEoJ6lUn7+jUs0qltt4OCzZEGa9YEGpmzGqnHosTBh1mN08Fq3ruhXtTBHgjK13pm69lWUOeIX
bTmRKpi39Bfj9671Ty1lRXGryK2cch5LgLUoJJ9vxwjr0rYO6m6Wd9zscTHIDsrhnSms0DUYLaCp
ZYLCoxY8Mo2nyP3FVz30MxuitpBnz8+TBwsU0GblUou5S0lQOlXI71Xwm9jZnqjj1qahW8xOumG7
6wfMEO9twTeq2bE7llUuWiewhtwWepnE9tEU0LnigDhTeZteZSZJtr8H6wD6iPS1JM2YQjDXAKO4
oCDBrufEMDryzJZlPPnz8Q3KqkLR0XnsGcoFCDjeAT3GfM1wRVVhKplooBOGeR3S5hahy7M2InPI
7t0nAi6D1aCvhyYFpQemRwnBlfw8DNyGltfqAkYHT0D15pJgysnOjrRhf+VlU8kNFcH4GxYDIMdM
+TEzNwdTDxQSgbgm3vFrmvl5DY4lj2uPSuHdsTrvk++XVuyDHueEYbFWKLVPRV2iHDmai9fXB0UY
uhTd9SabzR4sQEJp3WTxbOJhnAv+ri38wsDHj0MX7qX0811ioMhgx0j93WGYedEp+Kv+RqcnocJA
w6OK/evZvLx6WDyGI48GH/PcnDHosTjC8OEOLnx9lpF6SCOY0b67KpchP4LHmrxaSZfmT3XdmZIT
73adfsdK0Tgb20Dx8L4AQ+MPI0RlhkMdoEf6GU7sq1+XMkw5v1xqKQhmaD00+3kQMpEHNYNBo0XK
SzrO7rz0bB5eLguhCk5M8SkY22/tRA2mtrVU6g3KjFTvduayKp/b4va7c3SeyOlyvjlPF0f5xDu5
1/8hewaZ21dglN7dPU8Hd+EFagjrwNSJsVY6yIJaJLrvrMlajDe7Pycp0+zox7tUXYJSQ7qBjecz
I8vBiL1CSBRo4PiZipjDejRZtxZIHIjAI2fjJ2h/6GNN2rZXLfFT0ijE+q/oQ/Yj5d2DvcRCAPyG
0VfLuEbKUMKDm0lH+33FJlv/WgU5KzZESrvu6Gpj700Pf9/8w7k5rGBNT97r2UnKdBSXkLtb5dEG
P4CZpcicmqyy1ReOOf6XW30eesrtUpJyMKdFkJIHfD70hTPgykJo/RfkoXX421zcydAMFoQgIs3d
JOKRjip/jM/Ongg0pi4bcwDovClfPul9jZfI4iuczrRJtrkaWMrPQYbGpFfzZeKL9yfdrEjAn4RN
BasxASxWDE5fdijb3mWI0lrM1CNaWVRYPv1obqEBfh9XeU7JAKqmHAJHsdKExW/gu2DkviUAjjEN
9mGzO1f/0RMMZ3BfgK4IkBDBAAaDTsCGycs9NwrgQ3/L5c+JOl8zQ106EXgr6URORiPUX71o9CAK
5ikVhcIortXYGmG8s1VfOaXsu2+DbCqWO8YOPsfrY96wc5/zeyniHq9HIimnnjRexCq9ZF3Sbpdm
Dzj00rp78dPUTPzD2GILtJc5KP6sNM4SSC9my1T0qnDEx85VOUwv9Zi8AnFtrbYz/vO2503HhMRW
SLxqVH7Kp21mhn1Nn43VuBXkCGaWWrxvdrhNjAjdpkgCE2k2CVsDAI6gnU6XB/KFaT/1kYXkS2YW
PhGJXZ6QRZAsGo3/D4UT4t4BT0SNcpWRwvAgtSybH75rdFYD6EJHrcP5SsoAp1LdbEzjy6cN+/W9
OGcCZzVBnoPDo6HKloPG9dEpMWOUuIzeGS8Oh6p/NMhHwkGBlH/anZdtNCRDsC1DVrxjJo2VwSAQ
PtnSUC+ILxv4tzlIpeQWoQG3mSjlDyPwm0/CCr6wkCYkpv+1wbKyAGeCnrM2T9wSXyyS0EG9oGRh
8s51ipXS7hN5Klc5L9ZfmosiRY16lz7Ng4xPdS6XjCUeqigVjdWX8FZWi4w08JXyVMf5tf0Lc7oH
Uvd2LjB+v40M6IE9Wv0O9+ZwuOvrQuDRc66Sk6CRdRVMdq9fiWT4pxhBcLdAYk9bCQoSuzneOUPz
/SRjT2FsfL3+TfnCi0Fg3e6Ra8/c8QOg0Iw2VyiuD/zsW4uEAGv0VbBe2aINuNtiJW6o44ANeVqv
hi8THuQjwGTBjhZDc/dE6SQFkq9Jg7YhaDE6nQdmXkWjzj073JqAgh6GveVBZY2X4ptMZ/2vrrS5
awFe4a7HOcsiYOMD0c9pCOMKwTvTh/myYYYOSOjyyfn+IuLFIw1OVxLaag9OGBpEAXDMRuZwA6Iq
BxYCrFOYxw2sAu/d7XEBTMVVkLNIWzovsXDFPaW4nxSlAyiYR957Vo605iUN+SYh5xqLOqumKtmr
nIYENRxq5ygLPEA1QyzI3Fk6Lj1fZKArBP1dK5n6O0amOQul0/TpwDVHOE4EY4qRhxjcHrRw0Vv8
OTN/Q63vJDNxQHbHiXvQdcFAc1gK3FZBNznbc03oiS0JYo2Io9UM07qS1H4LToC//PzxdZa0NqHx
nJunNn9y31SxwTmzdRKB76RqdBrrzGtv9WvQTKtvp9FKwa9ScJ4vv3R4n5DAbIO/CJbZVCfb4Xpf
6r6nGuKBWfYk+pEQ+PmwvFpB7Yx9d0n0RahUobfhtDJBVxxAwZlWaIDuQ5Kf3PKjDy5DiE0zqXHS
k47yrVMvvu5LVj1c0ldwz0xLFeFXKBMcpIwHPjlIYM6oSxwL0CHXvBCClbVqRaSE7NY9NXOjCCt7
ld2tkNPa8Q88qnS4wPJju2/gEr0fsd9ldilbPzRccpg2Gob7o2SCoyNPCNNIO2m51+2fu4bC9lQI
xa1w97bSRzP8DGXUL0ijxpThfkD+NRFj+6FDNBoDPJ+ji/AFmloXnMaeO77x7upXcGCDItPJs7pa
Yaw1k1WRkG8T0kJq+ewymfmDMtFnysGdIe8lDCTcW1A6mYMFmE+QlUk1oRLHrY6sHFVya/ITYSXi
O0DzGPetHq5tMn6IzgY3nCdY6uazKO5lvnW8PV8imNMVJNMj7Frp8Ai6DG2Q45vNnIJrO5sF8Bss
5WZK2o0w0M1oYFmKOSxsh4RrlaPVdu+XYAn/b0dewGfZ4iyPK6u9TNQKmLlknYiKQ6SjhnAoyGs7
weJlmAm43lzhdYlYVIjC5ISy1wC6dcsQaWubTCxHGwtrgeAPI9yT6MgRGeyBmRC2tJ90LFqMKcS+
gb4WEj4BtHxqLuwh1/TShS3RMcGWXzZPix2r6Cf4/Ixlf0WwqTLf64ithdXUPdTHwLZ34s8JJYLS
kUZFtBykk2t4/NMU5feC9tLaXYSi5jU47lqWgtMAYzY8Bflc2kBR5ostcy0ZttxfuGtMcR0Keq1G
i4sMXfv+SZvQw4Jop6Hm9Zz0Upog6xNHQNcV8oLmOtT1UVqNm5YrXBybvn/0kTHSVu1qJPLsTz7z
mghsyLlGBksH9cS9oVeY5/LuCez817g82rRnDOLW3HJmwQCjQCNF+Fx4ozVgcMXcTBJMjjFRbSgw
tytV4uUvzbK7IRwZVaaF5KiaYaax4aMR7vCZ6bLz4XpKtX1X9nfGU1LGrF22UXs7Eb9suWD7t843
L/VoTOK2W2wfXTxe13Wlf+Rld+Tdz4UEhxoOjhahj52m+bV7kfvJTHPZ+CvHNCu/y0CYdAhdq8Q5
7nr2wkS6oqU2H5ZCMYYv0G1WxXN0Co3htX3jpRunsbgh+u/iHTgb40xMz4RUXsdRbBeHW6BuOQJ4
I/XOzyRSocIBkM+F+5Spy5Z8Am3MJMUq0zjKyq3bU9qtxeAtvXU32lWkzK7vPSyB5qa6Kh8/joII
cWoPFdJoXP8kQX+Q0j388HZ8pud+SM5QEL1KiiLprQXoFwsMd2aUILLoOHlYcbD2HJyCwv0290vj
x71oWUzrZrUIGPwxXWa3Qhrf4w49WyK24vU0mwXjRDU4+N0o4OQk96go6fDGdj58lrVkSo/3f/+5
y4F6xFYSCJb0Y/WxSR/ypVe2+BW35U0gQ07RIy5kRDBznhGAwXJHGCDC98Ox9gxnKa61Gpsc2xbV
KXKgICax4hABgsBjT7hXS/wvpwXWj4YwwFkkj4CJ3L32UNbc6TKkoqxYgj9ZYutelayfG+zXOCO1
trzZqvpaRl2gve41AuZxjkVroF42szVBjOilRFMl5OVQ76JXAci0BnlmKtrg2HlDH5xtDU/OoUez
UrUSduWAhS2poJLIHZSDm+BKYw3zcGZe8GrG+IM8tQmP7WYgJ++PX1nTFeIuhbxBfLJSVqSgyVU8
v377sYxuYXZYT7iO0r1zdlZ7A1v9aMzYtVnLHesVmRAUtp6HIePM0ofVqdBOdocfZtMDZIwjaCZU
IFaW/Wykizy2q/RVX8Qd0Vr8NuoSFKLiFDf/wD3ClGprQspuPt/h+iHOZKyC8gsAhpyZ80UfQsBR
H5qKHOWV6zbrR7Zw7DYe0nriLCL5CzmBiUJcUbL3tGKBatIRvq/11pZL3dGNjpzqWAb7T4zQa5TP
ktnUwJpzd6fXTKSkfVMDV83DNo+ToxoSuJcksf3uJiWf+XXhG71xQQhfNMaIc5POL5t/+8x3JSnY
PbXI7k12+MG+nBF/vXr9ww+0lH8P0trK1WLzVz9+wkuC1Kvqist3hXroH8vexoc5bb7ooR5HHvLL
5At6uGUhlEkosZf1q4HKvZUR4PRxaum8x0o3GTOX3WwX4qvx7GGaWU6G+LaC5ufg13+/ARFjLaP6
Qr01P68/WnYyKmgiedE8/if+hnvf7lP1wxJSd/0QC7osw6HbentOC0ISgBOBwRsjfeWC4+HsJst7
dHJO3cvZtzOgvoRbQ6+d4+ezrjrccG2KOb2LRwCrcu9h6gry20rhMh2ovL/0iN4kwlIIpqrXZKYF
7h7BWKk5HYtjcSkoKWw5lc+S/kZMy9UBN6g+9OGf1P0TXcrwsuG7k9txSmrZMSe7940VOSUUJiZP
tnJx7GxmQx40Tb1XBad3lw+sXTNIzk+TVv5/k0e9UDf5nnvKI6L0wAlOmNiI3bi2FYn/lJQrWL5y
C5XVwNLkcCOBdLJldBKrPvUZsd4/E9ZAd8uPmqhT7e2RaNEH7xciv6XIgUoM8jXjkjawywj+XMa9
CORFTCOGzH9nljgowDKGS36SVQP34Hu3CZ3na/fbpxk7/aBC+9XCDq41tQL0y/rKrYW0T7UaQqN5
IY3D9kRHWtAQy37tV5qEadHhQbgcB/JdJFD84EMRzNHhINaoejEkpt5d+ry90hHxz4Xnpthnc8Yj
qW/3nMT9bhDbFePUvCtPJK0JCmlSkSFByv6bz7oIxQeH09eC6GVttO8pQQTAqq7cSXZ9vwBIV4mM
T0vFwtyAv/8JZznWDa+iDnnokfN5DmkuQxK3n0J20mEEi0PSE6dO2dJ9S/UaPNoOle7V7hf5tEGr
eyzwQXgjfBmNC6uHWBjbtyo5e58n8t9JWcojbhi+QjadRs3p38KgO9xLhUsx1JgjaU3I/+RPFNZ6
E8GmPe3uLzhbNrrfLH+Wcbr/88Hs0b1AuHG6debzF91NmUp2pihvKh5G2qAN405zDN1GoW3yOyDq
5nLNERsCZI7j0prl0GGa4M14OmuCLWESifL8OAuugh0xZyK3QdcHQiwstu39jpywG7hT+K9rtslp
8BKFy/fWMX06K6yySgHjMTvmfOW+hcwBkMm2Dd48/luQCXUQRmpzkLlGt7D/O7mWejIM8f0VuxPd
fCrJiFUjB3t2cgfXwqeXlSecKo5232+H6nfsvmWnet+fM1C11TCKukL5q34F6cbyHseMthHaNO5a
SfZfk28fnE4vD7K7GhGNAXU0K5Jp+dSYN1hzjuJr8HTmxkzQPgHRiB00fppbfc6R4tWE4gfKyo30
VVp1gCOSn/CQ1c/LslnX0F6w0AqJy8sJ9ZiMD67y3LcuDDUjn7I4bLBxKXOL84bJrHchDLLR53vc
LLjVVPsnJu2xX3Ych03eimAJbJFxzLStxQVXjk5yIbPPVHYjTcxVgEWtkOXapu1+mOais39lcAKs
N1m6ITOgaZI4XPWQWmxZPq84cIr6jjUAfei/ubrLrUZmz1+erFnAyYbEj6QYKIccsN6PnqajYRKP
0O/hGmAVW/2xv8+H3XUl/6rdtrvgRJCDr8366D3BB7MRoXlzq5H8ptwOAhIxDjpU2oTuYq24XjQm
NU+LvOBkzcOnwfNO3d+mKM1DE7MbCtfqNUo/w/0oKeT7sHJotX3g8LK0IiUxYM/RNtgl+q2/AKtE
NClFSO3BHWdM+BtCRJoKfSOFzOdrmtQrsoWT0JUac4dzfY5J/RKK0I1gpRt/kDDsXm3ml4PMrGc4
TlRD8xXKKDMWzHXsoJyuOvu7F9O6FCfa7kkjfkgqrWLYw4de/1sKVX9O9EEGBkVpFTw0vYdOlz6A
SzeAokdkjGl11LHJ/VH3QXSdZELGvIjT5tWnlnJ3gPEmctZ2PyOzWIVZ9irgbfFuGFRi8ak7qUqM
ZcEnunj6SyS/r1K320bJUDDbVP9EauEW6y8R4sLKxELg6E2a3rXI7HAU5HcVL4/UyrHJq0jgOmDd
xiSizibmxuRUE/nkLborOSP83nfKTNsGu+a+keSC3O5kZemxCT7leqVSA10nZuVvqOJrQForQWwA
9DFsU4MTXaEHohEW1KfM5hLWJCpyjB4k5Xj6HdFCKT6hw04l1L+Tk53yk7n9C25P/9vm7c277aWo
uJ370GS2N0xSY7WPlYVLiPQtxeCh9uN+wXaxyo3qpMM3OEmIUl5FkNUuFF7zylaY4JuZUCLRjh2S
BwV6bOXEL/QnQqTgZo7rwc2q67WXZGelQcXUyUk7WJP2noY7I3nHnwTfxZu5VyTmrFKbcBhat+1M
geziNgIF7NjPgpLq+M3Jl2WIObZ/iNfYDc/urP2lMZY3OKdrwUotooHYx8C8cG5Y2ekcjTlo0uVZ
B5UwQDj9ONB4oWwku6xewGtbPSwq+SXv5yDWFoAQmNag8su9/Z4pY2rCESw6en9ZYQdG9b4ZDOly
WyrpeGP4FzqZtKa++fjKFN1u/LVimVWN/OBZBNsGvpGOGMW7nJ6+fpd6HD6pUybRPkZrAe+/fR1z
bCzsuSP34CVFsMOg5eiVcBM1Z40iHTsHKdSTQRhzglJF+CKQ33FTZRkJIpv2M8vJWvjM6jv/7cJr
cjunuVVG2tD2y3yp4zaVGJCQbzeyr1BEN4C5MJk7g8NKdVb0OSbkGfCwmBsb9pZjf/wYZYD3t/S2
dIAJvEQPUkSm9MRgbNVDq6tmjE5ccjUu9SN7QSgj8Erbmvyix8hzDIqugy1z6fjOfeNszekfTWbH
x/32+1EiEK1tyE4SZbdNsX6d6mE2pDUx50EVxchyESizALOd+eL+duWa7JxNJi0GNt7OJk46QFv1
8sqstqtYTgTt3iXPtNZH7wV8BOU/b2xANhl6AaZsFMu3aHgOPOjcdkRes+lmbJylbvWvDtvGC3iq
bcrEmG7Cc2BqhbKcB2fP2HNRjGCmp/G+pHXfJeTPRnz3hMsnqqPKw552Y+e3hnvmh9UNo7vSSCf2
wS41gpxMSMdDV/ubxEew92e75d0Zo+k7PIRdGhG5pNoamGgAJ9J9H9a5w/aCodCC9iK5Ig==
`protect end_protected
