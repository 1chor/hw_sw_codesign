-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
nAmapBLa39XuRr6p0CnievVoXA37DKKZpC1TMqavrSSeeQV26dxpZlHZOQGX9X7x
vbajNcq2fxUgAk26QguxN4VjPaQphFJ1TTWLPMLKGP25v8M0pr2vyW3ac8Y3ELdM
a6+MFktMXD72zdqK55cwk8faLeS0d0TrY/KTpDcKtgs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 45955)

`protect DATA_BLOCK
ZlWTNtxpYuxxweQHMce5OPfl+m/aGbxdYqM2OC4PG+LJzt0eZIQGqO0WEaA9YMwx
/BAvqZn6DPnFocUeKV9KV84S0DW0k7np075OOEWjt1TWA7mbKEWHAGDr+cifjZCM
bzgNspw7ME43BooCH7YVroho7l3jnpMS5sFFKoMoOicfewdn43foeIADf2cPjaTx
FwBhn7cRpoeEGu/arZMLaFavZD6VE9jUOiCDutIIaOoONTL+NZ/JXOm6ILbwCawD
zGkfNxurNekzepnPo5BBK5WJwSQC9VARFSO+s8NTJA2/b8b7ADfhGyW2r3zmWMgr
QBDB05NOyvD9njYUDlwHxcYUfwhJ8vwigMqxMZWeyxUvghhKXiyeHa0P1MvHd+4Z
DULcFBl215hPZY/wMFVl7XKTwtJmMjDGEjb5ZfhpIlOZqGDORzUD7UjmPRPuqwJ7
tZNFVHbGLDZR0Gut64e3Y3eXbmIwRYwd/qFnYbrRhvRgXScSRCna+iIGGmk27dOo
VpcfzCzX3BM/rL9t7tc8BVePjM17sGgXo26BbVA+I6WAPAIa+vuVvpPrO+zaQCvq
slGgC8PyIWVogKoDzVFyXLx/5WIqiWljY4UjonLS84jPgSq3Xzm/q4izhUQAXyWZ
0dQi/2m+KFEuybcPQNYHKb/vHNIaiyqYiE85NOLjK8TzVh8CSxmUQmwvhPWzXHY6
+Uq7PWOwmVazcA5G+X7O5NpUSaMFX5CcZtME0zVErXfjQQ+EEQLE6ArdkMML5O6t
aaZA/iA23wEqv9c0fa/baum4wUdjSE2RGN1uy/BEOzoEpyK6regW5t1E8brsu0fT
5zWoXvBalOPSv+YtFONgPWADYAte32hf4k+HXQFTi5BYJsJpf14I91gjpjxkmytQ
CQiJWwX3AkO64g3Bj+Qe52kfqtWnR7z+Ula5MGErx8LH9WcSk2hV8p004jY+7D7X
cW7BEoQx5NEsmi5wRU0C0rKs/CuqM9cDHVWGO5Ft/Ve5pP8pVFZwjWF2o4rsxkFk
2Z7Wkupjb8TC6CZaGkX0MnnHTVSZ7LqVqvw/bIMrqdXBUckLVZZszPmQt6H6JODb
L+m4pg5NjRRtKQM/pxYMGTTvhtlaA5O3gEXLaIl3ggTXG/FAstvaymbdqPhaAtNH
o5F2+56kE89r3rZadnUxVRxC0uIVckm4OePLVdNjh5dXrExVXQX2VTzDS5oUzpCa
r8cJP5YNRaljeXWUXAGdAYXEqxacluj6nYfEWu6x4fs88CZDj/m0ESPE0lSPcFov
UM5GDKLTYmaM58c0/SfQ9qZQdhpobjDPtoOZiuuOablLveuNNkd18jlTY2eNiKYY
S3Balv0MVaVriU9omXAUQN6Ps/8juxaP6PBhnr3pi2TcvC+OYWxzuLJGQqrSIQPZ
rZdM302THUnbjTQShEcn1k4KS/NhKOz9oUbcFt/F/3y4HBxnZhJxRixCf7t+Q79q
ks0AiVI7CEk2QtftCz7xyujdYvOrVt2VwhrKz5Vaug0o6HEcmmP9Bg3dOs/k2hEf
RTHCgj+9z/qO1gG6TSssZSKSphiwtH6P6D20tuk1m32x/R2B+3RF+nELo1F56qZr
i5wY2IWeEIw5Dwiw/eD789U/X8cxoNe8jfNp1OatVCcoTMyiAa/dniKTL01yUiaD
zQHlG5PKwNy+5f+e5Yi2X/FC0BbqhscLkLobP9CK7QlTj+bbfIBt4m8oniqj0dhq
SpAfrGg3kfqHLtLR+2dabWffiMJTBC3iH44GkG9ty4Fg5eq1feJfs3m8DC9C/jHI
SwB/At5adFnknt1CmEQm4SaBvEB/GhVfWhBxH77JacNPIq2AcLAlVGSYovXxIIaw
oQF6H0G26N3upgYjidFTLc+7qWAAkTnWGI4Gg5WdagEvVqYTBwx0N0ZAt7sLYkv3
P46RATDsLNGnEy+rbP9tVfYmtFKzo3hdBjd4oOwsae7nFzBjSXEUTKNXrH5UXTfx
15m0V/PygtwNkKwzBtktyPtTiumNoNt8AVU3LPkzKOVNCfm7ZPsaRQ0GvZDYNqqy
7X+jJmc16IzMGaebWmo48/y3cFuuBjzqce6epOTfTMrRBknpps9PVBNFDISeOzgZ
2vn7klGjcRWeBg50oWa09KNNomlqQqpd7IYKz1ACPX9o3tWVpk53jErHkb2i9ykj
YJZko4X+M2rszmFSSUTosgEhNOy60w+A1f/QAhwpzSfUOZShKQVUZI22NWQHMhKB
ekiXxyu9FY2L+bPzbbpww5rt+cZ+d0hs8lJhGZEO8VjyMtThgMVXA4RT7Z2/lXDg
jZ3Um7a2JIXjhOxa8kDvivhHvspKawCcwYIN4lo+MHA7n98sERAL3KMExzCFsL7K
vyFYCkxuuSTIBpTXCzfWARqhsG5bGsHRvU4ODBkFLuGW7q2msdTlTPKGiDzVR16y
ar6mcg4jDPi+92xJ8i/qT2k+REaMbV5thyvTs5PW+0hdPr1rHq8U7avpebwmFtS2
lSOI9XLmYX1Nfoi/1JpEvwYJC81pIrdt2NdjXrWQeqipDg/sWvgy7r454SkrlQfY
E9FVH42O+Kje32eZZ988zTDflYvYJX+XpQeWdzKxDyjbdjBr8Q1FlQTnvOiSRtkE
jHXo7HqzySXivXcVlA2t2YzllTmre98g8ilvEkJVWu0qS2agoFhZnt8+KKu17lID
yRX7U2WCMuktzKx9A7m3zxG98IMfa+2gP41WgEQYRrnfqo3epvXKZ12pIm9uU24o
MQbQKTV5lLK5sWwILRddwRW8mzbdEEJUvgkybkYYDpMy1ScNhfE2XLIzv/3fWpwi
C+ufKA4T1GqS21GS0HXpF5PUkQbE3zZmnNVBIXh/0p04TLtL1QGb+SFrWh+dITnQ
NB31/lUkLVsqfieHgCEvyTZb5rSne1vR30mUl9Yk13+DLdrep7QuLj1FJj5K4pQN
M6SoHP1jaGGWH2VGBqMhaPK7kRGpPN3MwNUDHg21MQ4cXUq1bboSfOBkaUEj7bC/
6Sor03Mo9xZ7DyD82MBV+XpUO0K65ZYJTtT+hO1ek+oybe++pmOAqPHCHKGx/M1w
e+MH8vDrU+N10/0uQ2ZiDvPHL8CPX2RESnPJhCBzQnyGP3Upk7yXQCMYh2mU71VM
KlrhnVrhYp2WWi5feXCKlDw03y59gEJhi9Ws1klwc1mNKrq4FSFruQdrV5/JQ7hy
t2pl9Nnk6lowFuxWgu0Y3z4bHAwZcL5IIZ+56xYMB2U3Cv1COSpGCR2zT5Qwxog3
39KSaomYaQrfJMJ5uGcJ2beJ297II5XC4IDIuir2c1teRHOJQav2+vrdiZOryNPb
yTh58EuqJmL/ZpDMNCUtx45zWxPW2wd2qa9/SCRemsSHXugQCmttInw6LnlfV4Kz
NEutHqlxuOowXEFPKDRUaPRZFIMhA/nj0tamgXKk5NwQjwqGyogNhn/vtz2WuxIE
98titkL8Ga3JB0K42WPktVayhCCcw3IHrkAHFllOO76hvAo4Llq8XGYPfYabY9bF
Xx82T0Uh/CzTQD+8YLqoZJaHPq5EAD6UPnQKkIkT6A/v+tnTlj4NVfOsSiceXf5O
yFi2OYhVmrtcDvHAUUVFDhGGO4Q4yOWXqLmgcaIQQCQsGxj14iqE1Bk4u0qQzHkf
Ls+wDO4b/zf4tsR+pDQgQNi1vKuKynUDeC9HOEEaOk1EdMaWU5jJOS5z0qS93PqT
bRrXr3Y809jnGDWkZf6z6TyD2epf5lLc6SlO7bnjxBCDMCPMyZoN3g953vumFQmV
65OOqbGVnV0l/ApjTvagdhs5tQxMXa6z8qq/G9ubEXmtb30jG+TRqJUTMmpM97/5
uSBdvu6Xo9ccCvdA2jM/PKUztX/8q+UoNOMjtqjfFk3KYMzFAQXojqKzpJP1fz4z
tb7AOMTvdIVZaJJhy2DNlfsgpag3W+EHD8qgZWLqzDGOcw23w1yEJPm6DElomCDu
QDpqY9NlqMzL4EJCjNAn51JAvBzlOEv/8nrs0uPs9NfcvyKaZ/tlw00AjD37d7Rn
kHg7eQjEia5lDnsfSA5LL0h8+LHU0iugR3dljv3Iku8cb2ZjMCsF3MZW3Pnd+jDm
H+f4W+Nzcm//TdC5uAc/qo1vkOHDmOSTXBNNSZOjntPSCcJL1RoSalROK3Myy7xE
as5/Go3Sb1QHFnjH27hVQnWV2ECNoCW7AGmi/tSZADtR833dJvkI4+8DwQnyk9b2
YlLfFM20GhqqUZZx9Y46tnE6ViUN62DgQjDnYP4B4YV4u6Qc7c2SCPGxpZNsqr7A
/ym4wQcFmQDmqZrlRfrteP6EhEEBTlviEFn3NOp6+SvvEkIluKZEQNVWMb1a0Gzy
7mke3xRozBzFxkoBtAtGuFWX6Ct2yGAJL1A01IaSqOZ0joNkO2VMr5LKMYEZf9OF
bc9d1ytEcspcYHwpUfc9YFyBgro6vioWfeyEdla7fwwXAmb/AfUpTPyUC7oaw8m9
orYo5UOhhuPo0fRJzkYMJwL73jm0HlGTUkqg4jxAf61nJholdi08FZUpaW0OV/lq
oP7+Y69xYiEhAIjdLf4xixAY5shfTKp8WUm35EYGKtMMqVRULtDb0cCjSr05tcc2
U/rBR+r6EXaZhwHAe+870+Y/p4E/n28S8khtQlIsZtcABCB6VSMQBCudJIPvcpPq
2+FWu8zqo7i/vcJVeCTP+avoDk/xGCtrTAZR4rJZ/Ky1wPo+PTgH/trWenE9kjon
Ib8fcu1TguwVs94NYns59prSb4C8GaUAZ1iHE/zR7kTm7aZbrK+JCM2XKiCzQlAG
ZruG5c65cy/YRx4x9HkHIJGkwcYBJor7ao2rr+BNyr+t9qQM3jQMiuJtqm6ca5Uv
n34sMlMQwJzSFS3QQRtRc2RXc3kNj/e4aw0sjIOjPoWmBft7HVKniT5cdRE38ixy
gKPdz9zsfQtCMELpttMT2Pt4rfTwSxHfu1pb/feOyK2lXgLdGr6p3o+MvxsqFHuH
1/USWv3LJGZuWtBbicbPRsHMbv5yxlqLjuhnGfgnAqFBMA86Kor/TbtY7B8NCKsv
GVK4Re4IUUDcRA1IaXJM0MWYumPKnYGxf9Ehefqoh5sIAfDpc118hKl13EaCoHS/
qAxJzeRJcG6E89iGcg5iI/tsx45hKJq+6G2rrIwtXlb6t4/gM6MXAbKg51yxQ1bR
f3e4u2Q58Y48R+RBrMFVSz6UyrVHcUM3DXP6cYDCJ8wtIBg5FSxhGVhR5r/bCz7L
ut4UiCAK2awE2SXnVuWos2qeU6LFWMKne97HUfryaDXb7Mknr9u7/oiC21dArnxx
N28WTkjFQPFGhpBx1nQmYcNCBE/HXA+D2nPR7mwH356QBkeTMf4qo/YERbBxFTyG
JhbHZix3tPw3vBiBddkyZfWalcD0iUAaNXtB/RZ6AMwqAvlFJDIVBkCsJQsV5WEU
7WKGnmNlW2bhUVqLoqBngwzbF1KZma4g7n8WtHg5zUiMK8wkSDGzO4ZtS5pRnZDU
zBRd8NyzDRw33TFkSGZ6YRyH2BWIxQp94DXE87bu1eiVTE5W/HXG82BqaDtx5FRw
WG+C0tvqXGu6KElolvUhrpQd6T65LsBOHgvnDO6hlUPAsN7SYg0A3QV4mJeyiFu1
v+t0E+EKrA1E0GBG2tLy5Q85KUQos4Px1DVHc8xPhg6ks1f+hK2OaEUebUR99jqZ
D8LRHErER7NDWPQ8VgB3a0HVL4ldkur4MHI6xSebU/JTbhnqIGpPsb2G89wN5BZ1
4T92BwZVLZ1qw3sD8JsJMuU8NHy1E309Io4nBd9ScKg7ai+CTyhc/YLwx9AL6hP1
n4qI8UGbuhtS1T4bO/ovozlyriRhY7ZJsqpHkg5ugKndvycy37zYweLsgMOk1t5v
Db+muwz9M1obKjgB7IjkPIDxZYIHssum7AqTzUwugr6tS9Htso2e40f/cO90wmjj
OwjgzHdYWylYJLnmUFYzjhKSSdlNcRDmtlKKGc3WxLhOfXCOoozZoMHO0S51JwuW
2zLiUV4zCHRse2H4nfVnFKcewdwnarGmSw447TyUFsSnrkVnCY068LIdT9Q9IL6L
7toaYLhmVjosCFTtp4OWD1nBp5zHYjJ0L4FRz3ZXI2qh7vNWWHp5H43hcwWBOQKQ
3WJFdUH/2gSjTG15rN3fwKnp+KLZPe9sZCjaL8QDR96EL82tHXPSuJoip9I8MTKz
uApUC8j0ZaKgTbQimw83MVxcOETqN8AYgx0gnuyFCVUBIgPBMsVrBTtnQMDyXS1g
xRDzEHOoiF6z1vnOQv7ZrfeGQcmuzkPv2uYPkgs1VNj2/YpWXO14VnS+vNDBZJYw
zNQyV4UAabVEGtZo1bxPnonUnv7zd3Y9EAMxFXwXrmRH33/gYKoLp+bA5mfDw7WR
XwnkpM7ZDaIbAynmq16x4l5LsL6RXvabOSQpir9FEqI0Th3SBfEhwj4XiiLvcIPz
PL2vNR20FDcAof4YEHFqn2Ht2C9X1nDO2puSULlfujhQLBgFNyoMIJVCQTB8Z40+
MSFIwgQmRLDnCnZVjIPQf7suYx928XZvKexF8blWpbkbmHODlPVxEzhJv1MLY5zj
b4nVvUjhxBNX+1l7mFVGkfMTpaEhZWy+7L3PSkqA35ul5Jrd5EJ/GBZtDLzyqe9e
5B2jBYmFkEFFtXpD2zrAghFKpwWgd0GWDI4JU2DB2i5n0XB5Sm2B7xFzIm8LM53H
RDN8/rYl3uwCyAoDehweOZCM42k9ac47K/fUnOc92Z8KzrcpJ6ivrIX1EO0qhtkr
SJ+dTNmhWJdDE1IAkdFSIghpZVQslUu77PnFJBdHW8fD8V5qGbZVdP6qTSRIJoCl
HCDnXbETwMfBNKWv6h5rZkovI0hLJkX4+s7vUoe5CKlaUr6ne075O3pCQDGjzykS
g12omNF7HhClmmk469niA1rTFTzxdkLbkLvxwyrBa49DWc3UQbRHbpRO07lgpeV9
GJZ4M+Anj7bOH5uPFMWaQ5o9q8hrUCuGo7goNEj1vlmIWlaJsGmVZGkPU+DNM720
/0bIJ82Vy1wFIasb382wn5dTaJT7r/puuDv+ifvYN0UBrA7zpUx7zh8nyKf91DIC
gNYEhXeANooM8UEFGq930wevtHyUfW1EBTL8Dvjzm7MeKSxShLz8lmnbA/MqqPLP
sEmql/Gh70gT4qWd6PVjNKzGU4v1fKF2GdRSzT42TlygNFa1z7QOgu2KfI8HPU6w
r3FOw1yvhM8NUnyNdseOMIFjw1rU1mny8BjCmjpHh8uej1DdHKeLKmEpbe0Hkt3W
KEESKOw7bPJj+HKvg0ngtGrb1DqtC1x+PZWF0RpfVtbBxeJRnPvr7i6+NRurqQnr
OMXYxYXv7TOH4P+9oEF5+QZB9F7oJ9GTJHBfSqzZIQ6x78RZYv6Xump/BgcFKlpF
JUPBDRFTJ0w2s7XIa4vUgV3U3Z33v+WucfpHghA0XrlLmrJIVtWS3/z+Qs5pKgwO
zgLPTKrCFGzxyTJlUbKAzUO5X11m41Zcu0y/hcY+aB7rQzuoyaYV/ViXDmrauLWX
jyYwihcirSyRlf/vdh2ga9zm2nX3hDdK7fx6a6BKzR/JvhvcaQ2oAHAQWCy7i7TJ
ozishTh/MvQ/3OK2wNaE4xRdWd6fWRKkJ5HuyMIfBzUao8g6RgIHyxp/HwosUJdN
6yk1XFDZLCPvgh9PFzfv8I2aVrZDET1oASmfKXHFlsVYvuVObVQHY3RlKIs9cJry
ITWir87GwSleY3UmubjcKxEHKl8aICAlzh09leG0kiig+F/7J6n7ITqyu+6P0yEh
Ga031zL4ztTTPvRQz80x8kjZIdyO8rya4z/rTppPV+2pjXkcsQFAWZzFzXpNSY8t
7Jbk1hkdBSO6Q4mgexKrUufzxw6gdgJpzXAs2UYpxk36kBWAw3sy8LeenWlOaeSl
yPEi+ZEgg2QtZyCLNxokUjCXwWzaqFPWsVR/AHEVuJK7RfAfbbgijZVu9ykGv6kJ
bAYeMBb+bbx2lE/Dqh+AqX2eg8miLJu04Ty1vSmbsWSzW+PobVm1orY23j7J0H16
yqMbYOl0BlQKX0bYlLKncJgXWWVD5I3cYK2PJh6y3fhcRFN/XXJlAOLVNU9h/6Vh
932CxrIdAKCnVhmv57yz3BakC0q/uWV96a8lfT7jAtUWRa0DW1sfdnKmKyG26UbE
3ZnzfmgbG4H8qWgkExap4yyuLuCTgZDPV5f5rRQrnBt3VrkcR7Lp9/WwAkr1JhXW
SIDebZqYukrgOt9NDYYWIXH61ep1dKBTdabpI9X3uwhQ4HtGCE1HEInoj1vcdrw7
+u6JpQiyRv1ricZ0d0YASSZW9sMYB26yVSPjQWAmi0v3aB3T+Auc4eq4gg+NGoy2
uvCbkxl+pl6Oe6wp1SFkxF3jWCAb0upRX22M+uPz+wQjRlj4iW1ZI3oILIWPYrf4
9ElhCmhfsgU7a43u2F0i8TjWkt5AIHk9ueiQVcAJQx/4HF+ydSIzpYiLR9S9gIbA
a8C3cqDO2eSmqLbpeC7Hz9uJaDmOLKaLYEIUG6b6vi7U3VncOwpHTqTs1lw7f7m5
uCst9+EIqgBwJ9YVj4QfcjTTuVTAIj2CFBlpmE8HoO6ur9U/ZaObSKQRua0BYero
/vBn23Ey2bfoLYLjpwex5IsdWHOoBM4QcgCPzNci6ihXPIZlBT+ru+c4HD1fVuz0
/Xgfy/xj//ka9yOu5MQ1RQANSEWGee01FtxJTUA5wEqnhRvxl5tTgQ0Paekauu1D
mc3ubhwRhnUHMUnT4x2lNUzi8UfvV5kZSMkr0Ay4D4chpfBLslgOq5rRo2/IiLsM
KKLTWKppQyf6ENCL54n5+r6FhFlWozVVrGSo941dazySava32N/cOr4dAqanqp6x
jKWYoF7H2ZX444bh1+lU6NDza0+dDdcbYccdNLUpo0QXmZF8OWiVcYqEsm83KElz
Lw+WtBTwFRi0iQEIwuTp23tvecVH0kCsmjOurv/WtJk5CdETji0PVDTuvKr/ovnU
GGG2ihfosHYk2NcQOVMZcXmylHtAIcVLJAtcWm53nO9jX17HTUpJUnqy+7r+kjUn
/V1E0PEekMTVQVje+HYidU4D6LE0U0BNIgwqq681UG7bu6ZM9oy2oRMeF7fusNV9
WlRjxe5syGIibRhyETJI4bCLWz1c+pqUatebZjhwdDUDRo1A5r/4mYIunkNIxcQl
u9uVKvtt3FYFzgTgY8/qNwexEyUNK7woUaaJV0j3XzCtS2kHQxy7a3v9czBD077U
rZHU12e0c9lxc1DaI2n/bny4xsrqUHl0r0JsYTfYhFu8CZ9Q886hlrS2/Sf8jBel
/OieydBSctI4tHSAZ7hLEX4pNjTuUPyZ/e2uwgN4WAG6cSlez0VUdN4ejaVCquAQ
l6537D6sClx5zUQr+2po9fe9YbfKhIe6V6m+IA51BbiSdae6fxRR44hpnPsoDl/M
rjT3M5bnxU2EWowe+O1BgAbJRYP+bBkzXwZs8Rs9Dj51jL2F7B79G6Mr7/Qm33sK
PZN4a4/a0NKFoqHzIlHxUzAkQ6xnkvwpFDIbKxW7UxtGB+JZxGptCEXlfD7J590C
gkTt460BCES8b7RP1mc+Dex+P4U+fApFG/jBI5umYLKYDtKrXNpFfzncSqoq9Lk3
5u3VKtlEEVAUR5/XWLdRBh/Ptq2apyBc/96XHjwAJWqhHjOZo3kYHuS0pERp7jSG
pvWnG2WGok/YZpIxrBsrmoE74sZXh7rnvWUCEQNKhtDxtK1xwYkRBRME0GWIXpXP
hQcePhHoYKLshGc25HHPQRwJ4TU9kMFG6S8HyJVWjUJcRXmJ+flnbXRGFlqnbhbp
7SRvM++/5v9Mk08Isoh9AenyZwSHjKYtJ09fz6pHBn8mwcvcNHxdvOJVM3KwjvXC
aOV9ai9LwxixXpWtVxo+ZPVLYbQc211FjfSAssgfDvbJwV1oR7U5mS7ilSUeKZP6
L5Yo+UfMX1lVk6TA46PiggTcczNMf4GAwfn4rlRCg7E5tKzOpXs/ZrQgxDwO+prM
Ox0x4QwJqYXqU6pfGrvlr0DhweELKvFBtnxyAAtfRrqruYZV1wJStpON/FAudBtN
t16ZsjHmuuktDGj6SGs/LM9I+vy2k/0RvU6EYmZ7IAEZfoDkgbY8SpqaMAA1tVgI
PoZLH47ky8t+CgLgS2w7eKrqk9SPZKkIfgAy+RfBbzyWkuKYgHy3TFR+M62sVCLn
ifXWb3DVRbzwq7ORt27b4cljibFowaTkdxifhTkD7J6Ii+7bfZHSU8crxFfAb1na
L5iKZkbaF2EQQPZi5Oqv1q/3kr9woVBLLfwwSwyfzOmCjwVeYAcDY9MYIP9VYOTr
xb4c+vZxpJGalrdM9LFB52IU10QSHf2t+Dk6Mc+LSZqNi8+/dTO0oS5Dr7iacwS6
CUjfTrIngmUyRW1D6iLpHUZ1p/bmq0lGFYevnojVTGzJq+FyYorj8Xr09jDYPqDn
Y+Co/608O2FbRRb+F08A0e3RRMuz7+gJzWk5HYwD0zXiPmZWaqj9G2t4aPvPJ08B
+ujNTqPPFJ6Y9WqUeqWKliKlSuGkkhidjIJYPEKnZWtcQJduyZ06ORXWeGMt3m2X
ou/bShRpyEUsEuxJ/AFWBBF3smppfc4BJk8uCuHX6aHhkQQWuMgJJS3u5WfBQDl3
j4A0OqSFcvK9dmjr/a4UVV5ghrmpJ9n06iTKh4lKiBAKnOe6NlFLfjZI0ZPDvZBX
/M/XMeUYsMl/Ql7yVga5VI0fFjVBu1h3uDwYMSg7gzdHI6g5PMUY440U77tnd16z
UsG11xfX/zDuQKeZcCLvxK5zPX2B3/Mbnx7hjkBePvwm1Ql0gJC8IMKd2NS9N9fS
lcF4Di511iM4xlyTdixv8hXIfSGQkEWMq60OwxTKoM5uATcSP4b7taZiRduTtjkZ
9OF9eyDzHRHlkUrh4xHIOgZOdvVfgG8u+0DE30OTTgJ+FQUFP5OSgQ0QZ8210/6v
VdHnrPv2en4rOm5CpFDYyBnDMW6MQ20cMKLmlQjgNMRwk+YzZlkIkymQfXRQPJy/
hIezDhU41Th+qWhnacEEDYra5gAqVKzrUXvW3NCpN7Ado1nwI8MZk/of7fYCCkgx
BNGwz8Cyks+OguYgmX+xuZlvUZFuTSli29S6MWIYqm9bBhq54NQWzmME0H3X8v27
eUnkkPV6Zxe+ktHHv8fp2fdyFSEb3KhuChRMSqGaihlsxYa7Klg0e/+rSikYOCKc
ZspUnqoR4lwN+RmgWeWM7ATb70ku9p4T3h3tYN5SYcFeNRfY3tR1AhrPO+IzMJQn
92qiJiM/C3T8DsuLSvZXWyrf6bL5dFGzmehsLbIrSYk1my5aFlu+lA2Pa3whS2G8
idV2cZxsT7/KmVl78dYgsBpbRV/RYfwGzSOvxwyJX/fBrkrYvESQL+h2NvBt0767
AmkhMkpjDRx4qnnWdoGd0TNFS/nG5aYp3n5L1xh+bp1r4s/pvlhcUeYHBL2GJ4KF
HdFcsd4kzQYezi/JHRSPxycFRXKo1wgtbFa4GJ6FBhnCrgy//ihZGNgBpB0IAnKQ
/qwdPtj7kaQSpuZlyd37XbL1sHX1ROTfGNKKn4HewwYk6Ier5zgt10crnEodFfrX
l24d8oAGOVNOE2BNW5RF3EkCyD8zB3Id/LKWGsqeert+1ZXegiiWif07zxVgbWWb
4RZC+ZuM51ygHv3wVjc0RIH/521vpQtKGUJ8rK1aDIzgQIUhgZu6ZGrEmlh+j6bK
20x/4/JFRwoxiGw2BabKs5k04RguuHlWXvyBEpEiDwq2Rg1dghqdy+BfMh+9P4IG
KhrKdwU5z6PvAv3o1EZMOPBKPjrbnNXPoYyoxBtrfwt8EGbjdsUL1wUqiVyMPdCm
PLxsxhVL/5wFr1JMA+7fyzCpSIhyjfCjLHJbgW8t4ZF584eGqbJizPfEu3SHF1PY
/i39yA2HWk4dEfOK5iGcnIS0bRYIP1ZXsL22Q3EjGLx4N5pFy6CTARgo1IavKj4R
dhidr7tZIZ14CKSK/eFBZVjaC6P41qPqjcrlEoj/cYMk3o64TfKXXJj2u0mSs8Cl
Y4ddiHa5iYHbbEhM5qaFMO1Tkz3CTp13F1x+AFlvP85o7/JjGECoRFXf9MUAS4cU
HbEm5ImSM95APS5+IQNShtQGSoJdxl6GUBhXhnAcT6lwAjEO61j+paVQuy71ltp/
0l8V/S612hEpjrTdvrOgcqttzXxkrSn0MITSfU9cJTGlBxSsqIGXEBaCbU/uBq3u
Kqy2UNQW/ka5P9oPTnwOcXK6mmKnJXTomXRURpxACW1IrXChKuxt40/ddgrAeOUO
9tsHG6LFxd8CalFLmRDco8awbP8zvpfGirPjlwL7Jl7+xFQ3yDvQnH4gGBMeWVqq
mgrApdH7v5f38jZjDmRGi3BvLsM12j/a1qCOom3LMZE0I7aIsIpsc3DaN/IBGgju
Pp8LdHsLbwBRB+xdG7sx5gf7i+bSQrmS6BhNRUKDfLEsyiJP4ou85134sXo3JQTn
Zfw9t9VhDeOf31xqKH0Tm6v3zHD90NMk8Y2moNZs/4BKcZQLFIAmlgHHPaPiUkak
BH8Bx7sz6fWYWTSy3JfHeNa4909NGq6f/hRnSTAzVY+PaSZBUjutJUVRKlFdN9TH
qhnLEUTZP4Ymz5s+UNd0J7wcyEHQe2FRRTyeuaeutzR+LaZdHt2wRt8tqxM6MXmX
oC+kpYyBs8RsQHZH/df0SUcuv635of+8+d0zhV66wzkZ1+3M/9SztRqUACDZqrWA
+HuWUVSwPSXtclkK5u+FocVPVu0uQzcwwVhTU8CgXJv7LZJojXYQXkg0MJWFI1b+
u8ejkD7f8qWsFbjkyMlVT1zKVNmgREevyAdL28GMbkXG3GFI5bF61Tjb97RFFigr
l12B/zdEAFZfv/U1cMZvJAztIVgF1OmRQagfokr+qyiaZ21N2QXaJbFPAOFnA8Vd
m55oBkriyqilD6upEL1hivrQmyrEBY9KRkSKFOcGjd0A+b75WzbdEwx1hounUbSh
GfiOg5O71XXs+LvdyIXGL5ctw+52uvOZqGci7eolnXDIJXwrFTifS2ff1hiCJRhO
78MdE4XfIrWQCwCQM0BP50y0GfuW+X1z5JW6zYswRcefMTW7VFnJ/O6JWEamh+cR
LvxrOh0u7byHQC7Xs4w/tkB/on9KM4vLVqU9ttBn+kD6lfWdFS7Pg+/mXB0BQCfP
pQoLBx6vnoa8dkCyeo8xdemCkP5CK5o1+vNDGlxBk/ShulpXsis6lZU7GNcH4y3L
MsvrN/1fG3CP56dHlElfH0zsH531TqtBmJQaAu8IRrmqKzK51hZTHZbIy1z1qB6l
rcZpH8Y7O3XhTB0vuTuS4AVbKQvG3xwzhFguDQ3tCCLCEeyk0RUElHQNPfxkjZkQ
2zX4OeSR6TzSBmRBPK8XdjVPM3Y8qfxeMrsBs28WkoIIuWnryrLBgyDlXWH6M7Cb
hiyUXKq5idIp9B9xRZh85DlxTeoyQ3/r2KsiJh5lScgQmGazfTEhxkf0GBjrpes5
MQpWp6tKFG1xae5Xw6VYa7q84V59xKcdfQAWZl8lPBPlHgJ9M7cWiQg8MK00xTgv
t1iKtC142JRRt2PtVpO1KsgiIKu6DLWzBRCx9lwM78dRsJebGR7IFC+1OWfmrGmF
ENd4YCEpvlQBncV147UFBEP7G9LsyJB0NaDEJsOe6KI0ANPW6zXY/CTGARY8ENZU
e5yFifAkIdP8+M2LTJrdoRk0XbPT8zaq+cPYNYi23zLlDZm5fs90gwn6K/0PW5mK
rbWBc+gz9U6oNmbYCQ8k9jmaBSURupDdJO/3SkwT+fZEWGv2+b5KQTZzm7oqvooW
bU34WoE8tx2Itr7ewK/S6swJ58afh90u8vaxsEWntsFTKN0LTH7ZmB8YLDGADtLI
9OOnQTTKbU9LqR2yiU0u0E4jU3MD4eib2f8vfKBj1OmILCRRgWe2rnKBQcImDjBf
EkqOjOMXpr5Y+yRNI55IhecZgx8tqTnb57sl3jZv1BJwjk2txZZPRCzPtcnv6ZCJ
fQ3zNNMh5IuVvTxvH8WrOZxLWR1IQv9z1S5EUFKscxVTQ0p4Lrk5xHBS5sRrKOeY
ERMaEYYqIDHKXG5FWEETKF3pPWpZzv/wm61n6YC1JonnIIYhvfaOXRs0EaPOCt2a
cPOAl4ZkS+NFpWVcvIOsBbp/0F+MGroTaIysMByHRhk0pOuEa5Y8I2lCmapYDGDl
0JbWsfHQOoElh6etp/jRgwwiFhvQ5PYc80S5CNC8+RxHrRrhSxE0T+6wmnBs0x8c
ErqPX+THW7wLpPMFVF5hlSbc8KA9Ir4fu/4HbPLHeJ61aaki3FxV5uQNCWRz5fAC
jaVx7V7G5iogOS25s2S5GJASbR0lNKBsHXZ7+YjMaJxJP/NJ1iE+f5A49d+MweRz
4zqlLc+8hc7I64Ov2aCqAcCOPDh+8KSptdBj4fq6dm8DRlE40lmPYD9tKnYfLDBq
mpMSc2dUpFIvEYxUJsAiwslfcUDoCSPazH5CAxm5VIBFLBV3/oMbm/J4blfh+2qb
H/wH0A10AW4JFDO5w0fYn2wOvHLOjm6G2fkZDwParfgalxWwZRVERn0s8oswdNtB
nled7AAIHqhE4o8VB9kvm11uVewm7NFnfO8WJEuFdIwOhcyF0K4X0f/8rjYTdVZU
tFi5dRtmGHteQWxmQcljV8V4BlEDN40Ld2mfCRKImBfnYi3Ih5Xexff2QaTk6V6o
NUaSUtSS6WPGndnbea5pd+v7lRqlEg7xIusZJLWPjWgEBhhtKcBfSgo/uS85zQv/
LFNC6dJPhE2pNFvHEdCTo4KtSqMCTAl8/tAB1MwNYHOdWr8dtqQPuqicBuiwcHF5
el3u9DJ97TMrMGt9kxfZh+dl651swa6Vt/5VPV3/geXtiCHZV0GQ4AnG/ALEdxZa
vmGN+UdrzT6RAwXf+J0CJ6QFbdNNWP/7KZTPcL+E6XVapyvqRJqSJoApUS1Slhdn
VVVquBfZydWXRW4fyqehrlmezw07YpbtLl+1738LUDjtN3o0+bCenkLNjYr/hHxH
ocsdi0zqbf/OOeKfPF6GMr3XnS2gFoMFvHrI/JUgvWzLh016cJyQzBgTyfXh+aFs
rmIUFXFlkZIXBJjLovAf9ZbeEIiDNoLSD4eouvRwpOJsnhUji2xQfEF3cJtk7DTA
gsAv7tMrrAvYjUfWGZ9I7mW2KaT+BZLNU+kcaplKS7hywJ2LFwAPb3HtNokzCmUl
tsM6ImqcG5HL6ay4HTfhea5xWgLJD6u4FGZYU2q8vXATkwHkArXopvTu8NwixjsO
hjdgG+EZj95ETbmOdZkbCvxkCMcwifKlZwYwtHO5tMBYbnH8S8TzeKZJ2NTPECEF
X9KNyOdWbeKIRzIcmdKKfVfFeRxmszURNJUwCku9mAM5VnIBTmkU34KkUCYaLrpw
s+KXBFonMQlzhDV22/odUV2/IxAcXKo/JWntFcf59jVHF8htlwU9ktknsfao7yGF
I+cHXCSXJr2+pqcuRtbnwLobj164ztFFADN9LoSUBhT9Wqs3ytsCgnnRPS8tSo/a
afrzMCDhq2e4qluRkebmzebB3ksIR8TdkwAiv9+WVjDlF76kLSGJsXx/8ePTmpDF
pgcW9iL8x1UwaY3RmNI6+alF9SR/FS2+AN3OZnZugE8B6zXCRkVoy6Da60IQbiJ/
mmYy0CyFhTxPwak3DbZa7ZcApfuQ52dUxhxUxgK73LlHZDp+nGvMNZqmstXwo4x1
V3pEgIPniqtYDHy9efTm4ofI8Exm+MpHcS3uyZX7Mwmncwm+v08NF81TpnvNeYPP
7X5dm215cOaAfry9+5gyjx0YJzg9jvLFQVTlJqNBdNla3WPSJTz1nJ6iYkFGf/0a
Q3EHlN1/a4JmVWN4FXtHN4qaD6DXNvakcXCuPMvL5Neixt88hyb1gT/P0ervk7rs
lEzJMIKMdJIAKJQ+A/6+YAjIbxvMje0bA/9h6VwglV/T25gppBSMpgDpXddWRkW0
IqgXhwZLeqJ1Hemr8PIa45xClyuoqNfFbdIpdltqiDBsuj3K6XQa4IOHYWVZbySn
Cl7dAJ6rTk6lnu0EPXHmH/QmweiVd0pqVR00WzG7fze40DuThQfUGAsnI374pOm4
9THQMStsJhgNb4VMY3l1R/BhZp+fQAlC4N5KEWHBpg6P5SCu12cgCR4JVfLYiBuY
TTL5aoOZ8aIoXda6P9RXqbW/MNAm4YM27KPRyzxBQJUI1mii+ZAmaG2Mwb6iNKrh
Lv0DLzjFgqJlkW1G+8toVZbEULKurlpuV4oX8e6/ZIcopKhTFBXifiTPWuj8OaYF
hLkjrAhcQaEg5Lw4rwUpnYkyyuGwKvMAAA2B2BuuwzHApR8xkZMx493y7pP32XnM
Kwf0WyaPi23X6PLazQ66zvB5qs9F7/QzevBldoMqC4+FCMUOaLvKGA4sS5zanTZm
20kKwaDuCAVZcHHWgsbAN0o+RXbRqLjPQ1Fh4GltZkcOego1ssXQkwIjX4fW+ZUf
D2CsOPy8J1yyRXMn5XuER5BYuNv331/DY3ndSJatPFpv62C5CpijoIfoENsheFbo
rsnLUbMpa8fLU7+nf6P0OXzXuuAbjXm+dE5n9BNMoy/qCr1J83MYK9/K2prjUfeL
UywKhyhGtqVZKzrD+oueigmEzqANmQ4D4phwHd4NtabRCvyjOatTvhH7IdyfMDHH
5ZFf9Z3cGOFUtVV/yRFb/wWJUox51hGkruhk1C3sUdtAe01bp0ZONmgpCWVq+j3d
CVmITtA9Q03E55zIuJcaAyiD60kbVIQ6Gn9GG/Bl1InocIOwonOPpkWdsI3QzdjY
n30H6v+zBP9t+bgTZQSMl6K6iC2Zuhg6oY00ag0iJp8+jSNN/EbvOP2WvglZPiwz
PurCHwp2jP073bIqX9FrmJgsdwGMMn0uMdN7j+t3u3AmJCf5fPGlO9BxEy4BGgms
NIsbFcSHVSTO2d8Rs7tlzOrXCJh5uf1g9pPRQjiNXQJYTdPLHdLE9zfyPcXu+maT
+90WOfbW76hR77LxoDRXvKZsiC3m1nkRfT7Vu9CN5J7sBVnBOUWslDNPtHWqUbWI
pbClpcIJf0AKMnOEN5H2TH2j2ONTYIb+4RzdXq9CNxRTljviu5jfFOg0n8ey4KWR
S8iuHSYauaHAEWh/34gljV7SIkVyGwdE0srWrGwLJayJwFea4PRdmsPRWLXDk/Ym
U9y8mI5xuiHet0OA5WyzqQVZ33C+MiHZ15lwmQwnsKjjAuRrPhH9Fwva/4x4HAsg
zdVWzR7plJv8dQjH+5JwXlfCuBt9haNm9NYI19iUjOZ/dXrDrgkgsdyBu8CQ+caT
D2XmNeDK2wG82ciz2fXcEOj6We/m7IOmQ2iMZDFB24pFTnTD2/TUmJXAHN1+VpiV
kaXBuAZMugjee7/ZAp74J8StzHsGensDNoNox7zR+pr0yB7mRIUwSpwc2LKPaZZ5
YfsDhDQIuNYprAOpoME6so1/jWqiOJfb0+zDHmQBkeRq0btsv+VPwbVB/sc57TaL
H0EzWTfslCUtSuPwlHPgmFZulfU6Y+qRk2bLankl3fZYC9SITqlMkrQ5WOdvqAcz
rnoPr/BTRxP/4r7SaDTMR7xdV2xSDau36kbjr0OPAwO55zB74VatVnUwl8Qous9Z
fLe3Qzf5MuFzGysSnwQTQp89pi1f+G/F/3qPFn55gflyxhe6ummmgdMuz9Hr4qRU
g3PG1NO9D+LsedCNcCgnMb2aUV8PhHp0LS/WQ2uT/VjCFvCoWLlEdEwbhRJ1a8Pg
SJzGRoq4wps/8lnJG+DgV5BoazxUiEovqzl06gb8jXSPioC8+NtAh+hHzRMm8JQs
kVnnOd1AWL/Ym1yraoy5rXn2VDXer8FuDqShIOQZNoOS2en4t2zsdJ4TopMDGqtl
bBlt+WIdReYhjBWopVnQ/+jM9RuP10FqiYB5tZoyebls7U0JtpXCreIUUTvZYFE+
MSquemrygn1qi1J68hcXx6yq6jrfAa7NRXqJ8gv0OUvHp9D+pqqANUoVIMrWdUBB
CfOJgtbFMph1+K6vYxXkMP3NTvh8t7E0kKx0xnoZ1LOrQgpU+dISfv1qkmS2kx3e
fPWVtdZBpL0W6DLK9Khs5UTEb986I8t5eJFPyxI5gRbagnM8WNvBE5vA+6qy/Nvm
mnQDBQhB35Cwv0iiDXjNdlEfigc5P3HNg5J+zDqHA/r//94a4dOXaN7ZBmm69EZ9
OgPRMswyaiXJGnY3JYW65hsW/WpZME8TCSwj0o+b5C1KW+woLmDFOQFeZDxwoCGw
c3mmq0Fv9hiYiXoxnIMnzp7YzekxiHdxzn00i1DcAKFuBh3mNg8FIk42TWtponOR
K5wwZCawrMpO3qxMaBL9kVnciaoeS5iK4f8a3zJU24cppKyWxcNyiHitrSMbfwLr
5vHQamnbfrfGyX35sh+SC7sorW4dM5AF3RGHBi936f9pGRsWq6edslz2YbaOxaGP
P22YQY9e4gLSv3UxcI0ngrnzWczyCOnWqkV51DrflE/c8IrikEOwslyt1ETDSR+O
EtFecHSpctEQxNg6ppKG3Rkr2npFaxJLuAsDqH++VvixkBGM2GYuikj29dtr6/eG
ellWWWMnc9fl8nd8fW1K5x/K2rMtGDsIHy+Voi4+2M2hyaBvqchDz+RVvkvQM6DK
Scj4JsDX7pNBMzxi3Esw+A8QqdUK1wkUfRSG0OhKWRG+gQ6I3Qvz9FgGD89eJEzI
mcLMsDRfZVHE0ttoZIpC3JTUUDOXL9wSWsQp6NR7fPIGdycLO63cSZvBu8kXNeG7
pHIaNxIpJPC5fYAd02vEKs2K4LCH7jiwaRi6715BOZ/z5mSBk2aP5s90g4XXE7cm
aNqMaq6iGtu9RJ38ZLkVpfR523mtqn/CxuZyBtDbnM070d+VGrw/CdbWegeQKGld
P478yDygfJCV317LQrhZJgchIgF2aldtdUjEwKcghpJK6nxrUbRNYDMxusJYW0+W
jrVJMGKOVMfv4R3iBhUCSo9yP99Mi0UFe/Bif1kUy/HeSiX912pECgyNpWHmEUcB
ZCLdDcWSKyk0mXj1gZTqdow1Sm1a3grzCw/gsATxdjvE1NPZ87GbEa/QZa+5B7T0
+TUG+/GaTj3uq/BaoeOieVlXKXeouupT0WfbySUd4L2Qsc6HA1IBnz+pk7DrS9/Z
+ptYFYgVTIWJkQDliHgXCiHmy+Z4/wQfoUv9bJi797DPh0efuMjhAKBK0J6wDo3R
TIhoxZkrVcbwytvIFCnRh8Rj8otArQ4tuEEyxTZzGiPXzPdDIV4EhP5mWPvpTxOU
WIfHX2oO1XQIEYyWznQCxfcJLOXQFdy00CKThp6qqDLNiRboPBGPi2JaRzRg5GFX
uBg1s4C5u8Tt82aOah1M/Ez/s8azjYDpSXIwfmDGgIszJDk+PNeNXGHtCNE0nkyx
qxNAmkfJjK3Kaxii5zGU7u5mGKf63yS7SfuLKanniRROGXeFLsfqGzsFcREuZEBn
dSprKR5rO5UYZTnMKHxpONFTHtDg4GJEXMeI2QN8y9sg3JRwJwEgS9GDAMLr+nYe
X6nmQTASdTh+TyhOEOuCl8yqCg2yWR9llRH0cSyKfaM+ONbKhMHXOiSixjhHvIat
ZDpfj3vc/hmECR25fuVro+M8j5oVlUHWRQY7bo9L/f4Kvn2zTnwrddEe0Q3djcrL
vgrZkz1e6Yf1LakIey5UE+esm5dVMCZGe0kos1mP3ccJzCC/ATfqyQvDN2qomzBx
GlQfJiyi9el6z6nTy06hVjQE9jF1nYCtdF+MHaEX6Pq+Kv7yIZWjXSDDYG+SmoNo
M5VQLo7I9Fudw1Q5L4n8h2ejdQ72fddBIi0Hdx19SGLndCsKpeJoEtpeabJXpED8
tbcaQ+cdJVDDqCQJdXlgTEG7hMcEtxvlxfITNZhGEaWgHSKsT7IPBGkjxIs/P3xa
mSbEFvUW/HQRAswp2akmW3OT2tV6K4XwkjgonmrJp9DfmP5IUqkTyt5kCgLtvsDA
/YHx4XScsRhqofRAGO7arX7ZrGWa+Yz4gMP4snMkNGdj+jVjsG8MBQ6RdanDJWy+
MGw/1uOy7bDawCGC0guqSY5pHKVv/AESjMznVuh/87mQ6lGZeVfjwqWmggxwST6l
m8WSUlSA2ZPPlzGrzYR6acBUz0TkkT38chQ55Q4qh1jctgN2iNRN1LuAezMaSAOI
7wpn5SiA7kiUukLHhiml7Q9Hd4aUyvMpWYoCRpDjLKMeLQtT0v9Wg/MgdniIKxE9
XQvmkOPK4867FuAZkmr0p8fncnAVeXy6OYJGHnVFC98Df0ndzx85IZUXxEpuGPK+
6HjhWZw5R7AFhEsk24fI405Mw0EqqpNkdn4vLUxyJnus9JbMc6jTbVKGvmm3k9Ne
zFwoZg+veRJrOSL2Y+7T7fnKIiWlJjeGb41SQtCauXb1BsDdY569bbVSy99z7aqV
tYy7tWqPpf84CI+c+xnM6XRq3wpo/sahOdXRF2XHsqiOZ/5CYrZ6HpQj/f9itIl1
2Qq5WWUgwXyxDAu9t0fd79Wgy9ILQT/kwYQRiED14Rs6/czPVzBI05EdoESYpLaf
IjU2blRGi7b0JIFY75hTWZ+44LxYAryP9O9Z3nY/rIAKhVkRdVka9lWmekFuzt1c
/+DRo0CsOGgr9U5KkObmrnNIKj1ykAbqFrWvUk98ctudxOux/Rh0xDoHl1iQq5wy
ErV7nvjOREEtI+XvXh42rzHt+Nq/cI+VYWZ1QNVr3Duebk7syNd2KI3FD2Qllf6W
3Bjs9aCmYfWeWjHLZk9AuSflIMd6iGlVzFRkveCkqORiwwTeGUbRoPagq2l/TWqK
rW9QaoiTdKJbOyepwqcKIk8zZ7rqhrVzwgAJ8BTRU9wyv7+oTBKCJSvAFb4nU0cx
x5bTWLR5ztvx7X+jWHbaOltWfAHz1Vqvy8tdjyN9Sgc5S5TLa/r+PwVPva7213Cs
yaRluY+YLtUs1f9HDsUVky6U0CdPh0Tu+RVlPHLfThGJ+I5jlIPsSoilqfVCRo3g
sVbP5eQJrS9bnarIH9gmKXYjaSpDKjgumksKxSITSFURW3mJbCT2JN6okm5GBaEx
2Xz3ml7EDPBnMN+EBVsY+BG+4wHJD9C3Unh04LG3j2NMcm4iHA0lnJao941F3Iw4
zuVCPQeERVTnuTzgcNJgHXCkG0Q4WRhnLje3jYMvVSt96h1emoKoM/IoqEuHXu0T
PIxtrmPpQ6TCiQsVmINzaUtZh7Kl6Zl45zWvLiy3yjqAwTiTWE+rqU+oJVBM2QUG
XEM4wEjmA7advLqUqQbuyZB9bbLW3+AdAWVoLfNm3n0FP166yf+XVBvSmHY5WnTd
nXMRphMc4XAlN/JcRKfkFWOiWeERVY0YdRxa3SpemLWrrCrdefZd5YiO/l6cDur9
WwU8zcIpKSos+jPDOMTT8/AvIvB1VXWtcfM362fRYArHqP8e9fBvXSH7qFIP5NZU
onJsx5VB3sONmk6xbuWyw/zJQxvs9aaI8Apn93t6pTEzDuMVHsAWax8khB01wB0f
THx00ZDo1ARVfeK1zjtj/mWxrBXyTYW7a6bM7m5sfXEnde3dVz+xSj3lLId1yRJ7
p3KPn0WrrMd1TzFq3H4txTIt8stejJ4eW1IjcTuVzPjk3qm2KwklHxWUnAYlbsQX
kZfcqvwiLQ3qHvGhW5jfDJteYYunNUoYdBpuDlinRLidqXR1kc0rJp8p1HbUFBGa
l0lJD0oXYp6DUSN4T2egnqC43hF8voo7L4aQnEskR6+/n1/GYvOj8qM6KfDnFpPQ
SmTLJfyrIIMF8efA8/xx27l6rsqF21jOS0FMhOMQEJL57T4wfLLhbiE33j8Jebeu
PKRmUsIMv5fSuL7/n3qCuOK9FjwKrZwlRkD1aahArHTbEdcdRtD+f0kuI9t2eFOZ
z5xUNUdKkbJ6MSxpDXb1CiNZw1KPqwq1qsAq4DkKgfvtsKOsiAKF5aVL73n4Fr/A
ApNsikkn9jJBUgfzj3ub/pwK+30kqVCjycdv6H6UYsMAUEefTkqVq/mfugkGNt01
KMyXeO3XkKUP8uElC8snWRbdGWmgHJx43ljbOvu/7+bFvS09zsj6ZsktTwmLmA0m
E6JbXyE5yLdzaLxaEZBcXM4yJFDUYctVBffNn4MuiKtDS+imOqeB7DOXLq7dGYW9
7BVK2zj9yM8/mpHBQQekWheqdu4ckoZ2GYNAckigxvUmtjW3/JsKhhlOlMUMXc2q
PAjYkjr9SI3IZ7u8WGj1yk2UQOPZZb7jKfljH67qmCWOtPSwUsQvMECBy8qrTR3c
4Vm4JxR994d69652k6tfxGphCIJ7IVngdPHGlPHdJmZEHRXkh+9TAkbJhYmA02mn
KZrlQv8AxIx49sviqkGa/9L8mVTECtDsguk1ov+ZZunAiIc2jAEmmfWJelGH5Og9
Jcdm/pS/uHnn+zTJn+0+QIaQ1eqkLFOl74pwOYPxVkafk6V+acwgIFJbtcZrkvQf
XZlpjTGCOqel3jcj7fSslnZEVzv28ILIMwXF+glber7rjm+ZxjK5J08qmR5cDPoq
LE1RA4WLp3wGwPgdHu+oaFRodEQiI5ENlsqEk6okTTGDr9VIAD+W0aVTKtx8oeuK
k8LvYhCoDhPuwp0Uh6CDc7pBN1n4F0nIC3LN5j+nGWV4YoLOIMllGfba0Sazny/S
YAQ4H2VdO0bcGXVoOiqF5siATuFjaUonHQR4J7QTa+SAWaXN3pxzs5V91Vy8WY3t
aid7LPKpwx7Db3/MM0/xeSA0YgHKEpe6fCJe62h6Gzo/vdD0Bp3YPjJoH+xIDX6u
//epCcDy6ytWQIvrruT3VqHXHUW/KFJnJ2ndvKs5vIjLRrTYx5BvOVD8Vhq30bgP
BK5z4ZXzC3qvb81vVSu06lExmJbVpcN1vy+HxGw6SsWhB5LGfHouWzwxUJYsUuu8
nm1CAS+rqHP8PcKvFUaOiaaNcsmiLEgX5+nLXZzAE6UvlR/tjzOaxvzNMLwUifat
Sw2UhbIeOcGrwCVLQBWjQzt5rcaiEScz99Y686A3N+IcNfBJ65zITm2pQb0l1GgN
aKQCr6xrco91bDCfsc6YeFdYSonqNVKePWtN9SgLtjh0UkPOWAIpXKWAlMZI0r/B
v5eLsjUrM/pUW8ZX7wwswe+fN2Fxh/rd/Ntl7pGECIzoCw1z2GVNdPi3PTC2dsse
E097SAaDsRxqQmFrkydkCglWAGy+sOM8roec/KbOmYu4cwAxzcttj1cssRVErnkx
NztSMHkjGp93rBHoRGjgQpCWAgDmj/hnMp5gpqBJ8GJSsaK81v0A7NyTztug7Ude
03MoXV9yJR9C4FC/qdyvuWKX+5e1DzsxJBYghje6wbbE8OHYg0pPZWcpwe2lgf73
YWFssMurZ20e+Xo5OuN/+vfgO3gRCnPh4vp5Crc0ZRkiPyZxNwtPNoJ18FI/slQR
qEeP5w8C5R393F7ExfkO0X3C1dH4CigqRJiyVtSCY8Z4GdAnb6dkwlY3JBT7l1+f
vgvDE8EQwz6UzG5MXnK87zlBQq+FPvIb2N0Fdo30U+pPeM4kvOF9LTx8dz1xarJc
/kEAYggCwSiPft5DFIKxBXEPVJ1CUsf0LaCOaYW759Km5VvgcGwTgKl/nCHv2JG4
zDMCnndqtFTC0zGYhYZHoVNC/+Xc/pU5MPOZpUSFiZZy8PIn1cdSMzxdmpxFA5vu
HQY62oi/L2tW9E/lcwF/m4lUyVqCwEEkorl9YBed+pKC2CYSPfDzBFwhQWA+NJJs
9O4D5jbKEfFVGxqaWYDBkxCHUvCboFNct+sN/mp1Pau1iyHICoC7bYSg6N5u1asG
p4XI258it4jlXDeSyZo5ET62Ab4vh+Pi7VV4ZHsVjnrNgolPvC85p06JoXzh0RSK
U0KvB6MRQ7qHuryHKwBZLHaa1aVAbrJgecUL0ynrVxYCxQX1MRH7FebxMzjj6u8u
JgmMr9IAVMdjTDGnmJ1WRxrpitjN2uxx762xY7rshag1QIjAa13kTJU4kBYTa+zC
rVC3PB84CnpidiMM5RiqknudLXlS6TWA7rE0z56H2gPeF67b6ZvWFCmnsot5pqH2
RmWxKWGYKKunZ0ZpBp5Qxo14uBpJ++d0IaJdPIV7Yh1OMqiZ1FBCMvGbXISOsidK
e8FhwscdXAfTf4cEAFo+Duf9uVb3H2wqBc1rgbnR36iMCrvpWdHfxEJZOMJNCzZx
XOCxAXj8DbkbfQ6nlMbzAyebiPnYcHiMtmCu9u9kqdngV/4QRvWVmJpBn7sOQS2T
STRSElBS6Xe1UO7mneDZ6gGutZ28z2ZnIr1r2ZvFVPVSi6Oug7hM8ywiyANxFtsL
17zx98FsINX+ec0/XDYMz6mhD02wGRCBShDsvCbv/Jxjvlx/V3UMfCx6Qy7L4FW0
1uo0g3PC9A9SfvztedD8GdJ0EavD1VbMQadwNRchHfOlJE6xtcolB/0rnQvOakus
D1vtXeAdlnRVzV0ZjCM6I0IcCGlimVc/qtLgUptFKyGiosgk9pMhXlu+OXLdhqHf
xxKqF7nLRPfWcwyONo0TjKcgTUuTzizsdjrFtR+X0hOy8tg4xCGemY/alVdLdQ2r
gBh0tQ8VBSX25E9iz9OVaFgVtTGB2oj3Xs2GcGxCKd+Lw08dHJ6U8s0pqePKzO7p
Y5xyUD3RX+5Z18++05BDJIcCTCv2ePUyUjXVNJokSm7Y3Rxb+3qDwrTEnkxf+XxM
qIvz4/0Nu7F6rJhz0U7LS3D0l6E6L2FmQS9cYGduunYMgUj+aL2RKzaz37fNQABo
pUAiYKI/r3wSF3JKdeeTBKYX+z+fWmLkHnqjhjcyhiwT72yMjIQFLUEAiKyTxvmG
Olnh6+FPlbsBWLLOThzJlB5nUweEbcoJbYDT6mJtZbnBpc8GEtLrf7bJp/7hdAU3
xcF2rqZGQDnfPoOPuMOn+iHzYXa+d5dvp0uxP6qv27tNoXcdqddm0zPn4d5X/2I0
d3qal/wUikRODQjPK0P+3OEi2FJ7J/ros5OeNnqWZqie+XqzNi9NtUiPUyMb500s
6uUFLkna3RvdDv3xxz9zCOB8fLpVc7LbEcrlTBeswExuaw6nqX23LyYVoh4f9Nys
f5yMqD4FEBHjodvd3n40kLS0ptMaY6sM14c69um3uJGV+b8XKqdHh4CEqc5SV8Nm
eK/lHLpuKJGGwiC/aj8axTsupXW38yGaVFBTeE64ol/fvqTjwSzmpz0xNAQ3tv4w
ovMsXKqP3u7SMRlEpk+fyW3EbZg937CTZEQ2f79IeZaFJKIMJPTaSvaWxzijLZ87
hQ5ZTnJtGKTNZEFVHRMYMil2vJn0OZvB2uHr0Osw9spja8D3QSmWQUqs5J8QYQ/y
h4qBz3hN/8A8ufxZMYnWZ8pYfhLt0+VZva9wtFs3YRiM4tftbSusZddNX+N65vqt
8pSZI2eExG9xLlhGrAyxDkYPAuSUvwzgtiFr5xn9M/E4sLCAKsrsbL+qk9RTxeLJ
lvJuw5q+BkMb0yRN9kq0GFCRcM12c87RD8I0cFwk6Th6wL4uI0q/q3LoYEln1A/w
e5HYoi2WUR4s9pFSnAGRMHucO4VRvbnyR/onQcrik8+gCc3+O6yGSk9mY8MitImJ
IlUsxXPxJetbbLNeTe9Mvss07PuhbcSCz9BOpUDjUQFdIasNb+zR/GMOqLIf+mam
EPzwIayy51sAHDvRqlVfI5ZMnUYIY2G4ymXZrkdyNfF06a7oxy27O+8+doBB61Pz
duMzoySpf2Dyy+4CbwXWp2s06eu4gcN/A17Kf8cguWeQz1+2/TISUPH8dmwA19lv
UQg2DWQzGCmNRuTa5Pxqsi0RCLdpe5V+znm6ai4Uwr5sG/iy3NoE+uYBEghInxK2
3B4RSm4YNNcXxJjq1FYcHwz+agc6Pd2itwyTFJHcLtOW/uVqc9fNnPC9Xm/qtFyj
wXbR/33ERTON8Iyahuyi9IT+enasHfpq+qSVQIli2MyMHtwC5LntCmKjxjvKaKuK
Se5bW3O8Yo1W2e1KkEW+3uky/ozTfccF7NCBt+rU3vVwxISgoxGG+AtLkMZxeyuN
lfNSN7vHxm2Idhzn7Wyap8IRPaRP3JOX6ApCBvUs8HuAUEIjaAa/BaxesgM4wopI
z0Jlmba9Cql2KL5kv73cm1CzHrpU7yeGmRrfGUkkMH4LjYahIykG5OPC3WvrzG7Y
hVhLHNhWzYAJB2VUO5xEn/bZR2OW+zun/WMx8H6PLsgMY/9M+HA5uyLsoVwvg6xd
UhldMSPP1cfATuOnf4XYbjoUikRwh+dDvUzHRxqrKL6QFscSJiMZmf7syQzfohgk
WtA4d9BdQLNmAR3j2zGUJjDuGVmSFA5tvs7qAH7UZOitQafehDpZBF5ud0gT+USn
pdleJtCobe06KwTRBUbaTTKlfdyMNne7cRD3+tv8hU68eWvOJaHMhFeJ+gKVdDGo
gTyNiKyVHYjeWfA3jYI42/8Q7mla8hA30+bEhIdlzmR7CfqKxqV5SHy0GyC4X2LT
3+ZgjMZ55woSKkoeNkUydR45U9Kgl14ZYYobcvYWs+tJwLef/AYDO+HT+RqTuyQK
KBeOE4Gk1iQ71fFGXLGb8fUBAo6WqXWrheg4WHnAB1SrIb+TOxtGbrnHN6cdzuBb
3Xlrt/1TIWesMaA0hLPr29S4iqLPtiFZ3dlvyxZXIWw5l5d6wqu1TsfsLA/qea6E
NLTMKR7dcDhz9mCjwd6efK2vC6h9doAUkSaZ1Z+OtmxbuoWNg9j/x4Rzxczla9hn
aEApMuIAyTEgYewLAXZLEX/7BdbdilegA2OiBOoPpb2W3wf2CkXnzrUG9v3BC6kL
OW7kXq5PdnfkbCZbc/vT6CNjI4gD/3uiRPQJ0NBpbA8pEhglKpU/inrhWYeK7a3k
JRLGdNM9lKENileqfdf5rtPh+j0NXVBgqbLtzGZ2n7iJiKGPIpPGh0RxpVWdnBVk
jXhe4rocA0D3l6MRT4t6LJxvdQoZv/4Yux8XZRWGSg06B91oRcFeKdyCUOXRQ7uF
bMcooj8nwTc6j6w7nSvu41ZJuoJTnIBEZK6+qTb+uPWNo3b3IFw4xZj2NOkJs6YH
MvX+tW8jVLb7Qs1D4BRDOHjIe4fvBfDXPknSRsvnGLmm4r9EXW0enseH7dGzqlM3
1F7Bh2BfuRCGPvpUrgr+3aO5Sc/LcY6OFXNYBP8AzfZdqY1NMLiPBLrdk0PMqgQY
1LxpgD9Ry7M0FH/9rAIDPO+kVzx/iBtkWJ8lpKTVQWsGEnNpHEGaPsfW5lW73MoI
JWILLYlAvjnApWsRJUwm+4PivENdl4rfxXttGP+n7/+1n860U1US4tGC6wG9XL6E
DiUb9gO7imzWEHmIH1Ejj0e1SWocIIejBFynuvKYKiPKEwGPi3rulElYmtxzBdII
Uln5IWXUn5tcCRhCcwRoTctaWUtcjWxc1FE8s8rsLe2oNITti0SYUeIWbm/N6eNU
xNOQCDcAhAeCdEHqP4iSdh0QeEUf5qyBz0TtnEBIcwIR1ZfkQHATADo+9JsnrE2j
y1bE1cVjGbhEtuckHW+Gvt90q7409XBI/lS3d8K5wC/QrxIN6B3bpxVtHEJPGpwh
Z6+6QtOGuu/nrOxPfyXB6m/rQYLURi/NoYCbSVjACXNQ85gKuGAQkl7EvkEh73/Z
fFHyc5nsZzscmDrPHwCXuKZkpWLdoD+tDotGCHQ2IWyEo9qzgXeiJcjZ8QMF2aOH
5f0Uv/dzisSaLIf0SW+yGH3CpfOZTUs80z7BGY7WUjhRh6bii87Xk1DxN2HtkNbA
CYuIUNTidK+gqIyTMDerKwh9eCn5vIwVOe3Hxz+3JXUpjq3/t1sC5gY0+zJX/1vK
LjVtWv0EUCKRauvh3DzbHAcS1pWAcF5SGME+Q0SQHc2dfsUbqvoqacuXkmE8bzwP
6CGlppAo4HYZU+7ijjRt3cDGvy8rUwbKVdsalv43Z/aoytGsfQTYx+rJoNx1D9dr
ek53BJvoaw3h6mH466Syb7HaT2k77ScRnR6rn8h8twNODIcooRtofxiSCfEYNU0W
1+RdKzqhSWBdffxyJpGTa+ODVlUn3PuC8IRdq+wLYFSKWD6CUIeFcitg27QO+b8o
z/tJq1zPm4xBKtDBfr+PWPKlPdv+3z6DjoXNPjsKjq5OQFobhBo5Mz56sawxS5wQ
oCjFAxpsxNH3RJaU77mfy+r8o3bC3dKQNKgmeoQbpg49ssK2D3rEqYGrPfPMLLWS
krssfsLzzJJvizHbu0YVskpudcxbsv5o91/wcYbSgB2PfYrZy4pg+aqQm4C2Pa/C
rhD6aEt902yPzMkEKICHThfT6zY8ciis9sJQ7hIQ0A3f52gAdQi+gSmhq8duXTK8
glXvfYz4Ukam8PzOWjzPA1m+C+B48YnpGDFOvU2jliY6nWIV1XdbNmD1TCEBvc2K
8NhPoO31mjWgahu4SbV4kbcswICxAh6mtMUybLMgTHIiwTwll+5qzuz3LlBxQeV7
zQ8Cxh9mrxa0RCQay3K2GP4k1XCoKZ4LEDXjHGhRuDedvY9jIxZoLNP+ZZUq2fMh
UvB7uMaWtpIpSwcxW94bw/cIzlqxLdLjflCpL7D3UcRnR2yjuP0vFb0OAdYF1Vvf
mYMCppkhFGM+7FNGEsgF6/sxjZc8AQ7BD/VulJ1XJyXnPGo2i/Msh2ITfBTgC1+m
W8AXdUO+asAG4y4oPZg3QngRluj2LPBDUOc8FZ3RLA65QeJjmiNwiTqde/2nWClV
QT0WdVGWOk4WtvZdOg3LJeJ+zlhie2Y2AvGa7zFjWK2KWRccnfavsvbSrxKTIDKD
4AEZptHsguSg7vZ1fsG2rnpYRAqEE2wBQ5yxw26uvrezbXj5xp4Iusqj42UFt8oF
ZWWnu3ZwrJo3Q9boeilkDeZ/9om7DGOtkeuVOrCyA1r9E9bTVzOHi9tCkPS7NyPW
xVDzkuJwwySgNsRe7Uu02ysoTBihjc+CEzLH/35xVrlHh1zBgE+eMeqG60Txow30
z/pLm22rsmfjbZ9CsWsrznoR54WeCAIDfsFRuZGatJBd1Nze2McLdv7Jvr2oEYwu
7ZCNQwAJAlqqzwM4h0mJMT2hRJ0M5ndCn2+loiTJNjhLFqBNu0q1ZVecd0JXiqzB
fhz7ihqU9jwbF8YEpIat63zejyoyGrnfyFJaQyOjJY2Cu2pugBudNNopuY4HKE0m
ZCE7Mx4biF9HxsXMhIObW7GYjJrQzm9sX4KlmQ1CiQBBYKPccQOxxLw71hVSpuME
/4jFLBWoq3FJTua99IHzUQ707UN/rxywQ5YlEK1iNiHYEZXUA0HMGR7KkP36ODxu
orPayBuh0B5IpOLarR69EA2vB6vTsR72AZTw/5N/hWweJrxs0V/h4FnwrT/gqhAj
bIe5Rns1N5l81Qh0GQ7LzezkrpTMl1qPmdsx+3kUH0JSGruPxx35FH1MoGkxSpKt
6pqa9mtvLGUWej3uJC6GSqpjKWF9w1nIaRLfm+1vqjZoPAII6UnOe12NXHdEAowz
hWAK5GNLZefWBWk9zXhGvFJzVmleSDfclCP9irF2JCaHNqU5p/8HElFTZLaCIKgs
yUCd+zgBAUNmT3t9sOfab21QTc9LToh1VoPdLOZGrgcvQvZa3DFG1WcDmTRWyl/X
NRdgLu3+HIuPXYa2G2+Z2dV0bRoBIZhwjcYrKB6MGJtWXoWWpbGtPe95zjyGZd/f
3xDFr9lusGItui7Dz8UvuBJSpZYp2QvZnAdLf2+cvCeaQdIbBxE9te61FC139NeS
IpzcKioD3Upwk78PyDXuQvv3A3dY4S9StKFN/odW3BrlAqpZ3ozyORjI5/ZkCrWe
+x46eqhc+yvnQXzxIdvrihF9y+NuixEukkmjZ/IbL4/fOr6oUwHIKchU09l6xLW4
hO7Zv93yo2pR5sKDNsETgx2l/KY0Wcv1FdaJJPwCGsSbcW4dTH2+8YHyGzKldaXY
5vz14qUVMnG416209QE1GLRLY2df9VFxkXpUD6Ci0mls1QyevnXRhWCj3yem+Th3
y89CShL8AxFbrRZEufVkQTgz9wcwjBxcH/MxNTDJ2jd4xS+DQyn0fTX1Gjz9fitr
gSj1FOV41It0FwNPaSPCezgzahU/HmmA1GVM94d+WJx4BpPbGOf3EwEsnRjvf0Do
hLhL9xk2XjN+lO5Y7GVsR2ZLHXQ6FAu7rL/PidqyRmhy5egu3mjPqi2KQdWUrTei
Lu1EOJklCnhyKBu2YRjt0/kGNTBDAEJamL8eAjVJBsjVIXtGXIlDrkZ8u/I5s3Wv
hnPTsSyuWlJJ7POGEk7P7U+bVlvP8kBqY0GGkTwwU6WC3c4eoG3CHO06HelZVhus
nVvPKcKpRp0sZjTFbS85yj9Vkd9eOWlhdpO7lr+IyRVgqn404hNayvXGxsal2F4J
Ug6TMWwvsk2xNQDX1cePeP0Rm0BAreXboULSrYjzNDzTqKk/mn35IACLCzCI87ET
fzU9GtE+7bOUMG/hiktCGFI/srylUApYMhv/db69whD1ttHKE9KwSuZwQu3wHfNS
QmQzGaMtG99TD8vUUnUgIN2oQw50NSsb62t8k21vVgtDpZgQ1iiNwXgnpZi2X0Eo
Nt+rnsh1lC5Nt3jRCuKYMaIN47vCHS/Or4VCEqxiyWPIHvO+4OFtR6hbSja+lCM8
aYDtp51BMJiX49DN2Qhg7T0XVoI8m70wgG4i/Tc6wg1/MRxvJPE4VK7+KlMIu+Wb
esJLTbCHZnBVBgrTDtMewBSHfbespgbkIgqnKrTZSOeDTivJanRGbTHNq6HcbWbn
qNzklXfzsQTUC5biokUt9HbJpgtwgHiipNZPsXdfFn8zsLj2d7n+da4aa6bXRwVv
uJVlP2Kt12NJd6CIpebbB+mCpHgvHkh7hL8/WHgG1i7AF+cD1pjoXsANxjDcNnyQ
HnFdNDztq1DHBRKngr1GSASKr/ImjDexK+xsr5xTNCRmlyePMqzRPk4e8FuT03s9
tgtkTt0EO9Ghau3V2S4RX65WhFppRrp+GEWmm/mDS9XAe+9qllsOa8G+cBBm9N6A
IxtIswxXHJzBpk5+b7aUqVOkfgxmr8lm0DMAsf5jo1FjNWDkZPdJnUp+4Blsa3qB
k3D/0IZR9jj3SQl/csql08aSMEtZAugf9QY5HRRmXkOwyH4UO7//NBTh4pUjyBf5
iz7CDCoYLfyN8SU4NQJRlkCR8U5SJjLkEPnBFKxVyr896WMjENisF02I1glwoESB
JvyTYFg7/CpKE4+SxXaTV7eG0lL7HUiQCyDUaj4kHYBSrcFZyrRxjH6PPMqYv0xS
e3ZSJY1BiVE3jtMuK+cPEonr5HEg1+GYQDoM+YMaxQd34cYAHY/UfcJUMXUKPO95
YDt34cUE4RQ6sFKIxr+o0O3kvU/mp5vlYX2jY1hmvK8yZ6+BSFIy/CB0xIqn31Vp
bKLfN9x765dC3X9hZc418TErCTnf8vZmQ+HYZlPGQHRL/fxkLla2K33qDQ6Ltvy0
AEcsEWHUwUGz2wR0M7rNr6fel7WTzukhkcylhsiFMAEHEUltn/vorXZy9lcFMuxY
dDZ/nzmV7dRb4FA0EXjBNv/S86LarYQFtbh9mQlEweLP9pfFgIOFG+5CFPtGEZUK
C4zKg84vMm5y/WuahBVEz6D5BZ7KU8IgxnGjrdQ76aXw+2RYOQnT02fPOevO8w9B
KgyA7ApjSANsuoJIvArht2PBpCEzGmicwPUyw6pXM0i+kSZNMt9ZX0J76a9wi8ri
PK1+rOCebn6HV+o5THmYGe5R7GtsTFhaVlJupewxbyjWVHGzoMNT0wL696ZAQaeP
7917dL3LFGJUnsMS7RVChrfiCIbrJ8MHnieHAkP9zlVUbCPpBTWCp1m/pRJnuR0a
wnJ7XEebi9kbmy75hkiZ73PYNn6I4KqODUP8dfmb/WGVBmRMhLGPlnugBNFf/oH5
Ko2l8MTnKibj0Uu1RTqaFx+cKYfQT422TIHl3dSSsvvDCHzUaeRwnwHb5yLROlTe
msmFFDK+ofHZF3BGqcWdsPdsip287EDOyy7EmiqRfvsGiqwWTOgcC0RoLQXr2cL9
99efnfvXfS7KLlT1vUzAfjz7+rRl5FRRDC1ourD7zMFZC6Ry0nM0npBFeohFNoKm
CtrmlaKlyGQKkEjNnEq+dqDMeVU7j519hgcF80wJim3bM4JGsPGEbSy++bXqRQ6x
pTYh+cX/CtSqFUJnYWyu+hZ/Y9qdwu7BlBeS0JYiFXGmxs0eBbGnTSdNkzOKFUmv
ymPuYMZzAKLaMMIrSQxfrUeV6UIlpH869KbX0aPlTtq07XUGtZ/jE3i22XQHfMLU
tp30LpNTHqCsHlfK6ctgIRW0eo1DIw+krO5We3ilUYjZ0wCFUJwEPUud3EH0bopW
Yy6oNfOcmpISYfk89sE6CRztzgYfNoTjTxQgZ5RcBDsARkN+8mOr/uGv70eO8NxA
n3splpRUwfzp/xYgpfLOEfi9vtsF8gpQUWN8Fyqculqc5f4jIp6rEM/G0OOU70us
Nn9eQ9YV0SNaVQU+ADBmKvsy2zUIUM6+oFx+95jDqvOWXtI1Pi8GZiqZAsdt79k7
dEsee6jU5oDHju36pm+FH+4Sj7Q4qtPEKPQECtrtXstMQ+/TpMNVB4mKVXV5MkEc
aow0AP8Z0MN7HumeRmXdNGrnWWl6GECX3g8hlWSLPQ1nm23GBmnWv/CCC7pdZaG9
ocWBXaNPpreymIWX60bV2/GkqiYQTMS1neZSYSCr7EX+WNHPNMVhSBRNVDIjxaBu
nR3nuUNEYhE/W4yoWg1jAvtlteSXjknbupjgJxtJExGwcAfstvvDcwi7TsCOI3Kh
wGZeDWC38OZMrn8sOfWtMqp2agtLWdhJJtpay3FZuMNTYSWy23m4/RMrVx/ACRW4
lXfCvajk9N8B8sCrKXL1QL+68WclBQbfFgvKPZsZT23oolLbLxdaI/FIEk0gZchZ
1yBkMjbw8s+Tely/jFRIMkKuSqOxlDPbxnCJszd6VsJF2Wad5cyggvynXSlyo04x
J0G8OzHuIA7j5mZp87N81ufF3yMBtQPwpwT9+JQXmK735ljYvpsY6QwkZpZ5pzs3
eWN+vu63nTNrXXPr0rSjN4y26vF51TkHxgSwNHb0RjcEzTY2nxcUsRUTTy6+2rIf
gCXwgG6NjPIg2qXMY51F1JlXJr5221lGjbNMNfIHRihV3Chpof/Yvkiu9JujITdE
kQSg2Yw98K1S2YOOmYS6hFhKuvWfCdDzwBQ/htp/lwX9S/bEjIVf5xfQH7uRtyNF
a2WDVpJLQA6eaZobaQLz73QzrROoCesfg7kHH4zcHx6xxWtjFzbVSYpXysD14MSt
uRxbdsy0PUcSer1GWVClMb6fCuZsmFwDR14zaid/hhlRTlEXg1Ew3vE0m1UdMIlv
ZryEFvwdNwIp7e1hxYo6ijtkC3KybOqzn2IXlTeF+dFPlmgZacMG4BK/iZbSa1lV
Weio/8hALpQNgCpegeVmfKjNku7Bbjj7e7/9rj4ByHmqMyniO+7y7w8ts8yQMoHN
nEEVvPMbXofvQP+HyxZ5hLpAGLRgyRy3Zx/pvDMKTHfkOoRuM2P8drptk5nLrPyv
ximY4ClMd1+FWIAGZjW2AKL2l5Hmd5OwgJ9cTdBbyn1zMCutAvpOXcsQOe3OqAqD
61xS1mEX15mOTO57j4BobO7d0euTumkoSUFouJAcM0tBE6M/+s0YOjzFjCJZaNlO
75RrxzAZBuoYyifoGVFvZnzAF9ABD+iH35dj8YYBbPEPjXatjhzOaSOTwtwyTiix
qUML7pONnEzjDO7O6NCynA//+sgof2vMAnPgprgo/f454CVmABO0aybPVxtnx3iD
EvxzRFTHhdfgK5aYwXM0P4uGARrzzxoNk2gHQDa714aMAKpNRYywhkh+mq5Puwfj
v4Wi881LAZb5Cr36q+FJRgOQxTQxm09vfHX0OhU0wTsDasOcMeZNrW/50O2k0UgJ
K8Pl4ug2A+MMxRbOlQKOD+KRoC01hYN092VEKvp246NUOSIxLBzJWg62rlkamPhU
36DGfG0hyt+WyxpBix0T6Vwyv4Y0xJ5CuWRH89DetwTPXYo+J6jzIGFTkB1vv/GI
dCZ1+SKeTgs/38KfAFzbz0j9UI4xZPsRZda6ivXEJo72UD4pZkp8U5yXjjsXUPyG
0bl6bkRFrqpGOfJxyKfqwpJpChEze+7iws2TS5bHiZz/njINkppzYAtqypeuG0nQ
WAc2NcO7+LyixLdj1mUg4uTUI9P6doMFt5iP5piT04tQaHS5Z1ZF7sZi6fm4lM2r
ulh0TLuy2GaLOv8vHNI9ggXO8tQEWut8u2DeVknpP7Mz74NkzPMliWAsMrYLFf4F
kxNrH58mwppwplr3PzN/d6HRIWB0+xaj+l8r9E4hw4eiPzNUGH6mSqYY6al7+ixl
crzc2I4oPBO+lrANYE2pmKP9R0OaoHxMmidO6uXAFCEjxek5BLN5s7OQE26lr/k8
W5TRLrgOxnmCTNYzvzSPICBcler0QSL0h3U1AbO1MdL8i5OO1UAHr52wIjp9AVNN
gYv3STTQh8exhLkb45jsv2Zj2Xg2+81tqPRONgslxlQkKw2xjotoVr3QCC076xEN
jd1slS9T/9PsJqRRCx8nP3psO4DmBmFlXsS1tdkhPG6zr2WowGdEApp1U5sxx2bT
OqXS4sp6TN33mej1Vb15E8fQKRQe7/sYLXB/89fJ1CpThZME8KND2tou+8T0Fq7Q
qI3Tq14BL1Sxh8Qnzx30qnEFqboskuGYn12qejuGPVwM/NrVomuQ9KGaCSYF5Po3
+9ReaPOmGepyfFdqYEtalR8V4XGtwDJ4nLhD/7hNW34A2GHp8mXHO7pWg5xsamd6
y7yUu7sbFg3faN52WpcYeyDyonhJLYjrrEA5azOpIcGlHUezHzEImFpgCa64gcwU
RzEZBiCkAT/1mG0Z12YJDZ2iMDQ4m8yB5wHT2Evwtu+S+F9grdDgJjGN5eYOAvIQ
G+4kyB8e4CGw+9lRWIINv2y7N0lWzX10NF0DlWnQ62XfKXW9Kt6zDcb80igzXj7R
lDNjcmwh1EO8Gq0ZpG6oiV+XWCP3IuvaJh64fpobhZnBT4LyAP7QvQzxVi+Xv1Eu
SHGyUw1xFG2F1yP3Kllb0nh3Jfm786c9dp3HUa7we3exP36aW8SIeXmG97ZJ/ugA
vEzpEoJuWUAq7gFwJ2LMqz1DkQds1Yqat2shmm84Tnj/ky3ShWbiUS/pb3GN1T4p
PtEjxL/Ozh/8yx50lSdYXelPW4kkMXcKPBCipijMmLKuKApIcbymBgU6r07dIaxC
eTfreVS813YtH4Pef7J/IhqR179tL3HLiO1WyyXKjpYJa/Z+G5BBejZKn6HulXAK
m/LXDko3QJupbkKD+sSZY4zgLi5DuW8gRIRN/0dn7iiqfdmNFxBu4ObAjsoyispX
OZZ6hX7q1aZL5om/jlr9cJS5lQqm7DF34tvnhJSOCIawRsDdiapAUV78TGK00hoS
82/qpfzTAMSkaRT/yGc5zZqsqbiwXahOcYICkkaL6URU+wDsm6gSodmpwd+M/4dO
i+dOvfqLN7oRanhckcovG7XMVEh64/UCLhgRXrFQng8esMSDAjvxWP66jdyOW0BV
73EplDrElKGhtA0gChnbJY7oRVTuGoEDgBzXs9ZOw4sdQDIWrjH0p5utvWfWg+zY
xBEIDeGMIxkCM2/XSD5Xx4/q0I1qu9C2NUQdKFTATnzo5WsaFGlrbV+ZTTHL3/hE
1OIxrZGg2qqCB0MQMteEtpq6w16pPurO0EGWSAopJAAAttm62auV0r2gkx647Can
+XoM+iJbI9S5aymghgQGD2Ll9aRbj+NUuDr/kGpvuDGR80Ah51eS6Bd7kjLq5kKH
hvOcUAU4dW9O0rUcrR3Cqhoe+9DTTWtMYca//Y4gwd84B8nek0x1Q6k+9SUW99Ke
KKDMuJP9nyZLHoUPnPV9WGd1rzL7UOXHcPmtQi3E+mrTq0VbYBA/vPFDyCGDiiwt
gW9yt3w3rqQl+1InTc8+EIFrfqbN6sttbmByY9Sup4vfkbvCGcGRRL/5Gp6d2xmb
Nd4c923TfhsC1BfFhS9hZ7ZF2N3DE+7JH/XURdxz88ZnWnG9uWMUm4YjphSouONv
fnhgHPs0mZiktA2ZcDjSVeGkqxpQDIHNskeI1v6nnQSZsk7EnG/UEPahcC6yuwin
2WPG+2gC6ATHyHBlM88sgO9kTA7Bw/AQlhP+qOQaayKlwWKkom1aG9T/1aj5sHt+
9bwBi5DA2f0hOZlZF2ItdFi+WUuj6FFx9L20dTCvR4yCwfOQEmeyXS+Y0NS9Bcwt
X/siIQ/sG1VSJTDrPGZyTzD/JXfInZJdeCFw8TcJaS+BJmuipNwimwvTHv244k4U
Qh/C35M5N3p7C37AfR8gtpQV2Ccb0W4SGl0YEIsBetjGje5lpTkSaNJ73iYfrlIo
JiJ7AntsgX/hTB9D4+j0Oj9kSAd6CTHbeR86k1jfDHZ+nCPQ7kydDsM9F4MpUQvt
LmE/BqU4Gb2tpP39vCNIwNAJ63zJCkq27RepcutqfsgYj1d/MDvGcMDzqP2kp7qy
KJFbem/HGcck2jLmCs2po1IVGKAqikyvruWJ3waiGRpaUaefucYjcTN3XkR3zYvc
lCU/uQ1up2Gh3kfEXygpoNqpLwRG0me+nsBJ+U2dQm9mYFxU1BK+DcMe5FlNAu4Z
4sAI8jlpONohzQDjeMRhTNt6Khhgf+PxkhjUbNKwW7aMp84A8svcc2ry2GN0q8jC
tfRFr/6Twu2whYpqw7apEZL9yUG0mBWtumwviT359sl2TtpGHu1e6w/83/qtuzQB
xAW1sXHS2xlNAZX0xPkhCc7AG9717a6TFi7EBcXNV+tgru03GTL7x4KUo8Rb7k51
umiiddjusrINScPd3tRfmML/eiXp+f+w6rwo7/mNm7u55TinhAWAeD45PuzR+foy
p3X0+/CHdkAoMAoV7I9FZ87NWXEPztVItMBDXUYUIUgLH34mxCWnS6s6bKVNl8h3
hr+R1uHzJUL+NrhBNrcSBm70BjblOOYm9uaMCBIYUiEBW3KSZw/nuy4Mn5bOrVsC
vUkZhmrQ9yU/3NFDuqu54NyuxSeo6LB18HD6OVduHJGZyvOefEEngObixcsEMdmZ
jAptQKcMCTgF9xq59IlE6RgHMBMdsAc4r7SwivQW+c440D2k1bi3zdyWPKE79rJ9
2mv39aKxZWyPho0dIVM81TIeyMmjrTYlqfnePdW5m+YwVeZHpSHzEsAJGcwqOYnd
vsF0R3JMH2wuRpV/nlPODK30HncGVMZqFSYEDmNSrauioa2mgPFDXW0xvLE7IF7c
Yso99zjASkA/h3YQ0H/wwk+JJFvLSGN/UxN48g/5tYna5YhY/Lz6HqQTe5nmQsEb
IJ/p6mnwoTFpBt0fUlVyOnF6475i5kgo1G1fKk8yE2dE+uQD/IRMtmYxq0/WBIG9
sd+rBuxrBi0UGCZGjzz29hhrzvIGDhUUZI/vIdT/pevIndJiCPzNxSaAfEUd5lC0
gb/D2SpXeZcN+LpyJzqJNjb5SdLRaSWYg1DsvVKmfYsrD55/SLm95nFuMZsFaPu1
9z6Ynf2XxJpYLecrzPjbipSNXM9MjSzI9dObjcWiyXdVKVRfvXonl95zOEUsbnY7
KDSeSusb5pw1FOj7cbAAvcRwGXAdMd0ChCs0+cpgMoCJ/+LShfhKXqToNHdbY77/
p58QhqCHT9pZiEoISoB7FCAto5x2qOAGDWkUCSUKazQR0lgcVtxuBNBwg2SLLL0R
Fp1LOpy5+WeRmppSzKpDXprlCxb8LONZcRrwAuCJX7DjKxMhN43ccfP61qD1YfOG
7qjc8K0UfhTgX6duAd8BytIjRxhyjA/1ZiaAEeBmRqJcyl+q1arGYXxmRr06VGQc
0gVEyJayNUivawcWDlUpmHdQHFQAoZwSAYkXtpq5OxbFfrzinjwWTCFENTjQu5B5
0sasBvI5DKm/SnKDQup4waWPWVjfPIsQLsWiCtO7m8U3nR18vCleFYqJmhjYUJCb
U7js3w9nh3/BC5f0QvZy3OqoV0JvVWlpJV3wRMSqj+JwBOPVB9pjciu5mdV46osX
QwdHPWD0JQgmGeiKnShKudQxcVPOU6yYaA9ITGEAdfLY8L72SVKE1ri4QwYqR8Kk
EDyfvXJqh8hmMtgQw8nhjGd/U2HpCywQr2aQ9Iu0G6HhXXV1KmKMbChN4cbfK8kZ
mk91LPu7qMINv7lX6by/muLG0mUjWN5BDld6lL+BaRrUoAx7TqZ0rokWsfRFaGWM
h4P6RkkRjkrXmDOhNTG9yClIpIpnR4VsLrbjAv7PA8NUzokOyRScNJLJydFRK3z8
0UOZxYB6e/hpiZgYrO3+Aeal5bu64qdD1poYqpfwY/ulU9VW3LsYBia50/zFEWnC
3Tddq7d7LYjydBHXb2leUCtX/FPCyBIlNsXBbaf0Ns8lFZC2xWXnN8da+aHnxL80
Xnw/feFkmC2ezIGUYMjK3eWLGkz5IFNMinssuZEkIdsPEmpuU8FcgLCOfFrWDFp0
I0zBvbWhTIyNF40gNotrAaZl93+PPg5a7WTvCNswxHjVkoV4aos+2ydK7Vmu6fuh
bvBnJ/euHdZxbDEjfGmiPVEgcR/7WsYSf2oR5lz+2zMfJLhUZRtqjrMG+Z7lWj/W
J0y7xZcFUD/vjKb6dxhNxdfSPzHvXa9+h3hQJn9FeZRwKrxCYqed3DjXD7zXhxnM
gBN6rLI2fArQf2AxORj7NmmLchj964WbzA/McT/nkR8MJ85+cI5wXUQg8Iy/c4vL
YgFxyGC/hC5UsTGk5YUfmuDP4ouKuU+hxwABRzappeJwJDS++pt67PObvaKDfpaA
DHJ3Suif8Nt3riCQfjopSADaqefn8p4/pMAfOcixqradgLcGZ8HRJ9OHGn44KwcO
1xiXgExPzln0pY5W8evRYkNz54ND+sw8eAGo/qXjB9NFOZzPz7kcSnnI4DB5th25
AwYnMTkzMyU3TFokTMpIBrv0V03u+jrIglwkdAxbzgEinI1VF49AjhyGECopDX1O
iXtWWsSu8aDcY5zE7BSj4EX+ITs/ezTxDgeu0/O2cyOu3ggn4B3rJmNT8o8otsXD
1ebBl+hVAySquizlTFDCrutq3RxYN5TFCWJBLRjNym5hMR5x+I/8qz8qTUw8/Yo/
O271j1SfJ8A5a52CfHyezH0z/Tq2Vco67nsQZk2VsHbwdOp9gHxy2cLXbeQ+A8iV
FGA0LlT6/fSIR2Xz62djkWdRoMfIDc21zUdcGgrYE8CCKwpE8gS0ZincxAxLjr5k
k62Rx2UCbPNVpwbk1c1HlWf3JDSNOhZ8Ir56u1joCExAJBNL8QpW2HQv6XwGQohs
rUbHqJaQDW2FKSNKb57jV3ZsmALQWUVc6PZUdbSUz9TMTQSLYXs5Sfm5BK9f+ugH
P6tzX8gXPFm9JwMTywlYXdHQnn7zavcVxaIzkm0uaY9IDFwHad3zYg4bDPUZO9kF
ktCF679HgB+nUWEybIu+oA2oiEl3Jpgt1bQpmcAi1cri5M+gTSkjDn2jxscTDAZg
TsCGawE+GfeZHafrGR0fH15Ge0isZMiIg3Og/zEntpBQ9I/A4zBkZhy4vV4rrVK7
Y7A1WEF5VZ1kk2j1nd980FIYoHTnCB4HgO+HIR3efjh3Zb3OBvGiS3W20tk23iAD
pwn+7zHqdujvqZnwjsNRS7ZDXGGCwVgPztApiWz1YdJKVSH5sKomYZTOIXDpW+tO
yLhY2zg6w8idi2gTa5k+Mv+OQU2q+l7Nv6vERIGYmQg1BH5IG86OfVYFPWaEnYe5
b6ErUFMeussXeo6uurmozidug1+BF9e8C0+s932KnyVIwiWXptg6+RSl1HSuHoQV
5SgXCG1eO2kYwAUqFvMiWd9htCGybv/s9f6INoVHMDoZHDuXABcmqwxIAZ+1xH6R
tq51eAurB8NckCr/c+eC6aEa21wFsVqbXeU6hGRllVazUjVVBMxIa0QBBFEnzG3R
Efy2MMuBc+tXMBPbNE8jdgvUdLwy1fGPSHjqTKtHq3TtuLv5SPr3EZqvD0Qm8sFG
T/hK9gEjCwvGuCL/S0lsTGc1LiuP5pnoHr3S5jYyehCYLDcDgToiWxgZT8GBOdYz
dUysWhttb4wyvyS5FnkE98MAZl15eHVckDh1nGxpfdFWTiWWeGEB9eNnEaiZt/fe
5CA+AEwTXPrDnGWPr8NNBAOSy2HMMwJn+QjNbtec69/SYiRFn0KN0/n38FLWxXzn
iyleXTumKY2DSf9KkKiSo7JEKEdsmGAEPOBX0UDcnUGEkV+1I02tkzuzpXoc7QoZ
yM1gFWcCCqTqWYcIeorf7Z6huRPPmXQ/BG+JEw3r4UbBIJgBHvXBA//yDbL9Ju17
Dj/9v7dtxtBebbk8OpEiwFUlxsXqxe9Ekzxuo6h1/grMsiC5BFrUvrjq6O+AnJk7
Wz4y7lGQeEJ7ZhPp9xDHZOnawlxctKB1zvDyEnW1WTmLQnGPUYzPXVyaaKZNo1m2
oAq+umhaZJEUNGHBNjcTU42w/SFl3+9djEzl7AZcd4BkymveVKcAQ71DXNGv7ENn
OvbFQFYtaNz3Y197A5skaF+yJrwJ2nRd2V2etDndkBjrsi6mSMoDfGJUrs/GhUcl
2GsI1oR+SY2z8trgmF28AUlLKi/B/6KydQEPSb5ejGfvglYhrCkNYoXM3kyTfLxA
Wcptrcw0nY17fHX4CifL8N9DKjsHbk7736BseV1J2rGBDLp+XNSbbSEcx+Ojj0Ja
pJzkqM86TVrpOq/XcQU4Pdg+vWVEIrtPGog8niOP2Kuso8xttOTXDobOQn/BTPnP
bqoqq34LujdExM6QLQclE/jrEKil7vElzMPRoLVFJp0iTB3lVju9Vczfa8DHGTQt
d36Mxol/uHLF6ColE6y1PqDi7coZl9Q7+621ny5lmbznDKMUtgTv0u0xwl3jBAtZ
++6JU5EE/rugM30SOwyTaKK/FJleBFNtUYT9gXPRsdYjGUYq8iLgdGJ0TSy/nzOV
stAOlg8Q61U35XbCl4dfaaFKIF1okYk4D8Qn4Gr0wYjcnYTtwjxrSp1RhPcMZTZe
nxr36+OwtTbnGqia5XRq0yjw/RgBH3B5P8LrqBrenPXWgo7NXN5Iu4Ctjryr+jUq
bpoQbO09qUKvbBeTz3JdqFcT/3XmVE9im++pQlO29YoFZi0BbX5+6ApHDb/4C40F
7lIGwlKdq1gffqNisQbbGLDaoxEskRPp+buDUtGQXbHEjZ0palvcZYSuUjqD243m
+xFcERXDgwi4KVD3q/cQmjPVX5CLiYei4mKByS3fChjb/X4AX/S7z/0rLZP5tus2
MKJxJx2C9n79veLEkZ9/XcS+e6pf2r8Ne7vJYB0+knU+0743Nv0ktDssr66Jl3+E
GrlNe939o8rp8jZICe+EC3hAnOy3784TJ8Tvm7dAUzxDLZ50VNJjeLssCLfdz9dN
jJbD6jCRxk7y1oHiGvFzvRRn00t+PWl5gVCMm36Ver6KAdRjlfslNK8FtWH+MJ6h
Gf/6P+mEyN1AxsPDoHkfhn05uxt0077kcTQCV92ZS+3uFBv0CpD1QmB7Vp2nRpB5
Lk/LHgGmZYpHkKkHVLNmlQzqTDymbrGDoz7GM+OpmKGP8gss9HYOTncdAT0rlShT
QpB8uQbwMEPDWYtw2EI21OStFtFgOkIR9YT3sn/PDGFTkDzt/PhAj1bE2X1bf4aN
sCaIrCtQgq/iILz33Q2czPt77NfhemB2SvqgezIltLOKVQ1RiczhOUlL+h0vZEIW
XLHZzpISgzG7VKsfNWueZ1osYY3MGsynCtXbqL+5K4oQk8Aic8aVdiBEHBX/vp22
b3cZekSNC44hT1YhwtnKjqYvh1+Nq/o1VcLq1g60yXmkg6KNfeq4u3troW9Fdf9d
WxzsPH3ODRH0192zfGK0YeCwXRI5bNbaH9+E2T+VvFs5JV6b0528DpQhYrj4WG/f
QP3kR0ZmP+S4wiC4usLr8ELHwaNaB4tUIT1/PNBk3F6tvQKZHJ+DAaDfDPHtSghr
zhBgwYpwzpAt5siYr2WRRRSW/Sq27PO6vuUzAd4FSWbPJB3k9O5E4sVIut+FKpJm
yeesOE9ZzX/buP0VNzc7BW1SF5wIKksvkQII6YtLuQ+ktk6WhC4oAAZIIYqdRNpT
e3XYBeCo+sF8ahw9N5nP0xJLkmR98RB79zlrz9zrgbgOOO0rCwWMSFZdoe2Pzt7r
vkuOfdrmYVHTXKBURF7qwY4HseepDA43x+MsGJS20z9r/rkFLNb7YGFI+Xp9gXi7
5lZ2Igs1o1r357IAE4clhPsJm/B/takDobl0AGOHUug8sW9RfQft98qZ9Sdj1G/C
2tWRAWPFbLquM4Ud4x9BIytK0WP1y03NqYg8pL2HiFCfehgRiHkS4NNiRnfT0q1l
9OcBs646Nia3fJLZBqwVdpJ0P0JPk7kIKcDr/W51r0KcXgpr4fFmbUf8G5XWQ3RC
otCLdKGulKtiK9IfoB+gF+ccgSBGgOh0vg2uoN08EoapNTzEh9KR4J5E1hfUZm3g
xtOQ1BN0JYOh7gCkAIJ7mcb2UCr+c/j2Qojt7pf0i7NwrytDwB+SnljUN3taOH+s
JMg3AUwQdltwrPZqm7TtuqvtMc1LLlStEW+TZSDDrOI+x4vfNghur0qaNEA9fwSv
sFF7N4cDN+O6orBQorP8Xu+eWZEW7md8gTFMrcDvJe9lip7klQuTVmrYVBRyTW1/
PsYjeCshellLZB6CF3DvC/E2gJ91nwLmlhCS2kMGNQi+ROeBGUfB6XsqjSllWGag
J89+kJsDKKN6ucgcgH4GVlDrtRHpfQtT7kdKKB1JawANKzSVg/hwpj+1i94Sw541
X0GpS2V17c4qa7T3SKoXGLSd85bf3fkRBCLN4c4PgR0oDxQ5QfSoyURE5jXJBdkP
vTR4hLspS/W8vjgRA5In3+m6BTG7WYBOT9yrqtBy/pwZ1EGDkeAdeNUj/x/BhaC7
7za3LlhkqEaj0SQI93xfF9xhY5ChK64uMnJrzeJqDFhHhWCD4wXK8ddue9PyHulx
Nb6OFeYWGN/U8SgB2LBgAmu3gvHl9UUbBNEhWi/cwSCGaAZYSJC9mYdG/fFfPjBh
1pc12gV+4qv1m0c59v+QdsXwNpBfuMDN2HskUj7TWxu45XJGN4ekYySqRWprpziS
5f8PzO8EeELuuMszC66vrsn7l9BWjrWlSTu7c272ZOrDeaqu/CG5t/d5pPiUo/Aq
iGYEW/W/9zUaUY4PKkeMvivUB7PBL+/+WYjWHttbdJZz5MVL5YnT7xuzLkOXSFp7
BZm/cCxtUrbvvatnfQk7NCHUqGMZEnnDKBVhP5ZI19XCc8SWAwXlTjdqrgzcUKo8
NX8QBV7oJIYq+jJvL5+pv16vwPkoxpcZ3iaMqVT61ydrvMVo2P1MbdEsdU4TFQ5a
/gGKGPAj8WYyWWcmebGiMpacATc/opKWQ8tdki6OodmBpX/bA4r1QIKIVGIFr7+8
ex1VhR4VEzVJ7P6R/VoYEg9Qjrhq0K+ZW0KIGwCLMNdpBgawFwXBmmIU2X10WaJS
OEk0QESz+0WJPrK+/TxKPpNYIBvYJMEVpc+YisjAI6aERfrmf459nAQKoth9h1/o
4O0wRGzmpa4e2yVUCXvY/lOVkPL/NHPX0IXjyLZA3rrmykuaXbXBZXw2h8Z4pALj
AKu2Hz3Eu+j/88xrm/QbQCjfN1zAu+DOU+hwt9HiRIz18xwMwlx4XLgmI+usLLCp
C2/mos9kfA01ibnj9W5Fq7IkuR6484w1v1TFj+SQyWQ2rBLpvQrNLY2Ot4JRFaQY
5UlGTyyF3k7Ar9QLEokE+nw/9Gjqx0lMwi6zCB3S7FN6d+y0Ff5S3TTIdqjxkUo+
RarYv+KhJJowlIZs1ib0P5SXlyQ/Whuyz9AAmC5/R+me/NEdZ0V+rCPsFooXzQ86
vLWYO9GXpy6b7oY7AcCrLHVMSSSR/Dp9hVZlWqBkOjmnVYQQ2dKPNnxEKB4aCwzF
EOn7cpRtaxYevL3MJhgBLXKsoRroXuJTGRtn0yifRP9xiXdGP/QVo7CVnV/ke60t
pI03/NO4CUl8iyFUtdEkTyJo53RhVXqFeTONS7Y9t0tbZ3x4g7P9HrCcYZ1B1pHj
IJrPCnuw46Jbv1V+t0ZCPfnAIuDwEZPzYwUWf7pgyBpFEOjDVYkFsLSp3lOwzIUg
BHkK8Tnozd3dNdKpdVWfYuC8MDiPwgVd9GYVRRxe4Xm8sVzB6pikODsZVoVeG0Yj
fln28EaW162Og6KD+JRB7H4CUvOFVyrsbHvrjuZjaeqd9Xm5Zb6A07eZdnz4SOGw
CrtyADZTs3GZ3Z4OhRewI9BGqhgTgAg0zMp3q8vjPXuLCEUJY+CUglwI9OxBCL9b
lwgMCKMB+4xKKd2kv7B7u4px10/DbB8IKMIuw0itQxqKkRpX2/8jYQ+64dCVRbOR
qnmOYTPzcYfeaMTI+s1wT3YMcaFka++4UvjvLOMhuG0gqw6/fLIJzwW0udvqCX29
bgFtPb9lNJyF7+pIDV3ap/vPXqr0pHLGv3JkcZtSV1yDEtr0gKehNCjWmktVubog
f7BDd3XwoDpqa3OrU3U4dAqG/sRPDHUEw0yNRGFuRfHV/zx+gwW+SrVpS0myk9EB
4KjeeT0gJGiCkRK63sgY8Ae/kaLdVaaPDospgpg0SHd5ojr55PGZBfdfM0jAAG0q
KDhdkn1FXfweGbdzjB5VOYDxvY1EL7gleW9bLayq1OV1kYeZ5DPaHAqQUrMw02XA
oP3lv96YUzEzdmzCkZNcDBvuzkn3CEEDHEKE+YAv9BXvnTjtlrOzx4K+ZyDQFYYk
G3JFKYjYrYOiOtlrnupKNNZrrXE9DkDL5RVpdTuCk+Z+cn4FWqQb6x5DrCZIWbIM
WTmYlUaJIm6+FOYrOzjO1mA7jzPonGrONXlrZYQSHSFTyUQraQP9vT7BBMxpxHQ/
//JkLLM5czdHTjIZot1PmwbONCE1gwXs2VyGPESrieTa3mRwjX8RqFZ/It5iMUP1
W8+ro5P01XGduyh8PSMK4gN18QCXpSklTo8GfeBhxs9uPOtxqNX2VKj3QPR9knfs
gOYccwZdW9k07NWn8GdOn3KBKlE4AXqPM+9dLBEZtUhTurCM2nMbyHhvkdy9AIzd
UOtIDywSMC4etZkPLFyeQK3/pcaSIsUjpiIfwgGU+2gJlsvPMvotcU5X1PedvW3I
Ykfv6q+Mo+elZ5mk6+pUyKe2vleYcviQERpcr8NEih97ZR3/MkqqWD41PsccqDGA
DoDEws5Y+pd4mNB0S53J4ayCNnSKtJ+sgSeSGpNeOOuZgLFSiq75g7E8oGPBfWhp
qYZJGcB9T8bY/Knl/oVH/BJUI1dzvmI2WEMnqORkJFM6BFHy0K7nfVGvEqix0f/O
VATxFf/Qcb6ZY8iEDe3tkH6nSofdq+k15QkywI0+ri9/PuMH34cxQggSu8LrPlOr
rxCS/24HKpxez/ARdCzo0iM9W3SkllpeljiyH3xXmZJ+CYpGY9Z1m2gPqdwl/Gok
f/B7HxeSnWnkScbr6s6t5sXkayLkQllll31jG0T/H8Y+fcmBUNPOjUjx03wJSfe2
fte8Iiv/wPPAEtwyG0VWZX67x7DE3NGk7rcplPp3LqfltmF/CgiPMt7KAqZXefn2
q2yRMUFh/gw244xyhtoqVTe973tCJhBTXbhtxs1Fa0WicpJXtlE6f8FHbv2ziDNx
3Xjbupd9/EfEvQXfNuiUot2UYkdbbydR2qDuqQBcrE2WHVTriENT5JFrI02kiBCt
WhHjNhGJ+FnvFEpLDH8F7fxeOeDDCgsIQivTsBvlV+p5ZLkLBrRn8ti4QxjyaAaX
fbNcSN1e7YE0lA3fnZsQXEUXOqR/uod2qksOefjiYZp1wzuBTDXg6Xu3HRAfKbb4
lgg2wgczYyKD8pUcJP8pB1lJZRyDTFEWtTfJTXPMkWCDeU7KErJK9Gd/bh9TlGAX
knStMra49C9TG8jZYYEKh1gY4fUp2Qri1t8hv+MFViVcbuyjh2c7bBt+WDY7Td9S
pkS3unm88KmFqU7XPDsuCmOxaptihNsmPtwrZPejniz3vcj5zq7hsAVysZ1Bdhrq
ZKkiA/6f7u0UyGwgNCH5NkNgYDZId07Y6E5RMAvH47FeQvgpjBNLm1NHbY57H8ce
OF4KD38GwrmsHU8bEhcIkzg/aSPBDovHHno7BrfsztEM6gLMYvfPIHlLqP5V9lWW
jgIf5OunF9hLqmskDwjIHeCZ/Opn8qWqGbANROCCWgMMY3Bi7ppvSPhmBsiX7qoi
/V4Jh3MgaujYZIV97TBIHMX2WNEegd59VwgOq/PMOhjZDXMVEgQeGPQJdvaOE+kF
5KAFYIpovIRinMiYBlpWToDqCnEzdB7KRXcNNGuhkbGf4NsU+HCrcrPeoDwi68BK
KaKCAlwTdMGew7cT0kIgVx7ZiKxfVa9+jGVW+8MIZPkNvwsMKseKlWUSZ18ycgHq
iy+fPpXqqHHX1QOAB4jvK1zwtIiYGZOf1Xab2nKaLp9QAIjOCiJc8brMFSzO+4KS
qcScGr9GOOn9UYOKJaRs2geqBEVAGele+syqDTNf/CxWk+OrcFD58dVLGhEIQXP0
6yTqJee5v3zUSjpVhgWYs3PfupZqVCoFEwnWQHs+OClv/TtBbuOguqtcN2ycej9Z
J3qfwlAI1q4AEeLMLG+1pjaXkjbT+JP4jmQWt4krGqfVcXeCCt8HEFA+4vjqh51Y
WC43IJB7NWb7iC/0u2zfg5+QG+r08rY7YSyagrm9aOhXXR/5ufA1aRsM0FZ3xoA6
TWRpAU4PayY03sl/fKBrF/YQjQQkhOYi2BQdbtZk6XnLzShVYL1wIp359DDeC4EW
aufHWmTSU6TUkNsCIyWncOoklI6Av4p4if3YxdTDSnri0XrOqFxHzIJ0nWmaqWEt
xznoYPZLlZNyaPrwpCrIovF567py602HKrSQugNxHLKsMRQ1IiHLYQlaTsWvIKpV
e4uAoSyw6uh/ZJtErwHa1QItBC7iELMbQxnpSS8PcyJ/0lFHNh92QDUbMA3EIGIa
g6OFow8pdpdk7J+eNT4Gj/MfuM9AWiJTloDK46tCDiHXDiyjs6Gji05+bTP88qbv
LoY25q/OxaBFJVkZM+REJ9nVU2Rcwm4QhXQTyRH+83NSd8COJ8dHdBPoj+UP1Arg
Mtch6awdpLCK+MfcwMh4xr92capefCupmp7rIzCv4bp1s5W9IN+AOfHIVfNJKBgU
3mj/GpPAHPW6C72koi4ue+ce6EPgRN+7GLaP/ihxX24KIkx5oFp793Mns86C8Gjm
6CLDcbmrUTJx3XqYZJxFf+TuRq18HDlwGwmHJtRlKnAxGn3qo0phElTl405SvACA
1QrXkWFGCz980f/CdgPUt/VoYsjPke9qFBFujO2BqHTbzTxRnUtduY0CGxCk5Upg
6bJb6Nr2/GtPFWGFepZfkYmvLPG+4JlI/fvViC20dzi7O+04rYRiS4vxWYJVGrJR
Y1xMCFr0rLjUpswMTc3BK/TdUjCgafdWmGhEcJ7wiUYpA6TOWpioSjnid3XHuvQ+
eJfuAOOIjGbIWHy5ZvPt0Ftr7FX8HnwSroTY+/uYhfnKC31mlo086SWWaxQNOt7E
fi+aIlD23C3pimCWlE4e3p/eUUV+79PO2Y8p9OhHnwIMFfboK3gaptb31lW7oZQ6
waMlLfhV02gb6/0WRhfM+IzUaoeK7TQpqPRQ9omETE2ho6nMJlZ2boZPwmvF1SEO
yUitVWPvVf2gpszLVyZvbrUUzQoHnRJwKNs2GIi81qhRh0gAaKiiAW+DnkAh2Fcn
/QAFTSq1Akyd9hgWKyIwfThP8dC9pi8kMFWB3omnxROwdA7Qd6HxH8Q//eVa+9e4
gyKgakgoEeXYIJXx3KVA4w/HWoZusgVoS1VTtVSHR1SJbcEIKqGF/G/lDqT2Hhfk
zX3PtgZjMg7Du1e6JYpQMbhz6eDOdhPMzXDBWIRTteBCc5khkKZuAAB4yPI80eYq
HO+lqGvCXxTy5wUJct0db5SskOJPj9wUigwdrYgJgVz4vNHsBuLg0VKOp3yExaLA
qvK7gxLWi2ECCsmMDDpKanZzd11fZ+HY4KYdRjVgZV3XOmEQJkDwFogt7qcgJH0g
cA1C/bvxRK56K6iSsr32VTHSNiAW30qiTF27Ol7KKSjPpoSZ+SD+kEDGp3SgJm1n
P0EM7Yo7S4Vy+SP7AHtBP3uzfNW18jbgIH09JNFfglDJ8DwooAlLk9zS7VKmibvR
B4NgW2L2XLrsNZl1XkiEna1uZ0S1opCkfPPJIOuOR0Y6KUWVFhx+IAsUxx38n1Z5
r9DwUfEsYwo2GbEfjVTMIUtEGm0CI6lSJEgIxPPZh8ehakB4aCurZAduaCcZNMEO
jOe0VmUroVceySEuwBUhTvcnfbBU+Zt4ClJDDOI9n+SmdpC0BiDjwJMIY2CNMuLe
j16kZ7eCYOW5sRyiOFkMjO3f0ql83WN8k/wd9tTTzZgF8y2rxG3kvVjvXNqFrObZ
A+7LEKNoIN8ayZrXe+xUYBd0ZWSPAKKdwWAO7OOEsnftLMQRqxeGRToLYik+rIV0
L+UgJBoDOtd1aXK/rvAITR5Gtuj5wdxgreM9K9FBiSOK+erCHVqLBsgEpCl0K38Y
wbY7/mBddJfgLbXf2guHt2Jvo/8jJX0b8/rpfECryDVIQhJBByaYFqrJP8pzQ0LB
hpyvX/p09MW97tfqIxGhPMOyvwHSlqaLrHm8BKK1gspeMVwkNVR6dSKWMK9HN3wv
FLi9KS4S27Sl6YDlrgdqQz1o/Gqjw3d5k1vn/+4ELiACnZ4PIAFLJXA5jyhKK+yn
lvwqO87eNTupneth9R1Y5G9q/794Z81JDyN0IwTf1h7UntkeOSDmGIszYZEnEgPF
22AezuaIVe/CvSyQvtnt9r2nPbPYQKtB5YFAnEHbfYnYfbAznUUlxiqcYa4Cf7Fh
+kho1jDHmJFlRFls0Aqb3hcnGHKwJy7Nz+XJ1UVfWHVIARxJ4CzfHK2B2maEWmbW
Pi1ULZR2Edl99nCkKOxiIfOfrDB+btqcm8Km+J6Rx0Kdw9SfFI/2ZNl+WqW5F0H2
ZvbPlfUPTzpFR+qAhLCgG1wVjfLGFx+8NgwkWAeu6rqTi0rQ23BDDpXzRiHccaJP
KZjMGpSK1MaWhV48P63eJrPeCr37MktTUuXKF7qJVzy9zSp4ky0S18hAHFdQRUz2
dTW/6KbHowEnD+fg+ObZtQWkIEzeRr26/i4/P3F0ix0KjPRoepjd0QKy+U0eXiDG
1d9AsX3ibF34UD6Zb31EhxVCLnDO6o89sILFgSPVCeG8+mODNuP1dQj+j3OrEOOT
8tADQq0tPLqcI7uo7ge2il74tuziKZ3gRZ8iRjbD46AmZ4HHykdxILIjJ5qnAsoc
W9oKr0h/aqyoT0jKGUBNHgX7/7ZsUCUK8TS201MaDkeqyNCZYxypwQ6FxqDiX1cY
cpwmMV1fdlmpxSr7lhC7elyDTkFEjkx4QlHLkGk58oj+D/0KGZ1PmsL9BllXYfES
w3jFU259rdcCnWDaynKItrAWiB396W7faM3bIVB+1jKBFUJrHmCxTHeQLcYjqoTE
K4aOQrPrHprd2SVHcZ0aF0QeoQGTVSQvx1GeU94ZjeEIyfjgWTg6+/oDzDbhM6rV
LJpAHv7aG/sOyVvblQlHA2ar/QFV2DpKj05yFLN9d36H+pI2OsB/PR0vRFmK9Tpj
G7H2v6vkrxfv4n0+y4nG2jCqgcrSw7JAN/3ch6TTHpqcM39IKH97/9ugdQ7QcbGk
LWLtYBtwMGihtjkH4ATl6oZEK50uf0hJdh8ayXPEID+982WPNUrabWJcdOeglUol
i01EQbJBhSLvjN0lwLQQCXB2xx5vVrIwg9DKEoXnMeI+mYh5ArAAcu55wk2Goes4
haeK8PAJ4U2D2Ves2/ENJcTMQZMOSyWmM0rPz9ChUOvkEPrV8ckWbd7Hr0yJ33eS
bjNkrqR718Ih7S3dS29xxmI7boOHNO7jUW4xBJZAWraRmlg68nTmB0v64Fu8lONO
fz5TYP30ntqDHLSCsL0H5mOHhrgOm9VdCSfx+UGQok0k4hLW3Q3Zb5P3nAN9POln
JlwGd40bi4RWlnIOtCb6FuMz/yH0ntf06NQdmzS+nPhXUXuzrsrZNrEJmHuwEqOx
58lwWlf+fPg7A/mi+ECwnVyIYsXzwFEhCUPFBWhbYhYuQizcvQc4MspjJ9AxSIEf
UZVrJPSMtqt4ZiETl0IFU6FepgCQDPkMEQIg4aGSmT/sh7ULl0efBTES4YH0QIsZ
WlUA2jLnMBAinoL755tc/BPt+gokPy8XrSgeciU0QY/gnRnVaED4ngOqmkpzKOiN
WDwKCZYUHGwQDCBW2FI5K/o2jtk98JxljrIPbZY81necHXv2C4hjgewtzjZIaCu9
/IPnAv7y6PdSJ/UkWJVrZm9cROcCkRyBsMvgrYyCFRfo2U4CdEPuaaePZOSHMRVm
ooHPE2zI1GSmYedzscWLJcXGqtQyMGQZSGVIjCcTgZmMmWGsi9gLOpdYMd1QmQVz
i0MBDU+liQLgWrUHwrsOQty4gaNrxd144uRB2P51h1BcBJucTiosaHILYFg7nK3p
HKwq2z6o1553CBFYZStN31XmbLx3ngUSUOwDJm5rgg7CRcd2lW338cVr2dfaxons
FKagMdIX6eta3kVUvTTarX9M+bwcVpJLg7MYtY8J7FtzX2wjdXv0nGHGATVziAGW
GjbZEfXBKNmznRwcAq6Rc1uCXYk21GZw1zMdiAbxOlbKRu6bpAD9MHb6ma6NEp0i
iU+5jJjk51wO97AEgsEBB6au6lZlP5LgQd1WajjOhvbQipM7XAF+FuzpNLI64rTy
+fMVE0MZAmdKl+Ibol+SyWcv+rShsuhv41zJtaWc49InzhKUECWN7BZ336CONsq+
mmWl3k2ohJ7MwfowpDZl+PrH3q5X+LSDVzjPpW87n5+WAan0gCwPBQ9sRt/baLAq
n8Ymx0WSPW84hYfRFUFxAkQupsfjyYFJJX21vGIx3GOG7x9fDJW3q+pUUdS66afj
4b/FB8AG25cOG11EwQBpom88kSaDrz9zrVhHf8rJEL2YaGo4DTT4wCGKZWib9vTn
G/KLx0RttfFuxx6toIq9LC0P7fK8mFf26J8pc6tKoAbfr3B+JjXHj4KPvmY6KSON
HlNENJV5FkSdzxNWdEb4Qvpzq1KqLu/inDiKSoic03/LBI2FIEKKLl1VFhwe2WWn
QqwpsrZlSN5hqN9znULJOEm8B31lMt0WhdTuzvXHObN37iJYrPQ6NUy/IMo3Y8vi
pkkMdWbsASMJHR8jLXaZF+iGEO7lXMGCJzewUpijaJhx28E6OJhCh2yWC6SNbsVe
V/9lLBj6e5l2CJOXXX5tmnn0JwXlsJ3LFHdUbPwSUXLbMm2bRBfSXP4cYXkyNA8n
zwSUR+FqgWaPn853XEb8yPSJthwOpVZQs/iUg7s5gLR6i68SJC1sQalf1C1qJ7SQ
M3UES7sv1OxngOzD7cMqJRRyUGg4Ooi5Ytr1IkQ9p40rRO02q6oo+gL3QoUCvkAx
FX6DTZzXOXD3iCTeoxuFQ2piWI3/hAty+gK7t+zrOKPImQL+TlFPyo1r5dHsJyoj
pe72z6Ph8loRMGj8eH/U/6718WaC6tedXmO6FkfWyh1Vn0Do/YknHqGeOpN6Y3ag
WvilR5U+ZW6OIiFUc7ki4t1VzuUraRZAW+oqwi1KqnUN7dhYf5n2jXzjflmy4stf
Pu/f68VxxAMTWQUAJAv/X5WOAOQHgAexj2eI8y7Wb9VtUj9CUWvsDdqwPGbO9/dU
66FMPwo4sJT1UCcwe0HWAi8Qf7J+BOpDSz3kPX3Udfb2PETwPqu9nzauLmMbAtyO
IQDOO992w+iDdq0bM/zjDlxCP5YcD+rz/etBqTe0CL8M25Lejr7yw7bcuIP1dtOG
BKG5YRCnogRqSN9UQOlK/27ttDVkEyG35j8+Jg45lfkR5ITlxZXU3+XMWl27XVQ2
/RPc/8COkiYEHG5SQBKaHXp+MQ+dmvJ70sNuTQZRk9PUI9LqDwvag4fVUtycwQgv
ZRbSoMKN6LmQTLw5YYejgfCLwvVT0HZT+cP/3yEU5BIiBogWa3wyu1kuaAC2KUTW
bh5P4n+zwGOkyu8Cgztu7MaXBLO59qCraqYOkbfd8a2Iw60PbIWwnfX70HJquIoL
uKf0ORcdZBTw5UKERub80AOSU/vlFmefOdBQcfVUiV28Hv8TO9/lw7aUQcN1kOFw
iR68wRRsaVzzWungaFqtwu/sjW3G2ICfN7bx0fWN+jYbGAhUB4LuKgRandw0hNNm
LGINj6LpAptrCS4Pqdfvxv2Wo2UJmU43SDA1IVAyf7rj4igzD4l0/Z70iz8SDueS
F3EGvy1NCetLitKp+sKWtG2WyWn2mWVfvZaWKgxgiCFAdi+JcnLPsK0qJX4lAB4q
yBX2Szf3XYqH7Uu6z0Pp2MaVyL4iCj8c7MsO7ekY50o+whBXZ2GTdlNYxvtPyCNz
iixggfJaXFPmBUCP8GDNnOD3OP5re4mn4skhPiXEIHZ/ETA1fIxZ+sESFDo829E4
tmbkCcBEUQpW3xZMI2XBBms+7D/pDsGd7vJx7YYjkr8TWKO8zHJTDuZUGTI9aHRE
5ExkeQrlXLFoePP8alUrjOZHp3LT6ddQf8J5EZaUVopf3botrv3qKczRpJ2tDKgy
6fr5RlaZ+B0lwYZPNMfHFT7mQAJWGrx75c1qifLJbyNgx36z9uIBTfyY8G8BATXn
fHfmtcUpGjZu++I/X4xCmDDnnRJKLYRnUlq4BzOTEBmJkzei0tjE55dUZ+FaWclh
TjU5OxrMkX5POm6ViQGg+VaCxbw135P9kinwJGcmfDjNa9r0Rcw1yS+xbhASTG8N
zgtlrfUt30S0KSXriTVGjV6yXTtUQYWkVr+cvQmh777vo8ZZ3cy12nq6MWJJU9YQ
7sMFYjozHWxgZBHzCg0SZ783tFu0kJ1wswEHowYSTszUfrzlF4FOpnuOAOXyajMw
kUlgi3jGJBLWtgCqYS5y8uipVuLfJHMvXHNKW08SOPcXW44eobxfib6umPt0ip9E
JuaqMOa8pH0QcjXNBtU7DdNJa1aGvqDcQJV7y6QQh7hErrpWRkClejaUmfrD/Sd2
sOsxZjd/ntRr3NCC8vdAcnH+KmVvLNScIjhd7mBSB9CKhdVecoqHYarpl38ZSXjA
Qq9pIGH8mS5ihnePd3yt59+zmmUjYHjTpqVg6LBhw9iQz3GaUV4cA27mUt0accWK
iE8zINgACsmjAPYCXBq11iLuU8YIDH9YZadWY9JzgExGFC/0VS30heFM+UG/lBAG
Mri8rfI8mbhGVC8F/P+zvv60CHSDZKRqcUOtPP+2Mk+JaAqq+nTuMvfx40TI14Kk
iuc0bCFKY4MsnvryaOgOa9MOIcOW8AXQUtRL1pQVfh/UnF9slbiuq9OqmFGT+hmr
9WN8oo+XsUgXGYeGufl/E4gTvT3htHgW7n0Bnasu1DzVhiQd3xB1htFPUuJGl7HQ
dhQoeeZWfv8McFsWjKJ1SjrJJGPuYYJdogseXSTFOV64iYi6dYRd8IP6oFIlrHcI
1FNcfuhRx+mbDdE5hDBIjmZ84CwBtAKgEiYlx9Mg35CY2iWfgd6zrDsSSGGH196f
iWcXkJHvkl2NGyPVe42nO7f5RYOGwNa0CHz5HU0eeCQOLpvWcJFc0Sa4jrEoPX8z
xR5YzOyIvfYArK7a3GJqSblk95HNMTsD8uJA8MbH/WcrbhT8ALX7AV6N2/YWn25q
QoMXEwE8Nt12xtFO14wcyfocWWx9+bOSekfVGYaT25na6osqFBjP7M/WuIlg2Wac
0TNqf++u52EJE1oe93UsCqmSWY5MpFPX8LXj5dd29XfQXuV37i7PqnyV6u4P8aM7
SU8yKqYfn32+SjcDtB2v4W7qHZGztMZ0GCdr0VPZanCbThB/qynYMhndq3VXzuFU
lUNehwUG525kqKsbmrJBbKg8+I6eGRkeOoRB9CxbY6MiFNVZAUl+riZ0OnLN6Jyv
BVR/DFeh/beBIT2cmdMOcUTjdldyVfIfrlNxXdKNUnFuifOxRZ5qXWxVR5RfR+nM
7yidFbmh7bXz/vfg6i1QatvndN98ag+UtQMyWeS1XIHwNG6ujHp+9h4xotzAC+js
ckbBzq9U3obMDCiXZeLqLBR1+TG064jpkj19aCNY4u/TS6zVtcVhC3pFtfIpCTFS
9yZeZhZHSLpwvxmeQL1v0L8i2dB3ACnfRlH4Iz3HznSeckB99p58Z5ZOfMSRJInL
dAitoEK27YXfIEipkyQVRh2/WrgxLtdGFQeBQfKbFALe8hE4gOuSJoFSM9KAXjg9
bk2X+dnCfNA5O5JEZX0lQw1tdxB01vbNVheorxGtmrpPmvsTa9adNE392rDVlaCI
+wUwJp3OL1d/dglwmM6L+43A6I/vEGhKYoRr69cd0rUH5zgUI2TMYfHqUYXkSl4w
+T2a2EXKLdy9K1aZ2DnSWIXvMFIe/79Wac6ttX0U+je5W7TORMGzqZK3iJ0/+tv7
KvBQrb/KHg0brac3gCa248SUMNfLDOmcsKXbO/5fL93n/bXURtK4ROS5rSIxTHoe
mPrHcci+WVbjTMrEwVVSdXecEQD06Soh6ydqWhC6EG3GEHSnAT1E+Ur7l8908m9u
80Cwm8uuJkmPxdJqV05H5wnUFsrSsiYsIFYbBN7IXjSWx43jInro4evVpAvjfg2c
+hj7qBi5JRftnXH/X0wRSM7Lzkp7bCAwqnZkb+BuPp+exM9PpFRdZipmqEI1IDUK
SFaRkmB/8jHRbqmqJ5zh/4ROQ5NINe3LxAyOisUXlMcCJ0P0oWErUBstu1TAu2q1
skTQCoZKJkly9psfRUK+w7i/tth0m4v17CxIX4iZ9lgIuVozFLOdQDunQHED32qt
pSacCkoyConF7vJ6Iw0ldwg5IRpuRjaOSXvlJGfeTjLF8OMdB2m2EgQ6LmY7XCk4
iVsCJFbnNxzbIKDM3WoP26vFiSzGHGCUUiFeJelCbZlcRwKd/0sh119p/xHzuaYr
D1bi625ls1Hjvn9z4Ci6Gm4Jly+HEdZFkFXP81zcsbpGKfpggfSSMcRMec0WegOl
Ux3QZOdLy1SaoWdIVotpMBc8uJ/womAIIjRSywcy8/XfgaW7IYxUapFk+SGG6tdK
j7I2QTrHM9VrHuuXuAlvt35ewuzEY7IuZCMJWGtiM73J72B/TuWwW4851aAIMD0T
uKmIQ7CPrhGb1oQ6P5zDJUcPFlfRX1xYxXMJNl8Xg2HEKKFIajOS2wlknk00/xHp
8Gl4/g8Gwxik/KcLEwhzlctpfzovGdPcc7iIHO3yLsG8VfQreFfd+mvK9RnLhnU9
LMyvGJyIc6+6W2IixvGgX+qhQFZma0o2aMn13AVZZiqumMEqqX7y99rsZU15nwMb
f5JTNj9iVkmRXHUIyE9elgVvCQp93FuC2kvSf5zJz8K1gyT5BOlAbzViia1l9YMJ
lqhsfeJn5Y2VdcvBl5nwwANzuSjs+2Jl9o26OuoDiWqqrEwizrAneqx6WSlFp+Ax
ifUcRNDz08oBc/EyCPop/1E6BjfUtjpf1S9DPo8WW/7tOA74gBQWKJBzcj59NAd5
qBAy6Pz7WSOHqQ2JSdtNPVXl3Lje0RTd4mS+90PsE6sH2hW7UGbBl26/sckq8HJf
v4OIiOkFuI2h8EwOqYKdZ1XJrDUdOn/nqXz5NSD87/OcjGNwumIPQbzLbIebN2N+
IMDXRvrt+GBjIMD8pV9iTBVxXpPVsar5ccgfVnE2X6iAkWjwAv1OC6Mb7bX00b0c
ibfegqd7NT23wzEt9CNiZDAtuwgu73WTUHnPGRAhWa4BxSAZwj2SMFZTgnIonHsT
Z6dyAZbkqawmlplqxdNmtXCZkWCbmrVz1eaiJflfw6biZXY1HZZ41jNMq5pWA04K
J7tc2b6bVpmJzibul3jo5XDb8SP8i/Lzz9eu1zckjrW7HTpFHk1xTN4YfVqVzApV
pu3tsOZvcb8GQWLlZTiTSkq7e9h8poSHXZq46qU6NKHV0whgtwzUbNNYhwoTqEq+
sq6Go6NGfh47W0avuU7wRJIzU2fh5hsULlN5JXjnmG8n77sT4eFVX5Jrg1K6alUc
/y+ugYQ32IMPiNEVZIamofJJSla2icyAal9Dpaem5wBW0IfyZUHVi4k1aduCRSmO
iAv0tCI7fgloQSEklGIgXFWXL9vUsadjkcM19PCASpd+KCzqwe5k+3vCE1k7eda3
IhJwT63hh7IJ+Gvb3TMQ6wUooAliFCixVqnqFQprZ+xXpqesNlFtlcROr2msfQUz
Ak/PUj9fJLllZiag1z/iMnsovA4n3fil14DgaM0bY3X2w64wAYiU/Rkg3uM06saS
kGj5aXE1XchENhnqrxe8clhCvP+FVkROBA4JWhoMsQW8Lx4s/dQhrwKw6RkU1C4J
jwO5on1GnKmIHfjD6dGe4uoL5nnrVgkWIfnu61UW3LyKW3eCdVCRpqM6AUwv6mhm
F0g4PgS/AMKc18t6OhN5nZRAjKYhVzuwzHi4xln7sdy4pCjkt4XlN5IUDcW0JJUV
UVRO8XTKj+Graba2B6drRBrx2rxxM7RencuRMqMAoLD8JjjdaoRFdVTDQEccunt4
M0JGUfI1WWBokBDUpNMteTi3Jtu0QrtcF5eRYxoTbFJF0SGNn2Stxlt50+6t9wIn
cx5VoIwypsrckKH4uX3aQAv3uNW0BXsRE93VJ/fACkM58ojXS+/my05HaCw4iaUc
qAWyCJCqYy/ByEslrlx3hsZU52xkaLIwMIeLLDQY6MDTencz2pNro2vfajVUBDQy
5voI4MpDnV2eaPxepP9e7Miruzgtu39BZkf/RYBYyxC1rv43RY2sWIDnow79ynVe
qFKE/neJsgnxzJctguzyMsdA8yA1BmyUCHeC716KlJQaRO+XB8t7wAl2yc5rSvV6
dUnvhexmU5Ufh85qfacm64DNkodhtECgIOh4DbVPX9Q4ABJ0WPw8SeSe+QOWHTLY
ig02SHd/rOloM2H+jFt05fmLL/tAR0oWOWFBNo6/g+pl506Y1Nv0oIZjwHsIoZZM
DStq9UuHMcV0JpHBCKpNqmavphoQNfp+dTgoA4kiq4FBhppYcRXaJfcvwmOvqiO6
GQ7CIn9wOqSaORV6xotDzVhevbWEXLpPrXNURZfKRuua10bEGVQ12KnIwBJoCGY2
X2i92umdTa7iOP0k7IHWxY5LCsnQvXYOftwF0HzhMS/MaibNxO2GanAEkuIJPtKD
78FNaONLlRvZxTZy0WDheg7KJzCg5z1JQ3lpJt8AnDKyirMCaUhDoUkz+it6KuKd
FCZfAjoRj/ufB8MdSoXf3W53QnWqM3+/i7b9FWs29toMmxIZKPnTQGhor4bI7dBr
lZHegPiZw11G/GstjcoQHYNc3ASrBSF0/KRSZlT6Ur9v0oqesflY+CCPY53zwCL3
ws4MypXYz+bdt9c/zWhqQUo7qfH0oabZRFst9dfBSVJ9oXpcWuxcg5EoTDPgA62a
ZiK4gqblp1dYXGWjOoKIqrPDLCvKmhNquyBywofxJAQgkcgn7NWwYM2SHranynP6
tZFzqiLAOSg8IoLNEvhSlgA/jArfap6P31bSq9tHrPCQtQswLwjVwgDKKfolYw2h
KGuHGwK1dQMDBG1yLUcwMsHpr6XXzbrLm71MZ2Vnaocoa6+auPKIhiSnDYTPrqWI
sww0XUnlUh1wkTxjurixQJBHwLCxCtZQ8wx14+2a+EEyxayUJxXTC42LhrvOxISn
5g+EDvMzCtud5HC+f5TxWfjaCAcBAm7gx92FHeaFt0wkxaVleky+DmpL2CUHhuqY
zwbngZpo0pmCwaHgg0poTtUem5851Vitx3IRsmk2SIadO+5R9jkf+iWAkvz0KnbC
6LV6pOFHj3+0ygh9tRirawSJSwPNtd49PxdnMEeOAh/6rShYUdynzMSpaa9N4emy
8ocCTs1N6UXlGl2tLNnBe0gsrqp8PqYDgOf/apN0oD6vzEZAhHhf5koShnpqarfo
xI0fkvQsAFZmUb8bJVcu4Z/HIMsNdb4oC9ZADQ4om044zErd+xzXCnj/NCc22+o6
2V3IYni3Mi0wLVKKvhyZ0XDBlh5h4Wj028F2uddNvrBfaIzXa2E87o7of29He3pf
4dh9ocoleZCN4wNbhTG/D6OwyD7Ld3vIfheep7y47BAdQMULOCFy0jZ7bp1rrSmP
FqnXwn9bYVO/69kLWnaHq2wrBoQbs4VPCrWU6itH4xS4dPo6XEvzbCfHiqvEN0qN
xmZRj5cAg5T94t+CF9sWt+5WlJdwgL5pqwfKu0FxFy5v85+ruHMXtGMln4K/ZHMG
obavRD8R5NJLi3y38RVj3YB0nG7AuRFev76FbyNw9ljVIMp0UVtinCyIc8Fl11QD
Uaw6IK2ihLJ/Et2UEj7m+4CmCOpduw78NyB1pL3hlmJpb65hmehTb5Yu18hXuMAq
R3H5B2FfMysLCcPy7ctRxCHq/5B/Vbm2wRM2rFQLv+5xnwpkph1bEg5NjKgJwGhd
cSQ2spN1NibHFM7A+ZAh9bX1KzgB+6mk1Y3WIgsO8CI/3jYM0lRKfwd6ZAUfOQNX
LajoDBJH8yhZ2pB14k+3e6AjrU73A8Aau5SWHS7D5XfWDcOXsNsOFUNSK051jxrh
CjA703H5GokAYGj8GQFev6Z7731C9VQynwfBOF9I0MlSUicn5O7ooTN4mlc243+Z
WwYDr2ELaj/DRw7naY0rW8yqM4vcIbwb2fChcBcfBrjC76O3hJDtocGDzvgbiMGJ
dKnEeMp79gys0fDrkKrngmk1RIkg3v3Urh8wpkq2ouKBHJ8wPhNTxspD2YGIkHMo
WfTK7fxgbuLO9o1DfDOF7y26Wq9fxXEXn6YdCuKvVPZWvvIKa+nyQpcZEUfVKq7o
Vbm5p0EXnqQ87lkREbFngZaNI/kbanBMWp4M8fcXn/eYWxan6hcwmkmBIvMzEeMs
FlAGp4+Yx+MnNZvRrwQGjKhydJqXnkQK/zCglrU8CEKBYpmsx6dX5mdWUYhTcNSs
h14kGSVszxn6TbQugvrgW6fghOqrf83ZauclYAIw4GrMQoUlalFczEiDq+Csnusw
H48pUBLMIOiFBI2Zmktm8Wot7DS7/JZzfuNyDblMlMZTg+l06ZtGtevvtI2vqnsI
esp+wBkJH5D1SIIiN/clgEE4zV5kjWH1Ut3f7qW42rTBigddxG13UnZVCGIgm8We
MDeOxnwSycjozEJhYu6g4QPzZeb4JAN14EF8HZplZuGHHJZbNSxQ1Qoy/HFXh0hC
gecIlbMopbbyXsSvDtfiw1xHFgBQ32q0BHVj/939X/f+nBjpdHrCcWR8FzRTm6xW
Dpcu3qOB3QNjQ1cTxLYG04jUA2U/xsxcnko0jWUVej8CELFVrCE/ReCUDfSGyViH
NWFHcIdASJFN8GbQChEl2+L3gZ2NVj+KC5zVJNHkEV6+W93V2USY3Z/h+b/3jy83
lSXl/h37ty8LnCDCfDKDlqIh/tpN45XRqht5T0i8+LoLN+nNSt2EHdmEBB96Ywtm
HR/nA/EwG/kZDKUitYvQbbYj0iPVpz9wAXUUyheRZZgAifE4PawCZZ8BiquYDT9Y
yAJdbjNYw4bexMoLbiHdIVUC/97GdoHFuPGfrO6wYeY+75Ot9WBABGPSkJCX1RC9
paeXjD24sKwNr5YbJF1LID60vyWzzOfR/PWke6gQrGONDQt6A/kuMdXlbvYXHEf4
C+up5df8k09bb647hZlAhNVanEsRSZ4eMZesroapHce4gP8lVTUAi1YrkBcll5uU
4c9DlA7jW0uee6N1fq75dHN2ydxTVTrxRXqOIwVhdj2HmWjOO7X+MHShkUQBuL+k
RFjOFj0Gv3LhkpYEp/iymioSyPiGrvvQo3JQ+gD5PvmggYORzxGcIycD6F3S0lr8
W1FEFIgOAF1ziAMtS+VjoRq1TO5T5+USD0Q9PxeFEy35zwSnrqAzot1/yRNweYte
lgVQr5alw1WGpEWvZh+C5346AbSjfP/gdSqR7DAB0Lk82kytDRtGPWaeyFd7Bw1C
Bc3IDOC5Ykdb5LOxneoY+d9PUQn+6uUtvUBsEMpRQ4fxYdOMnWcCRawPq8sm3qsZ
7o49dHame18+kGvYB2enlJbw9Kz400LtqLWR55SdQBfOoJawcxwFlE0qn1IKXi2u
q9513SaROrJfx0I+HkgmcelQ/cWRPI9FqfnYw1y3ZPHgfVZ0iP7gN8s+g/i/6U1v
AbphY0X0vAA8rOVa6+gLlAXdrFjBWOZUdhP2bXxf66jkWIaVICzY2SYhJG6FH5/2
re0viBg6dFIQbJJRqU+Pz9DNNQw8iCrsJ4xOdF37TLQycGqnqWVJlvNsD5HbgXVo
SUcAQvh5lZhc2/ssXv3T2pDhpbGz/TgDR+wEBHMIneVvUeq1nBachesU62bIdYtQ
nQtz9DZttrJMo/muOCPvhnpF1p2T09FEacJ58fPNeeaIKLEtboMp0wKNAXFGg32+
xuNFvlW/4ZXbzvQxSzTaQ0sxsHiZXVu7VzH+mU+ZHWSSM8877t+wClFPkKjYE4nL
YTgAybI8Dcof51Ru7PvBniHYOzJIgSUidz8q+GvZE4H32TE11Bj4Ei3gP9c72buT
ft79+eYtrFhysLvzINKrRlVU4gZGxkjS23YNTQPDGpNOdGAne0u9iClKIQ/lNd7b
P7Hk4jBzoQ+KUbR8POjlNlfiJGuooahUEIV4iVPBNwXe/aBz5UOqXJ31Zd3PdXWv
KkppPBdSz/iXamD9TMIU8hgPMRBmIWkNuy2ghQ3J0ja+hm9x649BK30MJAz9ofNi
4DY0xoNBLSKYcRXJR3TZnfkf7Dtq9Vn0L32lq4UJf+wvi/tcAVdG7c+K+heqqhLz
YAVQYxCyD96TDe3lvvv727vt3i1tvzVd0dOzI/1OSKLsadOlQfSIQ8e7fPxaPkG4
`protect END_PROTECTED