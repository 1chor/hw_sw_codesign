-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
G1lZEzblNhCUd8GHDMtPOC7+2HeM+Dmu2cXCN947sYXkBlymVCyDJqZjrvPZCQCE
Vf3VjhMNsrm6pJJMCMjkCQQZeAJE6bHigEqU03lrpEW6pE5j8kJ6BZc1wqdu9kIb
uJyBB1LYSlwVT0Hlxc6NpGh3H+/dshDnDeBJcmJXgow=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 19885)

`protect DATA_BLOCK
YltL6rQ6Ca7TB1vvLhUrdA6M8LHaqE/hc5+uWabW0YufpBVIkaagQCuSUG/FVPwY
fDr6zGHbsmHiG37VY81rgfYIMpEVr4w8OO4g13omrQMzl7vLNRucHG2qktWKWVAf
udIChnolNWY61PajVDakbSFtKz4GUO8779aXgNRE2CuBQcYBouFo8n281j1G6ONY
Jad9HFVbq3aZLFliuXOpCStoklC3F/qLIrtY366pPavOcyHUS6eDcz1dtHIqFZ3K
jYQRD42/44J5Xny56ODU0aCWwe3gZTKiMzVla36ysSMCthLDnPpztj5Q63SM8w6r
4rjPM26HE3ewux7oRRPV0CSPNAQA8PxL4ohMDLjbxXRgFfqQx08OYEM4ueIppQDS
+nnB40EjWqb8fs4MvNluRo54wrJpgh9HnirGTxA9oO2TUhQOZbduM2XV6JH4xMkW
AWcB05WYP37O0UPQeUIv/0rMzIYkh+pyU45HQu9qO5l+3QKyycBtNLApjC550yMs
jC2ihd2NobSQBmWytAFvm81dW0euUOUaJK2taPwdxxQRZgpW41AFEfQmrrnzE8Lb
Lgvz3KaPOs7lyJpFrdsR8ddkg2yNr5rN6W1unFSg1lgjoT6lwAfZRl89bwV9uIwv
BglahLjxeSWEVporhmVeQxGwbrUGIhGWv7T53ou4+9+NzyCGHUZhap7wi23hjY92
byvRa0AaR3PaOjMzfpqdQOEFDYTUwtddUWcsf20ZeSKyjv+Ue1K/moGx4aMIDXs2
0HwRLc0a6pmtbKgsxHt0dRg9l166NLE85MssMecrU2kwTphbIBlkLHOIwWNzq+l5
QAhn+VFbm6nku13s/fXfVCLA0+bUYQ65SwiyGDL4YMhlObsC1qaPH6YyLICr6EbC
2hWd9osManqCkoxV1bzmfG+/YN8DAIPC4xvpuu4MU5oIAM0nEZSoodSxjA9R6ILu
yGRVYkdSm6jDErYop09h3dhKgyGm/+26d/D5DvgIcIVskbLHiDtQYOPXjzZQFX14
vO/YE1jJDdlIKidRqXfHQjDMTW0XTTSkXmNKnZrUgMaRGK5ttAHWDFthsb4t0DXm
vRIqzCx9KabrvSzil1kqFCuXDgIRg3W4P+w1Gp+jA00q2SZ/yFRwkP1hWLiB5UDv
yxNIGXhbvSSPHChpyu4kwRVG8sLXC1sCJiCNLKO59kRb+MwSd9VgGPoTU/nVFEJv
n9oCNyH5chyKg4WAnHIJpExLLaQw6FWS9lokUpLzm2M9m2WxHho4hAL5nVAxd6vg
Nvt1TBdNLIOr8Uo4jQFAt/t23QZSq1IcxpvZRGxH1LT7mFFUZGgEjDotGHKlG3Sl
jZrFVfzP6tR9DOTEHGoP75G4dg8Gcjdk4acSw6jkWQL5TZq60K+eYBJ4F1X/q0i5
SqsrP2HQ7ur2xBs//xt3AiNT/8lhZGBHNrdgrnk9UD67yKWOWiIv2fzQyOGmmAS8
4j0Rqbb7bgR3CopH3Fd4inSl+ZixOt/1duqNIDcFceqh9b2RhsQsBFScVBDGz7Wi
uGSpAENN3wrFnkzlmqqWfBaqpS3gZAbn7T/xbZQPh78yPIy+ksuXdFeCTDVJxPM+
djsOTfuczwA1FUafXVs2qew04UV+vxidImFDwsAY5beCGeVh2RC0iD94MixJ9N5z
hm0WXFKQsYxzhUjN7xmdG6s9M5GngkI4xBQlvpCz5d8/meeFgsQIagTqOdRimYv1
TCumjxH5ARm4gzuQyE8NXJc4+WOovu7Yf0XJDbUGVrAAOlRLkZPL4Nx6xCfYMadT
OgQZ3JiH7qeprOqDi9vlGtdx2RU4rxG86/YKYKpWzvHoCqg3PFu5jWo/aapGK3QN
bKV040B8K63TjXrXcja+oXOV+xjooZpV9Mh9yZuc/IsQr7diSulGVFgkuz5lCrb8
9NYTM9dpKFIFkZoy/l0Gw0/0YRehfc8TdW6/nV+aSJpSDlraOUSpMlkOtgbKQOGd
5LEFbU71YEYjG1CYgANFhiu8S2746Z+Vq1lMR4PWOGOw/treQuHXGcRoSjEHM7z/
Vdlak3AIwC5Djt7z4St019Gb18pkPvp6us2OQC5FAPvVkHAMhMDBecUhFmIvxsw9
0BiHQtkR+WNTYbI/vHdB/VnJr4mvNRRJ9qg1Q6zp21buqB63fJVf1MYN6DddU/Ue
rfPrWxSx38SGetANOR4wR0Nw4XHzg1M7ai2X0iBa1tjmc81VmB75uruKrx0E8rgz
G3VanufQMivYgc6RvaQfKpTy7CpwGeMaztvdfjt0zqfNHsEKzQrbzMLXQ88bP6/F
DCS7hIfLgm8kjibtUtA4WBHl20klY6tRLk7xh2HRTsX95lvwkzCE+Na3OKsgS8XC
cOcgSpe/WVgwjKS8sIYY5LcVivqg+JnKQ5ISI2D6djL7E8Gvu0K65keZRDatxAd5
YqU2T2A34tQZcQK3NNEJuSZSW3/qGbO7XcPV9ECc6bBxlbg8+JJfRpZaEXC2+XgR
FrZr/dcD5n38fwf0KlzlOwitvHTSMx+03VVBG/WAQSg1ldqGBYjtLG0CS+lSZGJB
Jeirc0AlLOkwNjBJTUbTUX3dQxi4AMQRSNjYVYOEBlUDU43csb0cFM4/JPlUkSMt
gCxPgyGLsOQpkrk8MMKJV10HxCrqUir46H4A6EufoJLonpAAeEDL1cQyhHfcDNw+
L5m/vBwDQZOGpvcVLVa8amCui0mNTBdul073WR/73NyZuoAp9vSuprzXTspJrAD6
XgsA65HQHa7q97IxCBhyhPzy/lkT7etuhPbytwrkWKTneXgsFM1CeNK9fev5h50Q
DW9zeXLhdKtJOLNE9w7cF+c206ZZ6h15y+2tB0bn+CxdWnvh6PnIqwXBk850Ldh5
7GBdgKbNChIa9FaLd4i/m5PWDOcz678UqnNShrwW51xWFpWz/Sn5ZtLRpJJTeDUr
QxoOOOmH0I/XReQDR6ATOdiyvQBmISzpHlMIZOm3XSPPE6LluLANsBr61YstzGwQ
/xqpOBxoKpQuExF0umOjJqllroMrU7XfrFBpGRvFouzJCGrm0lWlnK+JDKOuWwm/
+9yObGNphLWWJpzklBqhfDqeUWfW0XSHcRENDUzUdq8gQ9UllnFQc4jHatypOTMK
ZbtMArYrp33RVxwMMhhi9ueep94RYw/Bis9/vap4CvJzOH7tXl7gpNG9KAJ2RcI8
JQqakvh/VJE4x3t3pMzJyrHlA0zw5epFsQEpe8RS35E7UXVcvQZdghqFK2edTNJi
aHw7dXyT0YpQIUbWexx+LQVclz/rdGetz16FiKzkABh5sQZomnlIZKS9aOmCdKQu
ndI6QuWzDw5ukVZP27rXQ3WAfmpAg7i6ma+ky/3TMjon+FbmHvSeJhlAZufErNsc
pi7vNtf1XKAtDrJ8oVGI3vRKJaRAQWuMFMaxHmGPCMC9JYX9Kdgu3VYSUUDCM7Yn
fxGCOqO4o1ukZWFb89Oi0EFH5n2yhRDqZTjZEQsqXg/ZRpwIQZiE6SLTsaKowrtp
PEby8QBIB37Wj8ansmonsBCNwveS5E/JJqsPe6lkMZMj+CZXDiTf2man1ZI8SNvF
/cuCTD7+4cJ7KHkQAtU2E+9wBzteAHBZck1BeXqJgcelCUNmejFqulfcvohkFtaC
lTGaNwovGTg567P5BDA1jzAlfC065LHgGnipBzvJITs93GAb1GWhWXhq9/aYP5vd
mgvuZpA5jt9KJxyRGX/r6BN2oTMs+hrTFcbz9e5QhnrdxHYtdxjN6wlOtz9xD2n6
K3R/7ZbbuSyRActUbb7QBYs0BcS3PIVi05UkJKDfpp9eAtjW4OgZHKp11cPV59Y/
b8vSmZK9mgd4E8quU9vt6a016U7jafYVXQ8J66fsd9eFaEwWYYsdl60ye1VjeA4I
qw8CGop7zUB33aFOPicShYQ9+AYZMmPnszFwKQfU2NPKNtd50yiUfRdaFmuC7cIm
Q5nv+Lawbs5qO4XwGq2pN1K75czX4tD940G1rWC+I8Q3A8DJCgCXVY0NpxO2Z1vZ
3Lfz8K3cHvGrziEC24weHQ8TN2ARXiBk7Pj9q8EUwYNdZEXhK7THkMWjH5fuLG6B
c5Cxcp41gKnGmOnxU91bCDTVAnNekP1BKvBitSjJV+VDgN+pId6copZszjun/oUz
CBbnWsT1UIA/4TgBRmMIzqPDm31pEpBxc7oO10qbt6uvjt14WPJ2eGmbbIff+cS4
KSMY95t8GPLqj3E8dbhiVXIv4xP5oVc1qPAgq7V2WvqiPNUYe1oLWhf9sG+Zqqm3
I5YRNBM8i70uuzzS+YFzQlLmPNRc63kLWshtozKKmr+7SPgbY1TXWRMz6GGmIlMz
K02tkjGEb/jW0vm1nXi4UDRZBnkJt8jW9nCj2X7nBGtmCSneVhARHPjWprWsPVsY
FOnZcaUZYqVojWjz7Ej5DfhPLsx+cm3jcnSgPnZL/AE0JCYBeJbY80GwxKSyXTLL
0Q+Bnm39dohivfjffKF30L8MQTo9gDaAPaMUqytGPwlzQN2DG30dHPdJmkIHq7Qp
BYm/FM0ZoqwEffla1qaK6BGoZLjY3/V3kGAtAIw8KpH8breNxar5MzwQGqu24A3h
f8KeKZ2lETdXVkILbR9o/AWXiMYq+hVJQve2a2OLuvD1ExO9wXi+zTyyw/oErvZP
8FWwy8FgqQfd28FWLjGPNvKh+0GfCXMKGM7tSH3lNWjRCPK6L3VjNJxsKTNPjebV
lJNZb95DId/YypMStAusU8xEaJ1taELoLjvJM7L7UV+WHCmpmYvDON+Z+Q2cwoSr
vC3TSFgH+IjX5IQP9/9pzSfC0kHFfuVKsIiGaMnsdKi92YMev+XyLO199NrIoE0f
uhmmY8Jb6c6AustSjpZ49SBGp3g8EK7yk/VZS1IB1OOl3QPlKrzEKKt73Wt7XqDY
9vmYyQUouRm6LD48DuWrU+8W3T2p3CNFmcoeBCg7tSKt2Ci+56S8mY2lvuuD2BWq
zKQY+EmgYtUkXg383T7j82LgZKD66lzlhyJn4Yc9KGzzXTXw5/w6ReaNrk1uJGmO
G5Ma+Xj7Hf04JZAWlVXRLpfiI1dic8TKG1VY9A5OJ7v1LhWFce3BM1q1WBPTTawX
Z4zLTG0rsxKsUBjCRN2bygh1BJKp6Va4042ppBZpVfjHrTmZiOGn4suH0PDY/Bcw
aXFFAP6CTlsYv4B1xvgygO3VKYT7gxNOQmPU38G1XoHZRTeY1vfEjX5HUNFdATyJ
GTn/ZPfo9jpSy/FyBgLask9ruuFBsag2pUrenN8mxlNQgxmEhQwdHmwaB/mEuzRb
VxWjj96eLkZHiRSP/1Ec5jcMB6AZinBluRZhcR8dcfOJG/rjdl6hLTwYgDdSRYFG
DYUiTENCh0bL8gHtT2MEumXJDwEFVfJGc2dzEWwBiZKPQoeY6ZHA16bXSTo99C81
qDB1Cxf9DH0lqlhsAVq5sZc/xENpW5ffJDEgox9ashlGelREOAsA7Fai3pXffAsf
IgG2z14YfG+Lhm5Ha5FFts1YiWbKS3dTY2s5VQ3CXvDMTkfatvbkuKP/1+pKFMpe
AARBksv4iBlK0pqTGsWE2IWNvLjt8QPD8N9hg8YqFnkwZK364iM58X6xRqz8kv69
Cfql4wy7CMTU3/bGte4XSCZl716Pp4r5tB0Mr/47hNgfKqaMh1XqmQ8mHIr6sVHD
Y0BvhTqA3s97RZvxzvbpdn3uKdldU3h+YWGx3hP1Am9C1xiRnwbxCY1ZY6REf2+7
mQZkuhXFDURwF8gWg4kZHlNcr5+TfoloN5QzKfI3NcWRkg3eBL/6p8KNioq/soFe
M9aa4LTDR+KWYYSwjYq4mchTDZ77VwK0tv6Lrm/csOMfArCPStNQrtm4US7/JkeJ
jqZ3f2r1spW+8vUqWxOuNAoJwxkC/n3m9SbbIMP4b4x4zSEkBRDizpv04ihVaG86
lrX2gX/bT314iHC+Ft0qKh8HydgZFZObRMHVMhVEikNEcGF6BLt8NJ/jdOlqLEz7
IVCs42uwTdnJPHCfCLREA0Yo8adnEDnbG6rDCOpF0xaEamANxgKD+FewE6BMBg/T
wKiKfIGgUWMUQwGmF91MZKmxx2r7RZLfcgk0+YjRiVDAqg2mWrH8oGbx1MMQFIXr
8Ipx2CBw21+Wm7o5TvC0jUTix/oVmXF4x6vjo1r6c4PqvGB/H8uf9ptOKRRH/pVA
SAXeLpMCXCeMizJNwT6+uk29NBglx6iO0Dya1ARD5/nyZJK55N6R33YsgIcQHMD/
doZpmoDk/mJi8P4esHNYvsQnPNMckMopno5jF9+cc5Og05LLUMsU77z11xUZ1NzN
NZ5nOQxPD154FRu7S/Ywzatmf3GlhyY1C9IIHy5AN995oUItXm+I+oUTU+A770m3
2W3JS7AP91GXgaJd+xzZdv+Ym+VWnU6EPYf6LwvW1kXt1M8phUTQfAPbFnuxXAGN
qPIVq2kBxoEvy27ZWRze/ppMD3D/TLMPQS0Fi2D25SwV5wLpjjZ23PYOsuDmk+Vi
g4gw6Co7r2NQYjbgruuYSFiUgryFNfIIrUurK9F/4p9wjXRX4HO+W/GuPlwKki7t
5RWV7UYx2T8uFvlrzM9Sfz+KqErX9J0h/J9lOP1/CcBoUoIRiSp1x0HcOH/Rsn8e
eRT8N7rY0RB5aXfdUtaOhUKY/wlDBCR2F3KJln5gFDNBW1OtOErsvC1/BmzkxUeM
tIPoo4tyDFwSRopVNrzLNVGsWyrgAlUgHWleAp1JHZVRGigT4lFO0l8NutHzNF5C
U0DQGMgyBix9+Xv7YAoUw8JYSB4wJjjXsBKzi4BlMUCGD5hAfyF8t7G7k/euBkHX
w+8sCS5d8AbwDvb+oVquYoorr4NgCf+LWsldsAd18w7mUONryRu9XoxXw/IuEkqu
MlQm8tx0wIBUNH54ELfLsyIeWKJYqjD4KurNGMIOLsECuiDMgSr9xpgkIaxeLfst
UCGqXzmIeueyxTb4wrNVjG/a3sQRzM+dOkEutJLnKwBaPVRnmkDsiHXEMctyKYqe
eMClj9fYb7a+CZDkQr9H9k36W/U9+LjHHMd1hxYsYmzgt0PV7+hzgIMx+y5i1Uzk
gnReGXfjjcgwi/H0b0bzRlzeI7//AOzZYdctn+o0VwjIFhESFMNQ6CfEVpM+pJsu
zEZ8jpk3yzyROzRRRJKMtD8AKJVOFmi8kqjVBB5UpKde+FUjwFi8OVyyqHzh8azm
vYaRmEmqag7zBJXhevyuBpA4ETdsUL7p9TQ8MKAZUP7JKDxzRzHa5tArjmFTPiqW
Bqpn2aGUglrQFYfek4U2caau4RoHcRyzUA0mTqj9sO3LEZG2VpD4RP1V5NXvkQSt
v2x7/brOogKN/KOEeu8Uy76gDTovNcGYmUwtha5H8SqF7Ym9VyCoM5ola50VF27W
A4ntn98zUqMQ24I8necxZoRnzP7GRGtXepAfvECBr8+1LhQTgm/ojHiEad6yub0f
xLjq3J+cQLIN8U0rjq4BZRIzSpZBdT8dN8zqNI/Yr8pq+jMKW+K1CZbim4eY+8yB
RepT62gS48aEybGdTEw6WUh1JspiyHcJnuqR2+C3L58VVu6ii1lBGeboXC15KN3Q
Ghg5ffO2aCYmbuI87Am5a2nHMiar2O1yFA/B6nWgCf1eX3yZY54arQVKHe888+tK
lHLQuwQ5OwYNx4nuHLLVF2n16LBorJxs/0XV+1okMlIdoSKCVh0xNfA32BJfOXTj
DCq3uuOQ2h1ynQzrgNO4qKDi/ApniBb0QainzZTmeAqlAJQCwlN+IqVh2HwsYHEQ
FuJG3Vu6X2YGgIcY3+jzYMkhmyzSlnxhLCmBdo7shWtkbpclpG9t3ELGP1y18Wof
UIQxiihcI31lN2mbWnfnUjxz2mtQ04GgaQWWlFidaPn8hUk0Ayb/T82MHBP6iSx9
vXXbT8+IuYhPeucJslr3Znqq1A8zRM7TyicCZgfqMiO4aqQNGcbmNIUm3SWOAfKf
NV6EEe53kCWfFz4UoIwnmYIkIFprrbhuYn3gknmdb55W88Wc2AEGFmLRPuFWBem5
szL+CDfdBHveKs7/JsRFfol7djPhixYoYmduRiWJetZVQge+RQ9shz/C+IEdZSzc
RDLJEymOV3J3nzWdNsGLQpQ/Wbh1gjkUC73520/lvAwI9ybSdP2XveTgtkQXaFf3
Vp3AV/QTX9BH1Td2ySTFhLaEAyivLGovJXgpSX3oL0vVyvjFfV5q493BNBu74OkC
PVrq1BI/cXwi6TwR+K8mRVEwLet0nAAVw4Y81Q7GduHkIUSr5YAr7WgLTJCwfZeT
hHqrCoBhU8yUDRzM5edjzQaklAaVgdgQvB9zlCYyNL60/dWSju7JmeMGL8Uyn78R
0wb3IR66M3jAgniM+Lh8vmJp3zK2zFPzSyxeFQd3oWeoV81jTu5/8JY6N5XSu/k9
G5MqlVvyydxlzVEREIAXgO1n5e1gopTvVqIiIqC0Z2tez9C/taoinYAWoWkgwz5W
bJ33l1U5WAL8aFiMRIdd+74WZomaPUDThiTX+LiwKy99IfqV2GdHt/q5y7P1pUAG
c18V2ulP/ixu/AChTx7+yIfeIl+3AQxW9ShyE+S581H3/n289Ue6xtSFZFvc85cl
oLy2B8Xz8ZN1jQjTYsSfnijc0ne6hdud2837XUbxo1+XEu4f4z7fHOkbO12GOmnG
wyhxITC8GqA47Fkk8ie8P1Ow2kNhwkW2MKU4ibg2OMjbAKQh4c6qhYyPkqNhm+pM
yAN5CxeY6Z5f9T3nBeTwRXxO7EBipvX5eoW0Vf6Qvu7GC5+h7ob9bhNdRa+dWeRl
DPOWV3F0utZYQhEJE5c7XhxPzEYzXiqnCdMDH8ac/gQkBEW6fsBuO77xHgKybvS2
aJI/ZxR8pRpZSZbnrHDDbMxDN7CU5oUaLpSvVAG6sEJ9QyicmHjuS6d1YJxQN6sl
WFYl/p0PiF86+S607397oj8j+d8zvgtGALi1igCawQZvAyIXDytGa8c/Rd0kYTjr
9vRjDm6bdLy9LHS4EvOyClVsBqXY/PgLndn+2M1DkIjcPxII/eEUfzChOqR3lWho
A5YmGjIeuMjHXtg279tGSrgsMX+nzqz6TA9Z4uPmeYrXoxGaIzwiX7Ln0lggISFv
baxvVkWbNJI0x/199cWNWKMD4Wg8t0pWszCR6PVutoLWo5jAAt91aMCQ7L5ry54k
gjE0PgCkLsxRD5WiMlg+FrdEsvV9HfrOMQPXBarX9joD/I/gQY3YONZDYz9WOS+x
Sq6pmfbOIS9qTvOV7+DTf78H9liVIPczNqlsiNuIMUNLRyaZKUVLXG3afodIw2Rj
amy/SPYCNecc5HD9cEFtlFyKovi8Cy4Kb+7TAfGxom/YxkuxGslm1gSxVqoS6YEQ
JT19Fy7FLZb+FiGzhVXmqTUhvnlpG6+7RRHFE2XrD0QxNqBGPrpFC1z33mRLg1e4
mNrI0TSoRaz2tf043daxxNa/206KWMAVxO39BLIoj2JtQ/Ul0Fp21GqgIDoflGV8
4n58ol4czLY8CFU+6zkSwHht+WL/+e54gkLH9WbCgL6pTRcp/CYXG8Hj/9m6WVyo
4SRoEeqRg6XO5DZvpCCpdAZ26h2RerBg3SniKFle6Mjf/IRPfsxpU9hXzoymbdTJ
TBzZVplQeK8c1PS1v3b+zl6J/mdsxdCHJcQachIxpOvvzBn9jzDhiICZizOXM9Qf
idqaeXsqjNA5lPyOZbDTPI1IorvDfZga1jLwHEPCbQpAe3h8XYyKhKhJB3vqvhWu
jBc//rUq6x7dAMrjsSNn5H7OfUqzKHGCpAfCNVCJYjbI24gMkSIDOjgPx5X3nj4q
9TCzlrvJ6aR+McKIbMS2VTNoZoWVY9kaifVKzyPXtfY6fWKGTgCMqEFPwf4PP8LX
FnaYkEo4jmohnIALgJ+hnEdlQWtVzf1kb8NfaqPfpbPMGafgSS0kPxEkaMqQL1vM
fNBXWOn3CU0V2+MX/1epTQtohtWmxCDPGABGFU7YyeciTdhMTf7VcHZa/JVi7DsQ
3vYMmlo4AkuglYue+7SCycdKu4/YeoCfqRwLgZ2MeKf2nWEE71l52WbfFGOt1g6A
ZOiM47JqZRWkwAV3sjiAGKAAsRlufHe2VnLfKGX0i3KdtqUZZ7GhUidl83fo10p/
WuBvdqFnttpcUDnLWRbNLI9dbYIgG7vxGwLhb6W5eTmapVgBmAwqbeo4GJeeu0CV
TSNY/qgK+pWeAH/2wnN/dlljZ0ORSipfFE/Ruf6RfhR0SgpTp0PGY6bkvZ2ulfl2
L22z359U4pgr6BayY7Xau5j9+1ntsX6WQwH1lQZnhocMzeqn/YYmwQLA7OL2jvd4
IkxKA9vqv0a1JTf/60JZcI0gPPP78jyOQpXBgFK8e1MSbXv9aeZd38wVHlhO+N8j
geO9lZyAyabekaQrHtzhuBUOmSHflwCQulS4EqD3j3eK9R9z+ZP8erlv/Yq6kY0e
ont+2GO1o8lDSfSCNJhvojmM9q+nl+vLF5i9iHRKtR/L5zKDz6HfaEPK0Kly9uLE
fOslsw5MWLYlyi/1tM8TJr/ZULU2kl6GY+XspligLv975cW8uDdVnJbtT/S5TZgY
XzwNoMEy5foQa8RnxY6EtoQH+qjkyi67Q3wEaOwzjbOYiX1ZQSxLfpScKU3gTw9d
oQH8ZZWRrrkoOF9E4anFen6fzWI1JRN+EPX3I6KSPpzpF/eBDHCHi7n3quoxjEUd
1VB3Yvx0KjIK/qMgLQrPCH4xY2u+uKEOS+cdPerpchu74N7004gi1Tf/2gDlN78M
A5mMpvaGdP19L08rLr2cA8sMcCGMZ9ZL3izSVhVjFRFMW96505yT49dqe8q5rvk2
JDyBJ0cCT2GKXYghIiPgvY43RKxuvubNpuTYy/pe4mQNVCg/K3U5dgKYspkmi47e
iUzTkwdAGNGQ79qvcfMD2EKVGrZ+H9dfFlxM7nYfQLD0xI3w9pdcaSKHVFAWMIan
3VIp+ztA8dfD097R7GPXCEYfGpAqURgeo7oBsdNmXq8lfwfS8sVO5rahUqNqM7v+
0pfYllj+Cf6zx0v/BSZ4Du+PSaQ5Dusr/0U4UZPS6lCVjH192slNHKov11RcBuJ0
t5qN9Od1iAeyyPRit5E/Omqt7SL+lGddPyQ7ejiqUVXD+03xMlmLfffJ0P6CdXC2
bbLbQ5khJI9X2x1AVTjcfQhgg/pJgOZ23296dVvYvpFsTId1PDXZXb805cDxAfS9
nNNsY/dOL3dnl4oMy0vkjdkEnJpvE43+fgp+VrCWKPXk3kwN3FY1+6rQ6qTlHZYN
IVwuQUHOUOyXY9ezi+Z/ogLRF3UXJYMsU3d1476HenOfIMCTcp6wN+9fwCxyv/Tw
A7c2UDaw4WXv907Wrz1gC126zHLll3XomtYI+ZIag2XAZSpa6esXGiS7bN6aU4K7
tqvV3wHTWqHzwPTgTzQbJxpam36VKeNaniejDVYG1/hR3j/msM4q1rezAso/h8BQ
sME1YsG0m43k15vGqktSEz0vhaqhPtt5G4nuRtan8PPH0B4m9xyCSqv2WavIL4Jy
pu0SYmRZOvpRtQUpcxP3lIWtWT9u8NfqmiD3iruh7vsCMelNBJPNxX53JxaisrqY
KQtqtkC21htBhLV2r1FSTilNCKuNx/TdX29GdTg8m7FIZKvNlwHZy+NnQxIdUVxc
2m09gY0HpNvGCnQ6+E7E+zAldlQWNDxsH1j+3/iYTxO8kw+FLg3aqH56gvT5xaF1
uW/wd3MQpT+EiKFV5WyNp6UQLZ9CYxrhf/xc6PqIIQQlLUjOIH0L0b5b+QAIILd8
CBC2P6QV8XH/wGanHIBbNXUFNeEaaZkvTysOixQEsHwXg9GBgXLtfKgCVxZ+rmfy
G4fTAZEyB0LRK3Dv8BqtWS9baHpWpx/nG+ZPUSnW1uraxojINrINRldpqSdpLW0s
7dJOLZ0PtCvX23Ba3p/vWRFsSDaDvomY+3vUJV6pPIBZZ79p/wNRpFaV2SG4Snnt
aDmqxsMISIN/QDPzp+BzxlFRod/YjSxABsmku/blwRx2or2JgXF3VM6lmV0VKCnC
58Cfcnd4yiAjaIwJ/M5guvHVRIjXddfqBXuN+oAWChRFXlEg9zV/GMsrvJ6mjErG
1uC3YoHIONBIHJPY6Zg9Jw/5rR5k05RUjI1N89W00HdfpIpk3/3mCSi8aRWWajXV
sGF1uW1FT19t1fZro9pdbMaq26ddRv0VMKdCUXf4hAQdk84RrGLnfbmD1IkpU31A
epxmXA5NEsjWt6ukwJcrxoQlQA3eovMgNGX3m3nzmln9/8qUlUf7LhJw1iXenMZh
xBoe84jH++aB0p/uoUZFJoFNEgk2gC9WT5kgdrcrVuHMnnsQpfC/Y+hwiWCVdJ4A
durqpSfjOTTdl8SSpyOs5PECOH075iQaLPkWetUZGMq7EhoMa0a+5/hoiuMzxYFI
7tMUZ5/mzyw+7JaAMjpQP5YrJSRjvsoPgx9WXHZU4Irytvp5g4ghxv3DKTy7iRrA
RISbDvcWt7/brh91/aunn02VLwai2mpBi3lYAKxOmG3vRqP/1ZOseJK5yFABlSwf
Bq+XvLZAAV4zMzX9MHUd5Jb97KuiKRK3DwEhfJbleSjOvIe3P92NVixzlyjL/Hvj
WrGHQQQJXYU/kjebVEF1szWCUKSLmlBH8zG9w6H19aKVez51y7wrvwEBL8szRpmb
maoLd6JTADRUWEuney+tP0noDHem1gIhrDghBrxyq/5YhOendw1awUuZ5suOr1gD
A/g0rNrp5gX9622sBbOfeJxfVgQ43fWR6J8OmBDeGeQnAf9/ltbHQHtuZxIRDIX1
DkygSsTB+u5lsiTFxzCTiYlCgt2TjN+ihJWOjeUWqgrB/gYf3TVvbv3RpEoljhQ3
ob15Maj7CprX+ROq6H0TYxi65z3vi6wCJjQYjqJaze8pymM3AzXXMupJfonmhtWd
9Ta7ctMLQQdDoUn1bNm2/IZHB27xT9hRYcLnPCC30GsoFrgOgvoM4NdPJY+96A11
OiSSbvCdBGgzxMP5Vb4hX45HpVWJyuygqoIUjZIJ6feZPBmCGJy7HYBXO2gKBGQ5
af0jo7gKJBvQZxmd1i3UVcIj4vWq6/cXQWTNVMkASVevaoc/UWKBkCrra1iAKH/V
aeqlWoS8WtxL5EKfdCZoSgjXtoPJQXg3b9uQYMGqPVCX2PGp9y5wv/fydAw08dF8
QRJIeNS8+W4yw6yMKOHUG6qG+HBBSahxuLx3xCEpcZv/p8hov1UOlSfBssq75yku
Xltsq8Tht/30ittnNt+309WoK+sN8mzESiWb0jgb9LPSoRUAf5BJvT7414wOwvWa
bfxvmYimKSm071l4Ln/BOmgBWj2Ysar+xAWNgy4XwBso0/+R3lZBQpsvggqln5iE
iYg7ATDkf3JR1SA9xkOvBEc4C1QZfVy3mEjShgslhg5myfP337I3Zl+xKsgEvqlD
se0rbwlzGvC9SeR12sbMoi1VsBBpjlRSBvSAMQJZvVAup4zwjlyjprwp52oTb+XS
INM540Zp0USWJW4jTMRFo65P6Afuei79FseJawyeULdpjJ6AeOEBAKxAuXs/wrwy
/Vmvjwl8z+rc1y/2xZjllJuvua2oAJc/SiYdZIJfcVBeIYRFweeWeGZHsX+LXYNn
jrrOeAeYNEkyTAv7Tnw27lhhih8W5K8ngPT26N9GhnAQ04dZ6jWSOHcGH6HAzMQ1
qVUjbAAueGwJSDpEKk0d0GtXfZ5WWlwSIkKwdZV9BR52Sg8wQp20jDYIF7lSWnNW
VkBD2gYJWKZTa9Lr+IzWH2OnYaJiEBzIQLSkJgjG5CA+esKysfCuQq3pMEDPQisA
60De8I6fAHlz8yq1SxA06QmaAeF4ITp/sbIOGh1ZHJR/7CGoHe3kicxTPRgcp6eC
cV2e1gAkRycZKNP8xvdSAUu92ReuPK5xLf5ODHO2iP/wX/utR+kmpf3JKL7k/V/L
gkqIMSn4E1xzSq7eeV8lXCM9fYPD0LG8SgzeKvklGK2F9doWFXV6TyYqjIzvlJ03
KtxTMSpT2SlxeNF9B4hQzqd8CxgQyevHCsgM5+4q4TKhV/DteqcRrXERiVktJ0IR
1zr1LEww8jK5y1F7fOtGw7Wm1telpm/kY7fyeqZIVYNKyepLSu/p3IGUsYZOwHwM
+ZEXmAGSW6GTLDz3vExAG/3XlVvrbbwUrIbd+z5P09rh3WDa8mJouCXDE3a0j0Fe
UqAYDwlIbX1JARsoalqAh31kEDeaiPmsletCh2FUP/qEJJYqrdVu/Ow0+86oGWOH
li1cXkCPYNZPHldMlKjwn056bUVAB9nqzPqyDTnjx95QQ3i9E1llOhCycg4u5b6v
oi+vIyVg9M2hzbqWJK3CAhkwggipd3GrPsCCXVT2h0eeoe5Gyep99smgV17iO7iH
Y6eRH0m7o1tcoftWJvniHS+55h8ds6O941BkSTqEz3Nxoz3CDkjDqneRzvJCyVza
HVm3g8L0EzmTSI+L5zcR6Szq5IGf8aTnlwCTglAYo5cOsFDClOD+EyqP6tbJFagi
doA37ZsDmG0tRDB92vSwSNCQGux2/Ev0tzyEu3qvqjGM1mFKwWTefnZtjv8HYCRf
8gdSnnNsVIail/583n8rMFfzelVRGlUg5oxkB8ndWzwe1rJEMI1rK8JRJxceL5N1
Zc7xlId/OTVEp1gaO88xAmryDQet6zFoWfhObchv/GEXtuJ669zHhtgs8M0F+FLK
yF97VGiXV//3Oxca+8N1JAFqkp8/v3FmJb8o4C0L49rF1cptJVNnr2F7ZQaGpA1t
yS2wYKgM6OD8puoY4dn0GC1DK7vC2sSP2y0uJYlrrtoCcil2UmXEC2I1s0Ioe8Yy
UaS/ZQ2mrWfQjkTPCnwPYEd0KF6Pn4oRwbmYHgN4XJPv06vYcx+C4biPFvdIfZsZ
xMRd0zmXGgQxipxlLztWGX5Td900XIXfrdPem7fkBpyzYQtaBWJUAPv4fcB1pUy1
3szq6bs13gXH8WK6xojqzH3d+4VlyiYx6uZUYhSnUC0MtgrqENAwlW9Brc6TNKoy
hV82twsA9jRvWjCecrBxJA8mlC//amZkT7DVVd8KybtohZoqIcjn5G1GxpyLrdDx
6AfujBdLwWJEXgxYxihAuHDjKKcEFlEXyRhXKW5zQQG3aL40Q5jIVc0JAReDTIyQ
Tixk1yolx7A1rnV+lFqdHnXKUz5EIDKqVV9Jd9gnSEe+cACeh/FYRgZLqrbQIfOj
1orvcjdRldhqbQgeGBvC0JGKN4qzALzBvw4128twzKITzlW3bjFLuB24UXfeu07P
IEApI9UWKj0sl7BND30vKIaDmqlObRtONPFgZVjQ+q2nLUClrIIb1Hd57JoSEJIS
oydCPMoqgg0OAOkjJgLxcb7dkMeOn7yXYeQwokKaY83vCJM/SdseSAXY/kVJcMEG
MDuZWxO2enQPwjzxcaUlz1TTysWR9qH3Uw0dhdt9bW+NIWAIQNF0JXDeFxolmXmX
yEEha/U2ZJSlJwDj0b26Vle/cZzMg400CUpW+Jgo88pn2InEuADx2BtjE/Qq1SvU
OeMoh9knKt1uDmoTs/BlT/MSD2gN5SU5K0F5XREWBKeu1mNm6bqL2xEwj7eBagkr
EZBupL92P52XMGJBTtnbdmQLGA1iYkuxQNiVWnnc+PT4nvFzbZJ+TLgHHRSsB0RK
Y3BxTwl71vGGDl2UOulNBEJEVCmbr5+g/GDaASoPTbCmfaxFWy1SceQQTabzusnv
p4dg9EWeb4hI0vqEBwXg4O+1XrXJnreDpCzOzQbAC9RbRPAcUKUCbr82F6n2BGpz
WI8Ynmq1e2m/99rEZYqK/MLI0rtT9bkNsZijH1Eg22ti81AEyAdmsLaK2Oj6g2h9
Nc8bSBr1qcRzs7zcFYYNbGw06nt+vWUzbsiY8w3by5GSSYfD3mZq/63XSOaMbxaG
9ktspK6MF00IrqejOQRtsCkAzylAEbI7oIIh2k0OVcX+N8TgkfpnRFWQTzfJfgDb
OtZ2naDx2z1g3QN2eRv3cwCrkxOJ8mqqOGr9qc4yQhWR3KyZeea6bjPAkmShozb4
veiDKW5/1s7XtqzuaSofCMGnLyGomdCzChtPp7mGLv2ydNtVEi73N0tonOz7U42+
lygXiNyt7HwDXkd7amg2GBYEneME1zDuqeTALTTAWDwqIvw4zNhtMVeXjlv0m2k+
A8vQtzjrOpoFBiKVNTusIhXC06qLMHNYRIQX0KfA5NfrqhRABGcyAa1H5WfJVqLD
QYXEAntlfrzkGMzgNXhw6ingI2ix+t+c0a3ymQz4faG26oukwOytlNNm0TyaMLtw
HUk0OzKOaSg/HwIVqJOmsPZYz0PbcErQpJwte3dDGeJQmpVENzuP0vYSaPqkCZXo
6FgxhddznzrOwo4PcLquEsLMwVNbMph0z9g7VtWDRswCyydhLVfIlUNhCzoSmtuj
OqGKawVywTZWgKtofJxCwVBvMHfyhtAsgCUYeKSVLxKVlFhpOa46+iJapx9Lo7k6
Xhr8MS5FLSaoKPGD3zQjRlyE036aEsqkhQhB3ZLf6TcCiGTHn5TmaEY0oQdXt4+d
oujHALntwGk748qgAmK9pGARCNKbRJ85pEYAU6X6kJKAdlCIORUgyyHqHiR2A8ra
ab6s55Q3sfQGR/UkIoJSB6X6qh8IspAsbrazKcCch4R0tpPxw7RVyzUdODnMMCae
ta6i4QNDwE6wbSt8mdNKUPN2/54I05rAVoAmY1+Mejq1JBYgqmAvucrgCSJHIjVD
55imkN2sAwBJCljrXi5bHl6WYozTN3bzrMhDHMooMnMzqUOgAlgxBjY8e8Eq9vsv
WHaPubs9QTwNj7uLbhl20KTcbakOFXHNQqg8ZZhAnqlooZKI6uIVa971VuosdRdo
J/gXO7/a9ZFMYmzlAefk9FMMX1cg75MGNZ7ux8IdJ/gMSy18qNQwxwWwj3vfXlyL
T8A/kPX8BX9RZkyZLY+oPGjJ8R326TftIiVYH/vz6BSh0VnELALEvbi/ypp/pvGD
tGQl0fUFQiOP5793OMJRCk6nPPVXgXKnVxAKxtXg7xvRuAp1rxQxYv0SJ1LBzSs0
VbRZhPdhCNQNZIv9285mFpxy/G0wcccit+dcxIjB80K1PFC1dgSJMclP53o/MKQC
wxjzt6Dg2WOmVIm+VzKjaam2JSbUEwtFTnQ4DmV7m4pG9ShJHVTG0LtT2k5wzRFL
JwO0V+b8ob5yDhCVZwrCo+N5iML/4Ht5fJ9aOd3IGK8IoyD46Go2fF5UYK08WtG7
VnevZ1pqqp0z02ML3ja5x2U4NWgJpgh5cmWCRGy3rdZS4eGhygJw5EnR8A8psLaK
ylFmUN0EwSNXbzBZPVj5IFVtBx1QErhBOVysNN40CpyR5/Ivb0gypvC1ZCyswYqM
Ctu1W3DK3w+GK8CQK4WVB9W1LXSSlnn/J6dHcsZNNKoelPgPKotmmFKK7uPZ6Jev
oAt4/gDQguzR4f70FFHui5VwTUQTBudBd+2hwZimXJB/9HeIlo2kOPpnmCQHzH1m
gfnigvqi9c8qyJhRea7dVgpq5KF/Iy+mB2Hv1SNwySbtUA8FCmnnmJSlSANY9053
Wm2qd2n7NXPpNDY/jtZveAjyGrR9XYp4OhsKiC7eduy02u7p+0BEWIjohEUbU+zv
wZnN6xacAfkaSUyHk3Imq3SQpiEzws8CU2w42BFWlgAVgpmeGfbyboYD3iECw0H4
szb9b2qf8Hacu+24iTPK+tJz9rwd0X6+OXJsgT+IigOIWE7AJ685NgcAMC+0WLRD
RpTQtv4W6MEBfsdD8jdOhM9q2ZSD5m5XJaOlnZ307Q6bX4uFPEyIRLFbY/AA1ksl
rbyPxpkAGadhh77lvVLv9sDJxALaNFWttkH959qgW/EJiVMmJpYmurmwDO4qodjD
25+sHUEK44uJW2pinOx5PQHsa8PadEyc0fKnQGssV/e+AJ52UMKOeEXbahPvZLEJ
eIhZ/wVN/3Yg65lon9IhsV9anRghjIzIV91y1BvEJDSnLn2hPBYcogA5imHY94pl
CjlSmxmsgLiLutr3a1tsc9OKL+K7vl+acqm5c0rZPK/1UVxn5ihzmCahr4HbjT71
loStk4Z8M6+NwEGvzN8OhM/jRNgDTRTznFboWjSwbdbfzVBzZIaJJ7+n429/Q9s0
cPKacoeJkcVSQm0TaZGsCtVNyQ7BGf2bLsDJZ6rFM/jMVEgb6+nS7vsgDva9Ru+S
o388p/Xcxf8zh7H4iRZ/2LzdiuSYfzm0+YSW+c13kQizhfnpFY8aWDAJKK3HwN1a
oTu1LjOtWd09Po5WQ+AOmqEvfvPKHi/z4Vtehnk0UJCcefijCzegGkdh71NqL8me
1ZUiVWEt/Iz5TgpPKEDJaZa+Qi50FJNwQsoaG/ykZHvC1JoZ03ocbyHO+JGRuwsk
TYT6lh/pvrsmI2oFEjRR36iD1q66vEiBsuwwDzzeezNTJbmXfv20Dh1I/wC2dgyf
4NofXgkg6gs7xMwh77BB3MHjJVbdFfRg9K/xDcdoMCrU19heTt/N/gXcTTUU6LVn
pOVBjMsRPllrhgTRHTfWil6U7AtB1jJwVUA3ZNSwsvjJfLt2TAolR9BVpXTWYfWr
u+4vrxaH+UnjXgWic4DDDuQyr7Zu+3NavQuHabeQcMmJKnoOvkJd9B7irsvE7dr+
TXaX5PmHm1ZoH5oO4PMlYgm4t7Cff5oVN3xNJq/Kd5qOrYvTo6VUpKarD8mm+W90
CAKZIPEQYYJbHJGckV3lglY3SRNJ7mbjiJ1/rGC4RvDG1Rasg5wIQZ96fw9OKiTz
hmGyhC8B67ODQLVYLbjsa0qbvS3/uyD7BAWlzl2he+n4/9q9mqXED8zg0mlL+tz1
2G/6esA4rk9LVALkC6NOX+y9u8p1wi25BOQF2637Zbjny2lDIXVNocJH1fV8ojNA
e5MxjO+cDsQFFbZBJLNonSvseWs9nLM4jKFmYZEDn0AVvHsCvi6t24hYHTfs4rcm
939+UCDUVfA4HpEKdown8uGeOoLDykZ8tIZdXLrPrr98vihtVR3P0D91rtGrAy9j
fep+HocakMcfKgJBb07PyubK5dQgWp+oRZnFHPQcqrKDZa50g4jP9zwU4QnsnPDn
0I+jhOEElEDL0XRDiQBC9XppOc4sdVOZz3kp00En6Hddah4zABIBpNmjKq10BuZy
dj2NWLNLifz/uKgY9QgXqOAik02+WsmueIR8Q09+u21CpSY4o6D7SCSA6GZGlHXL
Z1x3gEpoYzL9wwXH8Rl1D9gGfMKScV6Wp8LadgnYtrpKTAwgnhlTI135oPyq6vWg
7EWg6TrHxG2JNTQr/Ny5+X06duLo9WWQpzj1Df0gj29eioJKBDSTvIC/Tgbb+Tkk
udKjrdjoCK7JVz7MjtbU09la90N/2rDBWgOI3klNiVI17FwNO8C+RdYCfcjaZiC+
fu7Xh6OLsmmbnSaFy4LJwutRxYzRyEG4+wJdxtiCKdKHXrG9bHdfB+PN7nRLdXO1
bCAXCglMk8Pd/75FnohQcLi24uqip3XjCxUrpaLZlGykkXCxX+4Y/YMldzN9gw2+
G/IS+QmbmuMrcBPN5LwJwN+SROPr7HEZE8Bkrlz8lg57qYwetf5oA/vs7fY2uwTj
A/wiZ8krN3xeabfioSGB2YxRiPHmmpJNdCosp0S1d7jopCUuezpNFzHVdHwNm6X5
Zi3XqKx2wg/fgFvR1xbgKeq8Uwa1IB7Sk/Jx8Cv/gtnnuTNB2y+V6HctV4xzqLsx
QZwcJWAWHubczjdCh8IlXMXRnIdhr2GunFnSAEPZrCUz/gcADIvg8TqOGVE2bTl0
vh4rn7JafV4/5LJ2zKJpoZqeLFx1uvQ4+5+OVbDX0l3yHOjngMhVPOqNftjuMZp+
0TjJFORuai5vksycTLWoqR8s7RiUSd76NexxEG3f8xnLrRt5O7GMDwyARV2ubZHi
2btFl/KFk47lFibJ1RAOsjVUeu6ToxwxoyE6eFvbENt+zuw4PH+jx6iLHcK+bC9W
dda4FL2YKJewLTGDIlnbxMNYtlPbGEXkk9YGM51WPP0KOkTuEP6tpR4HGxurrzZ0
+LZxkE0mdEhsGO3jeJNq8+dCe/u3el3DUniqC9yLf0XJLDBamgKL2ef+VymnwBur
pk87odMKANBcZqrFVbbU9nD9scpQdFd+JwnZZYSBQX1o8X4BovFsxOSkeS0rV14W
ox4kYANt6ei5N8g9RRQ4z9Z8fUO2mbGbNSsWirX+oFbO/P1dgHBn2uiJHND7OKwt
O6aKFK/3sMVQgC0F3COhfTNiytyKjnm7i2Ipkvapigw2hCHZn34EnCSa+7LLvpEE
MX5odpno1Epe65iru7alWnQEWFzxCZhh4qImeggNf5L6miXMNzX9AkeiYqp/FQ2t
5NAYdqH9cc/k+hWDTqjO2LVzkN0CCfaEfmLQ79LXKS6NzTI3kJt4brt2Rh0I91wU
NjNET3OvC5ftkEzCsxFtg7vCfRNmOQyP4VhPlxwj0d1WWDf3yI46zQG+P7JYFg1M
0D8Wdzb4j9zmcwHPfyI2aD0WQZCJE/kL+LrAtPOdsXFpsQG2uQDNBpKyVBSr4E4L
BO+KSkCi0ZBmWp77uFs+Wm8JRy068hYgop/5E7FhQefNXp2GKdqssI7RYtezpsp5
3cHAcJmVtDIlC/GT7lDZxM/uVVsHAO1BauF2rzcjZJkxGHTfJOPCWv5m8P7wU7pe
7fcn5RPCHuoJp8UatDI9JkLQHI6KvUfQaVTA4bZcwosnnzq78nlLDsWYsuoK+74F
awVU6/+9U384SRsvu+jQ8UEHZljhNtbwRThoHrjAmPV21EFrEN7sG8arJiJFaZ5P
zdmIHDdYK0H8LV/QcbyoSWXQPwym/VBl3v3UKYdsqpI6t/IUq1ZJlKymb0mVSRuk
22hejMqxYuYtr838FAl8/aqVvFxBKEqD9Ie7Ipki/XyxKJwTlGfwNhNJvQ3io6m1
lQwXqk+jUF30+BzQlGTjEate3F6RcfDsf/4k7pomKT3lCzFnId6CijvXZ5YMN/V1
lR3pAKk5E0kSKUofB8Du/EreBYDcKZMoHSjggTEQBXuFC4scKsD4P58B0xLl6Rr5
LQ9Ux/0DjXVvZjw76FkIb72EmOm3f9N1X5EoaxBoXJ11Gp3JZQSibIBtLG2lYZ6x
6AAn1kkXd3WA5PChuC88/srXVODccIHPhFNYK+HxDmSeO+4U/Sady35wsNsZktpW
aIKODuXIeVfecushT4YLDU8dosMR22d7HappSBCi1YTzg8BH8cK5QJkH64sI7IEd
VDaTP4nxbJGEgxZIrmogDfOK1BgQtY6sz8vL4ORvUa4WO53y7m4pYSy6dg4TOQ63
dpazJ02azuAd+ekZRfc+r9VYBzJCiLad8c4upCBaiubo4fhFaBqw5VS67U0NYzg/
KjVokG5pcNey8eZ1pJ8EXh9FZvBAo7xc1WATdpGnf0Tdv0wwDTQtal02jfQs1WfE
uxc7AGf8ywbMXVO9Je/LEOiRbKGlQrqk9+vdIry7Nb0omSS1ABsT4KxBL75v9h/0
lWVNCAwNKBjohbdbaacTfeaP0gCxJaRi9yGH8NSzKqqhDW4CAMONm6y+nBmJR5L0
L6aiBeUtYt8+TmazB3vPV3gKV/BJX8Z9jwEt082wy8Oce7+6Wej0t+05e7V/6dMZ
4DggV+RInv21TdTs66OxbwUy1OE/VVDXW1JhXSuhjvHD2RRsiOTY9tNCzjfOfhcW
FbHSN4aJDm14sQPzPN04DeQ5a5nTG+6hddD7nIT3a2crhSH7tvbAdmpZBkWRg1Cp
1ip2WJtrZJoeOwba3H7oNwrNdiYoHNx0RzDltBXvHvZz8wiveWxCxUjJVu3bh6ws
L9PNqQsSwYYIX6D2a88LlrifOKX7aLq6UdbIGW41qqP6p9OpLFrr0D6Xkxh7TE4N
NL+lp2nXHk3T4KoSK/DjmpdFA1Ihxo3gymyI1+okwmW9F4Bv8z9dokjJux6zDzgT
PDawfllvRUwL5hf2bFCl+QpkmztPAUAzHecvK2pMg8kErraiXphhPnc6l/+3Ryf8
2CG6bRaFJHKKoQwob5+rtzhoGBsDqPVOXe0ZMy9eZFo6XkPQw+f8WCV547V+W8ft
E1OeZQV9gZcXdMYl7O5028Wx4adL7qhv/vIRm9a2gGY0CJTXXhY6P1NSqnqGX23U
ofU2n9d2/ECPGziR2Jv+aQr21lUBd+SHuxLnPJB2rgPSaUS5z0NmooP7AdAI9Yzc
p5N9lEuFLh8Ua5DZeDq7x7Af0XaUn2wOh65wa3PQpTl20J+PfSGurCJJOwcAZmwa
KFGTRpSVJy9nsVZLiWimtfVe2F9polXju/JLDdDdqsRNWZ01xWm9JHyYUR1tM5jB
hmIoWyiHUxhKqOisyM4JuzM13HZ+yTQ9pVnOYsJOjZGdmscaUCEanwveT4H1RNhe
eVppB40hN8QxT+wN3Pd/n7qoXRcWfFi71rbZ0UB0l5iuIqRrfRZXsbsDYWkIzGtl
oarqPxrlA0wCn2y1sMhmALGnxqSm3DFu1GrB5TfhXqdrHNnGmU2gPrNYJ0WdBHtA
5LWInOMCr/lbA3IeajNsUt7CHEt3MVA+NhGo7gsBucIbwPxTtP8fiz4XWrVzPdmR
zHOYoPJP7tZSQjFxXbFVAzJFP6ykrmQmZXOfrEccQ5gnxtZBvhSx4zvK52V0Zm8T
Tt16Yjl2CTos1rSqSSYRa9vThgZ8EdgOT5QN7g9wtlVGk1K1kB3dtGK9H7AHBtkQ
XOhAa+fJoPnNIIXI/auZM5Jon68QSgmDH5mkT1f7sTXb5CHlAy1RJmbj8yqX//5o
VKHPNSiQeqDowBp4kGb2uz1gIXRKHSqQxmEfkfMAgGY47BWr7N0n78pW4j/ECpK2
Hz+ur66RBB92XDNe4nz2oXNXQ1Z694kb86rdRbpKTPzyS4J1przTayjOn0ulZWgE
o57dNM7sEYZ7e/AdarFR2GzFa9w1EKLqjtgHs/AieQHZXLtUjOY76hD6iCIeewm7
k8Zh4vPMa71KGd0IFrqxS4GCqrc89Edqv07JcsrBtrSugHWZ09Q7iMeaKAgG6hzC
mMkvvSrWadUSgDOpmZubS7jpbTmzxcd3M9zHz1zmLOtZD1wIE+wmSX6jCe3JE3qM
r4TWlookNomu11WIE/7SxaYklNZlBa4tz2uTytFleE616MJFD3Zamq7axGnGTF0U
H8WFuWyseY/1WLMJnjZOCV9iplFJ9gBHpnAYyiNaC4ob4CWGLto5FYEQ4BfUpeI9
91Yq+KYG3SFUp+ibyFT4mJN/XMBJRoAiA3Fv7jnNhUbfL3rvUVjH1G80B9cH3SjS
L9EZ9SGetPMYkY7p6Kt9hjGGRnU2Ziz9aCOvn6/D2cjycf6f0K7o1sYNrpKazD5u
sj9mQqHYwhn5WlZb/J5lOA5Ay3jz3ianyBAWkPgKpc6Wcg5ZNXhmIATt70gOF84T
Yn87V4DgoBtJK6yr/Y6+TseXmy9WMKPO/J2EUzKuEpqokL717KHi3Z7fEbDmrfOX
7mDBn+wudQiGh41zsV7Ncc2GiIya+hingQr5ZcVBK3uLRn0ApIUnxXHtZ4FCjcIk
1QM9KLAW5mJzE24xIRc+szwgBydwknFfJK6Wu8h4PdwBUphL+9Uek+gEOgjs482T
nTM8/ga/UqJe/CJV8RdOP7tkvBrbRfo59ETNAPzcZuDZsyVZYTNnYfA9oOjjgSSm
YO+lM4V7xctYPRZNtg9gY+/2KncXOtxMWr8LYIaKgBVOcAU/EiInyvNG1PJCt4QS
lJFs0Nc4En5Y9jsVfzje3DPRuLOTFcrFaIeur7VgameYzaDbugvXV2JvjCsD8deL
DKd26e1++wbX6Iv8lylP2tjmAmq1mcdUrlWXE2mpzzkEX7Syy8g1fBONC3Bk9U1E
KVgoYPV93md4MLN3Ku9ut9OU/Qc5OlyQRMGuDORzNAeLAZNbr8L9mvmwS57gNLPK
FSLHuDLX+8izkZrSmCmfD4g34M4eGftJjSv0s+KS82mk1B6A83OGS5cR1kO7x/ka
H8nGWhcFZMtG5Z3zEEF6mliwHTeBo1dpLV326baPHyyvOXyrDVigRYkEUZWa8bgT
08QQ2KCPRM8jr1r1BAY6iwFGZwRaPYKQx6cQIfdrCDkD1VQ+9vm8v0GMzPJczK3I
DAXmyg2PHjF6/be9kMFrEpryuPArBeviPtjk8H5GMHOotaO2OHF2zEq+Hw5hvXfm
RDWDbw/bU8DdOpaniFy6a5ZKZC9G3cBoyVJ4TidQ3rKNOlJNm4eQaQ9pMQgEAeJ4
J+GpAztOu751hIuW9zw+K2Pi9e6Et99RzD1ELnElgkw+lE1TVUJcPSMmRDyUCzac
s6PXs1eMoOZAEnF8npm8xQEJbWhRb1x8haawneQhucd+3nu90iAc89sVmAyp6lih
I5Yr6WqJcxttYduAizNjnrAhbkE0CumV3APzj9MuhC7ssPKr5VMfZbvK8Kt+Rzf6
VAjU9Lc2GqW/1HTgi4byAPkfrX8iwVH/TlTiE0t3tUiZKK3QDX+BHoAX5NJlcOCP
nGMOTzmWo1R2TXME1ZLjt3LtLvt2MLd5WnJY4mmYmQfdFUSOG2gDo9UrTnQEJqQl
lGyNM1Ju/Lpq+CTb+3h33prbxVbZVb1w/XuayLlDlYWKOASb+ILTS8Czt7OqBPUX
yrkmvMikqT+QOC6Z8gJYGcIB1ts8MXdqVAZISMa0SlRDi3RFY2z1ZsmxdZ8sbGos
All/3gL2xFkOVIq70hwjiDaSc8aeO8F2rDhJDQWk3+1KAy39vGSsojC97c3hAHnO
pR0oAz2I2gpWezChyyre3MlAw69dyOOUAz2tk8F1gAokR9wBepsnseyhi+rF1E86
XQ7IbJFMSxb5ShIgWbdBxINzu9euiL3DLSSKceIw0MbgXihmULAnKHpv5zyebXp9
7pj/eDIvSmu/2zMgZ+BLV3AqDGtskAQlLgag8mdPt2vj2exrvOpyCUQG5ytFeopQ
LlcfIqehcGg2exFJF+YuWzEuDrL6J5e7XixmpWx/q5aM2WkL37EqJaLFMvlLm+N2
uyW0tJDE7D+FWDlzhORlMUpT0wu+3Dnwz0fGbClaG3RFViXpw7DC5DclQ8edVlDn
RnnUvXNkRQtCvXqMebAzCJIa1BC8pAsR8pG9SN9levWW7Yq/TJrcvISSs+XfYmVG
thbtJ1yvCzJbac1qRPEHW4rT5A2Uj0KvpFlxbk2CLNiheoYc4uHVAg64ARJympD5
cEgxGxUKidIk2B6npLIyvWjeLAeEpKbip+27ieYoHbZcvIRWU2CyYzllWFR2Jrdz
9QppSyvwaqyGMO9oPSRZ5T5Enkd/65uVOyCpDWSUw35JoI4Vg9m/P8LdRoOzOqJN
xzrwTj4P/VeoIS61OUwEolz1cCqp/f3SRATOBfosB0w/FWGXWot/sEfpCiOXFfgV
/yC0rKEL1jCChhWx2Y1AIWVB0dnpKeEErAJ9ukn8hdx5vStIkzgYQJ2DfJMsidoa
9vfF0ePIv7G66B5rcpJ+XH05PQJnx5e/DrcSZzV/3eGFRamysNOZyk1ghnauK3HW
h7/GKizKgPMg2L8tm7hIca2Uz9TSHb3PeQP5DSAEkIRPG5EuWPSyTGEIA+RxrtN2
VoK5SP51PNGjrQkmN3A1GgSSW4kvNqD3Dafl/kWsEPWV9vFdEN6bBgQuxf2PJLdc
K4HGp/xmyrDudIWU55EeOo30oIYkBHbG+yLDKmPRfXgei1skeWVM0rtuV18uo5iT
gkoQewX8i+wG83g62tTOwuw1kO8NL9GOVCUhtqsrtBESX96+QpG6m756kcPgopA5
VFCyRy8MCmx9MDHwacPjz0rLrwJDl6vasCAFmXeuquYo8+xlPidX+colSyhPyp4P
4keJLao2Sts9QQwG3XImhDFHHW3je40+SWYU7LvZAxGJvfgsyJcOTP1xxYNByQSp
MclyXgUp2gka04KzYi4X6jJSb600kPWtI2gTE4NbtGn7zC+E2pRfwhmnfVlE8cFH
yzd1j79XTQxctHOUCghjWtutvIVTSJMqM2s5SGc8A4vI196WApItrkxdDGhaKzRW
b2A/TsS27FwHucKqInGr4j6jsWbl24+bpn3GpUd/izfkxUg1cvMX8j78F/3oRt6p
Nks/7R7Uai9a07URZQo+BVfPLqVSj1jpuEXNDL+rfRvMLWs0KWVUQnKVCmhu0/4g
DdmQF9c8bAshHivl20tL344Rxxx5Ip54bqK7a8fvJpGR4wnNAyi6v8brMvSrWYRb
tovQcT4nsuLMyPlQPxGJZooxZq3GxpqNudid7ESGyBFAjolvAGtX4TfaU8H7DO2a
cxbdKon5WTmLeXzqBrFB8RypEozatNowGMJIhFbkxsU21zoANRG0gOcgx1Cnr7hm
UHQqB9ZyTec1vkFdvsF/vpR5YPhpJru+eHF2e3oGglo=
`protect END_PROTECTED