-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
YKgH8gdkiA50qRRjJl1fULTt2XdIDAUydl4LbzTZuHhpwmcdBP7DHFmTtDlQkprx
mxg/ivz4wFNR/XybLgkvwDaltZVi/VhX/L9j7V7ydRfIGSgkO37aYv5MCpyibziJ
j3kI62bibadlFhO+myR5upeFEEfEkhN9IYT9SKZPHVY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 49360)

`protect DATA_BLOCK
Fs7e0oTcY4qYhbe2dqm4utvo+Q5DMASr4JKcxonT0OoZIJJdxd2mnjkQbttwYFEY
awCqOJPWNW78DAqyo7mLMh/holFXcDdQklycuXyV+D8F9l+8V7FenZL1/yJ5Frjr
DsssK5fKZrsfaqH5JClC7PGD+qACWCoqUKsc2ED+BNl1AstDQx5ZzlNYJPfTBTP1
INrEVBBmyj5SfZDwWDXVgLGJkdDsKm0mBd4SLqlYCozwjJu2fN8yZckep8jPqnj8
8LmQl4skQY4h/fDayjaHVZWNc6Ze5ofI267YC9e4Ai9JvFhT4djNBQZHJGuEJ0j6
m/sDrx59t1hYhWocAJkLDcEV49q90wEgtWegj/4d4ILXsmcNiP+nT6+nYzNNt7OT
UububdsdVdNxuDvyyAP8N8bLYEmZxm6xDlzD/Ln8XeKu5TNP/IlcJlmRnIgjvLWX
7UAAQiFau3H2n7rt5Pw8d+t24BFZt7UnWw1vIGtusouAfq80ki+OoMvnoqMGUWSb
mSaCQGxx4rcO5ZXaBBnU8s0+OvTtWMSyzRT5cm/7Rwgn6IqC/3NcGrSJRTL0EMeN
TxRSEBAaaEjhwzhGo67hYmYZXANTT3ePJQnnviTjkC+VrKGls0nCuDSeaV3v7+pB
6axTCRjmix6uAZ825D8WYDvBLO+/BfE4UUGLngVTii6AsO9kbIRfopNfgRFrgkFH
jpWZa+5tTjHCDFXquxkhmCFQPEeZIczcTwZUFJYhVRcJsoBiV432enRVhEJ0AfBd
QPfINvXWAegD+qVwBiwl2fGdEtmDSaK4lnSWWUmuB1ncbCGjcFlBNAPk5nRb1zdu
ZbwUS18zplCWYdonyNmNPwTjRuE7KW781D/a6eXseMn0mZKgb8vEEVLuFEkDlzce
P5+GCHEaJuodmP31F74V2msAxp7oPrHQMG7Z3lIwRvPCtlm9fDSmg/uq+5y8gB6s
tzTN+m9C5wSKBZv248xpFpHqgh31kNL2jsgv+3opEmUB5k64gCKrLRMYjXF4hprV
esbVe1v74+1L40g00N+y6NSgACk7jnwZiQ7fZGOVmH/2yngeIsO02FcmSjVphuUr
B8WyBkMr5/gitA+ENi7dvyYdVHXoM+6PrjAuHzxpHFfmqLsCvmbxxScv4+w679Mr
DKEBUb7RJL3TRwgpKTTyWXVaHtl2sk6Qp+chcV7BoSp+FjfrwyYR30IXUjipg9K6
RZR1/kOJLqXkki8r7GDUdGFT1XAS9bzi+oa6pEbujuuEhvV4kSHmcDN9mlkbYbrw
V4/KYb0vDavA0qqNyL88CBfebGhYbuUdDNFzsj0EiRf58HV3cvz0EL/xXC3Wltg3
2X4j7F1ikkbiVeu/IHh/JwciKOBIhyD4FnA2m5kuYIrMTtEeLOj2m2tYmMLFEpf2
GeYcIPLFPay35u8GwJkUQo0qZPTm/Wukk22+iR1/aCzeIPnkbaDxVDcUtJWgNW2X
mvsL3+aIDU7C12v77bZq6wokZEQH/Tk0/ZeJJKgzh6lu5bD4UD2MGcIH/yocfaHK
sGsZpJI8AdM750Sph0TO2GIIKZENU6zqCWMNBv+5t1bkfKdMImGZiuq6Jh5igNwQ
G4WOuHrCMukqWhaptr3HI/c+3BDyxz9cmaZI3aZf9m7QXfZvL8he+0JlkBAL5InQ
mzeObsCMceRejPg5ukhmaL6qu8ozYhR3qj45/uy8kBNtgXRXdo/7gymQ/E/RI0w6
Uyocnyy9vnf5N6H/zl4D8b6GP2NA+D7ddSfRRP1ghkmccRBhVz5gBvJRKYhREukw
MnW5oPp8JT222iheJRXrb2osese9Q1sDT+FLXX/IuadLAuO7Dz4niAEXXCIU7M1Y
t9aIwfx0U/8fIZncq3xuejgXuRgEvHP8o4RLfy761z/0nm0PYf5vLYCbENalHjQ2
nrvZG2tcnmu2bTs4XhOkJ10PGfhyoMKV5xXv+uM1pyiWhElZkKboP/nb2x0MH017
9NhLGJl44RqUana7ojpLx0OUJAsQOAl5rb8UebQo2fGMfQJWzJjjL8U5wrMFfGDT
Vc9iYNQE5mZfXf7K9EcJfVTeC4E5JnFeIOOPfDpgHyaKxteGv51j0MLUTKtV6/5s
Q68M4ALywc8H7GF0Z+sF0SdzNbpF5vqsMr8TRYK4ZmjGJAUGretIabgZ1Bl5dZ1q
TZJAgx191kSZiXR34iuVhUbCfw03mwRVxVatwFG68qtUaKv63gKNCHafXnN5RjxK
hfVs0rzeYcwbb0gD9W3DoZLIGfY9vjjUKaHbeHRJtad0vgxpJWKRjfvriF0om3Fq
uer5/Ke3Zr+uZPjZwI6/ufJiWEeJ18u0Uhiutc2GN1mCKG9fG2oU8ZIVG5IvSqbL
7Ak5Aqy4xQxoCxOf+M/RvKXIrKvyl1ZIEceuDILyRP7Cj2TwS1glM/ZFVSb8imsA
2n7Ix2+YMooPXw4plyZ3MAn/p+xZq4zC11BsmMf1i45S0DQiKU2SRfAbCZ7MRvGw
Vepjrph6T4AqfrQ4HnNRxrSIe2fvtAyp6cfeRR4UhBbzGn6LffSActot4Ht0lNQ7
d3RVFPJ/OXRShVKpn/loOfipYhqPRQUg3s1/qZHbpQqHOWrQ02fGdG3BDmTsHeBG
+jTO1wN99czPNe8B9eRRGjqpUqZE5TSCg3l4z6O1iRKcX6JBGrGNF+Gcq56qz7up
voQW3Q8nwUf1pcv6ppNjdb+XhCYfolZHxI0ZHheNEYxbpasp8DFdmXcX0YUj3jdi
MuugvYDMsXKwSdB/CgXKkJkSNOw9tzJmkWq5yQx87fCzw4R2e7AuqB+/eyvvuF4r
fQR5ThoV3FNZaAuF0Cblde5gOuh91Uk5GVHXpy1xul9wm3xYsEOmQ/BeyrWWQ6KU
H4rxMi3fTBBmcP8AsGEG+iBuMzGXmPB3AWV8E0ePbiEwGyw0HNEXgWxM1mdSWasY
O1xfUCmthL/29pQk+0mDBs3si+yVVW2Pf8IofRoPTfhAc6+YVrMR8a5sXCd+DUgL
fcARYk+innhgKtb3Lm6yU8S/tILiXfWGFuUz58ste3m64v7tCKROl8DRhglodj1i
ZKU8NEKuKi7Wa2mouWfQ3vLhiVqqTB8p4GygjMqiFn0ouMHrFdP4NIl1lRwmLrLs
eNaSV0yJg4R7phHEBYX9fpNb2Zw47OKqV5WJohQDof1LvzdDpfhQF0C+GNXmMsoo
4aDrwpVmeMhRSx7QviAy4bgY5CqNLGfsDC11x7dhlOc06RNd60myPRFrXz5XM8uL
cijR+7qZd/1P5aW6YjwDXrsAOhupYIa/8TOA10PGb7lTSLc0qBxYOE0p+EAja+rl
waI417Xn3MS5klUPf3VO3/QDBOGbNv2z8UJq0q1Obik8+lrPxfzAfysevLapLIpZ
HpwG7WfnxJjuwsiSlWudHK2BiWLIZ8Eg8IPXqFHqkZCn5o9xtpTiEmdbSt4gquOU
bmTdIfaI1OTJUpfg5FMm8gyPu7wExlP/gPFxNTycQo1dvPp4OPjIfHQ/iKE0Yjx4
thbeZyAM1k0rtAbUbGmfcgaGRWigef3EJy9FD79dB2HQ/MPRDob7NEP8YjHe/qBM
7GNa/0v+GtgF4yV0WnmlSMSro7dR60lRxp93U4S/VEVsSACllfK8hiQKfvzXOCKi
+v2aMm30SnloXTaun4gIVZrDt3fhci72Cua5Hxjunyx5ymj5Rv5ZD7PlcLGOhsUR
dg3Injh4kMID3NOxkQvJgeYojCILsO6ULlDDK9ubGKoWBOCf0U1Sfo3IdHqB5JrJ
HA9O2quHzLQjk+/QIEAn+2UZHEWugqA3sS9Mh6rFLsvRdfHUkHVT6wvxTm2nE6KD
2ArwWZhjPsdzb06XNB8GtY4tYGN224PD1PDkXV5JjZBl9bHsv0ZUjDt6kTtto41f
OCchMGfDMmlKjGvSdOxP3MBduZDt2NAiBAQ7xunVkvtGtZbsObIWlaqu3tavML3j
CeXzSe1u8zj9i+7EbzeTEECtkp6k5ksVy9gKLBZCkGXFTcmmkcRYy2Qb3f5WrZX3
fLLtO3Qv5WPhG7R5i+3NdS1vtfsRxSjZL/GMOaOrFIF7EqZC5lw9Sw02jFWuByPw
mKvfQwnNRRhEDHBxLI+B4hDToXrbiMCMwnpyc4F4P/fCfz03rWya6o4EceS7JKi+
wo0zpTwscJegq5iN+sQw5NCodK+QAglUayPUGljeoAboFmk9Fd+ZUltlrQ6CtDYT
upB6yOP7ULqCDbd8+0yhONTI/fZpEt4YAkLgf+SGHfvr7yjyl/myDSt8aca28bjJ
IS8FxyC5yf2HODzHXJhDyJ0gao+Zr/iaZfMqwA6qazrSd412TDNK37pyRL+pRFlQ
JIgAbzU0OFNph8KVKhVHxndfX4ZGEMD1XB779RPdVL04bcpBo3YxUWUsmEG6y9Y3
c3M0chboik/i39+v2Mx6Lxkjx4/TSTvdEH6+04neBHzl61QyDaCn9wfYehlzChGs
euM6Ah/3iO5FJ2+37re7agYowpJW7pUs7J2r+qFYJCx9dwX6gKJepZx92qa0tp8n
W4yRByBMbPElmg3Ow+5KcqDNRvFYDWS1a7mnRO0y6rE0EThcNkSVt/Od4CHsfLJE
ogq4b3XT+iPIljj5v9lIute8CBuKj1R8lJg5rf7J2Qosf2bYo+domRpEsvFhSs3I
EIlghnMgJm9pM86pJOBVzub+xJg9B8nZ9vmXjAOyNdok2OfMB7wzAT4zJRXyefr6
7/uP+CTq4+tqQyDEbjPZImhtX71rhia9SksWrc53Z4ne+LgoC1m6N+TxBrNnejOD
p+4T/nNBCLO4ovI+mvqc+BFiJeVSZRsF+95vEXkFmttMAJKrOdn8E0lbkOJ+fEXC
MuaHdTUx2MJorGFyWwx2KnyNrdvzs72W6YfJRc8rLexmFKsng8ROC8cT9VYKOcE5
VQ2AQ5TMnpPwL5cX8y8u/9jU9b0IfIZ3O42z9H6aWlwDaVacVU0Ou8em5mMop7Dz
hrKgeclsqSDeC76RZK2ADsm/R0sDPoCfbUKGJBxoN0oiwklSCAR80VpRIwUi4xWr
3wBaN6ryZ1z20QLnkZk0xIrT2bpKq+l6m0Yr/j5EFOuaEg1xc32cS9YYocw1WOkZ
bPZI4nCQyHkv2kCz4l3B0wdwMsSLRjLTeWyE9K+673hAysTIQ/KY1MU7zH2PuATo
67OagRT8Whi7LBZJl/22G5W+jJu4vGmPSeveDgInwlRyya2qSggnrHc8/TUsNlz/
9CKwgX71szMLlScV+RO6lJOB+vbTeGPpT+v2pU5k1xJ/EF+7sp0AgxSkuFHgCjq/
vLXFuvdC/ynRi2C+c7RNFS/xqs86OmM9lisu58OVrMo0iliizWkqMukf0PUqXy6s
hFdsRjAUJtf9QxU9w3gtepbUu9QmvhswGHV5zBlhz2eOFZ/mQAuwtAI0EwdNQs4g
0oZ7sdvWQPwMw/SQti/CYqmG5NXJGO+JXUwI6selGyV8qDc8wVaPPu0TVkOc/V0h
SodwGkEUnJhry17pIFm/V962JE8VMI8XQxIvg0Inz1iroqJXAae/Pxo6cj4xmJoE
z3XrPDKk3TB4ty9QECNBf8jaGJR99fvNigJRBZTHunyHUcSbVMjMK2ivAxiet2xO
xVzdES6iXJymyRxMElRL/mP50NHlCUMCq91ryIqZk9p+CcF0IqrpyudbRHU+kmhN
QVeCbAUUKq/NOyx5Ap9UlS4MpAWRXLb82F0n7Ds0FCQeeiKRFtV/F5pvuWeKJV5r
4V8TkEJtr0DY3O+Y+RxEcHVBFQ+Tkmvi5MImVdpX/DTteVmunhgmSkK2VblUVT2h
ITwSMps5aniLtNbjhGa1tawgKtULiheRGwVoe6kS7iqs9+9jx3+al+taONa/lsZW
ethn+J5dJ+nfqLR/JhuuFb9U/UKodb4wU9QvMuUw149PgkSzZyGZkHaT9usKiJVD
Ee8Dh6JjL7JwBfIaoepmJLjNkovbin6n6B34B7T9cJ0ZqXL25Jmzz2htXYbXrfhg
OF25KsFPjZrKTVCZiOpf1m4LwLRnaTpXlnVzxtVCt0kYgNI9f5iI4yNmYpfJ8yys
qvgAlChAToG+momeUmQs3L74iE08O5kFLCbWv/4vfuKZ8R2gycjv2MUBFf10ezlF
aTgLz/rPrPYTKyb9ryJiPXVN8lXcsGEmY2+GDeeyKdV0kdoZP4roExQrr3C9b8bN
bCjN3jLEa0Qz6NtvauBX7gFTx65vYbD+x9V9zt7nEgcIQKnMRmW39GQ87wEDhQDo
Wj3p0J2KbAbLHV1zZpaG1SRWHRXuDdh50UTuJfxUb8NM2XCoMbarwBAqtar1n4NW
C+Nm9sxa/4+ps4eeu3kDjpWatmbh+2yr+dgQrW1bZ6ih92H7SHGhre/UDdXmre59
7B6ZYLb2rSkJAySpH8F6FGY9i9K0KQUr12HbLwkhrd8sXbrM3O/zm2zTlM+mU86O
djF52xPKG+d4OYKkrvSoSEfgwmxTX5+FAT4NYs1z3pdL2WNhwK2VEreu49MbHfz4
/PbHuS+diXxCX9jVOHacV6X9rCnRU7T4y1d4Y4aCnv33P+mVa9QFESdpSKw9gqRW
wzPk6Q2Gdct624kEw0QsXKjC+R3Pg29HnfehhTRE5RGK2QI/PPfG+A3dCV6dmrw7
xh4X/yXRwIYetuA3p+pDiSNHBUt/8xq63zuw9IvuYvfgzUlLRhPERyBWTP+4taQ0
Nyn4KpYBjHMSjebWA23Ipo8gWP0LphDUgIEYQQXfJwnl2i42B1+E1GD+9f7xLiaF
qdPnkpzvkLKVdNJ42pahwKS1S/18dwAwX8SMIgOyUce3fDNDN65VWElW6tJdINuP
TieNOad+a6UUnUaS9ovwfRCagFk3xxyiMoLAtJB96t0mto3k6XClKy53LdXSOjZm
OsU3K1vt5bZFin1AfQALXBqa/+kWDvXjFzKD0XsoIN+KeDtg5vWF3b9qK6EIv5AK
B78UPJNxuBxbIpX2fvx0XcOFlxscr+4SiZNmgDW6IVzAcEn+M4ljonlK7gn2MJgI
6pfBFM2utjnilj1oN4hVYnH/zrJmS8ijli3DU5I2wKKiULl7+eOwLA3XuNlgSIzO
x0WvSxBV5KsbPFmmWszlaIHgc7YlaHPjwZbIUeuOVsEjewVmdqu4Ydn/FgdAQYoJ
H7pODptvqpmyfFNLKvxLc5CWGDrnU92ZBULtaJruPfuNDz89jtlsP76r/F6silhG
RteiVOaaUs/J8PRbMOUZLK9WWkU3C0u62P2bYjXoYSaYFa7D9d8sIAG4RZxvcCpQ
/tZlmaI8SwJESZVAnkbcBNMG5ximRGJ00vEHGDAbZIeR9Dyq+2D+V8nTcaHoSa99
rilUWCROuOD0knGL+t0vnq9Nf1f6djxBzw8Joi4JZcfFgOGZ8aqs2X/T8SrDP7hu
0mZxmBTKfE7bnHfwltk4px79aSVtXcHCPJBMgJqRm4AoNssYQcdAztyre7JHcr/B
P35emynSnwjamZ+DNvZjaICiRn+35TGq3DAUVo/VCt/443bZj6rmS5LWbEYhSDFD
5ph8hM6VxQIjNStp+nr+/vP0DorZHsQix+pg/v3wEKyU+xvBKm0i5Jd+Ychp5b5Z
Zo5V8zR0CqZGpUX9z2n7o/GlRhDnK3wz6cB2gr2bvMxep+k8+x85KvlEX/12zISW
2Pkp7mM6NpFKIiYpnFMmgtmIAv6NY71rsXmzbkaHrmG0O3VRHon+pQ3FCBHdC5oe
fVebsrXYVZcYfijmRSB9aep5FAKiibYBAW6FbpXjegAKOIZ5Aj9laYyH68EYQM2t
x5IEOUrsnXfUyMln/LHiWgMktLvrqjGCrTuMoT87aB+7kY9GUkW3TacvF6l5k3CN
Wl2SZE/VqgAANALzZ1SznxyYiShm+4vJ+cN54i7F+0QNwtrt31uDw491BkyxoOUe
WWbwO2fR2CCD8Z9fI5VBHXCCccKGhSAE1irNfOQShEHMIBGnbC5AnD/QErfOShCN
m/P2FVvTOvwDsI35fMwcdwBMccWZJnOcmI26dsxoIiwBfpgn4g2AvMP+/8fOiEgk
c5+/2J5KW9RtAMa14Q9Ize5koBbK/0VmvtCqYDgkkw68oNstpewBM4PY7mLKxlA3
T63eQRWQcJ7kLXKwaMtFkmUbqEUh5yYjRcHkhcZruA2oqUSso8TRArA5OHsCVm+i
Zsf/lYAnSRTjfEX2donKePUgoZDAmNOLSM+SKDy5rCj3cvf2nlwgyGS9s7ce2OLg
vefydXOfaJd23mi4EcKtnyg4P7wJg4nAxFZ/wWfjL3fF9KOw3dFSeK1c4P87Rdm3
rUuvxzuBpIpQTzxhvUTSekCdD6PH6hus4v6fwbomIs/uy1do56Dkr9VV0gES141S
F8ceTAbpErsbMA/SzquKWna0KsgTYTGObdRYjcCDe3kSasHxsHhzJNmLidaVdQAA
gTGviAw7I5BT6Cw6JKQKTmufUyRkQSDh1lcVAK0O754tPwkxEoxeJuwgVTqrpBi/
s9wRPY5ELuGV+lIzVW8HHnd3go3mcvfO7wM3COejBtViHJp4DkJdkDz9RSqbmKsW
156A4f2ZNE+WSVtQp/YqwuugaQ3aVW+6fJnLzSL0pYdmknSKTwNtSxmY4sAZj89G
yB+boAU6/KdYZKBuaoP/f8PWj2WF5BKfELGdLLcG1hitx78N5IObhhyNTbDK3iis
coWLyQrU52Zf8iGN92nGTCz9ZXA7yt3u7h75JqtFKjF7CW4z2RWrKHuPLIqDpU6c
j7EqcL8tEFDUTH86Jn2FwyhaWx4G4782CvFMeqJzPWhGga4eGw4Y67JDwgCdLBVN
VjwWAw+IU3F7CNOhkt0Pd3VS5pOaHjFP2OER4LUeuUmEiEDjZsc5QcVAnOd1OuOV
n+UhAgDanV/nKhxOBMf36CA3xQIhbmVsw/77NkBZcOjqRbnSlU7pFB/eVb8biRv5
4sDaZkKBrk7KKHkk/GBUm2ID/qIxqGizUzWgoyBg4p3wjPSnbc4Hc6P5NyhGV8Ry
Q4y8itC85fU3WWJ0wQjbiIbqWreuOO/DuDf4nTYnQJNw1weVJ2mj4581tK4wH8wx
E98B8/2D1TSkH6s6M0Co3MIfD4R+yN69DKUrlNv+LETX0bemKFd5pMlffsQJa6Qe
oewvDdPnmpLM5wc2d/MLGNKgSOc5UvMyzFC5wEo9IheTvoCoVKMzTpCpAuT0P0mt
77Oob1md9XVRB/nlRW8+CPltadezcWpEMy06UGD8w1vE6g5DyKacCmJwFtBkF0Du
KXj6wcpWlV9GQO1YrupGoDsOl3sVzyucvdu2HQXGvlYD9EijXaecBk8fphn6RvXP
6fJesqkks3MzvR910LbsP+kWj1x9S9RjE3KU2nf/oS5j53doaWHQAGXo4ncUnI0Y
7V+fYdmbLT+jjXgEbbWf+geWZWhXbEPJoMLCSIN6128aYB21CjLmdfk2tdU6AeQh
ckSt9ZswZ5JaumM6Wjgvu8HR/bDIuhn6tqHMoaZDFXL3qDZF4JNfsLFizAYiyZlc
+P93Td6aM+iGNpEQcfKV3QHUF8HLPHXlHUQwfa+9u7zYaNrMgwRl28YpEJHxiLyt
CwhcLokE2IEVbdodoy+bV1lJ0QXAuvmMQbC8EnmzSVi8w2LhifoDjfblBuQYii2K
t3gAutumQ8eMamMnrtPQ5xbjDBRVEZqEbKUPeP6B8zrCAZPL4wQuRvO5uBmUXD52
g/cOTIrhbKTfrsHIQ5thquP1BkcSViM6k8dXrIuoTrOMRXOh542OZ6vrPVrBWKD2
+iYzTT0fPrmKrkVCulz81CIJm1qjVtMX+vEYk0AQbYmAFWzyDejgqsSMT/cZ1RIr
WPmUksvxiu1BHCcI9DPMznQSCJm2oSpOsjkhqiCHoVoS6ZizMZP0wJ5fs6pSqEhS
5koqoFMYrilUcgweAcSt3l2n8RRW4W9FfcTSJ/aLrvYKtTI9BWGHyIJ4SHGXfUxR
kiexHSIVkPIYmectmr7/9K/AYlviRStHWL/Vex2QTPkvIuX79V2kB+pEcOWLVR/3
3jEwciOJxiToNipXi/mVfB/T1T/GDiXHOy31kuhJJarvzHYJqTyBG2jDpNiH1GsQ
IvaOF5HL/rwDQYfBOsg6VbrvP77bxwgeAnr01pdl7/Da+eU+pQLHXKIiXRyiRydk
qHspUxqIWy0WdOUyHdwcVf+qTISTHtEqR5G8x78zJUMOd3uyOErJ5sZyJIAb1AWJ
8CAIuZZJwM9xD3rFJQ3GoYpQlLA9Hm/yytQi0Ovdjc7+633utAB/mULEHF1Pqmht
r+RhlgiElG6JmLUcPno8VcDxwjXLhsyK9hsnD+iahk0/MuUVdmC3xqHtFyIw29b+
y4HZZK1VjDvHZ3PX2LNcLf7XA2kSKAN7Obl8kQ1HhEby9A0/xsigKGjrwXwSvn5h
8oTfrrAPm1zn5OvTmIlBTflS6UnaOlXEa/LS3sBlZ0Sa9GOVkzhVPiDe4YKOVqq7
1DWHD0L83fC+/po8ig82/lM1+FIQNxZ19RO0Xy1iupcbB19gYRPQegv/WF//j66K
zsiCrs0FkckEfZsockKyugIItKJew7Nt5vc9M+NpDK15kBqhmcM+0n7wU6pxYQt5
M3nZA5dAckt4clPjgh6APPSLgMTtbqgv8pBEJRRIJezCeF5ZrTMKOSN8p3my+zpL
rclMW8IE8X5fuJygYnHGjIrCi53emhuwqEIeLBEfMr700kDVa4oY2U/81FR82+5+
Fl9zV8BrCNakQIZJBq7qO4fTDvr/9HNnVzYlzA/isGzqOWC/jAXJAoJfuyixoKMF
SJEQFdO62Ij6xAYDwDMAqiLaXMk1DLL55PUZX5Zj/cSeCSAczM9XYL6SPfu+Dn7K
BKHc16KmBn7WEOAXKu1ycPzc1RSTLhaVYu27Gs36yOMqgYtznsTT6lopulQ26Kwe
I79WtOBYIdPbZXrFy84tF6FNc234oWHYNjljCyhzBu7wgrF43RU5F0zvg+KEaDpJ
dlerBLTJGTiDaN/uItM9urt7gQqpAwuu2GL/2iquyiVbsD2P8NypffRHgPmvdkYw
2OQFtm5CXJii/FiCeJMuPad9CyYWHpfcf3hBPYhu/1KeBVicmC0BSXj6e7v7QZoy
CLIFRpBMmEPlBDSMV4jO0mCiWbXXsWASr6BU0Rq0xZfaSOxeqew4uJTmT9x9BtH4
1fSoWGvmOnVjvb+MaSXkDLQ+blv6IqMeZ4ZM6wj5OKe1m3m29IqWFNSyDnym8+XJ
u3wfygV4jFrOt8UCwqSj/Sl+rtg861G+ytql5ESnx13RE5bxikoRY3njlwrHyvfd
l+Yf3o4oj/E3oncG37IbSgbDTnZvmc/aPRH8rU38Yc6MWQzFe4dNdIcDnr+lFCnw
l8oy4hCixho4P4BsvoZr/I4QHi7FjP4TEOakL2KmrSmJqN9qU+g0Ayfg5ZlNN9/5
GspsYCs4tPtc6CQdaU+N1Oai4tBEjsmkHcc5nPjUT1wWkFqmdc/HobM14E5up5Pi
+UxpbzVjKKphw9c0wlkQgT8ZEsjsozb7u2D4BT4sc0bLcJtjsVNnt2J3yys5waOi
Hw8PqFIHgI+1dX8pt1+B41jX5Brr93i8j4qla4zWzYoNPUQwYI4KxYugFkEkHsut
33uf0b8vMmvEfFNvG7tWkCMM3DfvYN+6fQ8jN5YwXUgYPs/z71K9tPQ4edum/1BY
TCZT0z6g4YUoYA1Vv6wXLE22+1jA4O3DRRhLyXHdY2ONU3Yzt6vnFmqt5tl3/R7b
fMVvypkvTt+m0TpU2GaHafPCqHXu+qe69Aq7SmS7zGtBOmQhl9/LUy03vKU++EOM
kud1R+b2xV12lR6Fwl4CXI0EqZeTIWnwxNvIoaAhSxV8GKtv9zXWWQOVKs4lzuug
un/tytOy9TbBmJPsxM/U8MYDVr7yHXPWAgEQ5jNdykAEl0yyNYIrrd8uT85niqrt
YJzp5r2HxHVyStjem3/l9TW9wQ0r3MyEi7FMq/AaYcB8+MrzhlgSB8dGa17t9Rbb
lSRjV96IsaPVnxql/jVCAcaffQ/fcBWT9b4wdhoGYv4sVikbczs/TbnpQQuc188u
+09PQZG7H9EtT3cudaFI5pQvVAVpHbbweA50FXhiVVX9bYlfwSw8nl/v/HWXJNA7
r45D0lveRwPoxzaMAfUXwEcRBnvoI1tf6hIN0EJMHS7+75T/fCSYmUpTVym2v6rB
dNtsM3XmdgOylJe1mdNlNWcZDuKtLQLGF2w4RIA9WpNWoKAFArREVXvwZlvxtxtQ
fdNVedy9Vpnouzo582CAkG9u/2U4BHvqojf/MClawSM8KhVr97dvPVg4G/KV1E3W
yYRP46x1C/W5EyyPn+6/VmapEUhXzEveA+Z/d+6uYrWjfGL1uLBKLrLsCGHUtMrK
HSHZMKbldsV5rM8wUqCA3fbpM+TZyoY7uDxXuIwY+ppLDA+jzvf563mCXjzQL5sV
f+k1CEybzuzOzi7b8iJ/4FXRS7t4jUa35CSL5sNcDdi9bx7fP49pbDnhtmN+jCGt
WDslUpWUBKv+Y6CkhG8lzVN2o0CVVbcvP6p/j2Qz0ZaPKq7yPAlTAmmwgz/ySAo4
4jq8AlhnB8+gIWpOQTULqPkzziXPWYthxLOlyE+V6qYsLsdNRcFTcpxSKGdNgOsr
RNyxaLmVTsqKoQsB94B5mQu43WEAzFHbGF/s/+IfVXA4KUxgWkKPUY7GP34YZNYa
j004IDGicKN8ZfMW9+ApFYAXUN71I8rAcqkaPuTPYjrN/9CNh6lGb1LYMs+IP324
0xmMMzHurcMTM+1pz7BjZsFcEuGC7A9FGr0YGvjtGge8JDKoBZrCNpWGb+/7FgCe
n/oZXywrhrQ+aUaXMZu9xQQYcCoO6v2MBwftYyqdsBociRe2qx1lPNNLiQPSOAMl
FtJyE4Hw748A0UAbRVE3W4gQnK+gtVg0IofCTgXS5HdsV/YSWZHTq1qK1B3E+E2V
RQJGGeSY2b20IjMe98isyCEOv4MF97BES8qJSN6PnijYEIIr+BjLBtEskrxyxuKy
u1AurPcfxFW3AtrcFSZ0jszbpRYEFpP523Xxxg1pdEdn5dEjLuj2fNDs8Ww2WLWK
B/+/+UctH5Ax6u0e3b5YrCc6ydxvSFVicOJfx8OIkmKoa1DA1GZM5E2AZ4tDgBhI
SCPDjElc4BmF8RmibZzQ7Y8BpStyEl/PWl3ZxrejeVg1FcCZVraC2ArIsiJ/m7Mp
ta9Y7TvrLcBeZkU6hIIgv05Yv77/n3kieEBCpZRIEf3Euo17lHnMyny56r3b2IFc
5CagLHfS1W6UdkpOUUO6fjb6Q5S1g6f6fV/4RQR2qsCcn3YHL3deohkaB8mow+fi
+rlZbNRo3WY0X7mY18hZTIAjBetZQNAs8VtfGUm+qKiSSdbwHtt3hi8LHVX1Or9Q
7pAORiU1S0uwJQwiSiR5rgP7qv09DIUo9GtXpf9+HO7cV6xzh128FXDq8dk9GKvG
gQih9X6nBYyB2VCcXKR559aFtuIxfDbRHePj3PIgcp6u7VWb6jMS6GLCAFzhFm4u
k6bQxWKXe/hg0deQP/F6MpTO1Kyl7zsaF7HO+mWVDWjw2zgmk9mirBgWp7mt7Wcf
MRgS+8dXwD8XFMXf8B9zTHLY1DA1ab3EiLETSXbzSJKNEgKE65KwPuy9FjfX7Qjf
2TO7KS38dW4oRZzMa4e6/qYymDyUt+9ROEB6nS+0T5EEWAOrfl9WS0ptDFF9csEb
q8eyK7S27JStiFvG0XHX4DZmRi/vwGG4nsqcPyG1Atio8DvJu9/Ov2iW1nJXYgrA
gCR77IBaQR8k3fu/CytrPGZxuF7MTOSURthmkKff2XH+fncLDq3tACaDbd5TGhbo
o75KM0WnLAG5Fo1Ip4SAABBd0CFb0IplK3ICBllARAdfnw1gX6JV2vNe1UgkVt2Y
R0196Os44KDg5D4XeW/9GSOznQajjoK4GpEHn1MYUj9NQ8W9mQH0cnm6rAgON1x4
RZb7R31hkU/ywVfpVFt1MTzGjE4EuJIGk9dOUE7Vyw5DyTbfcAdPBS8GDlTsTNuC
aFGHp3Y/PeJ0cBKjwSNKkyovDrilx88x6k8u0U+zP5sy+MsVfxtBl6ZyqX269B4T
CXQnFX8JBxXAS7Nf1UhFb0f+XG1ebiyOfZNg1wmPjkdiEu3Uk5hLxaiSY8u6r4Y1
ikttOrvHtCHqMEevqOkaemnK3SVRLqmV5Nc9gyaS/5KU6yZ0AynovdHdL7WP3hOX
axYBy0MFI9w6h47G6w1es9j/uyKgKQ+iH/IQoDDq36/LgnHeDsrQITamvi5KbXY+
f6XGJZ8TjhYi0wJbW2XlhOwwxeINL2rb46c7tdBvJ1mW9Iydi5KCOqL9mEwLybxN
DQN/dv5mxAwzlsxQ5HDu0kXKK7G6fW7ZD6FginBElfLG2uUR/VAm/yiaGIEV/e/2
hIsRMUbiFl3u2WojetWShPBIMH/EFUWEzJ3Ojau7mzYyisKHmljkPuWt+5XVvNC0
q6em4xsVrbkmXzG+AC8jMyrpBJUG1RdkWjfppO9U1LbPbq21JCley/yfb/wGyqg7
9h2bXDh4cXAphGgQSuPNwPq0Yn+V5VTgolGxG+I/3x7XAKufdn8Q089DtUkG2cqk
IloBUVML1ki+mghr1hK6ObEsoSJp9JnO7IZa/9j0e4JGaY4cPhRIz1FPwiSGCI/L
sbQW7LZMFYHHfTPASKOq9Cdm2HecXjB5+Bt2lAAGCrVXZ5/zhd9euJoZaNH0v+Hf
oNTg3I1ny+vH2/6dYnDT1t5JltSuw9s5AJcQvUnVvMQOCmgOIDEXymo3bVqEdOog
+3BPtmzH0pcGpEhK7Q2BrKppf7SbeTdfVCZc5AChEy0wQxOL7qFXQVHwmZcxuIYc
YMgsOGgDpzFYnKE2wPDMR5vJKAt/iZY7icXC9/vgH/5mR6KDFCpADqD77UUSGnPK
unRDXQ0rXQS5pkU5EmGSBEPduMGgFQ5M1W0ZaGYHtpWFlvaSecw/CzpezQUf6IQ/
ZCD7ObxdGDlXwgU/RayLUrFAnGTYL6zEkdYqInazxxXqFBc7i5xBTcP7x2MbqKbm
eN/9O+S26MbggyBJ3x6QP3ar5zVt1CX/BGbZlw3v8BjWyDQuYTKCPkkNBbT2gMks
sOu+YoWmXbonQobvRuzsWLY/yYzFFxl4vIBldUVSQ/vjp1ATwQl0QRrWQJng2ZQY
Sq2h/lRXhdetNqGswcVfHMAkkDCLzCZf9Je3Kas07bsOy7FNiKVg3dfNiCDOc1rq
8YZc0cIJEYWJSkt0oaznbAPgK9/XikogN47xtDkA8qi8+d/eXV7VRUuE1zDU/cFx
4tchu7/Xm2egPXQWexwM60k+JuNz1mtd6WfL0xZemVXOzSsEK62DCZ05vL7ult8y
Ab6UHD6n15tir4BsXbtILkOUDMzQ34z2WFoIdE7toNUZQwFKsQqHJtxBL7v1uFBj
DK3X3RvU+MqcQ7uYjqIIWtdSHt+BUyb9GM5CnCHojcBJ5JLwYEDDtJfNG9oDdBTh
93BuJefVU6/HtVZvATEC5EqBr4MRZDPa5NNexR4bsP99jEwtdkwPP2KHkigY6ReX
ACfapZ11iTN5LgzMzo1e3FQ/ihtiuBpTw9Aq7XtAfms6JrE1maAAvcT4I73IHl5z
vu8krka0F5SGH4yct986+REo9vxSQPj9gUTwsFggioR1ovJQXGpWtI1Z9Tdf+OI2
m9dHglWWmZRR1b0zo/uhtNSAA6nwrQI5sU55VQ1mOM+CJU7dHBs0L7QLHAWp8Z6g
7fWUyR5ioqETNYlTv2gqQC5OC/+L1CNm3oGOqvRUy3V0aKCC2Z/2lwUuwSEgoMNq
v6SfMqzZ2zfNdIDAmqg7gaxN2GOs4TKJyPwkqxhZXwpg999rOkRzT/Y/iwVdBboW
uhag0VTTAtqCyFH39H/9atqMGg8EGqhGDnQqP0QFx/x1+iW8OwbmEUVkTsHiLvzX
1R/skJaG90OH7yCGDMPhs3cxV0jNvv3szlzO1C9bddK5fykwHLg5bkxXL7/tD8nO
+wrl6jP5osqrEBzUsEbOTMqMc0P0ABn0lA7n+5vqy5rE8XmhDYWug/kaBGLo5cVA
tWhbtIDEEu5lQB9YsNv3Xup5R7sHmkq5bDXrTwAJhWYoETrqpKUqRdgOyo4RjWDb
e2UOoNAuBKTTOf1ozS5jspCrhUI1owiWSR9bZa9JsvtUJ+cdswBhSgcm3ixfA6Nl
8z/E8mvPgfomEyQcQVGG9QdLAH9d+mTuCMXW8a95QkMC16mYizOz/4Ab7jCE1oxG
pf5hkcw2kdz3fOHVBxMFICie6/NdW8XY9GQ9xekXvFwHLoHqfU3h5yeLmFKybsIv
Loo7iGLhzRYFzJ205autzz8m0zcj8yF8zl7wqrzx/8X2aYu2CRV1+wv7AYJjxAL1
z7Vai3nt8IqFmkhMvherilW3le2dOLONM6z153zW9gaOhFXcmGpoYZ7gnBarxIU1
dyEd+5M4LPksGcqOFo3V/a7l2gazFHP7RDWKU1wE3yfCVox9pL7fl8s2O/4IIx/s
UOo+EFi3kVJ7ZFpDPViuczhfcwnpioOZTd2f+X/cIP7Emo+SNEe7lWlMJdrRuksS
F11Rvka6xPBjVSq2LUN6LcR7zejK0w1xMPMwAWG5Y6SBuJIb/BVqW/fLjgJVrLUB
joDs1cagKPaWSF7QAEvUhqghSAfUQwD76fp0m4uSWEsu+yz0Hm5QpMsYEAJC+duQ
usvMliqgWGSBhxtCmop8TSSKh3xeprOOjjTYfhc3rfBq/sehMotHGCzHMlPo8VB3
9vKJn4U94QXsjPRmIFv1CxpgGsSyXJmc14YFFLDkcBH8avwBTuIkcBQXSDEbmd+Q
4LkD6AF8x6Ko3G3fa1xy4FVxszmLbaPBEPFCw/+Lb5VnrD3FXFVXh37Itn0EoPgy
L0xfLOzrOufaGpc3Xr+SsLgWYveWRgwBXitf2b1UfBDB4UaOtLB55vK8KKtjV480
ETcGqEk8EzUZFHYXCl4KTyK+wQeiZRJIQr1rSaBL+DSoTDsrzmXnM21KOjiSvo2w
fO8GKKBk7V59c9tEKgjIZxrsMSlXJU9T2vr13T6TQR1VNmjyGba729qZ8eAv6vNL
AueFOYylSDvstB79rf6wCKyW9DsklG2iZzgKLP/9dxCNY1lQDNi3n/wcRJ3Q2jG2
HiTedLOHZPRzEXpFlJkCdaDgrioFnuSURwcfp9qJC7I1P6hMUWRZHst8cvcTBGM+
VOqK+ZmT5km/8JQO1pYX22ugio9Nad1x45xiVuoVWTry1EcWcJ9IL4/FEg42mABO
0b8+sY1R6OHzfrPnliKf2VUgWtJESaADNa+G6bV5pKRH7qzOa0AXpkP/SesDgvmH
qYhi5WBUBEpFPsqaJw8BbS+Ew86hzeLAEcSn3chhU5ebsWpxz01Mdpdoc7ywMs0l
lsBsY8Jjw3FRzQjP9kdsj85ZFvMDasMkJC0zyWRj8AyJiMqGmJ+XY6oxA/smdBCU
aDWY3UojFzrH0SJMSZRGd1lC3TEvXs8JnMlnK4SqWgK8gdAZSLJaukvL9+tcZw4H
xG+0dN7KdvqRl5zivm3cDJ15cD9JvVzsVFRS9Z1wGKHTkvPeKc7A2bJjxrm4ELEO
mSkn7YYGwQ3kF52V31H7b0WVOf4zYNhHtlfoLKKtdprwZOoboTXbIXz6tT0YL5Hh
jKluX1db+3Ktmilk71nnbZC6m7bOZlIlsZz7K1Y5AAMsT+q7JevcaqDiqEQI+leF
ev9TsIoRTgOaQB7xCVt8GVj5g9jMJrwQ07A2dbkM1mpoLMpqAt5TWCDH+Y9qDrnu
J1q8ZDGNaXN5bBaQhNTzwaz/Yvl/SPyaL4NdPkZZkdYH3sIfarKYmuEEzKEX8KfE
HEC61ktXorjWMfL3N+yIdAx7dybDuXch6zYjmii6qMWTiclSqU33Pjj3PYWzwaC7
siYEyglTvatbuMr87nLqjyim1vq8zXzxe9A603dTGQ7DEAhIoWK8/WjmOoQKrula
C5E8cNypisq1D2h0J85E70nIhlJw5wx5AzujYrITUfyJZ+8cZIQ7BjpN+czuotqy
T3lQADBvRDKAAUqCRn95KvvEhu2+ij017YcQwNPL+Uk3tYi9Ird3RV1bIKA1J4Wm
9GaLhD5AH13jqzwdCcUK6aj3CouM7VGjqA5Jc2Rb4Rt8KXv68vj4XdeC10qNT5RR
v48wql9llGDNnYujh138Qtxw8/jB4o6mUdi+Xb6IIFtGvCw7AiMV31hvr8jcT87D
TGJWxqg1WHk1XOZa45OroQ152HBlpAmuIsgXhhPUD6Zmnf/IGZDflIMwE+TyZ5dc
1YQqenk2XC1hJeLk+HiN8O3hnX/9FyeIGrp8mvtMygOb72ggMTJQ2Ag2lTqG9cY1
KUmCbeQ2ZYQ8SQlFEbSsa4VkJ1TINNdVeadQZyUCb0SHs21nzgz3UJtGxV2jZagU
TMbS1t9BVoMpbbbXUFtJzrBO/nQxtWOLvvpCcoAuihSkjHiU4JG22lTL3vREOLXG
XTeScN9hu6oyIvWo+VkK7vZqPiNML5KbEDUxior3mkEuIo5UuIz8p9QOJI3Wy5vJ
2YIn4r1rCcIzg3Y91nZkKtjPxvvlOvCmRTO3oXKBI1v21PLMC2mxf7ag1s0oC53t
CRiL/sSECUZ7XTI16ME3F3K64n7+upW8fL5/s+z/Q05XOmUR7AqllisI5kWuQkG+
nF5HMc9LIGouIYv1oR6vsA6PbL6mNXUUT6mGe0ExXhT7UxItbUB3IBnMcJeJ5vbi
zEk6jLSo6PBDVcV9XSTIO3Byqn6pi6C+zKR8Bs9sGl5jUTHdAlQWdbv3Ut3Ke7iM
66u3fjvSWmDtPu14quVXakMhZG2ppAVJX1PJu8sBGaU3eg2iXii4i6agQjEdF7FC
9ScQkgddRqfNnhjgyud2dxCE4duxygzYxE+Ucl1JknYztwlC0sY3hpPZZDTJTbyL
KZ91/qm8bOdCl94he/upYO9vstLiv6vPra1z6c2eKGSji6h/Fi2WUORTHSKBllNn
5+VYWdOjFn6mY7DKJNFUwFM77JDHk2ySLVYwumVEAXxnCvnso9QOBpHea8vKhfkD
QpB0ncVjYZjUcrWqgEwcX65SoLjd2YSWY1XjyR3iUbhBVncfdVigkqIyws5Zguyg
/9H2KT1DabQZWwJmvproSvz3fPv//rkIFIq/lRbuBIJrxi7cag97xw07a51mlFEP
5frfT0XXqpBATVQMPwQHSP5SBOtufe2uSH6hLyTnbEOPlDDEkQFsqvybLW/PYsOF
QebpDkWBoFQUpg7/XT6u/EpelZ+sYoV3NXNhM5t3rVIoFqDE6e0s7FUjxYCxjSeD
k+S/83EAvml+Uau/5cCQD7DCmAobMxLV6UVLu9NbqV8TqahZidJYzFqWR+FzTw4M
I3+MtfQCxlyC6Su/k1pGXglg5PJC8CN5l2AuEJbLW34dyOdyXU5xp7np+HbMbFur
H1y4ounW1TWdkFRPNqDl1tfsnqeGueVQcg5qkJ48mc31dspw6EC92IqguWm7rhA4
cnkendDFy2sVKJudrKBcfP2qPLL1C67o8c4ilFNO8QnXxnXGZKcTSJUVGaie3yf2
3unXL4cyC2D8FP7Elhhxa0DpMXt0HYkpbprCo5d6FPoWJ43n3apxV2jkjEbVgXOU
yb7Ru/pI+2ZZNbuJRz8PHwe4TSB+h6Gp4KEeUqHh33gBVDHbK7g7wtLDwsAGZSqT
dh13LMoCx/mXDcR/+MKewaIqgdRrfDSLLnJLGnmXTefHVlkat8L5Mi2yFxpcXJiF
a/W/xlPJ0KzyR2lSpr88RQMfa6T4PficUCU2KsDHv5JZK4uXLmj7/CNw/xPqkG60
1ysye4QuEv0f2uiwSTPNDD7JT542IolotxW2/KBxBKjUkv7mUnTS2AOAgsGjHAxV
pAN9hkhUEiiQX8GQfS5Fl0T5yRwfraI4ZySs3kepK+c+M0FJyYvvXtw/LvX2p6SE
+l/zKTnziUj42BzX99IijvFGGgSVU1uonkibTWkPN0hPa7WGhusOTs5x70vGR2HA
rbdM+IfU5mtZGMuhQmrkP+gFc6VDSBmgh7a9wSpHxeY69LQHnfZxKTF7uG4HKnhO
4ftP33A1Ecgx5XwUveb4RhlV/nWv0v4jp8O27WzFi5xXYqlATVOqGtkXYqHBRvQw
xZGpTOc36ALSQwBAulI7Y0AFBJYrzAJBfsOUkW1AJizmW8YS5fO0zn4IfgYepXaD
Yucux0XUVqLmXkSncNf8AvuHxkPUDuTZrR0IdBT5eTVWS6cd1DNj9nMdNnGiiV/D
Kpznh4n5stxbLmXlaQrKa4DEzOrvKnRYOwHTJ7IHNSrsMYTXbHjQye7OsOutMsMZ
Gr3mrm8kX4OfxhSc+RuiMyhGfttKaTluR0hj5e9KsgwjKdo3I2aXv3q64kXP9Iuq
7AgLqQ+bMp9RW1QMRHB3uBYI3txN6ekM0fzBux520jSWCYgWMZMHCIvqse7I/GPL
OAB9HVzTrcHbAVmxwmN8h2w7vc8eYazKeaEJzTR9MnrELXgNLzkiUWxG+LEaP31j
+XS1rUIc7rb6GYt7IyN+Z6WqxdIPVzwx7UKlxJe6aaWmU09TnR44wSPq7EIUBz/p
I5cZOojsFVz0qSXMs1LO73g7RWDa+nqnRAtjy24886Gdpy1AF18akgiYHs6eLkPy
Byt930rU8hxLoUv6kx8hM+OSc7Kbu8XyYKnWsfglPmtpCw3sL8z/lIIQvgb2ttTN
7yjJJB3M37+Rf4zhhH3apg0XYsFJJkLaO7kVE/uUGobUtOZrPcGHYCoqCPmm7msX
0wivspCaApm4fBhx1uQlY1Kzzrwl1QxILlK0MW0CDzM4NeyTsHQqfNG9PmUzGCSA
X4P9kqBrz4ccWVNohFyD98BO6curDb+9ssDbNRTfAZNrW3qVfWpEGyEXE1EsHgsv
r1nzrf8g0lo3TcF7v0ID/K41PfoejHgwUtvLVDJyVC8rtRwo6AQaTYui21qWVzTk
ShxN2gMasCeGsNHmj7c28RmwFlYXhwbOROJB5s3aeyj+xWXYG5t55BFgtyowwIpG
alNyhdRFFukgVORr4VK4Z4mTH8JWdP8RJGeYsk0NsAP6Zu3AaaMQF9oXWb0dsjjW
llCbYkRhMYSTi5HuWZw0Zuw3xA6BSaT9KqUV6BTiZQijHXlXcWW73h8IysWe4mq0
jrx8SU7ZdNo1DyJPE3QamMVu80jnQ4XUsZaPiB1iIyXquMHhCxnJmtM9FrLsq6oE
c4Ssg/ToeQsyXZ6dZsfS75jfZI3m7xhwWUzGpvhASBJxsDPphdVXd6XrDE3zm5IZ
BWIo9dKSKoj8vjRuOKJwn6ENbgvQnpf15RlCWNzhf3dOnewCoRea6VYNE2VH+vEj
mbhq8fAfJ7Gj2qYYV0whzsFHW4RLRHl1FJ/Av5S0+VPy6utIqSUArPW5KddzbOSw
D7aFDU/9I/P3gfGT18ktgj/HQqo+nt37jzmN79SuUP6ORNU6pUl0l4rgfZrSFVap
IAF2psiKcQB4G56c/3X9KTJLkKBcrfxP+GW4qIO7/OA77b2MrbtAoVK+cBrY659q
19cfWJQOc5KIJMSVkYfIOY2zkQRJ+h+R4L/y52Ha5RwOg+AvRnY/soZU5BRW53bx
i8XtR6SFlIXWxneGkkV66oQhUoDxyPhho7Pro8Q2+YKCTMn9NW+PlWAU6GENCD6g
fgu1idaG35xZJW9zpgXKQbIImh4QjvArj11qUZ0o5Sl03Q7GMFQOSh7cZo+KKgMZ
D9MMfSqB9lT//r4KbLz8pU6aU8xMvj5ZDRkdqoG/N3w1cT1q6tsHfafIUANbxag2
x69cnbeYQUbntgszIBWInvuGwSN8iPkcUybe1zsQLJojBE0umsk9oipOi+pmxYoT
92qhLOYXC3eeP2XfYxfTLsY8hlaMlXjACdViPp1j7HQMZuvsZVgMkPqZSKZL7s0Q
JoMEawxD98wb2k5PHF1t4aQ/yV92SDHkjZnFxdRh5fkk+aAwEO6lqi03rrcBn/ZA
Nl38wwA1OsDJJWFqURiQW6prU7ZEmKc4BdrtazJIDYKf73IpeqkCC9iZU8Ue2t73
1LxCpfcEX8/+DXKch1ZRDhgzSapKmzzA9IQ0UnRNAHHPUJ9BVW+N5ieJJ06br48B
XWOKYhwhYRYagZIquC8SkuiWap2lqaPjx4Nb5tRbtKG8zAFMH9CPcWfBbD25nTRl
edHlsmxW/vub1cIIT7IMVv5Ve1GGi93SmfDgcfFa+O08WJjzIb4dIs5Tl4S4wZ7r
lzUeTaWOuA+LcvEgeZ7V7S9pDwD/pDsxkGPzUREPBH2aZuwfLKeG3KCCgUaSUzs7
cIDIvt6TxHBwIoYPxvSE579Dkbs7bwj3bXKyZM3i9xwk9Qk9hKPz+DX8c6jzAFfI
K6kfVa/Tl4Yxi6tatzVFQcKJm0MvTKduzgo7SD8jMXiQkvSJngHLgcGwM36ckdMR
7h/wLANrRg3rG4cHL5akmyWuiORdKZazTPUvnGR1Y86LyKc68bF22Wn2LPBN9N5V
ZPNejJJHrK2GS4Hy5FwYA3k1b3IrBk7cewezV70j445NzVDeJXLk4jwrxvdsZ5cw
YXdiLy+Fadm+lGzUnTFm7d6ivG152Fzijp7wa9oY+KQ4MwUB0ZZTB8oR8eUSalMT
kusbmq87UfRJKTn4ahQejc8EC1BzKy5SNyGjNqavNlyeJ9OLlprOf8YmmLGbqYzR
dlNmJ88vARKc4sA/o0D+Bj13BnflR5gtvyLJ/KB4n9lnbTbdCVcjkF295mpNzBIL
eCD5XGD88jgW9PdTffXOiGTnHQKncTucDrb80uJO/mr/mavrECxNhikgzfq0RP1E
TT5oiA2M2L5pVwXfXtRgd2RigPIe80soModgEkhkejC8p36RdYMJ/jcgoBP3TtmI
hH3JUZ9Nkc9RDOnV/Yl2yvC1iSl+6wh01y4hZJXbVRySm4wwCOeLDR3yXQ142+F6
k9E6z1cWpMGPZXUl/mVoO+oyr5j9FjJAwg5T0EeDrmJ1F1rqrocqkgv08H06HN+/
lRBRlkbRE9B/SEL1tHxG7GCDhPxg8CLsRmFH9PiK+4cu5Qf1rpxqbwkyvF5KH87j
mmMIxsNf098LHBdFFSzejon/OnqS3ddvqBy4CZ8lWcoTUXzp4NjwXm1m4HxW1ZJx
rBY1K0Vz9pjsgeiLlGAd9C6XEqdIPy152xCU3kk2lSRGF2CQUzI/rafFLcyI6nOx
jyVJapj23jJW3lDpmq7kz+S4M/mUYbr9AUm9/p+OfLYrHUMcrw+8P6G6uL/KnTvm
Vy1guYF49276PXPHr12kIiInC8Bh8VsmCPIPa/K2bp6J/spS/psUaamOuiaCv4ag
pza1h8jB0Go3taD0l6qtHyGOzlCpf6Q1+IyIpbsCo0Fp4Y1HNiIN3ztkSnyaZvQp
roiWTi7yrvtpkkwAjUInVSF1Emy8DbRASRyxBp4nkRIPOBEanWRSVFEyvfW1F+2h
WWhALcAeCg/JKwofDvGToHm+8rV1FlYWDSDtc2GnIQmtlWuyrLmNbbXDqUghH6f4
QM2USerF5VXET5I8dkBIgH3vt3fXOgUKTKjCCVSTwgNrAycDonlTRxd3j2HU4ELl
Xnv2kWqdzniaSO2jlKSjjzYQoFC9Y4qALnNUmUZdAwm/YyQ9ujG/+x/3cAwtUvhI
zmQN9bIXCe2K+DwaIjK+onNQSug8K/AdU1BxviflncQW7+xslJGWmoOz1nsSEvbS
gQesCuVNSpu3lTdW9VnIQarR6aV5MKotYjpBCd8xarJnZJ/qLQo01Sxwgft9ipNr
l71mvl02x//V743OpdbRl+xaBUB747wBjpvXfmyUtQdhiLxYyj+E/m82IwQggw/4
8gT+3+B8o51I4mE5SKEimIntM5FzS/LKvCWcOCq473ndvcNMy+v94N9C/7Yke8Fm
/0AH/VKTFBpdNjVUqUim4RXHVq+iVk1XB+eV9gY+ox1Wq3YDJ/ruqKGYQWitbYNw
VnvLe4+bCq9OgcoP0HVXoUeUyyGDb+sAnPjYxDd1K1YwlML/XiaiYpRt9ktB4fmK
UIfeUyU7CNQh6LJEHlfN63tVdSHtUlu+0ydJ2A9B5QSHMdIuZklxhtwLQjOXZ+kU
5Pi1AcFfBF0kpq9J4OGMXinoybtIxeRTFbIkExSFbiyHbpW618NXKgOq2pajCsZK
5ux6Yc/8PnJUjpxUusL3lXtLlG9g3e2k2YEyLB/gJp6oDXBXaWL3UtVzPsFoPdd7
Cf1DsfGlJwJcZ2fz96PZj7ex2XiAeT6LOzvpT7HR70+DRmCcvqs6T6puKw7D+d3s
K8gr+xNnv+Q5INJS/RPi5tI70CdTplV3qWaUQGYB1DtjvaC55wrb2SnT07H8NuFP
SCocnKWhksV2YPcyy6ZMUQg7d43dwuARDLwwGPSXTRoRn61Bgw2YPI3Ieu8r9PTo
sRnkxu1LHYGtOF04DQSOD+rnAbDyCWF5nQuZsyWBWbtfUc02g5UO/yAjNUmk5y3B
z0yjIwOVg6xyiWGZvoKR8wzI9FPNpLqglMg/sr9Wdpx32u692C4+yoAqq8orroe8
EO5xkvmcTfN4z7Mr7AvL7xEkhrAY3qPaQTIw1D8jv6g9Dp6cpWTWvjVMj4dt0jIM
uV/zn0df6CYAWmdymKU4AQ5GL6VJrOHSpekBjdj3tyDDKo/soDYU8alk/8XPu3bL
GUUYSjQ0AfSC3DmzBmDWe6MWpwgd6h2oaM773irhb3W4V7Yv9CCdTDyLjdnY3VKm
rl5tSILb5rH+GDUhYIP6bQ0kbCMAq122TQeAnmtgwX0fycpkYZcWWUaKZot+zuIc
2mgRaJKcJ4sEFsuqEQ948xJNoyd/L+rXCb2bmLc7fpAb8H9iaYWkYBKc69ntoAki
z3N7hWIAs0LrOjjlsnFb5dKPx+/OquGi/CVlYbZw/Yu/AM5XQF7b9yvtNyzj+MhN
pCIpEfqRmPBCszT7fkbf2TcFLcbBz/r9pD1opJcfb/g2qd93QN2dq0VkfFy8ATMp
WEUyyOhb0ZBT6zNqDM9br9Z8pO47Ls8dK78ouGttQaFwT1MuAO69UsW8wOV5dGpv
kpCDDeFQUlYEEmGJvTKOhSt4IL0Q9oPLhCMd4z4smiDt2AsIGaN35U8+8Plzf6qf
AlVTfzQPFU/K074ouFYidMtXQycpLkaEcUZsn0g7TWXFqiYMB6r/jhIDYOhB5a1p
nKEbyoUcexX0sZ0Hvhl4Oz2I/unTxzWCsZyfSUFUHIzRrW4J8ZglTTgl4Q2Hryho
7wkEnq4eIfvsmEQeKeRdsjbRp1pMJW3ZtvR1I5unBJv7+19/cMFZP5XJ7P8QNBwd
0MepSBkyx2rY3JaSGAnJ6R9u+h5kXi+TamZk37pkSb07m89QI8yZl9UxHKnSI6+s
nLOYaK/Z0hQenhoLjGQa7h0FW1BNEScgsYcqwp6lVvp0w9SStNXLUOD92Qrbue+k
l1avvpHRtAxPDD/jiVFjO16L7cZ254uWwzkS0QqOIvp3eAjdkJ7TTy7tCcSYGbtC
VEpIXNeA6feaxZJ4lRVDOfsGpsi/pJEs5xJQn/2TFQTkFtzFCks0e5QOY/kMd7rY
tsdPdO01ZIBB+brmwaWED/5Dtc25GIDdPWWubsKN6VmBe1Lk4Is34pY7g49FOcUa
rFeN1fKaeEDpO33ee+kpbgiEN6msj4eXDmaIeOCdkZBQJzw6lijRlDZ+4Fd1lKji
EgaI99mhSnDqq3aBt2s/210Y520a+3w747h0UAVxEw0o1z/BupbMJLl5QdUCr0tg
12zN83zrI+CvJTroXw11XhuXtc+j8GP+KGrJNbov7eosqlyGJnJg9Z5+voXl96+V
IOmjNqd8q/+mnyX1wiQOO6J1U29k+5iJyixIVO13tDV4PJ9uRs6/FSfR/DNiZEeP
kB/UwmAA2IPI4kSNX9uNBe8mmQ4bCbyRl4ec+cAIBJ0qdRCwF00luNlWP3Fan1SS
WfwDHnborSyEEhv9BvGivpfue0En4eJ99oVlJlurkwgtP6YbDW2LSMnKiZYkkZU0
btB6E9acOpg+lV5cbsYQtHQb7eh6r6YWP9kOnepVs+7USZnKjXDTZ7KQKcrnH6bM
0J1DwxCCMhZYR8WPiPKHNj8j3UZfKO49foeZzXPr5/GlNz1WZm2fOZ7dH/OaSr6z
fyLXjfYphLSf2V8Apm/ja1YyNSgjhbaYlSU6aYD+U47TSRCFLugoIs6P0sR+dwCL
R2xuAFToU1Yb67TsZ7O+lCO7rVvf3UAOkvQhAUOIy6BHN47asJ9hmNmRbTsUEJZL
ezd0/rsriBJT8H7dADFfjttM50P0LTN7m3QXiEwMz5HYjKdsRH5NLYlv5LxInxj7
Askez4BXw+wlrUkbK6pD9dxCjVJYU6Iumj1RASlOiz8r5A1WpSKX55Azdl1ZQhLH
nk7c0lCVHzJ8kPWwerh9tlHr9L3bDBTSDaYB8OzTJBgkl0ifAr2EkMnDhjp3f7be
2exd1dnq5FSRG03c4dRQk/NAqEVxBHW/8tpFfm5SOps6fHmVZdpK7StpQ1r3q91o
8GxiCyLm+Smo2LvzH4PBYtG8OjhPP1vaq5kFiybFkBmcoctZPyaj/yTnzAsE4j9q
A3bF2pmFIEbNYC27DS4o4hrvp5RHArVvuyFKN/ldsyRKSGnTEoe6BlZMWJaVq4PD
3wiNH05LkbLQE6dQ4rag86wFE/gvwqWtwxUYDNKa3uqaiJXMifwhRsR/QRbvxqjM
EUXsVqFiCBvECONSp18jrnm/NKY20wjtBZmCM1k4rbIdbBwoOL15nsGxMAG7RLrD
OiigFW6tlHFoG30l4HQst0rOHckUGVtCe1NBQRrJ7JTNG/TB+nWI48qiLsFT1OMD
56NYK/B7tA9xOdKpilh5NlwDn0S4hHfvYUoAVolqw7JyhGAVEtFO5CuuxtWMCtXp
ewQr8ZqaHdNX84IasHubOy438oUAKMLcz1R/Jk5AdnHpZHvQRY/P39bOKSR5stKu
KCchpu4K5K4p7HQHG78Bkc4OVWhjhBf2V7kcZpaTqF3cNH2b+eDKBoQ/CnWkOX2d
eAftXgj4nq937HjgggKaXyIW3vxMNrNI98/KO5snHwQCqNwA3wrushJk9OxIE2rs
Qc0yuTPXIfyG8/bHn8FzROANRNp5H85YKJbpIbyjAygSEB5rM4s0VDGnhPhyDlTs
KdIbRLLEiJKa7xDfcQvDyaKcBYrHHr2I9heB/Lq5tkuEJ2gPpdR7ip9VS+DdVsOT
0a28AMe5xcuPUj+bim6/nNeJW0Fc0MeAurGIqa6jN6prdnPhK7tLuJ+W5qRz8Z7m
NRse7c82vSKVEwZc5FyT/6CbgKaCU0PqLtSt/08jOLeDOfymKSWIh64wZiQoA/mw
sy46FHHTCgw73/WnSMGjQGLOOmqbpLzunQtPfVaDy7/mgQe73e8mLcM7kFb0UUkf
FmMc4zElzoQV7bwfqjSCFcxmE3UEouq25Sdl5OrEdnwIUS0Zxy/w/m0N7bVxKvW6
wFxY2ZfOWyrTsVWdnavv55BH2d2JXRvtt6tVhgpqvRybpkPN/mNqm8YIC2uMEKJJ
2zSSvEnRvlKl156aTyIcam3WyFP4QTuftV+mfAQQTPBG0wxEVXgJvH2YJYHsCSEA
WzTi6CuQVhcVwu1/+N13gEsEVEOwys0d9655FrV56Wup0AfsMc8vp2914S1Icokj
rEoBToQMBCoBOmUZfGabBmnciMHwGmnEhMVu60j/Y3rkse3HksKHfe2Nl+Ay4PUF
gpN5DRelhEWCnrLnQNjbzL9JNNtr22ux7NQfX9qicVQlfHntNYTysFHVP2lQcIJQ
t0cwP7hlEA+j5poVow8kQFKFIhuwUTTtwJtbJj942fR3sVIAzF83Oy5WriAI/PST
MHcGj9VvS1mJxohuflJOIDxfiGqfNLJOQoIqSxE7WIHxPdW4PbR8D3KqBUubqrrB
VkuLJx3K3dIJm16JrgKkVOftiSrSWDbPwDNWyi0wttjYiEDDTm284UPzrvJd34oz
R77DTb5dNwARlsbXD3TwNJVZ7d4TaWT4ju5HfccoQY4wKnL0Cr/07UMlWo+AEAen
BmGl2bD9ikuV/WWkTDFsfXtfHIP1sjMoBO+A7iSkSq0qKQyXcE5x0m4XaY9TZntX
WXdZdeQAeM1gq5uU73mEhwOCaOujz7rv3bRLyj0FMJeoqsVNmr9Z5y4Yi+SGKBTu
/rPjw0luqfuN8RAkEJE2w491/tSX809ko5LP1G3MyYlUkZfX/Y3hy5V+mgecieMY
9guAQAb3P42jEJqBLRAnnGO7RT+v5mKhuy4FHSVAHxQg2h2JEmBwZJd09Scm89iD
rEntMeENBva4tXI+HGeDQezHBwPlfRgrI3Sch5J/j5umXWvyDrpBVEfA+PJUNufu
9STJ1FbyUA4L9m8+BquyDp0WmJiWyESZtAhUaINDCg7adZIKcQSm1lEVM5d4ra2C
nlzjOcM+mMnbwHaVwpXiavBYaABWRbzv8O6tQOMMHYVBNmU35Xb4O7V39my3pdvK
w4Y76S2Zcg8Ft17btDj4wxe3I9UrNQhc6nJcLh3fCQI0WWd5GwajgLeG0CB6fju/
VOxhAAHhMLnmddwTCeY3/Hr8vBxEcjIR5S3gDreK9AuII9MVhPLTJzOAId1f1774
j5QZqoFVUhush/i4ts4tY6vkJHYJuDbFdLWqv/F0ZTkrNlsFy+/axduE8kvxo/IH
4vzFCo/cSjFdbfCiPmmjnLRoPZy7I/sHlIWUl+c78HeCUVBV2VUSzol+C5PSFVbP
RLOmVfoZEWrqd/LLhvM8QzB+Znr25jG6KlXlBIuj/wLmffHXiO0IB1SXXlYBhA8v
LdoLSRmqBGzZ0ytdWZnn0l/aRrTMOSwF7ET5hlJ4c6T7owXjmHGqmEW+OH75ox5e
HWjJGrZRdu4fK2A/7EGEeiFxq2Z+1ytI0jMrPoWFBQTRpygazSQyV7df6lAS0+k5
ZEeAb2uEMgNhenRDsNiC4fJOpPdcSx7gWw8Jye5iu2sLwm4mIq4Jol0iFKHronU7
Hm0A+WFNydTSrGW6yKwMkek517CCPKdWPF64BMnKefzlXqJ1JqGN8gRuUpPRqJFF
wslRdaCnG36c/+60e1rud+gJnJfa4P+dlBKFXNAquUzo/2bUsZxTMviwR4nhzfye
I+IL8TIDFZn/ek1ko1K5aSozhJqiRzsByk23D3jMOubskwAGzKYbapAXRrFQU6/n
PTSrP9yzbaZ6dxOaMXLyhX0d0RqZMGH2j+XcgI50ltdC0WzI9MTBYhVplGi9oio/
NGRfKa+74UZH9QInRDdpPcEOqzbBgZ6ScX0HW3dXDoghr+zECptNpCKDbm2z7+Ip
sCrs8CXB2ESc6XEST2KHPFapVb4NL1d4AHSguDpDw5DsNwRAj1wkgt6UT+rZ4afZ
jBXwEB9nzzTTTeo0AouIeAwGhUksxRc0cgoknZv8qgwHKD8zImpKGubUGAyIeP6w
O7ln/tfBNWyJ0cG+LAAFqzYtGjwEtGEnm+d56ym+dfLkrBwIaZ0BEO3Ir2Ev8EOg
H70B7S7xCxm8jS6F4JNHZvVMGgpIGffeOVYuUTbTWfHOO63gEXlMLXMgQJZnpnXT
bx/lPW47XeSNsfCi3Xy4nynFGmbZl//7HJfGQwYr7JSknfz0SeXgbIayCu9B3YLh
AJo5FNdxqmfPw3CHoz2Q5gitNIhEnUdcpMdus4PSVLBRxmtH71OilOdz2jMuVhpA
HvbNgQcl47yZb2fBZ6NAy4Aa+djagb3MNCzxhYM32hb+Nk/Cb7kIX443ch11Hv+0
uMaA6MC2X72bPN6N9mu6nf9CcI8HaBJYv1ZAqRFLaZ+tpHB4ixd3kLNQ1+v4nOuN
MFs1XCt+5Zulk0vnVVCZdygAL+7ooZeDIMyxgOvXbVQMchUoiK/pmqyfGo2jVdJH
PsJmwXdEE3Lu2k/wzzrwAfzZ+/39uf2EGWEJFisb1TUEwQAhIyNfTRM5XXaI/z0T
bC3cv/QuY3d7bGIKrZV1VHtdi6TPJ1dYlAVpx/7aM8Q2nBt1BUBxhQN+d1hF5XLM
j7HqO62cm3IZxzNQXYvP3Ix8lycKIsawrpUEvZYrlrgtkIuvA/X8tSPffdgcO6nd
MHjnqEd9o72SG/83/1/WwRQOlBDQ/ue2P1sSdiZ9wUY717K5L9zyyYfFIQWovd6q
NLBfUo4GnkArypfQj6KdDeJLYM5nYE81GfT+oxGnJnaDLde7EDJhWx5/QnBPeY+j
23gXniFyknvu7+dINt6qyrysrcXSnYUfKJs26O9X8n2j4epZdC67BmckFvu10W72
Mbmh4pXhlRwbh5sZcO5hNmVa84p+bw+wE/5SbI0jIqKpk21k6XHONuO6l7VgVXCz
J9yQ46Qot9n6pVsqN5xILdova211IOpsAfm0vaw0fkRKgYzt+O8x1OIffjfsQ22q
Z/QaF+8qkxaOQw1SE3v3UGP8ixV8u31qaMvIMS2dToIpy2h9iGO7lYqwnamfBzT5
YkKM3n/y0CScgHsbqruaQuuZlgCHEPHh7U8FLJckWY7K5LpOFBHNUl1iABFTlS/W
oVRE/E6+mAIo8B+29OhJ074zyXYpiR4QbnY1WsFP98xBOvnM3unaxQy+EimS0x8i
kdQfGAkNncI2OSwNmeBDqJoD2AkRWAem5ZMwHmF9/Q7wO8DppwEcHfniJadNYDDm
NQsDPnkNiSTGAlvtvn8nIq+Le3OxpKZyAdAIiF05fonzJIE5LTggig8AbZm5161W
mAGWbbeZt79g5AsKouc0nFF6J/QzDR32DMyyRgWeKEjHnAvOBiArS5wXU8y9/zcV
7pZUN8VXjnaKotJoecOjDqOOhvw32eu3QxoBOlwubNyvexoBmR3r9VoWQkbhh3Rn
9fvHDpgDjXfaxjJ0H4IppgOo1b6fNp1RGnf7jgCRS3R1XIVLFVXTZBJGSVoq+Eup
/JZyWVY726Ejx3mllWT0rIdjBRInKyUkZjTOqF1ZV7Y0LVRbkHxrjcmQs3z0kt3O
9O1ZDrJ7MG9rGLHuvjPlp/QQHT1vzZ4P0X1Q6uI7qyN83RBpaWdJegQwVhUkqLv5
30nzmoTurBSbg7kNJzwHPPRjj0tPeKLCsi8f7ySu3RFdfaZZqxbqXNvb24JhysdL
rAlRKkAJj+7iGdJQA2YRmP6ea5fQ3M346eOF39ur88aA3QDUfbjBFjaoLduMpP2F
rbm4X3ZHa4McYohuvMNzvTc/DP4rqmec0P84VNUDQlOFy+M/Kd82cXSh/5ex0r0J
5xezRHHj0NUgiqoh2kKJV4d/o8XAK5D1LYOQkMNAzz32mwqQCeHyQOTb1leRJLFx
6AcOQlmIm00O0Fm8/MrOJ7VDapMdBD8kTIlem25sVtz61+yRRoEaCXkx5M2HWtA9
Y7T1gr+y79c8VdMz1EG+2zKCl28lXX/MUiIoCMwXqdXPCU7WCzlZTcvPF0yH2bEA
2LlYIkECyXVzDT4AWf9aHLkbp+Eh5lL4Wi0VA8U9/EX1LYPFkwL/edy2JK0ZSm0m
aEtEsfzxKCxIu+xcmdja1rFArfE7tatV8mP59e1y24p5QwT299Af+YDp4QUvX90x
ur28ETLWIxMwenr3usOgpCUprGm/rutzvZmsUfB4NSk/vh7aX6w7f78SUQKWz8r1
NMVrffcMarU+Q7/ykVTKxKJrPC/lLIfUZ+ZnwqHt35tumWeH1vMmlrTDt0fVXpbt
v300/Rp7d0uelQncMjNHSek1GLtluml2OYxOnkdy41gbh4es8qVvdniBvPNkWgNu
xGu4TQ3L/72N9vZJT6ne2fI5H08qAywhiYGSW+sv0WvSg1UwTCgvuuaxxkvWFKfn
VzZB8GHib7pd0zS07pwREZzGsjXhQ6fcXiOHq1/cw+MPytO4+xUTMxNp9fcBO8lM
7OmAniNNP01cXyKXM4iEf1wufRQURC1RXcZ0dEUXPnS9PfVhvB+jGHq5DXkHCVx6
1IrFPt6I2LakRFPmhjKPlOcNcgg9AI+JeM8kRtMiWKzE/q3ltHkU7vnI8ykFjbG6
S9sBvlktTXjd8MiEVTrKXSWzX6ncbSK3aiL7zEDeKBUzGbXJDx38qATBbWFbtVuG
voMQm+uLlaxbuY+gF99HN/ltZZc1x+cjvIg7nCbGX36L32RLxW9NHTNz8bPswbcJ
NTOCVCPs+l2SVlDjrnIKpwaVZZLuKu0CmOdSgM+yzUllFnODlV0Id7wUeJzWsbHT
k9wB3krfkAHZi+t4ht6SlJf+DyKggUhOMv8OEuq/2oVojpTU8ThRWynDha6XEUV7
4V6Wuqry2U3Rn8aN5dbRL9T404o2DTs1iG2JAm7LKnfz9mc3mdz8u/u7QUNmTMkm
F32t5fNNpYoNXN3Tl9SBC3h4ZIIXaxP/vzcLR//MKx2+EojrGGJPsrK5gaoSsZvX
SblQ8rlSMwA9CMXA25ijQQSymc70Vfn2dL7/un5wINAZpw9ILiwsjho2abeuSfp3
Q124ZrUrRKGZ6rwq450U+0DNtnQkGS9ez2vdmsw7k/6uAsVRsRWHn8yT9MvqRWrb
3eVKVRqN9ZT49/Or0SlvNvkMDaD7yc1J81Rtap2vbwfvY29BebP/Um0BLp6vRVmX
g6JXMa2BDBflGsthNSsDojtfIEv/WSkImjXyyAJW1WwxzfJB0ReF7F0j3I0reTYc
1oNTGIvNbzg7pkiAAJ+UYiZZowsXXWEAP2tH/4GFb7Y0tc4qqkuT2XztDzZiV/qU
CkMsBsBn0m+d9P1r9yVvPxGeAWs7fuK4ueHPSh4Tq1nHQsstnaq198WsV1QFRgZA
VkSQu0gfKt7YB7FgQSrdNlKg+b8/kxiV9xNGOTepg8WH6KVke3rCCmaJukaFrD71
89zIGkpXwd6+VFaBa8Fwm1f4mh+Yh8i2DClEnN5kOFRqynelrmWhPvhz4stYtu/3
swQo631Ib/ov1G9c+Wbez1z8XJdkPICSbJLS/Rfl/EPspsCfD90aMWxZqPb13h/L
hdb95DCJGUeNMNVV30Ay6JMiwpji0WKmvi1i+CNZM8H/fyEIe0BBOROlDu5/BlYX
khDo1/cC7krRSnflbshe2P7fPx1LvY3cVhaU+m91WKUvFOyxmJNVgTTHNKB8/Hyh
sLSazjWeauwv0R5+/LShnoBIJyCQuJYZ0DEsvDVgnd1SA+77IMvl1r8Z7q5o9wp6
u90cmfQiepaZRXydRE9ddqaYSIDfsSpqD4MaefFiGzTXysek1jwbiO9xD/4zZyH3
JAAy762yypoEpo7X8XVmD02H9TzTthY+AoId6h7hoepgiW6j0oaA5OhkpUspCY6u
2cFUirVtNYUzk/4ciegYDBH3D0uXKdkCYbYZMCjJc1pxcyIIwR7LGCcrtzzpKDpP
nU5DRX94CAMMRy/2189JLYHNe8+UrzMe+tyL0F2SCKxLIpOqXMm9g8MZZTZGfDG4
TbDn9lBGVRJibQlwpUACyqDm9Ak2f4E0cx+tX26QaI20dIrpgCUKAbwlaTTNwufi
yniH65z2AneLHo+A9eDJnzk09y7Caf5NWC/aNFqNe5Q6b4j9D5lPN+wiZVdVFqI1
iNreBmoqIkRhlB3mJGlPAvIs3/Q9LkhxKaEQ0tBdHgcBNx9MvbfLL0iqhpWsCHBl
rThygtgNWkvXwLfw5jVvyunMNckzSPCAgXewh9zREyOGAv0LEzkJ3j9n13U2P6Q5
v2irXCUQmb5Vi9n58l9T8Kw9znwvUGDSEgocFeip0LWoBOlUA/zxl5Qfo9Iu2qF6
qt2svK+TPOT71zoEjxqJQ1MWrlLP0uWx89IJR806B5+nyM7LAgJ1ldBg0Q1jIlQn
E6A7r0g0jmB33QllnUMDWFNcOPQX1HThZ7/USsToi869hoI6n2lCWPMKB/okiMRp
7LL3renSoh4L6j+432E8bvVWefyGjwzfb1iZBGTrXVIo7jDofzaF5M/hPs1Cu1oF
e9WZwE/wqx2yJgEVqBEMBweBko94QUaEwKQ3TipVxrwG5YFZvEWMBghYuyCWgIZL
9pXWTgGs26YQ8PvqLC27T1kXBcn9TRb86Tqg2QFioYf6HJYU0rYJpgdHjBqSg+wb
HJDzxYHo72M7EKwxfmftbrdAuFYThPinUvnoNo3c6+2rsa9lI7daVgV3CoRvlPcV
kXdm3+5k1OPnYYqRn3/yhSx0sSm/9lDnD4sun6e715BI4FKoTbNGsSQv/PrTv9mx
HCMFqFTbHRffLLapf7MY6ecXdOWPLukthqEMODRLIqd5+b+Ypb/O5lIszdTgifcP
c363Zx9YbTv1HU/erHuIAqQONti7r9ohPQb2x25CSqN/LwEYYXNkkQndEJ1BVf1g
+MW6swjR0mODc84I8zl3xs0RNFu6+D/dHlLTUYvPLnNxpP/3dHNWj746Cl6vt0yj
h00Pn7sB+YqBlEpVb3KCvb90NM6YGeN1TF1cHgQM6VWrrGy5EyAgsBmlxZjbugIu
cW9qA8DsxGG7yTNSQj0qYfdNpiH3zZXGZ4FqXym8AaeRTC2d87A/7LM0XaUppxHH
iqbnd8elBLpKxLvvAOCMjpiR57qiuNmaMCA0MVtE1PSpkkst/SadMLXrfhd5fE/A
jMASL/f3ZxpnRrybGiqSBv4p6Za1eJATwHJBpW2Ny00R98xyPRrvesrlWQc3rGXD
Npib63qsGWfxb4Ckdxjt0HmHKnctsoOeSK6XGPm+LT5Tyc432nGURjV5xOwga9sH
LKDXiqFlHRvfWohg4GjF6CdTizD2EXTgnA8k49lUXGDu4mVx/X2GECwASJaebR2l
N5yx1oRI8YMUfaqX0tFf7coKRBCODqLEVP42efXC2nTyGVtLbwKuN/YM2Qw6Ww12
Cd63ze4dXZ0RKMTXIKSMobWoZertIShAwKW/UCpYYCNqKs8zeKjhxPfpYE7Og9GI
We/yg9Dh+AmVs2nForq25BAbEcbpkxLVv/0xlQENOKDbj0977cAkv6b590fQx4/d
abtfWUbqEmfVcB3GdVtwhLFxoB8KbGsoEjUf8LJxSYKpJu92VP5+fPH/hgD6P7mD
9MMrx0kMpl2v0Q2/ndioFSV1oLItG0/h8MrSUqRpHOnOuA3FbZ/e8vV/UBBv9T1n
RVwbM6h++bU05X3q7y3l1JYuhNBCvPNfRhCEOhqXjg7ubiQbCadU72Uv0EWMmRxV
J/tc1ZQxunWJ1gDUwYdex5tqWi6L6wYlrfOlLXO/grWV++WbboqDWKLOHYiVcAol
FVoSmLRHtI4MZ9CHTWS/+Hotq9JOrCsnoGw40FYYDFdzSpQxTzPHY9e+lPHH/Qso
BlTiCNJ7chstSODpX39fae6s2gloaw7qpaaT/v025RXzYboHO0wW4FuT5L7zKtoU
vd4lhir164PfwWWhTuHp3Ihfr7xhgYlS3SdfeQCPauD74AyaaZKpgpvFeUvr3LCX
ZSPop4KalRtSqaMW7sfF3lgH/jLv/NhKY2H7JdWDJXqUHHZ7/WjuBK3oS7DXGiAs
m4lBJZdfQBImrffDth6ZiThObvcoPhDWqDF5VlYj6FiL2fcHphBDdgDSM4CR5sBP
2nfETIaOWBoEI6Cz+kAY0tGpXHR9e8x6mZFwOrI+N6VmzgV87cPDMKu1vQTRvWsj
4Jsuzszv2kmdsMzhghm5IDQIlEPHZG3IIvInDaSRnFU+TgviLv2MUTkYRDxOoQOV
sg1gVLPq6wvBRWXA0wJpGOBTHTOrbpM0HXjOQt002ccugfUFuSBNwxJ7cb3gyqle
R1boyGb3jwXs55/vnmZ4Sgn8CKcnmoBcUlNKFCB9Rp9GJLesE67fo2QhFbVqw8Hr
eNzKjb6Uat9nPvR8MmY/2PaYTEhvzpK6HJxVAyXKJnAPoE0pNQNusaPfcSvPog2k
h0SQDTiwwkQeJC0fN2zz6ympLOl98686yGbj4jpdcEyVH1vVHb5ZleZq4buG5ASr
o6R9Aie6VYyWrr7xa4p9lFwgezwHBh+/qBOzQrvS5rWsprSwmPbiLrdudmLonkQA
3e6bxnVEq66lmrmjf0lPxl+md2ecgdhBCNAuu91ZhZKMufUnujUIgeg8iqoban1i
CMoPRUUp2yk55ld627nVaOE9T+1fE+u6fWt89euI/r7QeCWimGIoV3GRyvxU9dI4
20VPpFrrHZRtYU4Ua8gvTK5JFPeG2mZfojS/f0Bru/mkdE5zO3BJqf+WsNHEI9e7
YRDTGqOwB5NA6Qj3J8ijppr/mpmI5oE72MYKil6LXw8wyXe6EM/rPiRZzcv/vvLX
KzIg06WPR+MGYFXxadzNw3yRNRth8Z/Z3yAyKhGAzMOiUGlXoG+c7zvVVlEDofjy
iLN8lni1iWAKxSahLTS9cgYyJ7f9ktNPgQ2AkKS+xksN7+nbiIf7jYLoUg39NbE9
7w0Ivx7C+uyUAX3UTYinG/OAag4A6AYlvvd2u6lyFZJBOt7AVBA4muY8SAqOC4Rw
gdhNRYQ/6ud+HeTVLsE3HhbiGpcmuim9uoE+7gz0hT1tn/qHnO2Ant1RNoSbU1QV
IWMQJj0yczpFNnxqsSNcyXk5m1hrH/dgLdcj7WdnGzyVVqCJ/Ic0LfY1Z4PvUJQn
hCFjbzGVeha5OEPX8aUn7NGy5TszVvgYyyOI1E+wufsraqFuP+mRvD5KwtNfnK2j
VDAYI4+IGGXFQACbkPuNiBLnAu8H1LGcIU1+5kbL8Fry+YOcmnQosYKBgRc+39QE
XfXE9EAszQ3gFkvyxpd0Q/X86DIh1TOsO9/QIDsIm+xtd/xKKnBb50HC6BrheMyq
P8+jdfLZIfdq5uLDYsiH0plP9i9kL2k6rAHBVnsIfLGEmiUtqcYmN0s1aAwgHsbl
x6kye/01VIV29XsHc7kdNjz+0Bh/nzYV8ZVIFs/NmrP0+TFy5/qYXyAJeETvNa7/
n8hLbSece/eDPfIh5icz4Ivi5DguuKa/dIJA0E/sNvoJYcFL8Qo+FhKrqWJWN5h+
f2wkYbc3J8scC8/MjVu54CpyEGkUc+0Ymo+cPCTWWlc0t+6DRl4opu1qEeCRiVpf
uvMLJ9Alpv4p9UMXv12nbQVKzrUFlM/qjvUGObnQucC94ocliNfNCAgtdiyOQOw2
vgq8YDi1Koeh2fwkgoyOjU7Ndzgl3tZsvXyguG+WBvqLRW3YHHrCNjd2jCwNleMf
J0pL9wyqZgcaNG942PgKqliS5zmoeTms0fBUeCcDheKZztwlZjPJbMYLkLgKC7Ss
WTya+lcP7ZUxlfJRW50inXuo5NCvswVjM0HGfshbhmCjUMdOAh8l5PMSio2/jbDa
WmoLLd58F8yoqhNV/xFs5FKagvyxAAAtr4cOQgLqIuOVKFcVOQHlDAzoyIZYfijm
3S/qdJlZAPXe0I83BoABHEJA0/KJxFzclkY5u+qH/Ncm71ZcK6KX6eCT1mZMPvNk
uAEyqsfkQ8bHzhPyfo9Wc7IGQhgi/yQPXRJXfAVQIf+WnEEdM4f/tBsU8LOr4paH
mU74R0oNqGsidCGx0gBRrIA1BasKBM5uz3kKDi5rdAsCsLF4mDtRbT5HAmA36sF+
95KACrDrqtz5/uU36Ms3RJHd6n8tQt7SO4AVAf7qI/CGTh77Ch2cHGlfevDj33Rd
JnSXI/WBSmDmdPhuK3A2LDvmhINPbExmox5tsKeaB7aK8hZ3Ve14C2jVYDodOR5n
YeDzdwCu75jGJCXxXdhs39QM6eYoXTe8Ak/OJ/PjhORkDo0RXwtpzreecDo03JKd
nzWzBlE0/23kIxvQlULmQzQYQuXVwEkr6tgZqgIsPCKhhOhnpvdyAkOWzawnwrD2
qDD/efHGNaS3p9MWoulTX3BiZ1eGlkORD8r+Il9SPO7dLDI+afKI0CsO7rRpdf5Q
9fLM7SfcBkK4Y/mBoj5dkKMIW7GDf8xUufDAb5NZYAI91xK9rvpBbQB0Y1ALTz6+
U9Mf5ePVrvdq0O56YYmwYLUR5Iq8CgKrO7Pr70u9AhAY3pI84t7k1GnrEPholVbS
FlIHOYNWZRSj/CNaETrHtXv3BvjlTF3ZkgGQ9ydwrT6iLi59ODOCyr8z+JxYaeSg
qE7aQqHRpvyIjSGXIkcxn2A2AY+RhXIzplG0nXS9qAY1t2cnmQs6b++dAxoX+9jz
1LCVa+aZ/b2vbSus6K2ckbsk9r1wuikbU/8fBdUvP06Q8jvMC1Ot2MS6bRqHr/X2
7apIPiZ/th1wgFHJfiKWNyblLKjaeAnV3sL31ibqXGg1rS97+AYMKYSNyrAnIdJb
6Jbj8obXFZbe/BU+jmNQZrAA5YWRvjxnVU4Qh2iLHcMyCyx3kSGfwSCbVYWT2lGE
jTrZ5EW2Rd9l41p3SMd7H9DViY8ASfbn1vw1T+YZF2LdhP0o7gStkQ4gDzDujLF6
WlBNBLUgNKCF+ljms614dFM+ZXu9hR6xyaLqUzu+xNoAw5t8YmUGlVqK5irFxb5Q
DpBwUVdpxwxJCIjgeGSKywOoqkyViIyLLQClJQyOtBeiIdd81hK649s1JIVbEy4s
mXSt8IKWUYxQNPQasRMg5pZRzBVKpMmN9tkOUXjdJw/uJsVwHcZp8ipJu3FhZlBW
tSdOYraoHWW/VgB2ciO7UC/3LTL5bQIklYvLwjYzgSN2vXL1/Br4cTc312uwSvPT
zkCciquj+gW/slv6AQNLYk/CYxUa1X64nxP915vRg8skqOkzbPI9tZUPlAh8ZyD4
l4hXXM65qhQU2GGPhvSVjJ4J/a8UAlh6r1qvHi2i7t5SGylLzFHpDqoZJbLKnk8Y
dQTmmZNyS2XmOWrvsUzdVOM++a81jHmogg+6JBY/vymNv5rmw2DZVMRZycnK8YdD
YhNYxDinHhiB1fG8axz/Yz0qyhry6nXCyMr/skCEjBHgWw1PZEJnLenIflEtVe0i
NJpWB9zMPd2WC02fY8JNSAhigdMkwKozCTlcC2WrUnz1WEhErs14zOJGaJEn1+YN
sNmreAXDRxbeFI7VEyjdRQSSOHLYuRzlPhY5P0uAyoTNkbptQ0otxAJBTBbsoyAh
T2jI2MRnBmriplrIyuK8+iZbpBHX63LakPRC36BzLiIKgTPbBe10dGiPSPNUGL2O
JPyeFlseqvceF/LRjKatHhjdIKHZgE3bklvn9ppRkX1fHR6QlNLHl6MRFL+HB2d/
wtTH8kciZAJW01R+KeT9Mp2B0ZfLyDp0g+wTykTY3unHYZHz1mChfn33+hCLanaq
GxB+NksOe6zAOy3Tj6d5Mlmx7o9KGLw3AbRxX/aQAHhqwnYgEllAnKZa8vul0sgf
0PlYAzbjgcCLD61NbxaPT2lvYTEwuxIn9lRxHpWRJQZRUp1K/Q6utZc/UgDy5BTA
fkOaRvxqd6mdhmk2fgev8On7A4dG+mu/yesRbTzvUAvF6zuZ0ljt0SLodZP5d6EP
1iJX6WkCdJf4PPsrn4nGD1EMR58CrYQpsSjxryjF907fmebXd1gD87tFxn/ciCGL
cQpCoJzteNy9TKShBLHy2dgLbCPWPQMASeYBITzqvJ5kd6uDASfk3jiJQG75vlec
GHq3dU2E0EKmpMIVyrhOzH52yBXqNoKmNDiGGKi+LQbOEWkOsxKrQ0b4NJO7lh3N
bPzj78GJfN2QAqSyDEbRaSZIR2/k9ut+ZwD6RpFA6rh6wu/RbZ3yrVpcwVAxGWW4
eMlwkxVURF5fVQHBs3pLHW6gMVMH2RTFIwn6aDLio21hbvVR9D2MLK/BYrbVTX6s
GquS7RgDtjLWZnLmaNvpk6wj2lZQgaF5ujmsMlEvfeqxRMFXtxlpEmODBx24efC2
+3RgGYv6WxEbTgVzX3uG+pxZa/PUwyrQhQMivrxWrKIcQ77g32aBCEzeNZbQAQaR
9o/lYnHWeQTfpHCexmX/Mf/vAfZgtw20Lkns4CGufBzk1zRo3Gr4pqRXXQHycx8V
NLrmGv7QZ2Ws9jQtQoB5zNCuuoiPItltQxV3bcsQSh+azDQcCghTcbE+ZiHM7rMD
hNZBbTzWr4nFmKXX82N2be+03Lko8co+xpQQnjyOo2aekYSapw93BQvLWjbpitgs
MfZRytm6zPbGvvXJ0bk2Xw/+hNHOmjwfRguReE1WS4DubPuvwMjA5IGftoRscXrH
em+bzbn4ptmxKuCZaRUrXtL75jBS03YJBG5jLzxu5LsMGhsVUWE0CHwXmdjxfoO+
9RpY2vy9stPDBl56VXa+NT0JODmxpQqpEGvHpMLGuZgs5DRmIOKLu/G5275TJ+Hy
EFCWEvr2qFsJZdlZluLj7mP5sehQvDtGuXbMENhtcaKGu1GLVp3eteV23fM9UwJC
OFSaFw30b3ReB+3SxHcLNl92uRer/CwBRCpjXIWooiffBXFhGWwabQNvusQhwXr9
OK5JpD/7QdGFtXHBa6iIfNu3CulFyq1gUP/shs/2V6zbKS8heNy8qevwwTtu/nNe
5VWeR0L3H38PwjcRu3tVeCdKVbktjWzmmNhP+hwiESu48iPZykYeWsOYW90QGHO4
am+9e8x4uR/tldLzEqOpKYaGR+abB/EI7MO9OcFYej9tskuVX2KaKkWZVr+fTZAV
CgquFXGSCm1hFBYCgsYFvqO5VW3WshaNqadMgdDrJXTc0vDZr/iDrz9Gem4p8/tK
TiGMmtAqjFA3RYsmSspx1EYYH8sqgf9ob0jblkxtnmhj41H6NpVOq+nehTKGn2tQ
hDOY+0igCVOiaAmeJsy7dT2vIXzgjPpRoHKOayRFr6SMLD+76KvkuPKummXHJZIj
aOg9pChu/TYUVb+XUWu/uum2eLgZmSbdn8QKv2BQCjI71fHCe+ghLpYASbiSa+v/
Cch+V6+ntJCv9fKKURfZHsNFKlYGI/+drswMDzwu+RL3Gm71t26jJJGH1qCYX6LH
iGuKguGoQxsm3bnqer+C2T1vPZS5Da96X+NTCaFqqNhkXSi6d1BWkm8B79sbduqs
azmln0mKbnfjQiwL1EbTVe7o50n39syZ3UWY+bqrrpmmsyurhwrf6uhBeWKjUQZ+
e4VxuraVIlFXV2AGlTYFQsB8UnKM/2b1i8J43QwVkSb2EFtrUG9gMCuFmGA6sZhP
oS81gwSPlCLuK0ae3pu48756Yp0lPBJGftg6/LoWypq3h/NtqmaISuxC5olV/GW/
5mRIXWFPePa8iIXxejUUdKEBizwneUM5f5pwJatTv/SqgpeCAqtbyOA/cEgFEyrH
TdTukTZmru551KWAeMDf2riBE/Qzo1cJyCfk8TzAn12nNBWf+RWOjqT6xKEtpXhk
7BJoGm328zopvb6x4ySDWsQ5F7kwgSv2NYc+6RkBEcQLXQJMsSu4a0ny66wC7/H5
MD4flgRk4rq2EOzzVVlArfb65mjrkIOIny278jpBfLB99Y0CvNXbQ6vN9KAv3SQ7
IT0BYauyCl5S65GxHg6plzgQWrV5BLWT/IH40CipemM3RoirRLyJ5zsomKbsJFyD
SUv34t122G43UUtL0fBqaFTOagq91rqogL+aqQPAP+jPHu632UbTLGW03vwIQ5hl
5r0j0fpFrIGURySFJVE3UpSO0KM03rOD4/YvUQwCV0/dy433mfrQ2QyCz9/Taqwj
USByrPHoNzT4pNWAFcMskJbYT8U2Yjxvsh9RzAZrxLMZQ6xEkU93KC09or17tC2I
zIVYI+gRE1bPLDV16RqXYglQfAvEIqz9BfmazJHl/Q/k/6RlPi5/PxrSnvIWbDxn
CsjxQtnKLRp41wb3Z81SuDelXQF7qyFdUCXcUKwFgMfb8VINFsfFMFCj2WgrKrZg
K9NkD7uqbqjnyBY5Y7NldLIAymE+W+5iXhZSVuZ2JpBCGsJr1cGhX6l3S+dLoWp6
nIvCCFxbEUj1OTMApsdMgVv7qhoLfd4Q4myWCZwhDanmxFQXqji0Ab9rn9efCQoK
hr+X1wLP7dTGhaWOyCFT8hXC9S6tp5nn7QVY3c+whissrcb83D5zDe6W6aEad708
Jr2UT22zrv5fexXni/92siTrtl88ty8iaYTJO2HbU6hK/45GsuAGQ7BaewS7t1wR
4t6D8Rz9fySnfjj8xVoj+NpNoZoIhxG9LC7e6gVlZAnq7Du5LgvoFaz3pX6m6Jk+
vXwYDoR8ItFKZvTLmBeAFowBp9YkYtumQr9A7x1UEAWPuiG40GO5bd/knwjsttO7
KeTOQdyCK36bx+DdmdxSXDIdsGT+xhBqR7MrOGAj5wJhusRAz6QgUxQHaPeygRik
w21RpQBCy7sXUtuIlBx439ih/+Ta6RoY0hRO0XHQx4Zeev+bMP9d881v1lwk2iyv
V1u7nY2owFWhA50HAc8cNrRKBSR2rmhRqE/g8ByHCxU8YOwCyXRmOSgeaebMoFop
Itm1ekQfa7t5BC0oXAXoQzeNgie4fZVw4nLofD0fUCgf9cV3vSX4PLymMHYdP41W
pMhh+Gf5vMW3SIKLsOtOpkgLBxFv0sGVYUcNqTU1np55Sc3hWYaQp0LKv66r3Ceg
KtXLf1yZq95wgjSdfdcB6R3B7oAjZlxKIb7Zb9RSQKsP23CHvNkUUwippsNfOvli
VZPv8y6veJd33/eSDbL8GNIo5bQaTvlHBi30yNVJYuxqtnqmhcu+mtKA+HRQvoRs
zYYcfCRIDBrlLsbHLR5T/eXElF1KOWCHvTLewK4yZ8Iq2ZqR5SXeRj7cLkyroeXh
fmniqwHPMkG3Tm0xS49xDBKZRGp8tFkV6F4aCeHgoYDbroduguD8Lz0rYmKb310u
fbG6W8SX7woRDtI3zgzDStnKxUVwRFObIJrj9HiWK0IhGdT5ax77mt4TwwIkzrcf
Ln3aUXCgWDPg6Xjan2KRsSWzDRQwyU4kKlVP0knnytAxAU4/Um/X7r7YekTqvyoY
4CrEnH4xQ2cEQq9ipZ8HZbG1i1TB2bQ3A2PDkJX6WpkLCVoD+tfX4ANd2aRNGZqH
98flR4FKSLI8/v/a9Axp48HS9N/S7RbWFkS8GIoyBEDd4mNLbaudBK2K3AOcT/vi
RmKzjNZR2BRRadUxkj96kcW31Of0UhiRvLi9imh1+gXGGFW+i7EZxHJZJQKOdBHt
pdE/fsB0VB9iOANrJiO022kLW6hcy3jhjTCfXnPkUl9vfaUAV6OwyzNETZlkMtRb
wR0vmbIqR11doODHrQKBZTNVsXSk5AyO/GW3GlqFfZrXi2hlIUnn8siWgJrWknWa
rcWpFJvsDAar2P6G/5Y5bL4/9o64FC1I+GmGEe9a5PXQ2Ux81wg6n/SOzRHYgfSX
ziMja8FISQu13TvO4AqFoiwzSel57Odz73TesdkkEwYeEHnPzEXcJr6dlYVl0nOD
TdSIl6Y7YMsMMuv++4kiDNkuMAvGN+07ZWQrk4oX9JtLNyiRlTpQnsVyeD/6k0tw
gPUCuu9nCENs6YEgjYZrrSdb8/GcqUDsTFKMPXV0n05/57jCIY17aYQ9sm9UxEb/
Illrtl9CSyLwVUBisKjKHv4JFjEpyA34ZtaQhgS55tOuw/a2S9NlyD6kdMnHm7P9
hetO8mHGT5Umo5R7eJV8T1WhFh9kawu5Toaq/PG+XuOZ6GR4Y3DDCSFkHbHE5cZt
eGGYHFmWhACblIAxBwVwMM7q9I4vbBNvqcUKY8bQsPoJpiXu7QHU4RzisrfIEYTE
lcThjGMGP3J7K2/oGffniQescdxv9MRToseqRW1P40dwOrraNONVdy8j032qpot4
O2vrKGX6UdXob4BsIyfHAhCRJ+Eu0JoG4EtOp25g6NhuiTOk5cU1cJH2V56zkMKO
vSzWPX6zTbtdRWm+yRS/l+eUGQ2f5exfizHlD9fXwnzZP6c+j5Rw9TW/lRIADJo0
vxKsTC6GMCXBVIrVz3C/Nby577K55SxZj5pXTYcMmAdviCsXh88ndCyUDJQZ790G
jLZIvizoGLjnbfKXW6AKlQ6OO5LqkxaRcXfj1XZRUO9hvvnwyrF+LOtUbfztlL0T
v04/HrT/UYrnB34jq2vZSw+BJWl2X62L5BuXMDAND6+1Wje+fEN4jZ8lMyoS+SBx
L0h2lRPCpxEooeW81xTm05rKW0pBP2PSfD5Wf8jVgwNtIJXtjk+YWVdR3iXj46Zh
TR/+uKhBtGmJ0Jdl8SaNWZ7dfQuordd5qo03DMHILIKdvtMBUB7qt+j0JMQPLfl7
82HnyIueE77K2dDPq0ELFbONv9GJIYvGnUMJukXmXmSZoIoz2FqgijyIB99gZ5w/
wS1hGsdVaqamrh5uC0seOens1OLbcs+e69m75Daez4dbdBUNSjl0ivE7Elz78ISG
kw8XlifxRraRV1d8N0dYTf6VRuDuMjE8Q98tTsvpnb/vHPZ3h58Kk/wkTN/MMOtj
EhYc2mnViYUtkNU9Yu2SdzFTghFK6CqoMZ9zlsE1+/r2MdKX58x/l9ehDgUqT55L
O1m2uK8dgDgZvTEbEKhLFT95oVF2Wm3cgauvrkZtbeA5yeOwQGFITOflc6ZlZe+E
MZlVHlN+qz8CQNDhTEHx4PNNXFASs24eTPcgig2OcTaD0bfVBEKRgmmFp9AexabD
j+NY5BIHM/sL31RXVO44fYA6vxF0z+KIDxdYN9GTBHkm4agPwvMvM2P21PazfERY
pF54qWA+ZDTFOtpv/riRT8gCUZr9cu0PYgZr3qrz6xpP7LDjASF4PI4MgnazHORF
FpcyDZs6X+8Z3YQrlPT/ObCT1ehb4KSo+Xzoh+RlnTqd4hzZ3UWsJBJHTbcJyd3B
PQKHhh8im/ZQj37YvNSb8dSZ3wE6/KTrZXJxu/3XpS/cZAJpUu/3+QdAiJpTZjGR
7CNY4+epGlZm2J18f5S2BKS0pW0mPacfPuF86Jxh9w6wXkkxpaMyBWFALLBI5ebb
PvP+0bISXAzHyY6TZDyWv4fztJJNRPOF8Oi77q/FI/t5qeSqyVUM2pijxKx/qLbB
kgfGU+WH5+a7IyEKztmwe6C1TBzrPzVjHwDPafA6q7QfJRubOe2OpCw1D1uxTaZ7
xxadxlBfGP1qvzGbBFl7xJuQSLAY1E+1SobW/ZEi11eIyJa5VFH6Ip0VJcB3x79n
FdbQ5SUX8GawI+8/KARyPogOS4k+fQc7w88McSuzOkHNmTjrixx4MbBI0zo2fhcc
rdVCdhMQs/izyjzTr1FKuR3++qDIaT0X04AMIEjypmZW8M04S/OBI9Ee2AVuO69J
NnhLPR2YD5SvSjB8p9EkfYJQhIjLt1OBwKJrNVOyuLjckAkXYyN2EBd17BAYmFqo
xbPaMpc7syAB+0IE/vEIfQKdAdWGuNqbnnyNt2y2uLbmRRdNkKbyGFXy5teFyaoj
G3l4bx68YgLVzYHuweydRGPmzm06eOost1OGVImeiOPC+imGWYOrheI0gPMkKDQA
Kjhu9WlmzZbXM4JKRPnoOoKV9pb9boiFnncw9pzGiTlZQZx+tUotktwXN44ufqcQ
HyQ/vNPan2jVQLv/p/m1Nd+IohNW0Kp1sTOm+u4q+SznuAF44w2BLpjS6pu6fZem
8M+rWYTTBPaDFV4opHod7UrhfoNrc/bSDQuWoImQiOR+4faxrRO048Qz6IIKLIV7
ZoI79Hl3xExiI1jV+twiuiZA4SXkECqoEyAu5cbo/zM1PLMpqBeWDTUhuWVjTpHz
WoxYA5v9/hNA7hOhTomzmsaN7dz15trxDfA+ow29nDHnWjBxQwl55Z9pYRsfUGYQ
vmXv/pTl3pgl7DVVnjS8D9tGFXErMRAWUEaKFObW/dNEKHb4Tar2QSYLJ8c6H+AN
uDEBCuHSSnAyAVb+3aLbjw0D0f3abvhP2GyNgFF1O5aOB2YBm4zM9dilMqQty5BV
cARjqgQx7RgkkSghe3HymfRHI8mDf9AOpX5dwrqU6oMBakg9gpDftn3aCUpoyvoW
kcmHLQDlgM41XXK5/QqWix8Rnf/qNqxNgvrzsfUuNwMCUMyDh/oku7yBR2dMUstK
bkr+E8xPFIH0sp8UXlbhDIPSMuQk4CJAl51RzTkeZJPFB2tm5S1dGwiN6SeuZCoA
OurslG7Dc6MXFkpG3udjclNGVl92CQPAmL2V13JpHd6+ITZonr7/xiGRbWw+4uyT
SXspoyQ3oJPi5nigsZqh4f7abC1Ka4wXTgkmo9w9QaTl8rplNa17Un2MsproORFF
YQ9MeXqp+IsogjXW947anF1NOD9mrVFpU8S7xFel1FasIku9RoWRDmcbkp7mnT34
xQR6JwwLJOqhZaCiTxbJsiTXtHqoknYRxfhz8kOUPkrP/9SmxqMgyIPVPWC7+CME
EK56bIm4Ttc8mJkEr7dLUo839NzMuWlZrXzlW0GLo21bB/YSID2Qdo4xkowq8KcA
gLHYyQu/yKEhCXbDK1lZW4ggw3Ch2ILbNKqBYvzshA9MJ2o8lBYCd+LKxa/t7A2w
CL2ZeGrNomk7uzPnoV20Qo1uE4tWgrz+aLBv9UBzYLrHop53PuOHApp+B86pfDIa
ll7Tx/GBth4qxu+kBo4AdqjR9IaNqNSXMaIonNtANpGFlUla7riAYfwd9VQzRFBh
sa+tto6cDpeM98nZ2N3gICz3nHbZ6akIJvwSTTcRBItcnHpm+6lV+n7Q9+yxCGgI
C75GNA4jtGQZ+R8vAaawCWTeFJ3htD7yGraoHewdgU6xeMp4dr1IP2fr0doQrrxa
rzRPuFwA8Nw7jGC7mIbXb1oZenzQiAYEflIs032leMLCI65cajBGCXsyC5s/vk4h
MjvVldgo9gQxOHbkRkX2GtM5joKoMgiFOi6DJdSZ3aixbKkMXL3eDgl7atqGCKkr
3niOA7HPc8SdyI23n557Yd8iTW2hQVmkZhGHxI1XpPbPN+YhTurvG+gN/N8PXul7
96prbcgV0wcqd4/N13XRYLRpo7diKsKu+/rQCd8GkbqXylDj0MyTYVBp532dZmEb
Od+0UuSpcbRVTti9PguzqYqDDazvIQjtsiyMbC8iyVj47eWvpU2kLgamS7cME4Ja
yp4cFys61iUkkU7CCrZqnQ7uMp3U7ssEGhvIw7COcgQUeQ+X2ZXcqiVJKLN+/Hm4
x3Rlk566oBYoFsb/gcLD2U4Ge/n0MVlGDG0sXnC1t//yutqsq68oYx73SJXROcCM
QECWw/bl7x3v/8BqPogzB1T25G216oCnN0YjsXjWmPg5LcRu83HEtotAYIZ5A6xy
30JwwV9vWy0zM7MpHaoFvhNto9wxqMxUrjWgHB/DAG5YoaYJ4e1mLeqQutDI3PcJ
e9cB/69iDky9aUJnAfh3rsRe1IM8FY0+RTSkglicrNIUQT59q/gYeJ5ayhKlwuxC
7G69fXBoOp94xWlZ0J3BVUHuYXKhQG7gw8MQdrjbhy3XggNw/AKWpL3bNEt4GVZq
HyPln6/Db33pHKnsMo6W4vDzFo+LXR4cyrA4bPSsuLmH1eGnHGilyjA6g1RRXjlP
oL2PNWLbkalZ8YkpKlsc6yXwX3VQbxzRXxxRmS3iPDZwrt22B9Ob6C9V2pjpli9l
RejkIZ6UJBpO+YXedP5d7pA6Pz51iWw7P7L3Oe5Wa9INGdQJwZgvuOazr9bgCkXj
Du/fXz6X78XOHVUyD/XwrsT84vUh8jaCdEMLXCn7P577j7Cmo8LXyUvrFj8PkYd9
8mP80Wy1+MSCuECVDXWuxCRyCcHeBb7KkjviuSjfHrq2OMGlx1jTIbcUHazaYjNn
5t0Teh1jt2qJrCHdE2HuTaJqrEmm3GoqjCCSuYQzdODvDzb19tFLZJoL0wqqwd/n
x8NLKZHfkqypqKhiaWUkR4f1mQxuyDCrUM4wxaF8m5h0uqKrxFEaUOriGcN3kYKT
pNhzvjAjJGws0tEEU5sReD3ATUi+Bf7tS1gJqFZR8tRvBpKiO+NyTLU2DYScLxpD
T0CDoRN4NjrXoGHiNO1fW4mRZQMn+S7DNu2X0xogvDHnyvhPdFdDudmVQKR/oDq7
pOVaZ6PPoD/i/xRI2za6hsYAbgWBurFeACswSyyavywIUjkEvDmqZy9E+92sWviK
gal3jn+HgFAwCJjrnxLBz1W5ZURmjAfyiNYBQc3g5NUeQ0Rx7J2mgThoRg2iPX5k
XMn4DX1HYMSB7+6KQ+0laQ5geHyYRgsDkzgllLxF7MhhygC4CbjwXfqpbqPFybuz
u1Ezy8xTnBjMK3Exlb3v5bHFQRrHpKK+oQ43nO3HOs5Vczsl1PFWdxMQHji2U++3
F5oMtkXS1mWm8T5riLPQvBQ3si2DdruPNcCFoZTwRLkHqknl9/AWHT8s217+eaft
Sfcs2aCD62XLbSlSVwT3x6Rgs3/Atcqd6kRwV0/2AXvqOZYR92pZaDWf3XwDl9lv
6jhl1Nu/epX9eeivcy+Al4RVfLne+Y09W5cvtzXDKY85jUdMKG28e5dzdFd2oJor
V/lcZmFu3nYZAbd1D8yteGfm3vRwRmtot/QRefuHgWr2ucL/UpGrJgYXGPyEbccy
XavSREofdXak0d2Jh0FCvKVKlL7TJnavPwmgq/YTk3GMAM/QG64jlIX2TZRLbAhK
xbro5e+ov2+71BqK4VP7GdJ6PCdnCCnhjfWn84O2/moh/jtaHmwMNY8PzUjHmPsL
oHcfPIVCXhh5j6Rg12Cy7y57DwdtttKaj0bZ6qM4PWc5A6WU29CoVrrR9UQqyyi0
Z9BYxnQLlfgwk8KHKwH60AgT0Ts0rAAennRQGX+wDKXa1zjq3HLM/BvJQJiyKISa
gdGONRCLNT9V6TXbl3mUPQHm+ndpNmLmTXuPAA0FSIU+JCGoRUS+KLSnFdhfwTfZ
mTBI4k753kdD4eb1p2Q0ePzDoB7YWEQZBcGGk8VRUXsoHx93PPKMQ7U6xig6srV4
3puDAGX/oTe1VmZokvU1zAUfJdY1kQrbXOGdRhXcJmrbjfkVTYpPMb8OgpGjtC6e
yHlJaXcN+0ubcr3/4AuzXS9nYzaW7J9Q0I+m+fxmqSCpD0A4LeK/bK+yAfiZB1yR
isl57TiTTLkz0L5Y6LfXHmuCWTHvOeqCJ+kK+O0cOjRTFMDwvpRherP/9YAKPWke
jr9MyoTEKE3U3dThELo6tLbZBuaWCTZOFYzsSoAnffI5Kf4kiJy6pIBsNEa9dYGI
22yFnVaJj0iNPlRdNqOXoEkEHpwOCP9lH8RqU68D/NzRlxlo4G07vVqIGuBVi5DN
SiVDTwR+7lNTdKNqlW7uMClvHMIqflaK/KRWutNrMnNzxq+bD5tQgzCHYK1Npizl
Obi7X86zg3sYaIjWVFmLz/6Jvx1snx2TSVHRyfeQDXOaLinyF85n5h3jb+fzEFVc
W2To7YLmCzjxqQOOMgirnoia2WCSmePBwOBRC7wJwcZ1Xc/7CO1mlttpBnLumamP
btRAqJFvdjFuyOutkYvixelt0hb7DitA2DVK4xOj81mMD/yJYIK2NlXoetFnOTo6
DYGh6AHXLAsHyqV3fo9qD92uaGMl3meYE86zx+PqH3LR/902JfpI8/D4UgPvlSo+
utuwOOLfcLNxkapp1ADLldRaLvG7Rcr2jEM+bSHK/JL/xkDKdB8phH/aEtORbOnf
NYwifvt5AYfNg0mZBq3Lv39otZqwELKvVGS1GnTMasKSIPrxQKgk+cVxEVCrzUni
9zzqYI8Ad2AgVROFsk3or6RvoVLW9qY+GbuAzt/hTxLfXN5l+5aEsNHEeMEtOcQ5
XFqinbj2xwpO333i6T033fHaHtHQtEJB2Dz4nQjABJL2vjwTHusiyKsFkDWG9Chd
eYG2XJ9I3/f4Tszr4Xge31tKw/gu0VqVdVxfI5941vsS224e0ckuyj8Vv/+OBOl2
x0mRffac8mzTBJ/JSjuNkw4pRBuHA9Ug52WIcKYyX7wlvey5C2z3a8xDRtsFddm6
+assB6NryMK0FD1nwpbmWrVQUouSn2W9kAg6gIyYjWuzfRvzMc4CiuDxr9NvYsim
yrJ0QD8UI7+DVIsuXN5JEtidrO7lz7kQKJbONiJSCZtpm+akYvMkwp3S047FkzHd
wFMVV7AkwJaWW1Rl6v73QGTZcjqXbn4OEPpMGM2oJneC3MKzig57vAC0zEJ2fZQz
GG7H33FgZ8M6qcAHrEqKddLkyD2gu8gw09VTPyek7CzMh61K3ouSjcg/YSkUBaBV
kJpekgbB/zrv8yvAHjJuXo54r6g7auQHXTLDkHcet6pymqfrAnH15i0Zkuc+i+SU
kaisdWWU/ECpQ919r6czPYRhNgRAdUG8jJCQjEhqxj66CPLfaEzSDXOaDR6gwwzd
gC6ZDBIYhHi4ICLw8KyvgVqiQYbZCwGQFv6x2SRG8qta/FkIYG5LFiXPaK/cwl2g
Q2eKFmBeqe2fqT2+EUsIUzQoBroEQRa0wyPQX5E49l6ipRxLtEN71ZYTkxmI+IJQ
CegQ0gci9BHAd6JWm9P4VF8xRW0/X5Nw7f9aGuRxZ0ItkryEvJDL2GU4qAxVZrTt
bPGr20l7jrq27bi4C5/MR6+vS9RsGIzWWhFpxuc2SO2qIMJEsRlo9voXMgLhLyvz
eg8+e32KxGb8J1ZnD6b4q9IgOb9VVxhVlWKPZ51NNZpi/ACmMb4WkB+qFCvzxOV/
ERebL5yRZEvfdh430H46LaQRT2icbDwWUkP/0Zw3VZPBROfmADBOzYW+mNBKKbmb
S/TShpTxKJt4hC0GTghi3iAE+1VSr0xFVeszM8MqrjnE3Fj+KfYzPU1FDjAqce9n
rDDYmv4wZDit6bZbDXdR4sYeG6Xb3++BswgK3i1OFd3FaIII5simrmwAkYubARNE
UVASLZx5/RL1T91xZVYwbGiIpRIAHNCdrEBw//10DXf+Ik14FrYcFdJtcrhPRLnR
a5smoCFf709LYeEgh08GW/2hmHzRFsRVh6D+ssjaxdKnczCk0TnJDsSLan1F0MjF
Ba4FJCHrToSiRu+9HkYjaJ2hXuiur540j3La8EtVmJushyEuujcaCxsYmYMYFYSe
YjT9diHQbwJP8ZQg1wfjX96f5qTmWMvL1Ty7PEbFFYEJWMT087XwpBVob332+9iF
pl2dezxZAKiNXOAafdzrF8lq8yxUy7v7LdO6OmPngXZ13jv2mockcsW+541eMfYa
8tpLocN/KGlDP+PlkxkuSjKFrj2qZF5W9P9yPEFgB20HOQr6NljIlNfn1KjSnYWJ
ZK9KegOmoRAVGOOVpuI7eFVFz5hwFOXluhanyYBu43wLdFYeNZr1TuryFCVzhui3
rWGNslJbVTdbhU+ruLaNAMAtl29eUtogm1S0uCmzDgKyRKgyFEQOK89Q9ao3kHRa
O/IrgqzDp7UbRKexKuOraWGkp5ajBGMK8xF0S6djCGCSnk3dkZRkRzv0zNsonYDO
nVvuKN8HqtZhtfr8QgM7rVceyOlOvvYYMB/fD31bxfLnvGcNV31jwfYh7HI1eN3c
wNPR8sgzkLK/6szfuV8GnrycIyPz/vcWXwYY32NllEFALHbcEEiKi6CcypQ6/K9i
Ofc2eHjfniUWufIu0CBXdSsBnRbQRN8Bh28Z3pTeiCBXibD1tjq7E+AHVEBU8dTp
GtT369pLvsT47bQ7caitjIUIHroZ7GYsn1VKV52pE+TCwqF2Mu1JcjvrAxIWZA8Q
jb0pnH1FLIXm/97w0rqGY2bMBc4I8wvnoZm5VM6Nrql2j3Xm64cO6wWKAIZPSHgw
cgmuZ1n0CbRf0ng+hXaO01Uwm2p/GgazCT8+9z6WzvYRm/TaZ4k01HLTtek4sW6r
fhF5DxhW9HwefDetL7RgG1TPj5eORfYIX0x3hzsi/7VzDA4XhrnQ5HwOnian7z2Q
EFmbwwqw4yJWRfYhyBZOoo9hk3eVCF+0+95O7n3AInL/OrfI33ZovMQ7XguiDgkT
iZfjGeq2xOXRx+ONK3g9Zp/dUz0wa4vvGVVR5COuicbRFk/kGCxxywBw3UZHI38P
lZnfLM7tcgPiD5N8MsDs5kqOYodSD1rAYwv2TcyTw6CTrMD5EfneCtoT95brupuj
1AZhP5aNsGyyEI+5Ek8fnJkfEs2LgES2SHlqtegt/s8k7HVQl8O2i/xdz9NbF4zM
D27RIBCCVOJ/67ROcIBwoe2j5OUPROuiLYGxjg+fIqL2ys4cWvj6LzBtwx+BX+dB
DGWV6orRTvJB0FcPbvYTAS6SGEy4UZUHVpyO84abBtRPJM+//Mtg6vZv0mBWhzZs
WOVZH8pdPr9xJubQTBdMpLF0fxenU3HrYUJZ5Lw1d5V3h987JDSfv4fXKuyxBPr7
5zc61Mj+6SPvOkMkBEyOIFCPwQAJyxOJ/NqNdzR4n+fPcIIrpPP/DDE8Xh26vKCt
4suy358cxwAis4aPpC7Vh/Y5YIA8dHr42XJme6f0E8afu6c8syY8ObvwY4kdIMZE
8TfumBj9e8fMOaq/B4Td2jbI6Gi9vX1P98rETTm5e45L3RbDo1vOfsiP+EgJFW1C
0IMLcFndv53TU4DwezvXaNG4tZWxjgiXodETH7N34LPbIS9XtqAi+Rqrcct6gjN+
1y4dN+QplQRl+0UbDKDtdL9b6CXMZITfnsj9G1uficaxC9PI1I94RE8DooBND+qz
yyNGtAJ8hv/zf7qoM1R+e0Teuc+Stuo+0FrkvpDiCvN1zDmsWKm0Cy5BF4o/zpeC
xPRfo/bLWWuwC5mQJBEPVv1XYiLEsoUEmrGeEVtlIwlH7+nWqGh7MGwereaYeEmT
yuNAUouP60qfAs0LBD+wmYGM2EsgBWhMuXyFBYnoGbQoWh4j0QXfbUDQsikjII0i
r/Y4hgb9mhU1YpVXSwgO9L6MJgfIrDG4CoFpDm2X1TkHt1Mp0Ju3fbPrIK2uwSbm
hjpAIlZSv+yr2r6t5DegANF0KXOOf47cyVQF/XU8aKlKgc1mtdiuE7vm+csHzpwD
eN3uz+dhmbWXR0x0I5zcGP42LVTzRBEQz0V2WenWxn9ddR8SWRaLenwSzpizIIOo
zhZxO7wk97sdPmd1ZSB+/1qXA3i3QgmwNTdDkUKw38hkihkmX9wvfP/V3y0UiIrp
2JHistnrOXowjlPa+KL051Odg2Y7hz7h9eR+W/gISxiGQat6OzBbn5KW/QlMjIHp
oDYR8ESiEWOlnbsFSg2gelYGgBqBCaSRgwPY9w8biDGH7UKZjhVJByoZoGEVVoB5
B5mBQ6yCUIzuOYsYAdp+GhNMwYRZfvvXj5dCsMZdp7c71Oy0MZ+q1tCeaa2/Ht6e
mu0L+EB/gIpGhFUQSO91l+7+yhHvHzarSbC2xFovr6uj1HoYGrYvnOKPVnt9f8qU
I02cBIDq1DTkLoQMkm/oMF1pJGcxanL6Y1wFmvAwA2ybXoyl2m17CttsZrDKOoWX
Agan59wNkfE01qHwNssFKRtY83sIBwmKz2Hosa1VszElf255mOXl9S0OwxGrGAeb
dkd7aVE290xwQRdv4KKaXW2ElK75TZ5m7EzaIyP4/zV5uWo5OYhoXvFiV0b1FN00
QP4Em+RikTbI4xMDhhzjlO1BQ0AhZFixanNrlQrNct4qKRMNe7aUn2hVjOa/HMRB
u+u/Er0LDmB70bx3sMVgNIzehcz70dH13S4pI7xpccLFqwb/xucghWpk1eutOsB4
NMpNGgCcFFkHuhRibTw8yYzyQT0a9hBjcOjZXpD7GlS4tewEqNuXvM6T6uIKFsUv
3gwDpp9NNEFukA9Vwk5EUbdwk5YKqQJivvTq62SegP5/pdNOuPHu4leEKtLI4yf8
YDpMZdjAs9rUc3jSNxxzOMAiTN+66q9Yr1hBj0zc0OD1dQIVXbcsiJoGzJLN5sGV
ONgwP8Ga4p2bsaYdnJHPKyK1yIrR4IndYowPyMlmuEULQrNGIkiwJ7CDKy2AUNbZ
EspAI3GAmjlcHbZgk3sYSRdOfzkekb0v6AvzTJNmow4fPiWXyP4nMTa5Lyg+qLdc
yxVNEvz6b5ikFAEuXjqrwKlyhVFRJxNPRh9FXh/2qDDRFhf1l8zr7r58VUIlBr8W
oN6lpL97Q8XAjsLbyEfjyliSr1QD5xOrODedlJJKlBl5eDWSG8bI/mFxi7NjrkC3
u+U392PtxMae/dwoALjnm5Az69EWtmqVtf6X2rjURoJm4xzKp1d+wWd9kEO94KaW
QQRqdxmtSa4gak2PHDJLRWqSLLBLNTtOWYBoZ8ty/uDdV5G5EepRoCrZCOgPNTWN
vvoeU8f+dvWS0E9WbMXPQ4lUykFJmW/Jl9qVH6GjECwXS4czA+SvQR/+N6R0s0VO
UPqCcQzLXQhsn5FZFzIgmp1gh9Im4c04KJ7zowcOq/5eRTRj96UpEKuLoG/uiLeJ
xc3x/bakptppYTPDo40VTGu1C4skI9LTeaY9jCWOU39zmBrpCrZ8o7hbteNhkmXL
B3dBDrac6qdkolM8f8QnIvMSwk4WmD5oksJNm830j4q8FYLgi8+Q0gFbLUZFjl8i
qZeEzrIad0TFU3SLDTV3KyCfFc5p5gFACGPTQQwUjiDCwczVd5M5gTJ4qVUVKUpi
XC3aE97NziKyC5FA3FFmM6eRUANqKVwwmqHiXCUIffeS8UV/ML/Fh6X3D1oeuUQo
cyUhfqWNhYKZ67yiHp4IiGh2002CdhDxXzC/Gs1eQ6yj9tIwdQUuvv2Zv1DJ15q3
1q1/O+LtdeilF70fKECX4N2NKPHjSE+c+vSvDl5wByXpT3GG9DIzZIC1Ibw/myUa
TGDTYjQk4WuUwqshJiSuCQW7yAff/SH9UtVhdA268pAE9sSVXRMjW2/bOy6TzGwa
g+qH4tESRoccsmkYVDAeTgKAsFn3IgbQxH3+bd8fcPp9/ynk6iXwp3KTxdG8JIfV
EqJvYbf4oWUwge0BlOXHGA3QuXeHlyypqG6YNqWtJAhfB5PFX13Q0U2bD/xPQAu3
o/YPbgrXNC27OFAF9FCtKKPv5CwuMk6XF5LTwtAguT3IWd7wCnQwU6fRWpTFgiXn
MTx4p/tUEjmwnoikTtWLU2sTlJzNsxtEKmDKx8Uy5DVj6AzJFKBorbUCqJDeI3BB
i5oXPcB4RIJHh1PupCDKsvLQmzGYe+Cs873Ts3JKdVtiXsl/Vp+gZa5EJFrsWz/i
HAXCI9RZr0do/Scz/6kkeyKN5CBVmGJ8NPWbl5S2YBA5juA5XYDth863T5/H4p3C
qWWf7d/CSRP4+v9dE+V3a6vfxBvqZ0NACEhhSnAhxd3l+ku6xiM65TqkQTATCaoE
8t0t2HSv2E8HRctJiy0XwhLTEqcC7nmdrtM/VFZYnoinOKfX4PDwD+mD/oDbardl
4k6dIn19ZxpwFPmSbLkdJxLEPQzA5UBHKf/uC7WHE71oTbNkKHN8kKr01Qoz5Sbc
2nkxORCIbuYFi4z7ZDwbnkcyDWYYiMknadX+BfIGQoLe8IAnGMY4g/AIoQnvD792
O/kPasLdCOROJWZnTvChzEypIXWgt/a9mU7cmyKRAwOIVsfuN4Iavx04tsd+8n44
mZtTzzUsMrEC4VlJOU0l5OIY5qA/vHnmGbIlt+B/vveh8KGgouN6Bm1mmHl3Yiuj
vOyCuNSwW+hywNnvbMXjttqLgjq+dQB0XAKEXlme3sEU9G5uBxBboRIZ+2beT/r+
7R+J2YnWxg1Sndt0zKD8C6jMKh+sJtHBQ4aBo3DWkRY8/Mq3UZMe0jhbw/q1gcCW
BdSmiVkUMWC35KFHogEIOhkAtmpVocHHluYTj/7ba/hE+XUC5uyVeHCap2n+gGsk
NRLQmtA13Jk8s2iE6xGPlWArNHmhfD2OFd3T4Zf02c100tOQYmDLe7i02usr0Frh
Jh10qZ1xU4bfAqLcALobcMRjWDW3lp2IEujbvJfaaJHRrvKBnQhfY9Ov/+FQZ34X
sW1rPB0+9PnUj3lKaFEZoPXZAYztmfj6bmc6faQ57VacJU1MNDwva/r4fVkBE9Wg
OOM86jr5HqGvyHrJ52d5o28pxJZAryGF55I1IJUSDo95PJQ/myGUhu6sXZ0DQOKv
eXoKZaiaNg7DhZOZ6/x3Od35safRnIAhXutBXdGjOqsaV5s3jdevDJ4vjpxWlZYJ
X11hp6Zfrj8xBRN2raNveWMcL+K7QvzcWEktKiT/8oFEwVDt7Gu/+xb4ekMwViQY
vnnKD/noSDFXcFGOFQwaLMLoGW/sNbkyfyG0X84HcJi0+JBv4v/setbqB0xiORka
99phYOI1XQk1YMDACCcpGxNNREsBmj4x8T1SxLlZ8y2VRtbOp1OJN++ysPa33+Vs
A66kl7xOh987fFLIBgPNKy6DHYrJRtnltzKdQMKmMy1jPRmbUcT7qRcI19HJ/7eu
nRcyx8pKw6ikypOWf1+zfrB1Jb/grQgGCCxxnPgDWK0jV2ndB9UwU+gJIcHGc26u
mqBgIsdIBseyLpPFdtwWQJIYRwGNUYTzuwAtCW8AGjABK+LFxIaV22rPLnEQVT4e
7kmuWeV/Xu0QVTnJ/UVejMqsA8cKcqve9eLVxDu2EcQxwkjgXNX9gxrZ9/Wzes1i
2BCEwYNYLkXm7sx6VMgq44kye+LZnnt0/Yvrn+fr/YfXi8l/ynA5XVvxx+5nvYv+
ucB6fGzjg8CD9FpkIf5tIwJP9j6PAwmUReXnjM6b9j+gcJRqQX6CTB9AvFz1+P3G
YGBEbvDD888LYQMsWlp68hEmypJnJXopUJhML/hg7tmSgEAD4uBxarv/5zasiXrO
ZGq1V2fNgCjfaYAO8VhJTKhZcmwsmXUMhq1XkaIHtXK9K1IhjK7hlGPmNcyY98Nk
UvnYhm0tjimBNTiToIyXUJYyH2GtHbKY08lqAkwffw6zSg0fpE6X2jq8lap3/7+/
alTBTXiSKFkTVwVj+P7bwzGMLrO10aWkHOBD/Nwj/ElhCFtV3gBRStMSS0in4utx
h1PlBpiHewDwAy9nBVv679gXVzdpTWkk7g/1HPEaC3I6ufeKhyiRWX7mAbWl1xdD
CkaAGSaMXubc7A+ilADMD6A6jdX7fMeg4CjproCtNe+X2S9JJlfaND80QuHQIMDL
Ace2+OG73BBq0nMwppL4J6BDUqEaCxlb0wAMR4IfkS7xgB2eWjW1nW59aYXKa0n9
Ein9WdOz7348DdHCHTfzfD267Z3J11V+ifUB1K8MEEB3viZZe/GEoOvbNZQUxwXJ
Lsu0kNqgnLCGG0A6FqtyiSQUd3iyXCOY24IXX50kD5RkMNb4rEeHStgJnpJV89Xb
VcuAHHfmeapbdNEU5Zjp4A8zeJjkdbALHJ8+Zl7KWhfq3J9doioOyF3nRNrXuRLs
uxYYIDXyG8qzOTOlymtm9+JPPmWGg0urEnSgbYD7tfLE8wq5v+U3nWg8UZl9fqXD
JlfsFVGp6JlyRn2LJr3u3qLotrHAPk8v6xBtgyfm1ddA87fmcipxq8G8Y15J9fop
c8Je7KLLFeGnLGnh7DPnQ2mvdwIcl6EOnHnZJEJE0WBNRXHIIH9FOeRX7SgFFhZP
2ETV6Mpovp3OS/Z7vugDVBs60DpJLRAoCBJQAiuVFCIoVwStxrxuh2C27M5jlJxK
KikBm7P3Bu5b0BWzV/3lImpD3AfoFiZ/SnUq557iUzTc9fcDbP9tjcJACgFIC9Jj
CqTFsc98t/Ft6oKRDYTv841rEcFUD6fXrcqtt3XUxrAl6HSf3KuEJj4lCwbN/Uf9
TZxp72Lh9+LiAq5KD8/VJlDxTpUGbjthUlqm6LgemvLES7zA84O45KkU759biwKE
XA0tVskS7+ujhSYrRhQUUg6SEaxvoSajIuBJh4RJNuFlsIqwQW9JYdKUG3tTZCjP
wzWNgb0Di5YxQhGDNQ3tgOGE1RHcGkM6hGolG9HxC3Qvmsam4ow9yOFVBZCo6FNX
S0z+Vo1hhg8+Mk4IFy/WWHtOycAqXusiip2bpG5/ZVWMZdtRiUFC7rqvAEYCLNqs
UPTJmZOg8GK2N7dU6eo4mTc1ZsbYBdnuk4wHKpRj6h4SFZNYC/Zq5EXsMYX00RGk
c6VN7w/8mLGBxfoWwRL4U0uNfTEet0T3uiCGKEaQ/4JZ18N7Bqhbhdk4T9x+dY51
dQdM36j7fGEQs8Z/tF7SMJprL1emopn982N2HV8rWJmDLKGYTvU0NcbYfVm59r3S
HIoTLPnRXonNvVsUxc0wdEr+MLeMfEFzayrgfKiYFlRoZ07PjrYvuMZsZhqSjs3k
kWkEKWyomxPtg74EY6ZhicDM5ZpANa3FndHFpd3dYWkoOiAx5U6BAwdc6adWClRi
/5+u8LSI3iNKtC4Qg/2xbTidqOeIgxK58/hntBLHnxFVNJx4d2mntdXhLryaa7Yn
D+PLPVkPa/L4eaEzRzC/Tuhp+ktZeCEt0Ki1yvggQMMgXC1olOHCXVGf2E8dgVpv
H1EjC/y1qAyOcHXYAwirrejNpgbUS5U3BZ1LnBO2CluGZe/djKxwAS1gRwDTmWGS
Xl+j79hCX2VGLe360t/g+h7t+VK/4CI0cluoiqRJDpN+gZxcVL6vs8XD04br4qUf
YHH44wuNKgtwc/JflvZzOJchmBdxe3bTMBRw0qb0RU8b20zRm18HFK1fBaiBmLWd
GLFF7gVmP1CD0E/xk5iNvcz+O5VlfoTobwF+zs6I5fmRYZC4+pL8tOZ+2y8Oozj+
p1t8fsBr+Qv+lEfpWxfNcUhXiwfFpYW2OrNa1T0iYqoi2uSxSg9Z4yRsKb/YPTnk
mq1aQQlGgdDIkqgyL4EvKBY5Wiazu359+YE29+90wR84ptCUUG6yOBSIGR0X5gep
R4ZxkBcFhYxI2n4HMLfVPtQcATsEIcSvMDBTCN1lTW5p/WGhPP0JqphLIr0adT1t
Jl66I0lPg9Fv1TlufbVfVlaZPbdNbsUMSyUz4DlBtIcMF99OCYsn669Bm5i/sysN
IVSlPXUZ8uSR2FUmpnnZRrCdNV8pUIKUgSsOShC7NqgR9tLhe/8TFi/azXYt22gv
Qjv3JN9l4IWFzeUzyVIVZBx2zxaddJBa69GoAvjVIYKfzz6UMIncdTuCslvzmWQb
ElL3uMDDRyGwFYkKl4YCFZJ1lPNViZFdGPbuJ6zy5fYRSm6MvTCF5BGI4aWHYqme
JECnro0065XQP3eIuwQUrEZorBkny5fVvzNppSj66tXZZw+GFr/O03CInmEh/vtQ
KX/SltzGBz88zdPdu7DLLIkMASFJUu5q/R3Z3669+xqD16vLSOUvYEhaO/piLj1/
ApWopbRqeoCeroXaR8lYaVtuTaVwRnTHorCoqdz5dpCRkDAgKVEsolT7QPOjrmyN
7E25/A8aEYbcmFTaDftV0WNcAf0stODKFiOlacAXQP6Cx62jFlf3AgaFgbud2Q+I
M3syZMys8OeoVZUEOVUpDAkElZH0VP8gQalNBUp59UbSb+WhDFjpW/q4jZRUCIGi
k/J8BBtTSTxAgNE4lAclC0sMLWrI2THvQgjxb/rpnZbXdRDnalSP2/puM1Idthxu
9rVOqTzUo4TnipHjZKGnwsP9nIxN7ZbiH0f4CM66r02fXuNBqsC3kVv77Duhzrwf
coZWTTWoUpo5kEAtcrdScN4GNVb1c07B2rzK2puZYvE3H1il3ptmgrcX/KNza2rn
K12WTs+00f3lbGhE0s/77MHoynVD6DDa9MtK7JeC1Y5G5Ir1TKJkJvU0kZmgfn/L
V7XLjdvj3iQQAl65wLotp6fK3Szsq3wfpl5IO7ktovdJ0qDpz9BBrZLOpGzWrO20
YU2C5CGTDQGeMitjsVqU7TlGHmBD4rrAE419oVRQlC4iOMz8egKuZAwvOKogjnAA
ZS0r4Hyq8nEzMlxT6AJqk3c7XC+GUfTXJ1/Hrvvn1AM9doG2L9ziuFnIHn+CIfEJ
2Mr4/S0eqC4pNcFk+5VmgBPRnXAkMyyEJt/Ej+CTrkJOgg0R///t49JUXEpqewy1
EL4soJ6FvxmXwTivUdjjxiwAstE3CrInzhiIwJhf8iSw+gpFEdy9+MzHWdzyFYgX
ayapTiYIXj6nnjd9Bn36F64DpVLRlogog3eI22ToleCOfesMRCPqKEjVZmFF9dZ/
bI4OTZMg7VYZ/gbfdcxehL453QvMKOM4Z081MdmW93xtFoK1cW23A3RDuLhUXFms
a7+k0o6rQtcniQRCd0YP2/kmcfrrjkolAQKZ63g+CfIMQvJdDLIBl6yRQK87/UW8
OsEQIkW4iIgOFLZUf8Jgq4hPPU5VGH8wAi+BIS67rD+NkJHCTWVi6E4iliZ+IN42
RLIzdkNnt6mpXgVZb0jpTdLfODVD0F2A25b/dkbD07JaaxtGRkNYnZQB75KOAmYL
0Yr4b2lvLOxtLDLqkJEu/w7xM96ZLatJrHBJbEYUIiWtrle3lbpraW6zGKg9rYp5
fd3eGQaVrTSVrTQwPZ8MZz/nsxjaa/a4vEnmQgU2FAoHY0LDBhNuC6Zk0WKcHJYv
lOUtZo6cgmrPUNcxOv+nFbt6ucC5U3izRT8HgGD4eb92rVLuJ0iaTylyszHQXvVG
GESzjkJbNgJqUgvNfp+UAbZhFwYcdQCdZCml6VSgO5gOoPFwR1bKasm9fuaLsKzj
KLstqbbaMMQCxA2yeB0qedx5Dx+zZuqfl6/el40fGhShW9g1DtVUsJAOG/oR1Xzs
0sOmU/eY9oLWPBSmCQZjXpBdA8TqbhLBULL0YrNMtNh4EHQyxvJsZYyheFgDCBPw
a3z/RM7c3ebdZ2YA13fB6eF0xAhDSYWNkPHSXnWBSr+NH3VPYpX+FOmvfMDZjK/j
ncq9qcxKVkbuY0zoQ0k39jqfJkNSsr2hbL1yLqygWYJPgWRFEf9CF3XQvD4vnu/O
HEAh77YHJ0kS0E8ZYCsa2/KT8k7Lf5q3qqNwnaCRdqEdkDscIXWSALcarikuhxWq
vJkzZU/Jh0OqNjyy6Xhtgd0Im3hKFWhdFpcRNN2N7YLPfEI9F6L+tOxigO4WGJFp
z+muQzl0eb2yi4rsDFKgdXDlPI+Y0+0lqmrJpq0bkcP9FYM3VAAjIziAVdcGyg35
bqxY80OST0MGkP9s6Yew1KlBQcLZVS5o+aRxs1jA4f6KG66TUWuB36hrCDg1Yd1Y
ufckWrYgvqesvU6pD5IcPI+9cH0jyZYXaDe6JJhASrtLmzJdlxlUMnbamX9/D04z
QVa6hHVAzC48rMe2fzODLbOXJ7ZF/V2lPem5cz63LDb/vZ7t90iw/YYtLRlyxdNp
8l+zT3lJ9w6sA8SipI6M+7haU+3lKa4EVXwhyjjcRiIiUm8hi6P6Tg4XFyM+Jkki
5C7+6L9Sc+zRrkBPJ+0RmyyImIzxpjmSYZNccUifS5egb0xL5/EVIBwtMVfaplkP
SMP9Tw9kKf9uYH3lsiYED+e0uQt1aakTXb71VWXMntfHSC0ktEoeWJGQGxkYJLdD
TayThWPyYSDLQdi7T5hskJG9fafwwm0ctHIlhv8bbJ7l/noH6mfcQA1yu3SJ2S6/
ViQDuEn3fUJ0qkWdmp7L7mFjwTwISrCuApwrKjpXJrSMhpKIMgBf8uH3bzgUUUbH
/tWvl4A5nVteojSCGeQNXGR09OZkh49E2Dh6ikpFRiwbeoHX8gNaKBFqVnheJb45
Ygd6GRNtMCv+cqK9JLPwdzv/9TUKBdddLY4cNleG2q9kOlhoioKXJDpl/WyE/Qao
LPElGpfIl08C0oeb/YdUtWhUxMCgrLi+7FAMLzd6ZAzI7rpz7u7JiO0/toDkpQR8
s2ATgQRoTmHwMFYHBW5Gi88wmCYFF7m5S/WuVR0/OH5o14aFRxtqufHEug+9yh4G
WPReTnsUuALEcujMaHgSKWKyLj5vA60YpT8GN/iRLVbQxp5/fcLVKf8WznxLFGE/
adxUn4NkZtiox2ftLzfGWDjCm+4cWi8tgM/o65p0NZfTkONFBIM6eWWwFJC3BOqg
oyFvkCc0pC62FTHUTGTobXVDa3+9mZ1tGHG29rcbGOrAaS+pQ5AtGT7kGhAXILXy
vWQS/7ke82/ALV2TywN0jteUmqdP5W7g5eXDPQw83fZApWRXK307NYTb9TFnbYmr
4t6NIilGsDlod0En/kOW13tFEDDVfsXoAbudyCYKhQAqg/m/49ucuR16gPlO4gW8
4dV6tichJdxajPN9uvvbZHZ8mc+3xIT86SoGuJKfoVktnw41TvOalzzczsgU3mrY
Ub9idObYn/8DnVxpkZNmOhcyzTKekwAyyC01e2YIO9icVnO+nMTf2COZV809t2xc
ve6w9mKYSdGugLi+cErj22a5VAU4s8sHjTyxTLjpX2fTw31DJ5lEbA9RNh6255cH
V/zkl1q7cBmuYQoYWhmP5GFI3Oc8xDpZf11uOlVdtHjnMwFJYb+wsUw4S7XWRGvI
aFFt18V2ojip8l9z+tzDgGirO8bSpiY7sV4o46+O1Jd8exU/znDSJjhfwgO5X/ny
gZRlBhvgO83Om2C55WLDk/CDDAlPiwtuH20blwTIUk+BmLNS+K1JcTZ1H0akBufn
R85VbJdEd7dgw3STmuvSL1RKj4th2ZzeCtKMC1hDxvLNwvz7g5PfNEU+jfkzfxT+
E60oh2qDgUZbi7WpM9hHWq43vd0iFEE0i8vf9jiNj6w6aSelxrsluzSe0g5xX4PM
mSdHQoJ7TO5wcJnRmSMZBDRJf2hPG1E1ylrZEX7ttiub//EDV/kwp5cYYYYdz/ex
zNxlyn4pXcjmJRhMI9QJhyO/I6q/pX33xcjoQw7Mdk5jGHMqdL9ik2f8ltpB0VHy
+iSDzcZq0bYSAD7jYe+ioX7opx6+Xrw5QyDv/y+Z6g9jHGYM8AZZyA9/IhOtbwNd
h6NzQvaj7fO8/kf2THywumqjHWIFDasjypFXS2bVjUskDzzoDh9HxE7T4VGHTnLA
7zVde+u2Pwzy/Bf9TndzDWPsXif/AqkhLI9R0Fm2oVb0OsxOr3JpnQ28Bxdk85YP
F63RLY2CFz/DdUK4c34bBKuSQe/J5Rpg2IZFY9JPO8KogbLB2d1qrSevTFByJBul
vIDdLdi/4BlNGASXSpmpPWpyI3Ed439l8gKkfCbyQ6WMdpB+Fi0G7EVMNZqzR2au
zfjhWmRAK62msIOMC9PVEysACOGYxaRh8hrxWsnOLm998Ymp9oGtbXURZvOZBpmX
ftxdlzuo2EPDe2PqdMszd9JxMJvriTgzg5gIfksKBvh1F+zAcRZijl8JaAkHXRrq
kLsKLFP2NYhNsgnVBv6EEFcBgDLZJABC0nw2OdYOn4M74ErhZdvOkQ9eJEcv4RZ7
TdEoVrgQsKLHrx32BjRJDw5fPewa/dg7+nAdb0nwfgeolRtfdMUblVtveowyVRAE
kxI9QK9Z4edhTaX/hjXFcDJ5v4bfRXI4ZkUr4LRICEsn7qjSL8a3BIsvEjKBJFt1
Nm12SzsGn3P+hPPs6Z/FD820MnR8Q43aLmJqX1X4mZGgqBPOFeIE9Bb9rXQhyRlX
c5K2Awh0FWbmjFJZSvdbX+0Kt10wiCDG8Tb/G/NML9Q+9WH+fPgLa4rY7fowFiKI
6r4NL84afDcXeLxzHYr4QsLIhL2C47Ypz0CHHIX5em7LdSWBIpYJMs6HZGKyNVrb
MQCy/UE2W3RLTNL39LI0+JiXRgYUnXQE65EujzuxsVroWd8wlrU3OHO2oxmiMee/
/vTm3seIVDbVz8ik3Zhjs/ZBiM7LSIAMct73OW9clBh9nqa+bp3ybXZfL3ufypOd
bCIb9/9TpOy2kEkNDM3F+n60xB0+4dZGG9HQb1S2PDCQyrUrfDqHGfXqwkESFYXN
9/D+w5ab8uvcw883hXWTypRIkmK+hocxovYWGkqbM+IfKibTv6+Hwu9GlonC7p6F
LkzLbhWj5QveXpQNEzsyWc4ZAfG6WFSYdzZwOR7wfKAF5CTTbrQ+iXmKGfKuTRBb
ULUAqTFf6v0KhQf9DRMX75S5bZ5nfd6TRpWI55HUUb0poapUXleCLvY0Dcj49AQ9
ZOQx3ufQfFpi+wdabgUcYAKsQ6k9HJnsh6rwtMB8oIgxOHyYTNJBkIoxwyk2vlnK
7wAx7C8P9UPlXL4tBSOZ9mOLR7Ld3FBuP0DU7lgHz/6wcA2Fuiwr1v7oVqsLdXnP
WjsCAsePFkTU2TQjExLFYuPv7Qg63YMAeKTpCKp5vJQF8LMx0zYitnkfVZY39a6y
l7h+lbQ8WrbEmeV8/D2QOAl7vCKOQXg/9pHjY541hYdSv8eFfbFQ+r97nU4WYL0p
+3tOayKgrHDyBK+Mcu0dZyTMmNzFbzsjwURrYLsRHP+df7UTFG5yiv/bpcQujP7s
ywZ2vxGSMav2zOMmjMPl6p34lZW5z+FHosg/MmX45taS1B3YTPUZFvY8vItjlzkr
Z7u/uti6eSGTYa9faLjgT9TfeROIng9VDVXDTqDaLePKJCzlB2totXxagfwtoSSE
OdEQzo833Vu4WprrA4Uz7rh12+7zAxSdCXF3oGBO3zqLWRT4rmjsi/I/pUxWWOGh
paQ9OhA9E0L/zt2FTA4HjX/a75rcGs6QuwW0wtIy6eKfcZs0ij7bm0ptZXuYe76b
wGoohvdCGsROLLJQJPOO6W6djkdyeDIvFlQNunZNpkmSh2m2k2ZPlN/Fb+NgfRJ4
GjqdsvU8OQQ2HkufHAH66uomM4tFooA8RPRRFmKr2GgEkcPv56nykgnhUOF11PAR
VaQ1+d9hN8mo5inqRlW3n2N6LybhF+Wkasf5PXtfNhJmdzdlrsmJR3sVOnZUeB5R
3i9ZutcTnfJEM63zFH+gtp1nDq4rq31gNjVFEpsO6bjY4Exw6pDa3OTUx5THf7WY
LiXlsr0adJfv1kW4akn+cltCMtB6b0sdPYm7PnTzE7wk6e9pXknrYBn7kB2VXqrw
2W5x72yQkm2ILm7D613qoFRGf9hkz7+v0v8CWJLT1r03fTMEzoTF6oQtyvQ8EjtY
zid1+MGIJCLNU5mUrRnD1BX8JW3awFDEm8/EBm9dBYcUxwNbWP9J+LIFO61q7TVv
//FpTI56d+AJ60N05Ivu6bCaj4gR+hMu1cFPKKclJE0qzsjEcBq3+RUe9FZFuSsj
HpLemApN85KJFK6n31+9INadHr3nHJ8Xkwf6UPKidditjaAFEt61h4KyQYgubZlQ
Ak2z9U3P5puOMhNgvDfNgpp0TZJtD4474ttyReHq16OLOViAnkKEZpenRF3G79sz
5xiO+jvebPsg2dYrA/w9WZNapNGIQlKKQLhRAuBXDdke1wc9WU2h29ExrD09+ek5
/pobA2VsLx6zOlVXZGDOly3pDmlhQgktF66QgcooKWjmBj4DOPirU1JMDJlmj0tv
GM+FXrW1HDmLXt5IMotTDUnV+wE9oodoObA2O3kdeau7Sk3q7sWbkpTVf5h/R9dw
SRqgFjdO27+GZ7FAYW/+vc7VnQJ9tRDC1i3dudAQMEqlP/J+neuk7S5/KvzYJcXL
jngXu/69R57wLi5cTqflSFm5IrxzRCqNfAHocLVPsZryKIDoE9jASJRlLzDn9r7I
Gp3pfZCgLDyCC+BG9e/mygrI7NVoHxZA5DIyegDGFyvXCXvlo+ohPZD3QuoiJD4K
AZpRmPwXS0PCCblyAtXd+kqT4dT/27UFo7e14N6LxCVgnBS/c/jhzdS+81gQzX9c
ThBnKa0w9pmuOfobXeAxkptVSMy96hYQ3nLMlkSSQjmYK/i0lHqEVEkEnKbt7QiA
ZGDXgEbPPy5CByKt7uPe2qbo5PmW+t85hRX+adln6OyE57Ahi0iAKiI/9IzNqpFh
HdsO+DrgrlureY6C2nGnTrFmOYHziNV/VGZKhrw5N8BtspyJDEyzIkyhYKMqBQJK
7R/Orbt1X2tPSS5gXiAd1W8DkVvtwutOP5glBRrnK/SIwCLZdzzVtMRbgPhu6mqk
`protect END_PROTECTED