-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
miK6e3aYCZG/3cqIDwNP9UsYx0jwTuVSDzM6woPJ+cZWl8Co54SjUSOapCuFqzuy
JneQK+ZBeQvXFsFLY5SvhX4kLf3ovh6j6QCZCvHT23LZ9duB0ivtO44PtUa3sQ2k
ZzDWYQI82R2gfWGJbbjpBQBKqlpRa9PRncI0bJrQeAI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6029)

`protect DATA_BLOCK
1a/i+edEj1duIdxvuPQ+dHLPDOk8lSZvuCVriNwcbxJuAaE0WO/1VghPNwPq7qb8
nSzLS23bFzBgkHghU7gOsJtQQCUX44oJewdoARAk70taJ/ao3foKRbt0lZzz1iXn
8kxWXSQ24HVreocy/u8kEE5GhzIu0hfoENgS6j61ZgpG7gyD8mWg7HcBCXKB7zxn
2B5yvz1z6ZX1cYRSDuK3XuCfbpFwH+VHzz1OhYwK2v+eB5vF49wVyWOYXu6ygdIj
GNn6tsTCzzTkyKuxJBDltdcxHj/lEyQnCi2ctHUy8Br9fwSNOGFzPxmSIVTk1oc0
56bMvuhvqGj/+PhReR7L1ttlO6FUJoYUYuZj+19xuDHbOz9woPAqxmo/J8mXq8ix
VY1/3fqmgjrz4Ksgy87DZmbNgnIM+mPBi2SDvna+8HhctuRYwe0BXrZ1gQJfPxv9
bYd9CWqsA3rrGaQebE61VdIB+dOUhcNAo+CHopIlmPXkog5cD7onQnbfI5qsJTqc
FnW6fb/rCY3GpmNCiXsFtMXm/NYyxmE6DUGZ/mHbUWMW7VGPcm5EpXoBnv3DZedL
YG2MRxS/bNAbIplgCpGIZLLJEtgPNxqwPZT7WtFPj90LSt97hBw5vTenw6jd6Sbh
v84SaWXqwDRA6wtdiUNK7NEwGbnl328BjN3unHr9HkSJLLPdia429WJTHrzeCp7X
l5g2ndpjuicWPsnIF1kkCO4yrpUd5U1utwQ7Rx3GWGIatDk9+m4GPuu1DaqnEHrE
qPJTfca3XbIBX41f28bnskovYbUiZk6i9HvRkoSfzb7SoBEG75LvWzRKBzU/7MTm
et4eFNLrcQTm8eoidUuCu1PA5dxqQEL8x/y4xZSERdEMqVubi3al4ay+8OZJr3RD
c5bBCayl4EFYpxxFzvKu3yAqvtjnbda4ND1TCjd7e/ONXIZUcePYZEaTVmbBp8lp
Sl2rBxe/GYguIgy+RzzOa/WYFSdO/tTg/sRIQ+qjG7Yde8zky8weh0AdYrrNMrco
33za6pQI/YtXMNd+/esj0kiwkzUusKWEWV1vpacua90Lm+G7K1zJefptCpKBXXG8
7zygnU64THs32BCg/74B537/5ACrvNrNgvwF7/nUHhNyQDWwTZ9x4xt0xeMEeS4U
fiY7Le/gdtsv4Oblw4ZUzxEtLmpAJZ+J2PA2/CZmMHNTze1Pceybec8fHiUfQK2P
SHiuMCxG4RcALiE++rGE4QUQ4H/zOM0dlsg+AQUhYFsGccxrwtvFHu6i8k7OY6Ep
E1PlIxMweSho5vESWWh+QKFklfrCh5dAFzUfMj65UevdTtegKXwqlssjkL6xsVrO
5xLX6Y4coZ2xJOkOwbfCijYcbQN8LBp+H8UHn4oYuOGIpWnGNJtmwEGvNfeH+oFZ
i6TbzYl83gt1zWcW+oKtA/m6eCUJE4Cvu6JHf/MKBNPIF7Yv4Ca78p5gpUC+e0m9
u+DoUsHFx/wljjbmG0MRUh/zs1k65i+ba62Y88T0pZ62V7gaNFcVAGQ5OeApivQp
5v+85SGZlk18Gh2lm8g8KycWnlfb+W0LffohNg22zz6cuQRQpxcaXWzvcOlW/sJV
xvLiD13pl79744D/LOgymPyfww7bfgfbqtcFt0/3ABD2H3wnVtO+jXxYTqIIDDB1
xcI0ROmDAxBgq5hOJtwriKYTuq0ch+QwkSNJcXQoB7Af7tEtrTzLcfWDmPxekzGb
DCt3C38gcQt2ObAsyWTDcAz0pu7XG11bzw9WNxYw5YerJfnNXJwy3ndX+V5cXm+A
0esmmYLmGGa0rYFRiv/CszQSbw/2wdVnfucK/cgKVojMIJojhnd7IOZ5MF5jFTAe
86LNMZgwJswLpMFPXfxU9db/XudX38rwQp7uqqkNzrgfCRNCYYCaYxq8gAlLfw/R
NNMdWoBI5llNAXfh18w3rNsW5OfRijj4o2B2C6AJw7qOUfWG4eK7jOm4IZTq6dh/
gn40DXDrzsUjF2PoD7AtIuaiIQCqZ6kG4x4yzSg6IRY/NaXA7us6uzsleflsl23q
SfiCA9nPTEQmngISPV+k4e3DTyl99u+UK71/RFuF/ptA7HTOKDs5umcV8C15HLDf
vi0ALE9WR8m0pUaHvEvGQ+skJ2havOrWbQGcOzPiwqsOWZtePD+mtvff7kBalFfw
pNHwqu9QWD6BkcgGOOfuXKhxfQW78uvLT18bed0k4pdgALNu3Ojuh4ZAJ7+iACfx
19RxCSRM/WLq28MsRTj0/Ju3WJ/QOI8jMP+IkyGPtLxlcKKHOCbYpWEERBZqf5rA
a2cJw48VgWv1oxBtQrBtJTVfx74eNUSpazPNMsJgOL+fMbbiCiOp1tpiHcWq/GL+
2XWS8b7qdxHt5GRqUQXd3Sj9jxYpZdkd2NHmgTBBibqY2N5TtQlhisVhF8hHTnzf
tsRz8l5xVW3oV84AnEJjKuzAs2WFFgRZyUYixSQ6g/ivKh6u18vi4ro3zTpX6kjW
P0IE2LkIkBY9xkbxmqjYkw7fYQu7N2gqRcu7kVkO+5huvRtQ/jOt3hIa9rduCMFy
L3le6O1PAr3F9F9qEQ7rH460V1BHz9SHzuMbjizEJm64mefzgySgNuWSpYqNj/w2
++bZxdrLIQbYtdE09herD7KtB+7qbo+wPCSY/vmBFunTN2yr3rm85NfT/zc6cU9f
n8GRvJqZ9uepor8as7RDuQzIq7ncSWIp96lRegH1J1UnaQzCuGHSWUWAZ2G2TJ4A
Dv6eea/G7nAgZcQIyJ8DAVhnNnJxnF1j4v4gXLFry+cLxsB2540fLp2P8AP+9lKx
f2F+N1pY6zp56PgySAR3CII7nq+twjfLUyflVIQ0xw5zUF+dvDNw0+nwIGcvhL4D
qD+aw2+sB5UkZjODVMd7euyCf05LfANelFtv8frM+4nAs64ngpqeCWhpaFcL2vSG
/NQTfJkyRu1eVrEYbqAkHaJOgRq52s+GCuZYKJB5zcmKBF92gSZ7AGOjWMXb0d/n
kGRx4oWhXiosgFc2YwDG0xBpMprdUKR+wLUjcx8CVF156Z4uXhhR7+tEjSDvffZJ
cX6ifJ0Pv45kacgB3EWv4Mk3mZz92rRfPG3PddvS7L1x9e6woHkdzjx7EdChkT6L
+ejkBrmlggtS2rCC4PVdY+dEnNZT7ZmWbcf+pmWhCn0G2KA0fJXd7o7mBQl90i4R
MglY836KxHXIA3/ByVegUeqOtpP+andK+22xRc7rsbF/RqO9juVEQotbumt4P417
MmFbTF8jJx7oX3rfVIsxI6vT3dJLIg7ZyqFFsrTqNyvTKHxtlyj1dH9hOqqBCI1I
vEQA4ahHz8BbulrNbqaPtSNTjynR0HXXbzTdHProLzdS5MqwJEhSZV2xR0SEBQTO
7hq9ImtJlfbU1o5pajt7aGqQYaPM2SfQrcvC0mLV/XhKF3V1ncjcxFItNx0Ewe8G
0uMr63hNUFjZmSfX7AI9qVgDadmmAfbwKxCfrAbtZQFmutSlLJcOCiWqlHOSnmww
DuK+nibERA/WwofxtS4Z2XUVBb0oizaYw2pJSWnrUrkFYyk04tq3L0Rc805rVf1n
zTPu2lWuXj1ezLMNPDgSbX+JX4yBYkrBo9aqSOM+5jQ6FobhI2CY2LLJUS9SlwLc
UMgq9pY60DqusB/W6Mbd7ORkbjdlf5AzybRdTJAs3PJrhNTi0vJVeebcgLwgFjam
ddiGF+q1hytg8mqrSUzQjgXvIeGRwt/mtvNo8mBbb/v2UG86+m8Sp3s0kz8jXszi
A6o7JRTa5zwtZTEooiuZ3LJlaPsYbH1mgoIxnErkLP0Mr/oPFqAy+LqFwc1qA3BF
Jh2DkckmMcgYC2C6WmeYAx8csU+uDtZzbaJxEJ80l/xZzrAboYETSJ67fYIl7a8n
WeNQThoXcVdhZ/VB9dZahXGnBB+nodvCWjfqcr7CyL1TDSX/Q9C6+8H8GGId+w8h
QpBBWk75vRfHztUZlvjq/mEclsLyzlNUzHEStYrjwbJ5aSozw9uztXqxCONnJ/Rt
SWNRdogDE5widVQ3vcZqkMqf9c0gXlNFu9gw1oohP3wNBSjjW5dOQRB/pTZXsbZ2
SVNrdZT1xsRm8qujWVdLQ2DHnwZ/Lh6vPQIEMD/qQGdkdwdx/VZgIWE7KwUoRrN+
m9pQexQJYOPzkQB49/+FPVF0YuOVKtmbfoyymrVEBTwW9qhhNsf8MhYWJrxMx9hy
vXYoh77j/9a6IZeZtBi4NsSh+ReR3RhbVBie+INdDpjZ2xEjKE3iPc263P6u25op
ggJCXPp4ixnaSeHd3QdU5bRl/KrtxRz9iskLyRUzn1azQpBxyBtdzpc/jnBzMRNP
wtQ8duicnRhkGPyXREOfFVDqtSNHfJmAnEMocDCrqiCvoCv32d6V4cy5iNw8bUWY
C256WD20qDs/Z7U2NE0Gjlg6z0TmXbmkedsIVlyhi94JlGihTJ0x7djNALaNafgM
923tjmogKZj+uA5h299OyGlQYRYNr+OW+slTBvrQydGFKKx4dG3XxfJg2ZnhiVmI
lVSQg1YUUDgDO+Pz+bfUz2bz11tuQI2K+hug3RTw1gjhh5+rKdycc7AVo+dLqYe7
Qlk/EEYacQDBEY0AxcS/YAoUhgISjOj1WKezZPspEkoWapYIhUkbFSKDIT5q5ptX
HlQdwoNQJsAdpCTg/4jUuflCTDXCeNtSX3SpQCsv4z3d64owzB+ClcHRL338F0C/
I6Kt8d2FbdBgjD8doNcj56e0UA4p2TLf9MI7Mo3HdMrVzL249r1p9583/ed9FkzG
hApOsUySmWlvW3F+dzatkywBP59O+AvjXvpeRNkHzMdvW9JLdfABxbHaanHJ2499
KopMRzi0ZIe/s2Es5sr3xjsC/AAdtnwgL9E6pejZ5AOrM0yfg85Qkbna5ubiv6qr
hKawyGQjuIWVAvCeICtMxstpvH/OOHy1OyEt2/LPN1z9TOhTdH+p29Waf+5bC/FU
MCLwk50UljsVGLF8kelyaxEhQRCbE6pLxtVVDNWzA8TkmMIleg0bbcF1iDtg9nzZ
4oi1BKdihxgobf7inOA3rs3hDWVRMWtuGoY90zOJhbSzXoPSluUqxXz3xY7OVdgD
lO2R2CTjdqjr62oqvuuyhKF1BSZz4uQcBoto+asbZmNB8HMoba8wIHYXNjPHvknx
jPdgaaRqir9f0zULYOh0kUY6ntrSMxCiC9OSJFGx+lgNinq6q4GuBV66Y37pDA0q
B1hhJWA0Ymrc8c79DFOkRYNiqWVZ45i22CiK0TWsl+i/d5ewAomxnThpqPDRvMrE
6S0imoPbnsEaRsaFa/92I+r0o7JN2jkIF27jcvM64dzpoYg8UPCfq2ZhH8tQP902
7bjYGSUJ/hqOaH0HqP68RFJCT/E9Oob7gGzG7XWDbNZrXcnv4NL5kqYfiJeRp0Se
fkT0E+yJ5bQc7IBNtD1zfA9AsbIwqXmTwjkaodbcHWSIRor1VJ9gYfgebnksGdgO
riSxOs6sRpBmDEbwh7q9jIpqDPNFbAhcTgI9CvKFNn6UfUFH8nv5eBiJmGdk3T6b
t9cCGGBtErXYEvgkqsTSUx1q1XbTb1UPYZUL8lnfZEupqx4IEGFDyWzIwa67KwV3
jKEYPL7uADgCqk73Zm5I6v7x5ILMmpbx5DF3GejL3bMofSrRCJAmun2rse8Mtvb9
2l0JildNM/Wj+DDfj47ViS1oHtzdbbsJgt4cuogbj9GA/OZEAyWG5osc5rnbfME+
TsaSnF1C+2SBXLbZJLifbsJkqhvxfnhgGFd0EDBXYP5f8UCvruoyyqcPa7GZ/n0Y
PT5PihysC9V3AOnXYz87DR+hYlYOopdoZgvBqChETCSumEUv+zpIkQFTaIfLQ1fw
UI0IRKUHDIVrZ0iSnIiCfN27qSiBSam9atHDXDhSzFvXaWOLJYBKDpdo9uHqGQ+J
axynC+v4uhYzNoBC8GcbW5JTgXvOdScAmemKs0eCZkgDjSTvmny+p/vs6FpiMoti
3PNMNvUTvFQSVvqHnYTENvjpgMU0u/nJT28eNMSaavItix2/VnEKSTv/NLSXl8PP
HhAr7pg2534+5kCF//fvFT0PwZEAejkXmtR/hmIxl+hMpboFype/+wetZPBTN79i
4gyCKZyt0rGCqyyCumM0XsrKYQ2A++OccEUASm1BgLzWkjH4PDduk90yo5Rvn9ck
3SfLgB1Kczx11wu48Bwu8trkjVaSVCcOp10D9HM+1X+Z54Tar7NpdyWwe+hTVoRA
dPin2lVN1r35F2BVu24PjRFHUa25Sqb9Evy2n+YIiyHSoxxRFiVrL9WLw1FXv4d4
dxve4YlpbSk/9Bfeln7vVBy1hK+4/VK9n4g5RCMmbn3EsIeSdvPM/HnqCTSqdNQe
7tnfYATpC44qaS1xsY8tEsnPriLQ53IyxrU8eUBWOsw26w/kMj1mfm8thtb332Zq
S1rbcWTUvg88OOEOxCAJj3S/ds5F2/cnp+LWxIxFqfXZFDWFnCWIif9oA1sbqSaB
OI9imiVLP+nFCSMr/7fD0oaax86UvcxNqucbn768yo6Avg2daKVPlvCle+SjtyBd
s3J1ug8wSsInknqsCDX1mkNehDZUgMofRWJXSJUV3v+uAs3BF1abDEw90jyC/8VW
Jh8n8EgGOG3xcwTElZn+mxr6+qQS3gl2Ygqnh3h36ia1+APt5A+qStM85xXGxNdC
lbJvAARuwncawBZjGlTMnTPa1Cdcetzt33xIVzVA3utgbPBSyOG4Q5IgqkywOzps
aqfo4yZrYdCbxg5rfnABAABZq1BNsOA4dTPD1ZSbuWk5P8FoEOKA9n6T/DECMgQm
u6Z2LNdQlPWi3qzUQtTjRmyzstWWVK+Dd9OWI5e9rZgua4UqKry61b3bmNYOsBgi
voA9uSgX6YXXasL/2JjPp51YBqyEDaV7PKQYUakAt5BT6P/xFR4Sl/A06kpVJOBm
pXmnVYaGphS8V1GfAM9QcYKobNFpU0m/mDI0+OAu8mAiPcxBi52P3pI86INORcgj
60XZMtvDgtdL7yZKpg8woePIj3IhHnafRSpN6QEysFhy0N5DW6xrpxoh5VYrnfhg
vvJP2U0quBm5FN/fIba0QZiDoJRMHErCZTD9xtntHukFGch+32H5AyhCeRO0maF6
ua2x9uBg2IWFEohmTcIAmT9xqdxguymQbUIliMUncB+9fImE4e8PVuIKQBSiX7Ui
bqBqjp9tPk3JunswZuvdXENxaHUYdJ/xZtQjZfbUHtDWG18bqEOzMiHn6S98fDit
lyta6zTcHWdeyRbae0g83pZwER33EGIy9NvXhXTiJFmAwwfPvrZr+YGXNvyrWUA7
JofaxDT4+qy2WAUHqEEATUlbiMMmvtzt5fjzZBTUcbk5nDYGNjPvFTdnE9jIEzVy
jzCcGBKNh3/S8bt+U+UivihWeTl6g6m9ihNH53fvqXf0+UUveru/l2p0bqZWwjqE
HWdXKlueo2/Sf2UYbA29/Pi6Gf3eoRYISSXO8qqErcWgi38xuiFwjJEUfM7ndQQp
SxNHo6vWlhE5NYTasUAZ2IWLZnmjGVhW9ZoxvOv5bSKRq5HVhpt0C8i9ofEpuBNc
qMFzlppOoi55hWJUA28U8K9P5gytchdnPSyTZp1DFMs3l2mozPVzPL9ndCwI3Vxz
djo9LY/OB5ZB7NR863wVtW4XGwPIyQa+H0SphVqPooAFAz3JQZq3zXYe/FeL+KYg
LRMDFm2wl6cJo3nSjJmo6uMBELPQJ/LBrA0dAxPV1S/ySdowtVCnBVMLA/YEN1Z4
BBW1b0SmsELH/2AgevasBrVB2PMIeUHa9mRRR/L8hHDOxScjKqakt9wfKlppCx9z
aWwi5g6v0HG5aXSufysIfEDgM4cIt/D8ajuzVmh+iUeVrLyj4pFtse8Wsv2EieKn
Zbyc689YFoUa4FcAcTClUaVsEqmdDRkWt0IOoSUFovXE4kXPTDbNpEhC2d7I8Qal
8UKnVCIccYzP9WV2tcCg1CaF139178lwZQ3xvBb3/S/o6/knhRrt2JI7edz8CO4j
`protect END_PROTECTED