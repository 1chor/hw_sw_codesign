-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RcQu9AMurG9Bnqhk/WewD5RdpBIRfUVGP3mfsEaB3AtoZAtdSp66rdRpIbKDlcPeQ3mLifwPMh9P
BpL2xbxVNAwkN0XOLH3iweEoCN/4PwTFLt3Fo5RHAmvW0jPco9vWex2rCphQTMRPdavVwWoeRB1U
YaTm/XLmtrEbZlmKLXSNhdPlTv6IUQ5s0kwBT7AnJweBSYj7mz9kxhhUrWRwjAqzKo5A7EX1/FcC
uCswJrX0fJedSfrJb1G+CbqdKAzohMYavH2N8Ytk1gxyMbMF128R1tcbKAnSododu8Sm9qTc/zbK
XydRHlTkjWBHhbENKQL8Gv2G8mzEkN3cWOGJEg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49392)
`protect data_block
nozowNvP9cFBW0OdkdJkl4+N9XWkvn2r1oCcgMDTJK+pR2zZKV5VpJ2Xsw8/B5cuBk3qt+AH/+pr
qAiiYEo5/UD4EhdB7BaTAruv+bvylhaeuDpxOUY4hEEBqiFLnEtqP1+vkxvIwwjMocMXyxnaAgzz
oVNrXh02TnavNmYEadpmQjJcOLYH3czPAWn5rEYmRLedjL/EzynLiv21kTYue0rguEnjqrCUiouo
unRzJaeyUUMZJD/UGECyRvAKV5AysECljeaXPQuJf9783FdnuXM6c4LZMk/p4lgtaN//FA0vQqf3
BfyqCBKGX6Ei8omWMFXqhRMk6U1famnt62VDv4nGJRVGC/iLXVbXSTJccvTlnPqcz7HSVAhpfQ/H
0RHtMrweJTusKlrumm+/3aR2QLEA8n24tv51VoKuf47ILeL66L5k/R56e5fmrL6KeONy0B6IP5jg
zaZo1Z4KacjixQUFDgciHjOeX39a/H8q/vmvQ4egH0HIeQLIGGB7gLwF0VDml22ZIaxM8e0gWIZs
078zD0kX0FGKt81YOgFYX5thzAqyQfgS4im4HlmxS37RCCzknB+iNYGCMAGWsOfgOGSTgat4Zjcg
ilOxE/l0ZQYAZw86EzubIVo1GOYjGpMcQmkvfBSVKV29xeEalAMutYjcMQu373LtF08n3KT0mbUm
Ymx+oO+jn+/AMXUuxnSeFodiofpWR3L8KaXWECcGpSSVX23xcCzx0AOLI3QRW/hR9ICBKBAxoIk6
vF1widAln6D6uWRYlbTRvYWBYYhIW6Zs9iW0OTMRC3byExAAr54vvNq+GcBumxttw/84NCcwxAf9
eSipXoe09oRoXmbfMnGoiZ34oDLvfU6BlrYSNlcCEFT0/PliZigUaQTOGIysDLdAzWugbJd09ONe
UA4gFcBRUH5uDqn/8n06RjXtd42tUHCT1PkCTB5lCnu+i1X7g0/clycunRDRxWHtarVT46uyQYAQ
gzey9yGP7s20lScNf2uv+6pxw7xe8M5wql7sukKUHJADwxPrWOlBxORB/y9/+vCmoB6zGgO85zf9
2AzdpWp+A1HF30j8DrwYYwQRzKjhhy3wqvyZucTmcPfvijhRU4kKdMGNUcOvhwnljFgTPS5d5/Al
BxFr3WHLokkaN1OA5v35cPkzj0fWbaAOAIuxplpP4vEcNlInZz5yHBeU5xrWCiu9nByY0Kru+wP9
eJ6Aj0tr0Hzd+OMY/cWPE6+l0t5E3QFy5jSJE6+Rttkjg5rszRTQVSNT2p73JhqmBVzwlxq0FxNY
4e/vkzj/2CyqPJ0uOJPxPIrE8bjXxvrajmzZtHMebGYBV5yX46RgeLq9sKfovQsHOasL9GG+/3U2
NqbIQ3vhZsxFa9qKV0MhT5FjoTDVUqIx5nJVMQ/ZKYwUCdvEZ935YtCM1NEX0hlLOsTI5gMiO2ny
q4h83Puqcn4l8fqCQ2Z2VwwDNmsdMSGqGRBjaKOO1y9plceNdpjAycGUMCiTIQajcrClox5sb3Tc
fS24awU9tX/rwH91L71bQHqZDObpsEbESsDgkLj817p04lUZtA49yatzqcr462GPDkS9puos2845
T/zKQO2gsNbt1GoS1TBO92Tyakf0MQznpnEzgzonRzH/F/O18xqBgxOqqcJtTCUffShObVKCGsK9
yNmSZXyXWWiTt3jZO7o51Zo7tKN4Ubz14bxfrYkpawiSbFIk9RKwbQ5XQdc0cin1oWedju16NhMn
H9uE39eymE1tVyU54/j0gKg+Hfv08G5DIVegwDUmgWGXKmvgJSZQxfccmlrgpL6CAcdx0mraNbFP
C3ykx10IMGQDmP/k4HyRlJBvdF3uhi4iGVuDk/4ZZVECtXbXwqlzJsntACzTZudrfOIxqG7Unu7v
avgqt59BsJjos+LnBeRXjCSobmhS067immi1ztOdLzr00eiS7Qik/IGd768qpZCtGFKEu/wMG+lP
4FhO9i/mpMN6QvsnBtJsFLhkURIY7hs+orDoeDUEWQtZtxzmPyjRgoPD2AG76RFHjvI2dzd+hMo3
1l8Paz5/+IWRVjMWA10L7PDgFJFfQnREK/ZX+PLA9Li6bwFf54eQPYjfdC3JaPXvV/x4o4aGgF7L
iytIN32D3b34XLbwC/29K+SCkdca1LUSnZy10AANr7RYpJquGH2zdzGghVBV0CuEdlCIYz/ixIFe
VoLA4yZE1leoEuN8rvdixk+uVgrlNN9zGNGCu+a6gCXumEY3S4QcAZu2Hu/l5qThbP219wasTcIT
on05dvsmeXR3oyRSDfIy5vwLQpsym8Ln/LKlDbWQlNagkanzFd6qaTtVxiSAsll9Fp19VWY2VEXO
Qtss+ldU7O/zJ7hvB1TgEhbwGtnADeJ201QxbkZ6XCfyy581j0VMMn+4L6NZXHgSOJw+i/ptQ2Qi
wo/kJK0aTYr74YoEIj2pKvbrJsBBK8zp71N+Zhxv7tDO0N2rkneWXoyIaQFb7VzpuxdLXqprhB2f
uDX77lNP2Emq3xfVjGL1H6Mynm68OsB3h8J3J+9tSqztXrF2kDVey8ydA9XESc6wa+32n2xXGg9x
mhJlSK/ULTgETiu2/7SJ/ZEvmLr8jLi4dECTZG0/rHwhxT1uMB34UprP1zpyJ2T0QmNLPw11W2/r
91L5hu7kV7wLMhK+9Lk8vEMGSJ5J8CrsboJJzHevcRzvGY8vhxoLzOYkjPJ05F7gb8Id8BSUlSNA
frglQX65pEsdIhNw9XpsBxFluVy3egIhev4kJ67ENvuAY+eH1Gfzr2P3j+bRRreYfhI1TVNEdqyv
qeTNOSXPM4aYJLabDX5rZZqZxwGkxzi9VVa/Izk/rHkHa8U7NcumGTRnr9OxqcRWvnv3RTs8Ot/5
ADYqwA5xRmm1ngE9Az1wydEOi9/FVBFzP8mG3vi174Up19D5Ie/mC1UxPmN/YL4Wh4C3x5Pr/+xr
z3Q28hp8iipOAxrKDJtSsRP0TIi9GKjJUvR+a4W3H+29MLorlDzTjp7ZeMFEwjOKiB4uSFxHeaYu
58RMEWxd81RZBu114ChEC5xaMD4j4vxz1SDje3ec8/9QhykgBAS26uDyhihrF08UBXjAV/zud2ys
BuqG1oD7AbMLDWgeJHk3SxbgcK9Ow+pDJj1Q8Hq1oDC3JTDsXMDSBg3EoJfr99oMEuoBOPB6UVNk
W5TEJKRn5sHVpDAFA1VzflXzYze2aFLeKBH6V/wbiHmj0YBYjMtlifeodNSQS3vlptirQaXY23RU
+ggjiBfifE6Fl0vOkMpeTNdajDiORqZDbgm3FurocMLU61Q8ORywlKL8PFILy+46dj2Ucr6T+6i0
cE43/UeAAWdZbs2PFoOQUTlprWDoUt8aQwkJS1wbkA0ODyC1ZeueoknQgx+VnEOUCppe4ip5T9ub
VNyes7q+m8yS9RkiR6NsVWNzGu0h+7b0pWIdk8dG60tOAueuF3ehXtXIuDl+KdR86rC4XBfdhXH/
8/gyDuuSBOl0xVInFC+C7oSsfPTkd+BYIXlcpqAT3GYuZD0GiBidL8sDahmGyHHCqtg8XIQsL42V
goCSYgrt8XchGCUBDlNl4hbwRSS9Qj0y9d6/1HrC0xt77Nfrd0ij5EdqX4sEZ3kgZIu0iQUiX588
viuuqob0VuzAUKkPLdM72X+3z/UXsdmDVFTtR3mttpRegoF2j5kYIcXdtIalyvdwMAsLvQQS53yr
HqNQ+7YmSvluTvuGwnR7qt7mGP0m58gkC+HN8JIolDbB7G7DfsPJGZBKjykxuBuLA7BeDHwubS//
QM9qZnTISP46yNkvgQWc1JryyfJsYjr1BrCk2n2FcfQfgAnun8jlssCzpr6gFPt4FFUAIhpIMxNT
2h/XvFRezewHwI8EvzJ95+tjf/Sg9K2yHaGPpN6j9SGI3rHnrcTD9C6PYHqEIznlPZhpYGFfDXpp
6ql/uUNkqPTnV7v0l5fjEGp7GE7qSAtWjvRF7o5t8VEzSYA01XppcRIJEosf9w4uTf6aJwJ2envg
e0EXm1KVHCK4rzKdbR0oXz4Z/ybf7+Vx49lpd/OYK7x6DUmE4YM3GVFK3G5OQep5sqtj/BHgUyHs
iznOBt64dzM6uFHpjRDZdff/74/ZSV1Qyn3cM1SHp8WAbt9MkmtZ9bzPLCs7WeJb6EKcnt3Kv2TC
xiD97HOGEVIqadtZDHHZ6+0zq+19NUPo4dFIk+7O2FIy4LjPSHqcBKuyN0rCPF+jE/D0GIpAh6/X
69oBtcJeZGLNCRKliVRpjAXUT1fdRwCvpE2AO9dpwpwNcFfuwFbydxYJg1asfOZ89Fc3TpXWk75e
f19z01VcRBTubokD7pV9RPqrLV7hvtfWorOWJG2LS+i5c+G9i1kSRG5vgWYw7pF8X4DlhUc2/08S
n3/WCCfqgVxArpkSzkaozB5WdpilPLaEMK8W0LaJjiBljKmsn53Q6vkk5ITQKkTJoqY2b5EMIO9F
OsYdF4TGg5SrTpSfXAkiEepjdyHBu9lgXbkPGlCm82iZePoZEU+x6YVl/QY/1Tp1OrfuHU+WJL3k
xDDCRCdiAGEHK/kYjZtAPb+5eYTyWL2rSsGZ9eBDv17U8oxBw+Ip6wundNEg7hygBgVFB05CnBJ2
Miih7ywM3KW+Z1DFPpF7lY/WxTeAHnsD28pfDJYvQDGnCUKZvstAL9Ua4RHcF2hEWYJuViOLGCOV
3szhHoBS0DRKsmzypJN1UOma5QuLJFwu62ID55C4lF83omeJxDHKCDuqrN42izkANp9RIXvjb0IJ
hkkB1aAzlo27OXELY0SI0d8vR907XoBCJRZTkbEtdVML2oNd14yFQpyazi4dFx3A9pcL1dUMbje+
YWDq6RflF+Y5L5vQiv4fR87X4Nr7su5hoP1mvxLkGev/Jpgh5swiSXOdXiIHkrQtaQaICW2UyAV1
Q4PsyN50bfObkOPrChahnVwm/5L4NvZETkUkB9ZdSKL73EBL4M836PqhisoUz1W1Di1YyxIRhCi2
P2o7ZiOGkl65PCULZmklvKalIaXVXUVjiKxDF20e751g4cRvgWMQ7VbSbotANH6FLhCPSrsJvHNF
QuJJ1M1jR/zqzXrUhxltEnXk6FGbMUQ754AQu7eiUvWt42/JHwxwMsUG86r9UTT+pziMTqZ6XoUK
MnhKAtQSkmAA4qmtSjAongOa/y+kVpw9iZaY1BiPq0gQPTNXLFPWksnXUpYfQqQYp6aYvOJHbdcF
l5ELTsKYIipdr2kA4GPlcsuc/P5+IJz0O4DhbwLYLJNoj5oM0D6l3EVVOC1ROs8S1lH+pmODdI2T
z+nQNYAmOrm4JNrd1imC9TH5oL7yDHRGzSaLbH2Ew57lQNBe1XbaEa5+kfwwwZ3RivogXog6W7rQ
TyP59Z9Y17RFcPhrb9xSdwVMjWl9oALk5UbwalweWF1n9h5Mxdgwo1EY9lhzD4coE4F9wNEn3Xjo
nHh3YK7V2qrTuvAPFLJLTaJviNqLSzl5otHTzGI+WXvCVSXARMmG0cDBV7/lEQREAmNnx/w+BZwU
WKiNM+Qy65JgrxwO/FEOBsx9hikYOVXa8GDCjl5ObAn/ZMq8utjQ1qQz2pxBTxaamJWc11rj3d13
7LrhNscpuntcYCkEBE2ZtWEjJenjlvZS5AVkPmxEVQ5erLgehPZ1fA87+j7F1GiMVPtxa4fEAjCb
RarfSsXh9Sz6ZilZviGKDnyhRICkIwbx6SPyPZWWShJHPG1BimfpN12JVhdDjyXl8z9fzo/MqTho
JZjgk9D3jvrHf9jpiNyFzS5J7fj4pS0QpsoEE3u5UwYryZY66iZdHP4hDsE+RSZPP/eO0TiBiYLn
IZMhl6dKhlcneuFUokN1QLiFm7UjVxqd6jDSkUp8wy9AJ/6CHiObIyCLnGgwn79kcnz7KJrT+A5/
EagU9Mb78696OICide0J5j8CAGvnR6oNax1qwViIB+uTA9oYbbK9ehAIt8dpO4Y/05I7UH4i7f84
8jmfFTGBHxCQo5xDHieJbpsHZYA9c7/rb7jYY+1OR/gyIPQbheI8f5D4mUYvQ8v/eXt7J4qgOWzO
mEJsnVAOaJj2ZUyXy0LDrHG99AlEVersOkwsVFyUnatdyUVxb3P/HsLTk21O5kmpALblEdqm+N9y
LXaoosbuW3KS4KXYtNd6oC6jL3b286FEBYHarImO/8/EzSQw7NFeEvdAL6Qb4Np+ghl03S7CPc+r
ThoQKxIvEtAls0BiOpqnlnvfahrz0cO2lGU0/qlgU7aF4tOHcLvvPXAChEB1VroNFIC/6ekr1bxs
YcTuPiEDri9lErIaQV9nKmRDMTyG5C++SsoX1TLy6zRxWsHROQYLXqyyAYi1IGyhwGe1Nv6gEBJS
wuY7Wq1ki76LxQBm9XE+o8MdqSm0sBok8NuGhWVfvsl6EqVd44CiSM2IW7Vl9MFqd/4+CcRfVsbM
9WITDAzhLTmvpfl02La8MlDMgW4/CBnNcE3gaGkCLdb/twLEPX02qcZQlVqnV5zHBwYe7THRxXA6
3TgrQdW1vHtX4/ivmiiYFUiVngws7rtuAgypGEgVq9tszai0vrRLG21OOQ7JZ3HE2EBWIhkcLNKo
+fFPeVenWGWr/Iw9nslKmKdG5OsiZ3xPAih8bqrw4pcKUWT8ZfgVBJV6+ShJZn/zjlTMoC0aXECG
8HI3KO1g/wYom3XKXOrzDnH74/nMjBtwFS+9gRST+JLyuIQ19in0fJ2HNa5KRfj1dZhOOQCRwKxM
N4JL5OqKe4HO5S7t2B38XYL2T9+QCypHI+C1L+ULz/AmvYjUt55mOxfyRCP+pfvLaU3/82St6FV5
kDDcmrXMZ7FdtVRhzyFDkIBxcCcW2B7sXaUebzZVTwM9tNtyDx6PPLR6nZtO/0lVRlYutcOS1zS8
jKje8YcQ9+uVKRdIKlLBLrWaVLQiNbzz3ZLb9oknEjvDNCtGhkuWjMKFQdQmK5xr3qH0LlRfy26p
Cbah6Q6orE39L5SnYcOXhwbQKqSqB8PAWciH08DhffQeh+OxdsCQjvYmcJXtjaLY7vY60HerDPR5
XRVGJyeC/uP5KhzXG8Kc7zv7ka9rW2hkQ+jceucVRHlJZqqKCsglO7dbk0ye2N+HJBXg4O7eBFAl
fHkWO0e3MXqfgFkUC8HoFLCYhioc6svQ1NlMTvJDbRbtH2ALI1Hg6YY7aLg4tOLQbJ0Fcb2MvKPq
SmkIyhnNQo5v24QBODlK7B4mWqhubj+gWsnRbj2YuS4kjUst/zROerKAmdXZ2kHv6X3e+ro+IvNO
Dnp30P4RDmnW71G7fXYakyHMpUHop+TFlCtKGxwh6AZaYODnQ+yMH48h+lpicS/KuZehUiNgKM8+
hwE8554Hq/1C5Nhs8gjKJDRh5PjZ7HdQJ9Jx9mfo9fgzuFCh9gmUptY63yTX1HLWCHQanqoFlKEM
Vzyf3zGaJ14Kr58qmy4fKqXLjjTv8wZrCAEI38qKGBzrTaYabpNYDfzPPhg+XhWWLBnu2LN2744j
Bs5AGLgiUpKL4mSH0lv/ZBctlu1VuYt6VPpWhMx9ycfbgOK85TbkhTtqudUmvmkq9Vf5wdncUSP3
o09OVoaoaJ6uB9NuBEDwfg1NVdWBbRHS1ez2ULCgdur9fTefk8eDk4yN5V7LvGjTmQNIjS6rTnFx
lbB4YXiYRn3Uf9BijJ/eszz6QXBs/S33R6U5p5Dky3EitHRjcUR1y/dK7Fs6xXx/qc02URohKwnh
UsfiPsc6zF0O5rqWJtxRODpEnyKTArmliT3QapJ5wgxyDCHQvDwjjDFHkNooghtz2rBf9ysIK8/4
lUglPq+yTGNCeb1zuKBTGWznXl4ZJXtGTL2Erf0jf4opcohDF7hdN64KLzUD+yzIxH7atfShrUPp
67fCaPF0lgG5kp1vsSElEQHOascVgf4z1x7ftIHr45AQBRsrqO+MOFugEuFhZBCS6/VXgTGDhbZ7
SZrrzEWjabzN6yp7/Yoi3P98W2QNRGVGTr7O9qx7V241qItERSVkxY7HK/6OxlbsNEF2cSZQsZph
JcraJ0BnUlHo0Q7vgbj0Mm+5GARmizhJ9IKTh+NH7bJb9gGSE2a7DTnbHHP4MviYkaF+5+wkzRRQ
fuhRQRrRSKjHLjqCekPkImk4QiZ0TAgsVRiRwtI2MtCu1xH7udVtO0EWkydtmMHiskIKkUk1bW5P
bFLZ8ysgja7mCXR+87qNMskyjRY6/OsiWD7nR3tw51eYmiZYD02IrWbMpuIT4ugs/JdKWiKTXzA6
bh/X1aGGEdEiZyrR3DvymAYZhJ1AftgEb6HtqbzRZOVI7XGbmNIFBABpXxHWk4oMyaNDfj3fRrJT
xGFKDxsopjO6NwXeZFseiJ/MWmbarSCZi4Mt4inS6p4HComZ2nBCE53uCILIyb/W8m3rr92u7t8M
Y72NDiiC88c/5b2NfY1NoKR6eRlfa87I7d9qgFv4h4VUJ7qt7dRsDU/i6u4M191UKvaZMLJJZdcq
hyqHMWY+pjT4CDcyjXp19TUx6+M6mJvIMu8TmKOuDfHMkit77n5pEZa6/QRqlCyEm48TB6F25DU9
VG82gSdFyp7p6RumYZZ7e8ac4wx/uMYCuljHe1jlaU1OIJeYXLOJDgjgcsLl1Em93G2bAYFpdHz4
/Tnl4C2bbCe75hO7TtNLr+exvHq418HYvhcTgp3NCxp6D4Hmy5xLm5eRhLISUG8COuk/x7nbBNez
XpFE6Rm9Yf2CnEtEGtyPx/VbHOsx2NkCwzQdn4yCpVlN4L8wG6TBnOYM1Dr1kFsLLmWxUwkIDZxU
3wj7iwnOaQcWP2o2BkstleMURwoiI6ow7OWT8uDAcaMMgfoq7TzXOXf12+lZNUiuGo4s8ZgNyZli
2gYtXgS8USbL4YpiMwiLT9WLX6SAzOaPy7xD9MbucSSjYsIW+T61mJMIQcXQJ1BvT9n7VPHY7xHf
VWafFEUTLuQc9G3tt5qdpvrZaRXL1/mZUw90grQaS1tw2ph1kUv7ouVrb3w4VuN1KYc0lumUD2GF
Wc4HgMuI4i+SERF6VOEDveugxTSOcijqdOINN3rZJrOERzsETAxQq5Yk9gtVzpdPfI23ohdi4tii
Qm0/mq4ITeym6IcG0JgzMTtFcG3mwI1+PiggGJM5qvlGc+hAuNaxDET3qvQXNYYoDFZ6An14pE89
xatDo3oirid3kXVJMcWul3b9pxUAw17RgouiqL+2p1TV0ImYZg+bFHDs4GIIvgXGo9AKUFq5/vbP
DZR7OaIiFB5Hg0Rw5UmsHYKgO/oF5nYsSWjqsOjzR3CV/dAbVHHuGLjMElfRjkOOnaOwrfpsRbi1
dw44hV8QRKlRXetW0GugSvwYQfjyFHxwfCCdoCwTL8KV3Oc/7Dk9WjRia8/HVNvziPIuxD5/WVTK
fC66DLpe7gfiVnQ8SyRRjzFVvlFZd6YOQMwKZukE2vHuyXLEzdYSAIokSXGv8c9UYKejBJQpuqMk
3ibmm6PThzTnTCnpG/wcjwXR+/JVBa0QNzzA31RIbi0577Necph4Y2O3T5fHTjEkCad8YspFCaIR
Zq3qhocjLAkHakowDP1D57hJnj6bcV98OiO8Ci/DkHKvzC9E19IPBQvUEKXysxCwNWap4Xb18d/L
g7Id052ri6F9avxBDuMWilO47rXOqglWpQUzQ8nZ2GZ/YJYk0hYHgMY8TV3Dc6sgur4A6iD8cLo5
L1MaNRociqvCvs5hw2CMHpm0y5NrK082MFRQPycbvScSxyLxR8M5V+5osLC+tIYnKOHTamDRaQlq
/5X5tBdoTVx/1mRV8nev30E9A60YOhTQuSG1GMNT43rYMrgOgRqQHhkmBKKHqrMCF9nXywGQM8fq
8ORlKgMvu8MqNZ3fohBUY+gEePNCh3htNNkHjfnGx+hNjXZ4mxkU6DjU7Z5eKk3TDZhLydI9ziyf
q2FiDBN/UMpmunOAdhw/53jmNsop+Gz6wyziMZXehAFouHuj7fDSHeEumrZL2RoOiBFf2VesNyqR
PkiPoe9xsnkPjaNoJliisGumI9G9Bguo6O7dem7ErvhRRLyeorFW6fpQMtxxItETDSjwPsfSHehk
Q4k6yA0XE+WU6jw09l2lXKSHnh1IfCRq8aAmUpV3N6PgtteVnrEsTmrvqf0hXiyXFmw6ykxoujbF
f/ITqe+ihNs1InMpqqU9Ll4p2vsfKq84roln/DyprnY0P67ZkHe/WHq8WBkt2ckBeat3qC04VnjQ
yxVftP+UEJwoDQgb5S4+vMqDHVCMjDXLSFOAZqpZfm9RlL0cgqzRLcs3pABKmqV+NlTGrj1QaisE
CZ6u+enSRSGmrK3UrCmTXCk4TMVw8VPunyD33Re55MkkAToIKcJsOmjCNx+C8BDT1jUjhY8ELRSp
ihcjf/ZmwWsyPR88KMloD8k8oMTcevJ5TtTQRZy8ev9k2u3hKHri7m4/C2wPUQCDG9IFTUdNrGQk
6MeT2vIp+wi4ND+9c5rEhcZHyd4iPJ1ObYzSf2yhn/Iic8fqBGy/QfegSYI0UIeTAzaoX3Pjrwo3
PlUv7fcX0AQsQwiq98U3wUGHoMZbsXp2LKnxUWFe3vuIN22NNz1hDxgqKLgK0AkhOjTK+ijh27m+
NZxpTkqGV7NN2QoByqc24qfewQViZJr7xy67DEkF7G3Km19o4IOPvkSqB7lkpm/ZEC5uJtFVpM5o
ZL+vqFJ0jatVbhEZQhiWHUUEcAJfQMxHLECn5E2G2UHx+Zw7DKk2cy3CofirfP4ulC/1z/eYz3m5
8rPIqFiMMnX0rLA6xJn6rXlu2bmpktpPYfSyWxbqRdPvOoo12YNqaVf/DwSFofOV2sCwQ0uPXD1G
KM7X7SEUmWi15FNIp+GqmztrwdJC2NoSpZB121dKsyy4QNbaU6n4Z/UbjbWAAmwahJDLP3Os2Xsn
pRwNobu3zn3mkeRNvsmwNKJWI8+zf7lm9bkqU+HTukoJJywcZGTTswIbZcsZgcALlolxdF83WMqx
xWjPRHR0hV9jZ3Jhufm7pbnf1e/CeHy8nUPFd6I/u9OdEUAkPgWWWIDzAH8czCn40ydkpK0DZBwU
Pvigf3TyiR5KENz4tDEZ1+nQ3IQ+CVI5D3cycX0jQGFOqJwgWANOzDUiWQqTQM74Dbt/beNdWoIg
w9yrhjfj79N2YzYcipBOdtqAnvxN6vMf1tudmDmTtDa9ZDs6cJwioSiTeGKOMNNNz1m0t9ae4Dfy
L02X1obUYRiL+/4ZydT4/ciBRq9isOKmh4ECgT0OBGU0VLHkupvTeW55jJGTK+Rg0xvU+N/J/6bS
urO1Bj2NwyE00bubPTKcmUk3lFcji31Kwcig5cqjD9DhQx3tilSkjnATFd+0yu50zz70+Rs9ltet
78i208FD3a6haLgH+fnhuYGAInNo72jFQ1ov0xDvnm+Eb8D7jeUaY30BqvdCdxWUGQCtfOwxUa5s
IVnntTaVHRJCCRQEwLF9XnpNZM4UfqF+tPYS5y5DOhmSDTwK5X/dql5WMnP/p2pf7KiYii86k+L/
9d3GFJrqiwztyOUIBmS/mntaeOnu+QgVFGtV4U156+OJ6m2l0DE1WX4AbAUf2ja4SH7Og5Fo32nz
TOiSYwUPD3Lnt+zgbZS95d6G2SC4yT2BX37pIa1C1PNAbn2gPcYgehW68F3X+D8GeSk+tZ255L/U
dvielj/M3wH8fScpilsdkDYO4MKQJZDCW0C16moE4uy24SfiOHxq5uYSVgI+YwUP19Ucd1NXy4lb
SXP14wGqeKp93kZdYTw4AaBeO6fJ/wpyMcAvfkBg+CAwTMhQyEFYeFGxPPyOIsh5BZjBdhEo4XkV
Gsrfwkw2nH1LYbcyAkUkDsZ34ZFumzeksY1H2dQxAPrlh1y6DYxrC2kp5I+lz7MwSf6IJmETi75N
aSZlFtjYHnxYZxxmbxn7MG8HYL/14rAt5y9G2XTuc3a7XTPhX2l2DJrWV+yeAL68e0Tzg6m6iLhk
emvVGwZc1I66FQcbkY4jf9Hj2SLHUUKjCdD1jJ6YSrjt2TtflTZ33JbQ0hTxrLwrvBgA2tRNyotz
a6FS7ygxnY0LhkiXShoTh+0Oj86CVhGYuQMCbRoEkr9GSWCthanIsKnxMKiAaPLlaHp48B7rQQbD
VLAup8TFIVyC8Nyzs8FNU3+PbZBnTfny/VZF3zrU0FyEvnWa312GiOMg99AfJttF88mUMkZpCIVS
Tn9UhLGES9ES4rNQ4rIilzbWtYzlsusNPOiZDZIHK1UnQySXi6LyGC6fdoihQpTmFJHe8YcOqiq0
iZkeYN1HXzut0fVYdGWPUoJMuLEK4xrV2Ns83F+ji4FeaGLKxErxc1kZOJ3W2EfGjjl6/ZfYJDgQ
UR6tc0aIqQO2qSjyku1cmjp+hRaK3fxWiLRv7GRP48eSa73Jdj2PVugr+HYTmAI6RgWuUM13kw7d
gMbF1d3jxnAiMsrbCAuiNNECMj0UzLrdESKpp3wnKMTYk3XZ+s1sMEI7WHUzJ55gUxv2ChT9KGhI
n7FMZvcrGzLJpokG2dYynYmuvSFND+rvOtAxj/cZLRumI7N0okVMwyLa9ffUphxn709qWGNN2XOm
eDyoq1VAASRyXx+56INxU/tJOY1wpT2dmgFvzMZdQM9D2oxNsAFVrI5uXGFcZLcuCqTvd7omdZnF
ZUjJNCCvm8neAEP5zD7DWQ3/vbOHOy8A/K3yK/hqQ4eNEQxJSrDaS7EkB7kW/W3oon7Bcv8nWgBB
krGuUL295uKiNioZZl2caNi3w+AiYHTUqoSOG/30Gvpo1IEX2U0vq6+0l2hmMC8B9baxolP+FjfX
dA2dfav8+C1w7eE9EuRq03hlfRndzkAmAC7fTQAHmIkwVWl9iTM3TCWu4aeHE0RG+RmW+brCA2zX
hJqBY3G0EMALhpPxnhHbMXlAiQPMXtmnBkhhwsoD5d5Eu5QBHFgoqnmF36AHLw/6XpN3LYpvSkZU
VPjRPz70tetqc0qRJ4zKPoK9igC6JhXidMJDiOfTsh+4SO1IrnZXNiAA4q9RHIDXhuP2GSPz/Lnf
FGxhMlkP6a9kF6tgeXiqjCVb55HpxZcTalJquLxowu9g0T1uuPEcFWmlS1Oijby+M91C/pXs0S7N
QXN3kKpUuXIiCmD9DqSmD68UgJyDh8JXSxAReAhnRXIsXCACqOJgnk79JcTZsXGs2yAQRBDoA2nW
3aD+/89LCgJWTfO28rB6P3LNLEHbAp7RDGa+gacAiMNvlci8Xyu6CW5GUaOeku9A/voUrgYhP4rp
02je9KbV9as0UyblBkmyQIL7l0vHqlBMSss+RbuWR9CXBhItFPNqx4THWjCtBXNvy1nWaFHHo03V
qp3OAvIhH8YON1kpoXzInuVToaCnIkZ9s4XINk79RmVX0Anu5LVWgT23w0yg2kHoe9I7lTyg6d+/
R3izWMGMXHbR+z//mGw98evROBmH6RTDckq2v3sc6kvJM5RsVWzhtl0IuVKF/emhcYIK/HQBnaN1
BbGNOvfRwZuI3aoZg820RHZwFpGX65OGTMzzIewPJBBRBK7K5wUAbe1xqXgGaimX98/qseA7zs7X
8u+NgJuT9WdvWpCA04U/OeHPwD85eL//mM/WKuHM79lup05seZL2VZIA2IDs4/m0PoEvgs2pF/QF
7MRRYVaBUl6Z4LIXgqh3u6uwiF7ZWUqMsLi6AfDBkljjAsjE92kbmnUyKpCD2X/CkPFzYWWTiNHC
9g0ug6mXo0/LXZYtePGlS4sLxV/ZAG+6qWF+b8Rysd6gGiV6yODimb863kIjBC3hVbcbuFtsdXXn
09oRvApUAlvdwCzDKrK9yu6bTcsa7YCRVDMjFS/e5jXZZ5b+UQ9Q+9y/uw+6Dos+z1CYVDplOW4H
FFhhT4L4pGS6j0Zm+EpnZvo4MdpQouCGJ/fcxy2Juk3Xmq44MT2jFJcMVhb7YRnWFDaZNrO5q7nT
CnvNu40n8qVHEWn2dNr6n5DLBzNhalU37+9U7qzpFpXVdpHZnWtgh6JsOzvaR4bUtbUIDvGC19Jl
pLnlK1hRK/uxloB627EmxeslQeq08uprxKaANyxmczHBwZ8f7aveFBE4HxISIBbMtA0oGX0W+JNQ
nYVdSqMVRAuMOqbmdcP/c4DQLqgEBe/Ih5tzWMVx8uTemdNtNi8NH0zAPNrnHxr9NmLfbaXkMqhE
6zbqboEpMBSUueX3QSXdzsGnSeO28N7/vgMId6RYoUtrECssKZXbfcpVCj+l3zkab6HyxZRuToch
Ntb6ZiiSzAcwv8JkkEzk9FN86BgtUGyNh/RHlNFkF8Kx6AQ77Gg3vhYphSbMXi06l1MFrNCvX1j8
efpPC4jpO4C/ZqKzk3Ii7pCMV0q7j/i0xp8dt56cOdLyp8tp00V3zCn93F2xk3nGqIZ5BSFyQXVa
U45Ww15+qe58XIBTe1kWl2PRDmnE5yAfm0o3HtiAjxBiBHVx1hny5Fvmh17D/0M6+Ohk1VmRXs61
fftxDoCMFkr8971rl/UbBxfNeO301LKXSHpF5uE7CiMKIPm4uwE2L0PUfFkuCscvl923JTpUSrJt
IuTM4toAHDD6Aw8QmuSzA0tl63e76sFExu1SfNwr5/HLyC/EvnIabmQvenpLJL6Z8Us5/YpGwsJz
lLMCwhZ+sFkfP7mastK/3ZbfI2uzSmbVknJt9fwAAgt2qJkGkhD8QH6Xg5wxlDV/FPI8XmHi8w6c
TBF67VZXu9EImCs/aCMlEH/3iyWiygMykLA9fxiNPYAwL/3ISH6+FYrWaEb81FcZuxUJs3xFTdOV
RtMDW6xDEv7LyMlsUYni4qkQFauZWSfH//S+a6ilfc6+v8DPbEQpGl3eHL6yf2/weiOEjTk7BgWg
iXyNTQghSR45yYXsKpxZxL5cY//Nm/Xp0pRWrSlg15ewVsMjYGAJ3eBOzdhhwg1ASwZOYQ3fSBMj
KHhz7it9p+957kk7VLdmrextAz/+NoFUIxY+pmflMRZWqqISusO0eRd+95VxBs9+PvNeCMZxHxeB
fD5Pr9AoZNR9w40qizbfqcEbB3Ruj71+NWugrwyk8U1LfQSqMYZD4M9ac3EegHa/6IkAh9572FDm
eZyiOjhMzxYHCBh9ea5H/nPxQLi4eodSXgQ8SR7Hl333c63dDrprP2vgTzbB+IrZAo7kpUirqagz
hyeLg5lLQpXBtvZpiDxyJdmPQAi7DGYok3W/c3eNXK3fHetiD0Jm2u+hfs1XY2sjEmHhpej9A3OM
vmpNjL1ZclfFllTvpZxkynWhZZ36AmPmCDlnnsRvn2qYGZBnH1SuGwXK3l2kVtAkdTGPj1Ltjou2
w3Ytd9WBIaRGAJ/YXvbQnx75CTMbd6mVTcN764fOdP7nGBA+N2NLRqCrCAQo6smbjD52W+PRvb5p
yWWqYB6PGJbxMzolAz1GXMNhkVS53/ssk0NjOTxJfDHIzQYs70B+nfD2f5QA9A0go25vwD+ZGdjV
5Qu7wErgfDuFhNCwGzV8X1Yx+5uIcMr4aC9FrvAKd25YdG4VbVee76kio/snfIIFGr/OQktbZbVu
+KRbyX5DleNudKbdpordewMr5WibcphLOG6m6WHB2TGLZCmZALt9glJeBrLFy0ne6S3rllRhC5jw
wsohU8TiGiDc3wQ3HyOvxeZ+ebGFyKQ+LKwNGvYHlt91vty+JkQIbEkIBbjueNlPZeRzZXplCxUL
TO+J31VeD4JmDJUhppLEw8rKcHqetfijpuK+u3JdqV9NRLzpNSkCTKyLByQdwppH+8R8L/yVdUj+
nqIb5NoteY68PUS0BcRNaocDfuTb9KTrt22xcLt+OCOR2/mzTJ8eR750i/ylxSd1lQaGtsgdPDHS
qhEcaL9ObgklsLP904xLb0JoXOCRrBlJJg0I+2JsyFuHBzycBZyS4xt7xM3wu1GwN+412ktWVSuR
tC9cRaRzxHRN9Hloc2Ls1l8Jk/UMXfVE92UI/4pC8Tpac6y970Cn/+MvFwdjcZif6iwV/U17B8uy
omdj4QGX8pBs9fQQtKM1GZrVBDFM4vKET6aC40W2a0GnCzLf69tGmLOs48I1oe4cX+kPOzPXVNMq
TqOp/99SHy+Xul2h0rYO3ZLbEOmv/znWwL5GOm+JBFp2ofCi/jH1yyIggzle0GPTwh0FOSlRsSTD
GdPsHBFrf5xHyqpZ0AXZU/h16x4Z1qETqlODRbrjcSNPy0uUX3BKU2Rev3lCmalHkD7S90CFP27R
OdMMJLgm40Gpc2STB1AChH5TnxwQ8C3uy9l7zpHvqLkAk5DQdcAPtgeIASzKD5vISZliFjdClyfQ
yz6d6wKxKH1PgTGqpRzOMoXHPUI0S2wATMAMVNzNsMpyacPAJmdlJus9Syx2B5MdOvPfF2hZt27h
J2HN0FHb7DFHyFoCSoEWG6I7L+at0lTD8ivhqO+UaMy+vzCnG7KMVKEuVyUdV85/CXyaV9EgTTye
3Wt3Vu21m8Iuhzbvm/9nBBbSo6Ekq6D2xP06xksJLnKv5Tt5Uvo0WB5yxvjRGh7DXGkdyiw9gddz
TVJTBbS1jGqMB/JtIQOeZqg8IzBP3ytnHE5YANu/24Nm5R67+GFSmepLCUtZO73qd+8tKzoNV4+b
CCAEl3lAYXKQVfgRvMmGlJffJqqonvVTbzKaLZmUoEKw1FEoTz7T9O47KK8gA5GZSic/pHOGujxt
Lr2rSSe4gkJZotsnpfmifX8C8Z8uP7CIN9Ybpxzqc0Nuu9HWY/S/gPE9pDoyCDTE8Z6En2pevN/u
UgztFLYDySgnJgp/KKsdh0DV7RLDUCr5NmnMqrAB1hFjA7xEqpinBJGkI1s4Op8fqkPOIfpfaxez
rj3uCNd9mjwO4lIWPeNTPFp8XF7wNoBfQSO1pDVgu4K5Q7JExJbb4EJWVv9gHR3OSw/Ze9lH3Eaz
EcevK3bHBR78vSrP1JACnE3e3w4hM6yg2PtjW6Bx0RHCqpgfBijgLIwbHIgIsm0QmVgnQ7oCX0Vz
rl1i8O0nAeQCAlh3rwSCvNBE9bUtASNl4UkapnHbedk+z7buoGNEFy2A+HgnQWB3FccEiG0M+Va7
qWAkFlju5d0PJaWnCeYB+teOAXdy1NQknx/1yh7lNJDgypVCxMQwA3K2eufFzetX9uhhgylj7sCp
VI/UD7CTuhODjHvL3WrH0xVRsTAafXoumD2Glos3X5wjPAA/HWjdIc79RL9sUq7gT5cFEGo3zIVu
Gn9FRdxcRj2WZI6i8rDdBvpjBUx7dG6zxVnmE4yA2umoCJJro2D9hAOa68HHqm30edwl/7Q/z6t9
y9XXtxmOBglFVrKV0B0IEETfLyX/Ko/IILU7EvEyxmwqXsgkgnENkBlOqs6PfRBMdX/H+D68BzQb
lWM5E5tEGl+HemY44Ck78eh2RrT6Wx+1Oao4UziI9rI0W9AwNSb9piZLndAOkBl9HZv28fHCyuDk
iesU8zWJJUwNiuQCWWQZvpUAU35zhg9l/pqMil7uiv+zdDH+pa/bmmp9QOsgadVZIaS1SVkF5Two
A8CZqJM0JHBByWs6zlOdAi1M9iFpnhfMaXv0j3cqSDwj+EbNCZzLKBkjC3DwjCD/TWRWlA1wARSA
qpnpDoDlm837yMDL61GbDtrtfvcD11Cd2fBxwxITmT0mLPgl6inChHvMNLfVpYtUnoJPFrRmNzIA
8SHKIEL+elvcEGSoP1RUOUNAwsVjs9ATmgpcvHAJqJw8SbkyTryx03EBA5rrxesvcjwAnJMEpPGs
Tf2gE+c+iTzKrZOrGyOh8L5bgzc5quIUjotmALK2a9WtwLnqLRhsNMSKa9ZhtPGOoFMIVq1ZNf2n
qes99wuMroGUWySg3wNRBWuRZRXD+irTeS/4j4hDcSt+OxVhzXY7IZxM3oV8jEKz3U9j2s9RrIKM
sTbp+WwgsurcoFkvEs1MoFxYMSOJK1YhYmdyypbvaSKFgLET8XxA1vAU1ia7sRVWOSp78vWvL7DG
HGxsNQO2Tk/piJ2w2CqZj1r/B8H9ruGZ6aCrgHsTUGq0WC56kfjDIVfhaCBZu8vkfup/iqhnro/n
0RLjXpzQ5Rq2Tf4AVmkeRG3uaiYMscsvxPQOWX0CzilbVH2J6fq3L+pSM9V8DBMDDLRoKgJJT9RS
UQyLJ4JyHcy1+GP2OQOysHmFZzb3yHoTjwLKL7Bz+Ny4rn3ei9qrrDMcjUGX30T7BJMoomLQVn8K
2RJh6XBJNTkiuDlKXmiI1aUL9jt+zxDYoadqc1LHtxlLqfRcsiG4Cv6rhjH3JgKsjz38iXB9gAB2
gZ2ovaXebREvb/7gcUZB0ioMw7cVbh2Nyjf64QcaVWataHKOKrr1896cnHoOt5cFgP/9GgdljDoF
JVO/Tqzl4HPG33p0J1hRgGwVjjXhieEWwT+2fwITBPq1Sw7f7I1oc/YHC+0MIwDe0DgQKqNMhHCN
KHEXLhpP73Z8a+LeqEG16D0jX56e4+YqTSd3SGw0TtfnbReP09wtYPBMeivkYnipBIgbWsBFs4cC
IadsOeWzKSURNI7y0j8qyj4htzCpt6fw6GL2FmsjQ8QayoeqfumWbGDIEZLVJRlPtPcspg+tcPga
ccwZh12FGqnmRKYubM3OkA1788DaHcDUK47iIeU+GG2V0bLwaXAN82WX1BvcPwkIE/I8tQKFk82n
WiFTt86fD9w1rC/i8boxfc+vTIFd1K6tt6kbHn5UBFaBm//mUzZItA35sjzJ2b87vhjCnFZWNr/X
zk04F8GtlLpRSjNBXuZoVOzAJjavYfBWDdeNZVpivz2NFgU+dBcYHKSe8Cs2qJYTDUUzaz/0z2UO
fbIUiMmIluydw8moOial8+gX2tdtZKs7AaE5dI/ZxFwTRtITPSXK/5G7YIHkcixa+sgkWVP40K/n
5FfUvrqKy5/ThV5BCEXU9J9bE4uUp5goDwGzuXjyVoypQb5ARxPfJQsWvm3v1RT36RZcc+rx49CA
oI+PQLz1eFFy+p1Z32M5bNhIuWM4Gyq5qEdb6zENhFdMZH+2zj1csSprinM4kGWDQx5Dc63XlR3T
j+EIvvSB+Ad+S35w58GuX6mOMTmpqIYcDgHFiY00R6x5x64egxZOx2xWFLz4dHku8NyTq8449jAy
5dxa61UnAEcVmxANO+q9rWJ+QKoam5pd4yct0QFRzTMfCI3/UXyUVNazhumBTSwratooEy6Bdr7t
xcb0mCr8AN09Gi4WIuSirG43Jw3h8USUoL/pNm52P4qCzOozAHYBL7gNQ5gSNuzdv4qLoCv97FYW
DAv5z6BAMO2JjyK7ELbgCIYugB56ERt10Ny84IoF0w7O5Zrg3hmagv8Ckt6gYtXMsqPXBn4eQu/z
Wg/tE4A255pHv5ekTo1mV5qyt1mo6YIL0NKeiX4f/L/optSjDVSIfqJzNfuxOBVtYeb7Bk0CJvOE
m8XYpUbifWCMWQIlF9VRW3oS6yaZ0SSp4EFsjseSOTS/stJ/fy5mB2afKow5XCoDLW1JuLZ6jrKP
De05hr0vrhpPzi3/VSCiDGAAkbI9tqiPrbcR4fftwsviCm23DOXsw4k8p9+zXastTPFgwsoWpSyp
vtsGy3XHG7K9MvKB0NKoY1kArsClhUg5p5Q4lb0/E5COjmP4MlqYAJAARM0lx/Sou5dP8pfjFlQa
Qyof7+XHZcmo151ZmXOsT61JI5VhGxO38YVbVW3cdYXJCtR5Z846Ap1bB5aNOl08IgGSVkF1I/YF
xkRF+8MY4lZwPjeJng9CHjuHZyfzbppixswt/2jvNg8oKLXEzbMbErJHLz8GjFqeSZVJHJnTY+S9
HqPpkC7nJ0+L3xKEeflgBkQpYLAIRKZahj8W6aMjPI9FhHbSExq/EPCYKnL9ApzFOkj6pjJRJgvW
U4kb+uhbqdfuB7cG5uacbaVvgvM2CxHKXvnTRFYyf46dt+uG0bQY4VsyRmQfcTdjZT3imrYmE+cY
FUghbp4LugPoSJ/zqHK2bMYP9F1ADOpvJKDKbrln9j/BqSsXtMV3xa7RD0Nkq6P2qzbAOr1UHsA+
3pF3xcLMMj300OmHJTqmFdQkTMh1hrvz4qvg3Fag86+g5pD/uM/wCAzF3Yi1s/6+sdNXz9HXW258
Ho5zklJ85TT4tC2Da7kVEVOMDCXU3NmSu8EpzvW4scXmjjrJ5VUSo+4kaQDs20ko/GddyzZwDDJ6
NQmkARc6p+sCetoN1YITIhkhav9EgVhFY4IQN5gI7uMTTBF0HyWNUmYdIhMCKXMH9nA47pHraoh2
AZG1h5EFPkRMAiZuOH24GwQWQv+xotKchjEWto/GFbFCnkPiiensBktqhnkqt6oknyYiyP+sVAQr
BxpdVFHhMpZHT0cmLLi7JqRNGXl09SuUJrAfbu62d0ZVrXwtz5LPaZ+Wih8bvYNZE8xit5cmKHQL
FLalbQAkdrcxYU/vqFZhGzE9P9MKldWPLVh2+xFVnIXte7aYEGEGy2bivpw72PdHRfIx23FENLkt
xKOeqYCcSKtXlSEVkt11t/9O+7IonE6xIa0Xkbv6MEkcK2sBMEuzcRO05ztezCnzINE6+ubGdE94
Vcsrntv13j+3xjsEJJqoi46uFv01VjCjsxahQzm0NzhH6ho59Lg2d3pf6yuyvZWJOzBR1Al7wP2Q
l+JKq+ulA94UMo/v597QDzQXKlwmwAxrYNn8PbxShtxn+Aw9KT6FOUlsgTT3nnKESzadrICZ/76W
hU8ERw8+wdhw8bHw/zJE2dBRzt4qcgz8q5d9bl8kZBH/+6ChV5Wj4syhxcVc3DZGM1B1Rz+gLpVE
bHrkLtQIsI6xqyZ2/oOQa7r+qmC66PEXjwoig/FEH5J9NhzC1sEhA84v82vqt/7J5FK4o95kvIAk
yEqyDK4tkxu5eiFeySdjhNhLI5jqjn4/Nu9BAvawZJk8Vc39YtoMxPNb0RLzZ4RpFKyUuNBB+r6D
m1gDTW4XcTedxS5zI5F5N9yDN+BBOVe/74JqSB4F56ktQEJMU/twjzG1IdDmsi+7QU0tmpqsNOOM
pQy0tZ4TVJYiW+aCEDoDnRjiSU38zj752+jGY7QKz03p/l/Ony+nu8UQB1y1iFlc23mfcY3YHogW
lxZ7WKpURQW/y3a35EQqm3N7vqfjAE5+Ao6UBVLcz00GsPXV40SEUS7ugN2xrXCjk/ye2IDobjUI
gNIGHB9dgzU4VRf9RTmFFic3Noy2ArC2fDEO6EHchM1Y+djNRyMK6AO7lgdKIsCC8R+rd0e3sowV
Z5eWf+1vWnQcVfuVeYBpRd3m4IfDKBR2likZE9ZTEUd5X65guyXVEAe2S37nC8t52a0Q2GqVPJ8s
qfjcGTiX3H2fHJ9/4IfegWzjPNPRh3mUbxx9mUymqIU6/X0RFjbsXotljDk0Dm8o4PXonsij1Koh
oK7gOgjjyPn9u1aDzF4wb5UhaWLpY2TTTX0sQ1hYqhuaG8B7EzmOReg64+e0IxAUT7tZFN5cnYeW
cj1V1+lR1EuUh+j1oIV5C7IME06SMmdKBQl4RBNJoGAtOhR0UQ5yORmdG0iblw/Njf09v83r2Y1e
29kxIchsEaj1bnXFUyClkThgY7nKJyYxIlDSc3Vo9auX8OSJl/vt1MKRhYY8rFUbEeY6RWl7xpo5
UkdFZU1W/C4LsPKWVIN3ORrxJgraNwvcjdDb/B40K9fkwZCKGJ3zCgj4z47naFsCSji5pWy2iQn/
+PMKCIczKsyCZV/kd9JZ/olO0TTRbYZPNdIUgMf9nSkcsF7uZEXyrYZfL2Wxtj1AZ5VQ0LpM6NX2
ykMlcy11pqlhEG5V8y2QEeX1AP1tpjvd3PKZ8yeFYX0cGBDzh+mxxV2rJawAbSXDliVX6J2oekSd
VI9qiWKFHboUhGmg1ogOC8rwy0MslC0u1m3JzObs2urNGRmbS/jWzbo7lI9oxTfWkWKNkxmTohFt
kCQvOA7QFfYa3CeBlzExkgWvD/rinLhRGAH+tOO3nFlOH+1IyAEjJBO/6+Y8MTWKAe9DWNZf2kwq
JkfKvfu29I206oYAllmIUBOQE+AxwL8TlAGi/uOBWhX5IEzX1WCBZnq31SMRpQ+upSdbIVV1zN1m
kgmANT3nNeg59sGtKc+p9DTq1Yu4lkfFJNlNWUzxWNBuCBErpQ8CWmWMaPvuUDtm7JNqKC+4ZwDY
PQ8rm2vvvJtLqTAFDiuGJ+NdEUxN3oK97Rkr7BojgQ+1YufBZJzhjyVzzVyPdPf4RdiaMqfovJgp
3WTBRW3yQsvsR2F19uGmkB+n+bSJDccB0ypo3wzbtHKobmRbuBQPnCUAkVDySiRYyPasko2VzHIt
nMWn7+l24j7PLGn/UMGS6HhXb7kLfO9Iw0xFR6LlFx6JoeMLXPKt9Z/TS1jNNVVsraz8MuJYDFz9
LOXSt/DQ3uVivttuRmpBq5eN2BPMdEDqnYG/hyWg9gZ3TXGrcHURNNHwEtbdVRz8Dvy5k1H1M2KQ
1dKLzUusznqZnvclekMonwbI8k7vS1fpK9QKAmYWFS7V+EM82sgAbbK5ysjki9eeXAvMn9NaabCj
o7XHqXPiOsNi40FxvqhmmTsQDL9OQMWXVpzT/RJYA53VdhYzxLm4TVF0FuIgZTEBbxetWscnWIHy
PGSq+m59wgiQ3lD1MLCxh//jrg2GisSK9TCBvogJShIgZ3lv0BA8Me+Hdskh0zZIKBUHuw52kkQO
cmi0g2UVOSz6F4KEmv9Cj1Y1RVMBEkpwFtD1EABI8whxRlS2p4SmhRF2pRPZElZ9zGJqXMWADimV
SqrMMl/xylbhoR5OqNYmrOEcANVRR473qYFUy6QtZhjm8hSN+VH/DGo5ik66T0ZH02hr4Giujp74
9Js6cmfiB7f0QTEVx1yb7grrmkmnJwvjQai19jholTBdlJhFc3s7ZeBm/B2snpesdPhjUn7uWM8U
136i5ueQPOSHMUqcyd2/kCihaazPTjFJA1bzCHzGh/MzYFkBC4uesqlVj3DfmMKS087T3inOK1kD
vzHPv1tK+ryl6P8XaN+j0RedEQ7WEgmDsfsphuuyme1B4lW2NQw88mz02Wv4sS7cFfSOE+oE9xv5
8tOp2FRNExRf0/RZ0J4hBBT4S4MNNFtVDIwEGwDtQBvA/1IlQlmNuVKqA2RUf0ANChGJeWTTmIUr
7P8tIw6ZozCn8xomqixH87GgQc/0utUdSwrwzzaBSV1l1hRLmGGyOFvdVh14cN/tfJdQwU6rH036
Vj9lqqx7EhoZzvDM3JNg3plkt/6Zisfrz3Hg+b4x8yg2WMnjNPuAxJAmNvuYB/Mgx2tpjwZQ6Dmc
rJ1ZmVGQERLujwbLtdQqRrAzP1z6jKV+mCrsEAcoMFWrI1DxDd6bkB96Dv2czg/o6XyUVmX5u1/8
MWn70tQUMak7LFUOzolzlqonO34qDEznTjk/5c/BCj6JlWrvWBVwV1Dog4uQKWq1Ncy3UfqDG6XT
UZbyRD9zfR7ihP4SbzzsVMRs2t9/bhu7fs6dUQtIPAauvHVMtdF5zq1jLTrnxu3miuhxtxedXxTN
Ou/AgyNa3wFxtX0fhBESxJOh34vRKDYMojxNWqtaZbSK8v7OJcb17wVEpLA+hSwoc4qZGpwy5jQz
9XBuX7rB4lQIpowXHUo/l6OEODptRz8qXsvfzNkgzUR25m0gS9qgpb+Q8ieMRlndMrLmbq3sL9QI
6Ph/IRjfyrDcSYRPDl+pr+HuY4LEeBj0EaAqs8KMdoYosRdiZAm4z6x8bQuURL3Y4ybmBEWDI5YO
e1sCnVKnBs7O0IgYhWmOsxqtRyn7KstAwlCSPfua0ig7/Ko/ihPIQEHmNcjzSZBKFY32e2I7yYTD
Wu5Fw7iyeiyc2mWoZjoaRcCAPeZoVFA7e+BaguxdYdiciPr6yy9wbqMrsCm6Bx7zR2YczTX1dz0P
Rr9ysVgzyDgon5pMSx51Hgj8Iz1NVXXDhtbtFfMNZcTnED56Fn9JtySCxuNOkFP6Y8Y1FMeIgqxN
UmWLufgctyprwD/uFekaMPfTAv6b8KvDxqzsqxVfAfMTrPX/ZL3NjqNbBJRS2XPOMDUdiE77Fi88
LmXcsVmxtTAtPCO2odymB5iwOdRUJRpCQp6c/eiJ+Eej3OmYU4hP1GCZxTIs9xnowjJ3Ecd6cAdR
juUcha0bc7QpjGvNI97fNBDZKAPuwsBcaDX+R3RjyFWStn464SSOh6DhABNECDFxh23Crl/rwtID
SEJp/if87dCXrIV2KwUUBsWsJptjM2nlcn8uh7jy9uPSHz4gVcwvG+BvhWb46EWIGUc2CLbW7gg8
HkOYnt2XI4eyreIZJ3hEm37H5zwpv3KpBsnL5EPitu9B906FeIp3LKki93zPSIXuiXFwCKm/ds5V
MfnK6UB0+L29ft73eNhVscsg0HcU7YFM10p/x0zMTdDwms3qZ4oUX1jOsslUqr/hfM74niZ47wl0
CCRlyhYbgSC5qN9zPL+j/EyglGSTHXWE9Crd/Ht9oZVjai8mjzqh3tRRXsqcb7adn3yFQR5mWjiv
VxQnRQ6WrHJPfTIBgQKuaxlsNHumhKAUp9LgjjKocVQANQyf+eUd+qkTW+FhJJdjSzQ4SON+kwwS
50KJlPhhhsvD6sMPm9GY92GbbDuXRDX074rwCqZgb6vEhr+s+02S1jx6+EaCALpYQRo55A2OsfoM
VbbZEObFOnhl1esiwxoEgHIYqY+3Ym2bZtciQfKV5oifh0wyhS32fOBFC4o/l6X8JzWGqXYkMpoZ
J1TewM01+Pn8Shxa7TzB63ZQB3I2jD2xmY2gdogy/v0CJqgWKwC8VM+xra0PTx2BELOyBg2oopTE
FTsnDxbJauy3rrcU5sgoDhh0VCGSSI4NELxdvuyVNXZVPJutya11HDsY5CUSS9vOpgdy99QqNx68
ll0/AM8FAU/xVy0HAZL6MjG1A07Gj0clZNMptUdDflnFZl0KKZdyrw3m8q/FuotI1Y/m2NP/Fgum
Gg+0TwEzW+cQmNPuW+21jmCPk/dSGrS+Io+UhDay/GWsKZjO4ZCjy0NYKPulTf2FgJQ+AMgQOs43
kffqus/YJbTlCqo04ZRTaQ+bHGVDLVY2erc0q66G6qpFdNpZjkgr8AoZYAjl9tU1Twne8JBv5LqB
bqLbFfsbDiivM6Z2jqeB2E68lr5TH6I9OiZGYGfqW0E9xf5MR4Jm7zZXqSoCtQZHLwbREnrdhw67
jhXgtXuNPcUDCYkOf8pqKhRdXnGMAAfe2Pm7bGWx04f9kyIWyEhR3b8/3qL2Eed/mpOwg4mbTl/X
9GIWyVPgO6vZJU++atQXuZ6nfXiYuB2um3q6l764iOwasaBQGwynzGBsfBAjtCd4ImeYqHYPqLGo
yG+GuSMpcce7oBgCVUoVPtMR97AosmQ1jKQRe/9IS3XJSiQ29cGF37FeVZIOiglfCDTsOWaIgWxF
mbCHG7L0nMnq2I74unSTq+yZvHK4SoKZFzZiZwcJoBpfDIx3KJefWHQVSpKBD9XbXeYDiMyUWzXL
Pcxdkg1QhGmtmLp/wZKBKFiB4H2JXDv49N9sfmmPBpE9DYjFHiXkUp5ZHMRuORuuEHmNZT5uXSDh
ujNKaMff/Ie4lhYegWYoRgDwdYR/k2K0y9jY6Sv0UGJtR/OGQ2lKtFoQHX+Vf1CA6J64weNmKA2V
w2esWo11BHfwZPUzHzaUNOD4fM90CcaARo0OYdgAgHxBWWnNaQ+BjBBSZAtxHX2SoOJqFI0HrZJO
iHfuPQwVGHd5R3tElyqstum+7oyfdW9au95TmyBx0/Cm3FdzJ46veJDZsoN/ri6kh2yc1E7WQoWR
y9Ne8kOpjh6m8BUUUeCpujSWwvLB+9hG58vIfjinmtsaNkDFrXe7uItE6AnJl+IL8ToEIGhimEMY
HgRpSjrD68xXw24mzUEz7ZRUmqB41DT5kpvTMntY7VSnhTzuwPzOEso0aLxShetaUuQGF/znN0yv
Kym03kcAUv/XqmCxMLKfFxHR91iM4DuD5yTqFbd9xKszcZWwCghqk10qrbFboBf701mpWnn3B/9i
gXxvTZo8JKQ0MytC1CVeI9Q8JzqlwKCL2D6+fgbhrzTrirrG/lu6vPwOmq8ZlHs9UYEj4mijj1+d
RpfVfXsesSH+z6Rk+qe8RQdMYoZ/FuIw10+kvQRPg5+ZzEgr/qwqM/K2vyvH0LqsOdKA1+NbhqPe
KTjhSGmlrrtE8yULsTe6mLNSPzcUiR+WXEQocKcuiyBrTScE6txzQpGhaNYBU1e8vnmxrJKiT6bE
1F5oMBwBZJYV/im90X6H2sPFnW9RI/Eh67sb0wRK88eysNKL+yrqkZ1chGsXdRaSMA3yWxmh0Gnc
d5W7/tZamRn6cVvWuhMyxFE6kZsRjRlLDCgkx0MriT5RDxuyLxWkfW13V+ENDD3DsexgABrsl1XS
CJHlrGX9jwRK5ngLiUltqPr3HJrslKnDMV3OgCy7DL7sNJgY1tF3ZPmkbMqkW3JZYFG2qxQKkWFN
zwDbXCdTKlG2WRFZ2g2ggmfl5/nqIydHevUODKLMAwU/CemeSAoTD1/5yiKSQ/VVz6K4qHT552SB
/y73pTkSCgUsdiKHD5rEa2bVJQn2s90Q9NwKEzIt/OQnCwSXueX1lcWFgl+lAUlQRzUklXyQ8TKI
DmL+4w32HE6nyyXSmqgdlWtqBzTqGUwabDLuaEqCXVemmsYdOqcH9AQ0zXbuIJ3uE9M0dK5WVPP/
PsVL5g0htyP4Ga3qEusSDdJzamtdVmzPh1JoVw0ot8q89g+JdpnJAzoK6kHQA8FRFtjlJuE5LqT3
l8F+IaY5F8sRU1cSTOGTWNbK55rjtMzW046HjMCIdwt+LEuSX+SwgMvrQG8I5da7nOq/2OFrQCpY
8eQDvqm7s9qBZVwWCOES8g/TvgOdG0zmkfQH9k6RbiF/mOJNWp732xEe9f4Zzlz+o9N7VDGsxXKa
2abjT9U28caNOXbjNY/OYEoOHSL50ovOxXNBrzdXv7g8ImLNnMWMAqK3lrWXqbQp+mWq/am5PkuO
2JE6rn8yH7ih9ClQHJ381tkA1UwYlwg7XJGZ6T0qP16wETTM87oOBhceIJCM5NwxbJ6T3oMDXGUG
IVvfhaBjMTsdOcOtaTZ39SsbbDbHjkpXnWnjN3kqzBGQeVWP8Bh3iVwVe3YaHzdacSWyjMxEr1Yr
EsFrFs34HPbh6gfcsFpluxaSRD/y4FW6sh3MaHuQ9AsgfhKlpcy0hPqf01Fm4fvVX2bDl51GR0mk
fAXJOCGlWucrvgG934KnPAyMGzyk3AsNj5lkoKB9ZbFBbq9C7Xxn8wHZrhOmuXlzVfD6zgGWm5fv
EdTFe7fyxFg6YUugcpje9bUdptmxzsP9h6uNzm8MWKqjT6jukqXAopBhYU+OVckZyytm4Kv/KowU
yXDID2zQCrdteBMvIzOuRj7Q13tK4tAJtWckp9rPntY9vZINwzKRIO02mD4+6vWHJ0rtyQIiRPTe
whM/nFRz0u8sEfQi5MyFItDyZkFmjF0saU9uoYtCcAuAzgNaX7bBor71lwz3874i2Pd4vxW3aVke
j0RZE62brqP4m8cG5UR2nS7Y4OwqbAPrWzkxz9MVUuDgHW8jkgtwO5O9znY9Ee8Cm8q+10VK0Cc3
dBObOLkWwSmDLRBUGLxBBOeZlg9F9onSw9D816rFV27K5s85cm8CDb9Vow5VrZnsdeLzAODkegIQ
WmfEb7thHIMcawaBZA/+Xjgf450ho9apw5C3hXbabx3w2fG6eirCfpjR1vS86khWMd2Jmd5+PxcX
ZGTFS8d26iBkRJwXH+HXG2OWJ8Oz74dnw/3+oGKFs9rfFx4IHcvJG7Zq/rbOba0S1ixQi60ahNF+
XD/0XDG/nbsYB1CopAcGTw/HbfEpQxaa4+rfhSo6JvBgiYLp/zbM01jt114ICoif/MehToKpwIpI
daCP7kinTIgLVzbhUNgJS8hVWw2W8InO8YDY/4pLdWGCGbkdqhysYTlBj/nGyfR/P3hVDtsHU+n6
cGuLBJQF66mivkgn6IqC2J6JIUcG6Ztz8LmM7pdWnw38dzyNhJNUqduxjKKcvlwTXJSNipTgpwCa
RN8z5iwmm32D7hUs4whN2sOsHhgjS8DBQhd/xgEi1+lysRkNsytjW7YiFe2njZvXepJLpv0w6s03
ddYVP556pcrqKbvbdfwhOwJvZGnTHkvbTqoPMMhfEZnyrsS812R0WIPFlaYKO6P/Tsgh4pjVtDuZ
WaY+db+MhQx5PMRFBN7rTr7ucAQrPJo1I/rDNlPAKrZCoyWrcm+lOtQVwePG14DFHAFr39HLCg3P
UwiCsnpV03BK/1MRMdB1+yVHx3wGgXGUTwhWmilqZeubnjgqUlHMmQ4dsyJnsPV85CNQSQXM8PkW
UrXShNX+O+A7z7AKdtYA+AniQ91QzXgm/mt4k1uXDGOiSsOzKIUcgmARmHhpvichBJ3I464NJ7ME
jq6YISm4Ej0gm7A0jzdbupn1NAGWOc5aXk4S9qZp73qadAK1SqLI7YrN8p6BuYVWnsp8QtGriFJQ
08zNhjVMEog3c/mlcIkeRw07xqe8eIU9eWhQS++tSBqvzlvRnV5SaltVcNm9sJ8f9hpZjOOKax8D
IG9OmaCJ84GahlAVOksJOU8x0YH4GEfi+gsxpEpAGitef48jqijIEZnAa+NWAG01evF4ZQPn/t53
BWUuccZwcV/aRMk9MwF5mGd1JhtAHCt6IQY9CcqxryFczddiZ/h8ZQxx3qv7QcbYDXOnot3ObFHW
3J4Mbnbd2xdA3U5XkHgnD9coX/MS6k3/kl70CLI3fpdUYQCHpSnL6KG4msCwRK7/EsQPZojkrPJa
mwPdmnAqZqC6IqT7ShYpGbBfratZhUvdcokieoV5a5dYlrCd7ipvxFrShloBB/Jpbsx9N9Vsrewk
E9v/55lBeg9pskH9Wd603415d0D8m26LgFVrhlBrB7og3OYySJa0lZu8wYN3aRKwJJoDtH6CQtd5
KZHHB/o2A9jXSbOZ7VKHsUCltfMeVaservCJ3mmPPzzZzBON4Au6pNwx61khoyKXJ5PfhXU/LLSL
8M50ZVCiZFUblj4/Tgt7yy+L3HgOFr+SrV3zUfYxyLxKWO8zdLvqt9sUbFlFYvSW8F3mWKrwQAPb
RkghhxWZaqMFqQRhlGuPLQ5ggpqjx5U5lmpLjWeaClCFIqX/9VS78HrhF9AY8C4hANrwcE94TG5c
GdT0kV7eBN14ea24c/w7wgq9GObAp/kJ69nhKupsCuyQZuqUT5FbVXp2uCMgg1ywAxipcHIjFylZ
H6kQX1AXbLplUpQcL1wHnpAbRCjT1NWXbrMElcJYqbhlK9Zh9Ahpyosc2Pra+KxoXlMI9HT1Bpug
Y6aVDNMbggidObWORTKSyS6Jtzee0/DOxrYd/jBJHLKkKColVs1iEgj9akd9bIYJB4VXecwj4kPQ
Luj4McTAFndqYHTjEIDlRUBxpvFW/f+n+U3ECm30XO6a9x9Mj+Cb09S9ExCWSQcmbgmQK5wi/ZrP
trHgkw3LYZMHvIf0iR0fDeJsilHb1j1neiFapYflNPyWbysMuqOg+eX4OTtEZp4KNt1UBhn+NVAf
t9P1yyrwoJE1hm9ngsZvFefLtBXrMsV4XS4/U9G3kADlBxsssuRDttwhfsXiD7b0h4gzckvUfjuY
byhd3TqmMn94GdShM4c8L5QTToc9nO7cEQo3eyZbG08lWfrm0t/tKd2ZCIMJOvakFB+07YTrZhYn
jvFkGKkt2aaMp+/7TCYH4VRVpT1USjyG5aAMeXofRGgym3gTSk6Lbx9skc3ih9USzKiMg/84i2e6
WyJCLkZHUXxEZOgd/nls89ub6hAGptJfW0D5+FKSdUibwhg/mchHmTMUEfSTOSowofmP5bW5QXz9
om4LwGwmSYVrfTi2jcKnvi6+tSbstEU4K7jfocNeN16rgSsGqfdqFHJ/0CCBMxYium/fVgCsUwVY
wcdsV314QdMcbB+CQT0wEaWOH3pezT6lp/MPC2hyulKqsL933mplf9Fe77o6PKsm4KQo6BhaR2si
BxrcL0tvTVHTscK+PFg79+q+xZ81+2N63MUo/YF2TXxpSQUGWEKMzeo9rBkMaIAIR0nEzkD6k3er
as6DgUtKxzDmOC9pQTUMn5bFqLx8dKh3eCaXd0DduJbce4cVT8+ux98V0YIxz52RcCd8yyl0r5+O
WwDgRfGkgiJXNiV0P9DBVuSvLxAifaf3i4HPP163i3ww6O/1WemwW5qM7WZtkVkCMi2NXTS8Xq2m
c0T44amHn058wHonjW31NwZA0N3n0tSqNbTw1Yot6IWm9akLWGTaHH9SLumS6HWHqZ/GhkGSObcR
VApoxDfLkvhcXmyhsZLZblZOpl54LIeAjLQ3hWyUcY/ekT98/PW5VSh3p4brTrYv7oIS7c7FQGOy
gpyRlAsk/4dj85vUCUBLcbE7ySIfcla0NkBvvbzv4PthfA41pG4qMw3FKbhjoveQLjk+QzdiI3Az
CjAdrAZJHpy2iPyfLYwVOo2IdBBn5gjV0CTmiUEgo4QO/LJFxlyGmugsBcm8XLds+VvqMEHrTGjd
r+n+0Hn8pbyVAx28ZfdVPfDg93PD5+oOaH4U/xi/V0DZ5LZBYEioB8UVA2W0u+yYAkYtPDtwbp/2
3eIVSJnIDxhkc6v5enxdRPZfZlk4OqZNnBwqPDdOKE1ATFwX3/qAn07yqYZV0glAMjgWlfZOSInO
rpljbGukOe8CB412st9lk4sP3h7frAn76mhunTynZ41UulOrOi4IDp8CWGG6bXfF4mIkeacMMDm4
pM5Xb61YeguqHvFVrBY2HjhwJ5nu8uv0uVXDHvi5gHHaeFbdePsSuvNqUOALFxhTUHnICkzoS1VL
8JTIcSosj5gVMF0bNcmsXwJDSIP2XlfAMIobyQpPk1a26vxpQf+a1ekJafGmvb0WH3aJ0b7fCvcx
FJ8DEM2uMaNNIzJIM3VPCRfPCHTu8Rz6tEYfegsvUdQ8xK3a9hx9QVNgn6xs4Y/UP3RvH00YiScD
hyWC04xOyk3h3sn1hj81Vw+Uy6G85g0n/K/yv6T7WEkqfBRiWMZNIW+gIwU/r5VRlf9aoGIfjh9y
9OxT3xiCCuQTDU2B8ThRJsfLoFGK+Xkbj8BvPBljn61fPGbAhK8LQVeCpyUbyMj9fHpleFqeFTJW
MasEsfFl3SaeJyzKfnwei7ux96t8AiHjOTml9A798yvoNktpfsWdFMC8vm9/QYRwU/QFOjrzRndK
XagrhH0eYjZ7nLYA8nZXttCGgnC7WdOqCNQfN4tYPyoZZlB1LwsJ/yBeZqQs9SkwfoASIj83W1cy
qOMxZ2Yng1E/fDjr7pzD7dWJ1+V+WcDL+WbYoAoYKAltyUbz74GxpZG4MP/YLlftICzdmTH5qX2F
nwKAwkq06ryBMis0btXNbNPRD4UQxXsgWiRoUO49Iz6++WUYZp64Nzmym/+jKvxiPXbaUGZKroRL
5w3UQfxnUF16K113bMBP9eHIuWKLA+DDwdDHRkk0e6ZSgmsq6PH6rJr9VyGQb1PNdDZeAv2+HJWA
A/K2+CdH16uuzG8Ob4V9rEau2KiuTw1+/WjeBKz+lOBeJqjcGNxTzRg5YRgLqzU2iZCufv1/oM+G
emdJSnv6YWFZQZ8AbbTVkPTOgPJUzpI6wpa0I7/E/lhg2j2drDeRzVG8Mfym80/yKW+/IlAEIrF0
LvSyvjPuMztJRWDfTvQal/B7oL7iNtu53ON3000qHXOYMb5MMGacv0lfyTzNj59UnWbqJT+vQcN8
/GpVjwczAHzHpO2W5vZTrSa1RwKMiPC9GNxTbujobBtofomBrCs5eHkbjNbXHitRbbvfGftMM7p3
aRX9ydMO0CJsVY2fdYgac1JgGq2dzGvAQzk/dv6vtuF1oqaRtAnlDa8dek4sb3IyO6Oud8ewfZHo
nxC+stlgsdCxJih1mjjY6ybFjH5Dp5e6gAJXtmOoap7Sj0la1xjCNGHe1opQao1QhFUJIdYVhrOj
ALrQ5Tp50nSCqSFJZ2r+s57ehbEIqnqd+bh2gZCbvkGBicqlTtZ/Y0bXwDflKrduxFbVKnpSjqkl
7kp/ikCxXrJa4qSl/X6jGE0yQYVsqvQGcJHr4RKvQdGY5xaZegzK78D6qOzHO2M548mxQCYCqa06
tanxStu1pZTsHfy33863G9UBCghtL3RzZWwmsLrL6QmsiuO4qd0cPudaSUwu1zAnwMAXcRaAHsDE
WyZlI/BFgSwd5WfkET/T4h2CmE+8AYRGKvT9ndmSJUHZ8n8kImdAcDkkTu4Lrs2WnJCQBym4Q1g3
kKfV9YWoWCYWh+H3R3LWFn+5+zosgRzoPm9jAJoo1zt1D+DQs1979KUsXFHdbiF7cGhzwWsGChfb
AcGH3I5jtqv4pqU/jZiYWZimvlsp044pYT3qkvs/FbBKa0dc95dciwRc8CPVnFjRi+Yswb4Dxa6m
tcURrXApb+cSv8+22TczfOlxnIOHls4Thl2ajjTXG8srdBiLzyza1jlRxV7SvqELhFyEMFpHv6mE
ENLL5pZ0XAJjCyNr0sTGTfXnJKbZZQ78WQ51CgUmK7G790pXl+dncQ7BxZQlq6NGQt7yDdhxf7FP
DdLllk9IiuP8gucCbnNCgZISiObq1ZECul0rlr5aaRxnvbUNpAopgwT/ily+RXpWqlNJCICTeuCb
pzerHcZr9M2AozdfRRcadnE0ojFpBROIa9Tfp9jZwocZ4r9Fc5SoNsM/nUHC645MN2HL2umeULAq
ZooAdhaaRZCXBp/0LvQvhs4rjotWWtyJSqUH1ofqFcZePuTBaKN8MlaQPx1ygjFpi+w4RbDD1Oby
ejy0n2nbcyAiw2vX4ZywjNNhkyEffVU4OPLpJzNvECV6/3t2tuJuC//npFrK/jKE7iifmphJ7ucz
Hhj0i/3YMvdodQqReSt70soCqA21i3xNJd38UAZiWpIhMjEWQleFVn2gdu7Sr10gqf1rDtoDEiXN
CJ7LdmJKIkUIcPdWlyNZ+vrLa8hQj0nw2n+YEwMPsCgFSgrYz2Q94m4SBSBvyfY5FYgTjK5uvtDd
vUOe9oPNRedhAQOuk0sZRVcrQ6MzfPD+Ujxzd0u2nfTdWe+eTf9uQzZums3hqzuvLe8nV/yfEUnY
SJ2aH0n70uffTMgfREoCRk538XVm4afm62wEh9kOn64Y5CQdHhGsa41lePn5d4/Vq6IEZCwkdjN/
Cy2zzbtAcmcG/mYTJIYj8cFhJWB/2/AaQvTRxDjyTuz3Lf9MEJ2lXbaq3qS0zCalC8eTv+05lgB2
bN6gTu3uGTE6wYEk7ugsHYkOun+canOLqmgk49VoLwpdjK+ls3TD3qd6CbTVgoonL5USCNcY4AkF
XI0aClg7AoZ2qjb1A/SWZkI3uPpt+qWqLd7aVea+VGJzRuORPz8o/n+prIIMq2I1Is9SP3xrVriN
MMjgfA2YUH4iWChp2Ckzz0AW5UoLVOyuCvSLiw1kD1nFooDWS4FrQ1uiZlGg7xCDlxxY80cah6Kt
2UlkH8CL2D0MePFeq1STCCW6d/nmGBSqfvvrPUKw14Oiv7hhfh4YXac4TTa2eUEWe+xyy6Bzsq8X
banxABuxrq0J3glduJPAsU4YQavPW9TIDl6jqQfa8MUXCg5zkp8vQAZ3deVr7qiPhgz1WKjTPo0R
XDCVHI6EgMmtDux9ng0056wbvYVmFZL/fqeLGX4kNisznvKPCOauE2++ULif8RFKmvVrJ6LqqVsv
JjE+82FZ31edB1NpFO05ozjA3cAc8bSjRAT/kKn9t2xTFhguHs34Jqdk1RFf+9i5/KU1rJvJZF1Y
pH0DOq6YObRDBWZ8ithOGutT29/YeoTJN1Y7G/I1e2oSVXO3AfNZIL8lYA4jLYHUL+BqxtAd9WMO
05uHVHah5ZMwEeahxVSQBqJ0LAWcfBYabPCDGK77zjj+Nt3puEGM/dCeVJ1itUOB8OqXxYzPZW5y
aOvf6qUuvvALNdtvt+uzXgnvaTKRRRgzohTJxsniAd3TZXqYkTL9qizW3uTus0Twc2NZKrlz4woA
yXlBYR8stbdDrDyJ8aqTppEuasiTOE6HMVCW3PD6wIP7of3556tRPMbBlp1zno8rqmU12fPbYXTT
rgWzRGl1h5k/r4vXEHw0Y0AwOho44YvOxGxzgRNbLrI+HrfOvLKgy2nuASdeU2X3LZ95CtL3XPlB
oNOfw/euwK/je56ZDMojXHj/hGUXr1j2NE0NXityh2gWj04BNBMVVsuGGFZPj28+QWW/4tekO9zG
Nmthau8ik47WqacjNrAYRflLn07WtRrXaykoXYPNlpi/8lETRelttaGhXVEjkid+rwZxtNLNBil/
qBY7ktpsEo4BQh+2QfvbQbxB6R5YQ/rziK4VDLHkN1VBBeqwd2AyIo8YDSqUR48KeYIgHrRIdYSM
gUFwrw0yVbkat9xB5YfPtZISys61Mm7j78qjOram/oYPMnYFGNxcDGx3x3sRRVmYcIEwmMsASLBT
KOAee8VRO2mXQomZogruTB5HCqojhDF2a1mMSInoHgr5Ybbwrqc4NUo1FeKrBKBGET7ct6AQO8p3
tqiH6yJBYZ05dU1REXoWndDIqb5WZUCiwVJ/OpqRg4B6zANX1ouNv9E6nLwtnh1zabGSO+3CzKMm
IQMrsAlAK4HkU2InGs8Athzz4JtZDhLPpeBqdgwdP/L25EPHOBG9havbZI56gA1ZoK4XZ1JUuHVU
YgCqjTWNc3VWG1lyfGXrbqmcJ1aFrElLnn90APy1PF0ZUa2Me8hX/2192VQnVDq+EDMoceaPx7pM
2fx081nk+rYoDUE2YlIXE1W5LcSaH//t9QMsox59jAp1CtQCY2M0HcbQB0rsPqxD3Av2B5GSvHs1
Jda9HzTy4DUYeLNpinqC/qF0yumdvD549ScibCxR2YPKgI0mMRw1WqsRaULnfor5TReO/Py6p6n5
vuSyynSHX/av2v8oTYKMiU5zMIeh9FMWlh1n28k8+DmUuhUGSXjzss6HKk2PNMrgvlvQWEkEyhQl
PhKuNfzSfvP3tLR9lGhOqQbg8yfvUPrGdNONpyXqLCBMPmJYilR6Q2Trud/H9/gVsVZ3hGCKTNyj
aIdYAUWILUaWak0VpcsuoLvwtghevCVBpE7w2/EB1xDz/STUNQSOvINVbA14P+UNjKtJqalUul6N
n3e8r83qjgkepEg6WY2fG5goIV0pNLTlsLQzfQfiL6twidU+Y9ejxIPFCpZrlOJqphTgfeHh25Ih
kZXKca30g9wBe1iNAyRqs4ybJB99jhhf/0Du1Qbu2f04gmCZNwJLQhpKrSzX5ftZZcBcBlj7kBhR
PLFxwzcT3+p+NWNv7nmLxs/QYQCRgS/rsmfuavgPj0nbiKKhBkbNUiT+4LT0FyewnIZwfY4GNQKv
/hVdlsIyb9NrIJ7+ENLJbx9HnofeZw+zAGWTtxSDDV/EDHwmv2emX61iGaX8UchB86G2tW0BN2Co
ka7U2FgAmOqH7OLsWL8pHKtGaw4AuuCUkW5x7p+oMaGU11dhJXU+UAu1LCsvbGvHHmZ9a6JU91IT
MZNnWxCk6SKVnS0tsqt7gSI7BzFQsvVV9I2fT8PsrfZn1mRuaCFbl3Kk2fVsIDBcfqTJF0Di7ODP
AvN/QZUOCLveZDAnwC6y5ZtXhk0QLdUiufRfS5WV3f8SgnT47EgR4SKNW2zA+uZG14KuAb015pec
AUAqdg1cnJKGtB/G9xHrpdJcMgpGFT07mcQcUgnmEPOEgTJr32YdHKWdkKasImNopXEf91iabGzg
5uWKJLKG7QjiSsPcgZdu5VIIU8KMOlFnu6n4iKWuBs/INdEs1p/S4cVY1iqh160L8PFGwQon9qkF
GS+todydJXKx5FSwR0Rla9jBCryHuLB/bgqa4O6uPG92u1PkxsVudkTYdmCsl885war1UqhG4I0s
U4FQ70/oKakQhkz5VyWV1GFR3Xrd5D7IQsqXkvPycbriSUSHOzs/Ums1hyxS+vKm8aqrST0kqLd5
+fGZIEleKMUbgzTVfry1WEv1qvyCt9pHkXK/weV2qvwoGZEMUYf+L84rr9U2RhDKPuSG57e3TZqp
f+s1CMPeS5TtQQIPQ+86z61cph9j5blYjk+9yOm3y3S47tGDrerD8DAaE0GR6hRKl1Dppcsts9kh
H1TYX6sNgb3DhmbBWrNPKpljIPH5Pju4DLU1pvW/UvOaGFsz0ZMtGTXYl71oOdHfxiPm/D8Z9vo3
3QeAhxGzYdKoTgwQwxePrDvVcraUKmPBySuBanQ5t7GyZO/4djj8++0NSD/+7eLcEte8Fbstptlt
2GT8ZojlELC8X6voxu7qpjvjkI9fKKTtBh5seLVDFHkkyRUXkUNB9tsLNA3VEtpc+ejfFn2GWWSs
GnY4pQ4d7RCq3wKvvSdGO/dTPhL++2697v/rXMO5rwnpgcubAA+YXzT45K/6qRW/b3aeITyV49Bs
30GrJY/cbjucDxK3JZf6xbrcoW8eWaVx+cC7fE5E3Tr3uxtGtyIWlLot1EwUOK7ZBYXv3lbbB2MW
oOvKzhAjPwYSYZVgtSP+kxlSvFekzAalgrH/yG2g3XepGo4qH9l92CktttyG4ARm3IeDVJGhKBx7
msdFlDesB0ybqTDt7xcX1na/tjatxeRl8RS9q/QJIxVq0MHLkkQOwtmCl+b0nMaeYjBiWgAzkN1k
FTAEZ49VTSAge42wI7eXsfKJro8MA6OeOUQArEJL5wJeqPo8LQtbK7C7AaVEDBHX9GBBd9ysbuyS
tiQ3fAg7V9Z9R14rcIynJc04mh8/P5t09HT4XqevPTmmG5z94Vo/ky7Sq+CQISr5UU2MKMO6LFHI
n2hqowvt1lT28bKdwqVXcwTRj8B54PqPOc+BBh7iMQ9tZBadtjyGNxjT07xWhCVmB/9Qndqb0PQ7
p+ia1ZFhblcB/vINdIKfvxswL/dQoh+LUPTIzxJqOEqkki0Jq58447mtPq27RAAJpsQtHUhuaXd2
qnvacYby2UDQ0D+Ci5eHYDhrYBKc3WJMch4n16XmGaHoYIJDWIJwM2P9YGRb8Qea/sQzMfYoX/Qp
6qXXWOcRluzi4b6c5OL32Mw8OXf1AngypTbiZIwDul6D/Kx3sH3+wx3p3GZG0UJNZipXdhOWCTJM
+CHImEgRwVCi1rVlgdirxVN/C4ZMsQhZl96AhRDh8RHnuvTZennYMCQlL2k6wQMOlJLuOJYbJ3nF
qwdfER3xHsesddLRJnBuiqeyLVA0D/ulvc9sR58yfjFpRmyRprn5vrngQPmnP7M9MTyuPmH0ASd/
O8kT1nE5DYhVFpmG+xFDEjCJOVmzrZKWBvNClH6RwGnDmaFx8N9eiafSKxT4f8mEiMfqRsXiItgc
eYBSvZZxkw1GshUbZYJbRJeChLW5ohM8KecViudFCMS3h1PiHpzVSH31RH4QhCnc3TyiDaghgEhB
WQ6M62FOBNiCUwbA/qZjVti1OSV6EqsaI3akFEUHalrCD4snaWPDbYSU0NMFPqKywFnYoPOKfcyf
oYvklNb8aTqDaBssTrI4kn6BUpTxE5Z8doiWhEviF6n1B1kErZfTFDQPx/vwaGpZ3JdlKJAstJF7
ypzyCKNLvLMuDAd3kCbQRtqIifOm0pqEkW0iH+PfqXn6RBO0lP1e3KdOPRxHKnGoJz5HhUEzwUL+
6Oa3zPGDvZjm8/hMyrj5bOX1yZCogQWNRjr23sQ8VUhUJNpqWzLHoJMUbMR+9D/GpfzLFdZku0it
TF+4YLaTpBRywahrcs5P9gL/bEfKEXyk5Vv/TLd2ac/PdR8473QzNzDCfq1l9J1N2RyUTiYkgpG1
iJ9kopri9AJKhSgigMroNBj1TFJpmD/P0aTUwJTnjUSG0G2G4InSAujUA7DWX52XcyJC4WeKUFp3
9TWUkBLdGdVVFYuWTWP0Cg3WeRgpyVXKeu8nZCik2wC+qNWW4a11oqjpCij78lA0EViff4wOcIx7
gO8XQULamw84R66kD1zjTMmwHo1p2MM4CkdZuzr45yNPl05dpm88xDZtCRCVu8Z3RKp2jN88oLgx
zbI7XyhC9OhyMKdEee4lsJZDJecvoSCHVMEWU5g03kMrGnQpEhiJ/F9diizjd3GpKkA4uelHhHGA
U1Y9DH7oiVZqG+2OX6twpb6PabBPUX8GYGjIP3BShxDsh6FzCiHgwhe5LTRsygppGXtnnSTa0m66
fRwM8DlYOn2Tnmuvb68IBNEy0WYRSSCCIkIXJea2XrEOdbnq9/Gmv30qz5bG1BvzisRSKPYwTQ76
9lsawp0w/xMg5EKv1iPWM2KdeeXCipDeyFz9/zPL+t0/cjIO1nB236CwA5+s4ItjzqU3w8sLa78R
udCzavBnHnXcr52L9p04XcCuk/oTQRyYdBgOHO0Mprtbz5/DrAw2YuFAPYwL/IMvVw52h//zNiuQ
cHSM3xXA5OISKAqwY2llcj++KLOosE8JBgYOUuZbqXB0YZ/VS9Pj9PnDnHpOLbGpJY0nEnTVk8zB
+jCFkAEAAMatV44I6xa9w5ga4Lo8Il6nIcsOx2GsAPKErIr8MmzRXGzTUbjc+vCHfzcgngjIaAAS
VCwIXC8pzzhvnM+IAc6HYgF8zsTI1Xd0Zz91ATYMIhqmW/Oo9r3N3ELullMe+9UDncf3P20eYUi5
A6jLT3xXqEkxcWN8rk7GumAxh/Jfq7fgwc8a6RVuOGGDt8T8feT8CfYui54dt10V3TTnxAw/ZGGR
d3wehT+gXTh9k4bPfTI/ImP560jGkrupvNaDpyukuw9szEpm0XHNFAjx8KgLEwp57g+T6SBnAa/Y
KAP7gI23cgNHYiJfnpxtzEJzClmwsJLFGBqJ2H5z/Dyo3M3kajagv1qw7rbQbVO60A+7CNqGZkNe
S2X1+aHXclO7lWg8HZNIRf0s4X4uSt/1MzCjtqOO+nocxQaaEMJ/eY0wGwlNyMA4LoXUq2K1h/Xd
X04Ti22z6yxxnq8DsCBWklEcO7HcFjCSyZKREikfN/+DMsuPgmmunehx7G+ivqxdxSekr3e6ivhN
J1bIU6X7JubMQJoRnPR+PM75sWDe+yGAEOWT70jGI6djrlhki5K6B+oDVB5zt59+SoTbCl8l4hXM
zTpBm9R38vfqI3NIX6MIa4OucTTZFe7v52NcW9zbvwcBnV5ex3AClJjrreacogbMUG8aid1aQe4h
zhr6+r7NLbCWBopxTcQvHHswYx/bGUqjE0QoiBAiZOmJ0wV7L3doD/5IH++Ea6vP0tpo26cmiKUZ
fl2G0mxpeoBwmQgSlDMs8xrL01pXo/mk0YDsyo4z9Q1dGJvbmiQHaWUhiaG4rWWsrLzqXtN4ZtUF
SUJ4z10ZDSxJR5uB/IHq0a9Yey1T6u69Inn/A2sbZOROu9G4ydPQzpY1FNlggFdMawiYv5ql0QSA
YfOJ6p3kad085zjdaYa0konSCLJI1ijGFmTbc06ODAF4f8uwn0PWt5bHHIP5Q474mQdF+fRAuhEX
ucr0wXweJbwVvC5fNuFQ9Plk5rYJwou6wWtslWvGaJ52cpt3n3qTfB/CiMsjpTtuxMTgjaf+MdkQ
oRYONc7cGfjXlytvswmByf9ceU76zjgRaVhHfYecBb3jEEv0YbUA9UeWt4VlUZBBeV6H6r2lxs5K
aeH9NFNqtc9a6vK36HVRafdc3h35uc/VMiRx/lTbJmnlT2VYVP7Pto+p20mq4l3KGOZ9ocsS+jYB
XsjFVtsFUuwjuLqmulWWKYxG53lZFYyU5Q+BqZcMKBQcAMSicYjmNteTwXvF7oLV8V97ewMeSQAy
nQwIqSkOJGlYgBoYunsu3uoPdXR7lXqS8T55kqKm9gFGTOOIetIdewVyDZ/K6pLkMkl8jJ8UjN5H
oLjdWA53/3LtdGCJ5nIkJXUsEdO6WY3VxuPfWvBAvoO+FmxwyT2UuOTb9lALKh3h93RmZGXgz7nb
dgqW7qsH1n/FjS1sCKcMOC0ydSSXnh9W7lJ/YL5wJAhxf8foEU05DHRG4RAmisR9MqILhvLaBuuN
1Q0qCPOVWTykysZLhcVW7yXTe1jsCA7T1Z2kQmu/ciRvpPDv9eSMCwp7TowMY0Ln8OHGWH/3RtlV
IDghGEip5jzQtpDFYPOI6blKAT/ATqE4jeNkRyHbpQjsD1rpVNzO/qtto5DFmj9jEp0pov4+B5zN
SE4elQmT24WXWxIKkmy8etRFJQdGGbQyILggzYAFNzmpjYTRNz+3L5tFqcrkwZ0yqLZpUrbv5+uH
yXDX8Ai/H46wDDJEpjSSI3QjP/QvmWxn6+Hf1NEscUNLmumz8An5mvNUyhLONQup4AhiowLrwC0q
GXIJvhv2V7Jet1YKAg1nIJnfYHtiIv7nJYVpFk8Rmu+R4AsNv1Sj5Z+GNtYTNB5ggi4OrGPAt0qh
icZbv2pQo4CFDHYA2IiPzjzvxbhsPQ8z9flX2JopFfEFubPmy0E0M/BSVmpTwQ1mLd6mG1r94Kpk
nAz/M+/WibTZWKx7sLmtVm2DmnIxQHWVnxpO49/TwwYwjqWqUFTlEadDFK8q8D4N7j9oMyKDUZVc
dGGMa2rQvSbna6GCyibr19YKyTOkNvzTCvosGu3WE5+rKBb4/xHuY7ba0sVbeOxvMFTsAc9ufr9C
KnU5VCD6BPXWjO2aY+e+K4NDJ3o1hKxbunWDIf2jT3joajjAs+IKlRdyJSSNwPiEKi2sMGhrFZ0d
HjR8JDCz3xIHQMH34VkkdVkLt4VcMF2497TA5RjTQYkBWdIv3wfst14rTh6AZLwON//T/lkVarsK
2fUCOi2FafK/wZkFV58e+6qb8fWaK/eQCPH0TUtQUvXLtel01vr60JCWxjkfHOYwL3YtMBhBi1k8
AmNb375gwWG3DGaIb1gaYLpVCR5aaKsCtqINcs1qLOLm+BdfvjwbcYFmr4hOJfUNfwMCOVif47Hw
PXJp/5/GZQQeiTcXLKj9j/5vGCaeNbn+4fGB0esrAP3jdPR7tHU76i8G5MnDvjs0SmeijywIfPwq
MrNM/ero0DO/EK66BugDH+8mIa0/JXCSbzTeHtpaAUW9pPncjrnSnFzdqkuGPaduTWSa9W1GImpn
8iB89B47JlcAWXWDzm3bpmvKxnFKeZteiWdWkfCUZ1Z15qLisAJaPTYnP1Qnkf5Q2J92YuOaXtZ0
ZKtOhj2NzRUIgr5GwrRDFv715ktwRK7DZ5ZibgIUGoFZ0zFV+ioye3Pss81REyaVJv97SXPP2z8Y
7QCW0ZFX6X91c0O4qdIAi2waKB4zid4w7A5y3bQdqHMT2u+mwQTSmYW3sMGHZQpJju7jA2v5bxd/
AKRLZELMYkcwxrDVKpFXAeu7Bzs/RDVNsJWnk05eumeEmxU5Yd8UYgzpzvVWRUjrZSG7wcysf2aL
nPcMfmjdasX6d0K3CJgiIRHyKlYIkNSjr72TOAeXmxykxkRRRcP9PJG03m/QPMTESlgwcu2rXZy2
oT52dO3x1pPWVCOFGXDhEvwFbtRKlMXQCUbeJBEfBnDLIaq7d3x7WffwPbdlMTsuV+DsiWvzOAm1
e1b/Cvej2ke6f2GxdX/EKe91J9OvAP0bqsvtUd8sY2ImJ5bZVYWjojE/gZT66ISMnrtpCORfN9rF
hyXEakBM5nllPxdW0/QEobQ1a8xKMfykL8FVWaiiVfdAVG/Af+i6yNynPjSKoi1i3LV6+KTBwclR
Ds37MEnrh0SfpgGkZBH3JkqbtT8FOEVyyFqIysebe/nf4q2XQyHPtkEXkjziucU37HBWh1ZO6uQb
iRMgoRVV3LPdjSGL3fLz3Xdx0rwauawzUEB69RInZmK+GgYAlj7q/EQyvHsv0teCPDd2n/5JsA4Y
V+F97aJqWI+dsyNTlR5AWRwHfiQH9tWlPwX0PtUZPrAM7GuX8A2qEIo9Ev4Q2cGI9FRvvKtcyjCF
quDAS3Vc2Una9oFdtcv8c8Wwpdbr6oFs+cSEF9bgMNKkrFL0Ar7QU2LzoijZJtC+MllA5Lh8vnEO
67vxJzvwo7PQCYLEx1QVzPWN0SIyjS2nRyk0MJrGcjQsHAVg2bwrovgoOUUbYORs20qL22bTATJr
tM8G7lyw/DvC5w4d1d9BeBrnbfhh+UoulWPcQhsQ12hMbEx0QfabVbkMGIJZvzY+A/XBSKgk5XsJ
Ko4euP+OnH346xAnyUjplztE4yP/+zVM4jPJE+lCGEB2VvO5tsfpdz+PmPfra+W53e3crmwrDysN
JP5uaHA22CeL4wLyWJYyFR2fmqTPHHDYUwSW9flaKNeTKW6GeyfQ4CoojOAkNsNUszED6He6uNKx
q1HtEXZV0yrnGfgOzxiQ2mUoqEwpLyIP+LV0I5HLHGVTKV2TN+y6fflEPVpTozaAraD5VVedrVRf
JrPZsQ5DkJjx8t4L2QtA/8L2f635Wc3G1Y2tl248jE32w6MOXKfz73k/Is5gGupXgPNh7Z6wPc/W
cBsJPXrVLPkTGMQsPDjHj9TBJGjcchJhWOWDukHjgiwl/Ryuy9r9aDRTP7EMyRblOyzBDMrG1vau
hITo/ZcVhnYwTyEveQ2h7xxuRfunKL94HC65TDCLPS2r3sOpY0AaZ2BmxqXzE3SSPU87v2MviRKG
m/eJ7ItMcGmY6zGoAXUnkzCKhxhfZuN5eLZgVC41aY1BfQz9h+zp0i2UvwxLjBp22++qdh1oWtdv
f41eXY5IkrI/0Ht3LxrrFH8jiJVouqLnJOJBx/Eop8UQZ7UshcskCGRsZ6ibB8mQW6e5VWSnXy8N
iqzB3TnsAwr5fhqqWDj2Yt6te/9C3gGzodUKBJ/4vq+ufRJFNd2qV+xbeqRxjTgEepjWxIrPkSPV
+zx8HTGw605GIWhJSsf05lkbwgNknFU2AJI1/WjDdI1tqEgaY9LqUvXjozRyGBQn8aadb/IO9GQ5
KoG+LJ6RowB58QQYtV+xeukI5TboMCbqZ9yo3YOHVspULJLeG867ZHuLSZIs9YvrXryDSHm8UfZL
c2RHHcKSOcYe4PlKUTYYvzN6rfi864xcNIklev3boEPKhiLkpldPATewiVvt7T/kPu4cLLszz5Mq
iJVPjV+mIa8e1SpZ7fKiZQS6v0eUS3LNx+6UyzCoR27Iei3eHHF6ORuXJ2fD6pIGbkOWXpd75HmH
l4SmvvzNXn7QtiGDQCOOy+8RBLSw/RNqy0VB7FUY/KUAm3gHeHuJ38DZSMZNhrErB8Bh8gXDpI49
ASOEcy/pIG3LF3Gn9t068kQrvO+jy/DxzRqKUV4gZHcNDOTZaw1OEvPAovj4rsnWcvWgJQiCqIQa
vu9TXjN8P10cmCZHAuLeFdTLKH1voqlseea7MUAKJtjyQtpI/mAGoDh4fb0T6uWp1OKBVZb+bIsZ
w13lzYE+mbonzrwpjv/8uhO12xHjAwY/iNaGSK8nTqnYJwSoHWUW8dqV/nMZOhVItD4dnzWqgn/O
9qa44WsrAb3bhYQ10OnsSXXnGHhoSkoYttdz5onXkGTo/XjaTBPCYd6pMpyisn0bdPILe7Soq13p
5KTW3TXm3O2RukRyzcghSG7cczg7z0/Vcr/BszkLUUXC14+9dSjppEvNbxan1GPVgK01JCbiYxqR
FqxR0WgkVspiizJ5FKD9E/zXQcdLrOKxBSCvlJdOCsCjh5qH9KTIe4rPNq2UQBjSSLkwqWPMoPRU
q43a9kXN5KKY9O1akr/bGu4nBLMNcRMSzt2ijS9dlu4jbbbUgfz7RDFIPwRoCFljzoNwv53TdCqn
pffCqRRnz0i78re+rdjZjJUYTMo2ZggSygtqxVc2i2afos5mc947oB5ocW98I3gYkEdzFJXano2z
TIuu5ND0lxoozoIP796xf3Iy21u8eUqm4wzy7uVAxbofp2FUHEFi8FWrA/J5zsZZ0v7F5GdcDG5Q
BZL+8YlqQpar5ImBhgOwSjXj9PKrhzKCs45r+YjJZJznVXHzjB68HZM9L1SNL06oPH0sJ8TBns0u
gzJRwTTnjjovkefIAAefeo4Nmyyl0a9cXO5e+R9t8PnmsKmCWCGK4syEnAwg6YBDp10y9iXDoMB+
NUsOpESPHev/x7s1Uxz4QgPBbAUB1ngZa45oez1nsuz5PICrS8MsDxddRuVceC8hMn2NDwD94qFO
rGq0iEpRC9C6oAZoEQdOnnOlHPSoDgQvl5N1c2NGy9WcwjB5tAugJ4LWcnb8OIA5N9x+yaJUP8BK
qSegB2GYTShUt2KB01FT6Yyx3IOu/SmTPUCmHTT9WvDpiD2nPIOfSsCSjuRe4vybqJg7pkpSooVQ
Nwh83rPTlMl/2W4u5B8vqA/Cnpo7S8OZxS+t5v7TD63TUDpF40T6pMVO3Wn3Zo/ba4PYM9n+B8jE
qK0zfmxhIaiLcEG4PX1JHQMwtXTO4goYj23uP6gArT9ptyjyK8/EcSaJvTdNA3U9bvf7uw0eo+jS
FGrhGS2Q0aJeQ4znIw8DeH7m0BaCn4AQKylHxZ+LBYYCwov9gnUeX4AlbF0yfplLz9y6qnTYn5Vf
MErhNLdQSpKxxmESqRj/4zS+/SXWHomihcjX44eT3k5QiryT9zmNQKc9CP4uzVWBSDMfsmxstFYS
86f5/YqSicG48iDKP5bj7U/aDNXY/nE1aw70Fz8rY6uPr9ou/+vZTwxKN9KX9tnZ/UfIo7z9t/g5
JoAqin3+VmpMUkhoGeBBdwQrJjFXJvqbfhyERGPVtoHk+83iZxTPCJAcj9brnlOnpntOpb85ZxvL
UP7hrbl1nkoku/zTLZ2uskEqLzgbPoaPPpdUpdBjcJVTiJabRDfH49f8/f1p5gOlJaFwtjpCnhtr
mkolyN6qycOawCR6095tzg5lLx2rSyck0mboQ2e0V1QSBry6j2iGYocZ+8GL63XH9XHMWNCt8bwo
BLltDtFe6iQDlOfcjXsiu+EuiNGQU9hCghTqDgRBYwvC8p8g4K/RjjLtbILB2PmapZ+imYksCnau
VGP+/WVbYsSzdxjtL1RgZDREMOgh2J1zaZlxW3/9l3yA6Y6P48Q7SOH+E3dsFv/MXLCMk06lGxLJ
ox6BzMvR8PCWHz7R50S6v+Oz/3EBxkqrxPnx4wAqOtbFdfNJQKCQVfuxn2Z+FLSHWA8jrxVUoEhM
WPqnBdFm10uajgXTaLsFksZqvijmzchXHKadK6irJMLVw3bcIOVZ3rlu8JAvS7DH/1aFsbC/gScy
kNx6S6EuyrhNrev4i4HeVyGbreEW/5Ke/duUj23hgcIiPdimnvFQI6Wr2a7rVF8mPUAohFNuDUes
yTV9ZjgXofO1cHJb4eqfsVPvzMFNjCFyXwG3rD8298JyIs0/WArEdTk2CBz+BHyDzNrBwuDgZKzi
3+4ayeQXJHEQzDGuMbJk/lqtjqb8JbKyTpM5h5x3ePokhusg4Cwi4CC6BSRpDZqGC10C2ITOsTmj
S2D+Ouz0wBEyUaQjItWt31Hq6p9BDOv+CbulBEcqLv1wqFbChdUUXRRroencIyXAFszHDdBP+u+z
P7TTB+qZs+q85+fVB40AZQbvaeWd715cHlwyNIHCpwhYRdFiNfY90GDXJSp/kPxwgDi7Z+oL9QG7
r9Rp4fILNSVVYSBS9vsM4lzhN4PQp6MeXZbOE4Ln0bjFR5sJsdLnMkPCYbqsJuv9MnBYjL/yNWah
ez9pfz1+1/at5fVP39xdYuh0roqX1J+iogD4Orh2lB3UX4DLxTyajCrSgIFDBR8BMoap5lRwKC9K
7Vqg9IhJciQ58RSWiNHL5UsMmpntmz+KNegi4YxUBxrNBH+9EjxtunfKI+i6/shw/CH/UF8KV0nE
EqTW/W2pWn/MeEW3mSwj751rl7cRTCGJ/efBuI/8S5OmEQY6IzGc8BcJOZCxiVLmNUSYeWly/2d7
ASSWCThE4EcnY9wy6ISo49VCtnFKryItDEJvcltNAOmDIB4/dnlSUzhiQTqChslJ3e3otQCFNwHu
o2PSzw/b8uVpHrEq8ikpa+6trF8qdanoC2CePM8Jm3ufHZFZHPzFXNU1GMCnfoz3ypSZCDzWNQqK
4tH7b88GZRQwC3zITLZB1KpZLQ0hHLD1MkV1Iz2W1awOoOG5llFFICiCn/lpAsAEG/xQSems6V/l
8/lJ664eg5WyB6haWcsYCLaodjECS7KY/ioWnqzG2HlvGContl4KotFQmKzgyidqjLzvVaNR+bP9
Nc2MVLMxXnb0z5S/MBvKgtjKwmB6AtX4x3/ff1KEB/VTvU106K6gPd/XeGmsy0k0J2Q385rp/dXl
hANO1dynShZHkDqwZVapJ5LyEnmwqjCrQhvNvnk4tn/p3ttHyAVneSXDA8t4JdvZ/Jrokv/viaQh
0LdvSzMZKZVIS5CbF+Lcu7rKdAnm0yrazofRhxKw3pM7SsdumT1QcY0V1+5VqeymFNssBGB+KxDx
L54Tqv9/ZjBnU8sN8aYSwnS1X98iAR/E4P4bwcxcAZQ5YWw4LiMIVyLAGV3Rx1EmrLM2l7ptdvd7
RMnlwMqM20qwJHsroC8AoJViDAJVT0k/F6gw6HaNfOfDtHIPvGuiPFyS2cCmOXLhVvg6at4lww3z
nTJymSvhSsZnJR7664VvPX+G/sD24M3xSqJ/Uukc03NR19D3S+DIKUsVMOnEuuVwdVU/il9J4jOx
q4B/rSPGit/RWhdhzor2EqYJcx6xVekFERwf10EeK3EVaD8gaCRxtcppH4Iyj9OteYvFeWA6u6l6
TLaZMSK1OWYUmi3OCGt9yXANWBmW3e94CL/+dQDKnk2xOruWTaZycr6f2ASZEuTVpzamZMl0xhth
tAEi/TwzPIHocC/af+cspR6Z6m/YzJCgx0ga5X4Ien5FsA0EMF1yvnka4amfXJWgwW4DnPqpK4fS
ikTux5UQBCxsGoWYSw1G9Go6K7erK26v4JVK6+UFAreTLWW+4ErWn4zhw3r/BOPm/rWw+c6BT4vI
31RK0e0F1zE6bw1usLxYMsx3efMtc/twUQqc62m/RUIZQ9XMQOTX65NrdssYPOCDqdYadKKiuXsa
9resV3EP3XgbOxrmuMMaSzwPRaCplFeHDXkZ54LhQUMN5IGbkmxO5sVWqryKafDmydVaS21GBw0v
rBolcRb18CJHttWkS3vNSxApGwphCbLu/eDrKyGDd0lrfL4uO8a3U9yWqpB722IRlhlPsLLGcYCo
jO8bTIhW3WsW7qPqFHZwpS8+GuoR7J9Xu4WonHuBriiv5CJXKJ6QO8brdHgbg5M7/GnHJvhmnDAp
ceD0j3pHUIIw9aJOP4XQ1JtC1QL+WNh/68IpOoLsCFFoMEgEUixwkJHHXusw4qxhsgaJ0PLPi11M
WHSTu/hy5/VJkprQEueLO820EVPlOjPwccxcfC8vlaHa/wQP6c7xXE9b9oNuuIqu07OqfkZe+/BM
tqQ+YijmCWaNaRPvi0w7SNJKdXzvzX0j9/oYqZDtm8Jv/rtIKH5KcdBJz9s9IUeZxAD5hlhuDM1p
30S90Z6/A4EIV/7qJzq7R1GMhufk4ubjKwREsF3M2hj9rJIc7APvBtKe8auACG/ko/vD0SwWXBTD
abPfQJObmj+NBJWtzFLvVBKt3dTZD17ZJHBX4HFMhP7soXkmfL81klOZ/8v6mO5V3Io7WV5AzPtU
fPdvuMr34SklRZostKS/MeQzYUbYxFU8IsRW1fZax5NU7fc+vZ0tanDLNgsvH3NXL+WHQjs9oe6t
ZD9fIUaeXGhtXq2DGyXDBjx0vNWKGgnlrddme0y4PPnkf/0bUfocgJv5jzZ7AlIX4ORLwyaMH92f
XnwnbLjFBTi+Co8i8p+53U5t0uIxKDRTn10q8woU60BbZ6mBvCw3H6Bi2oXNB+R0IDrjseAwXDbn
rn1F+ZXiraz4E/ohK3cuA4FPnh3XXvi+4EN3TkNt1bjU7PrIgWSWMfbY9z+xD0Fy7TlukRtTA+J6
Tajwpm3K8WC9of6c+UPCcf+JRFwV7R/qXTipvT38tFqUh925eYkGGNYYmwR7BDRBu7OtN/um2WWg
TsWCGPX+pwA0EbhGIVsNbUslFJgLnUU76FJVZDisl3AEHmUxKMd5fMK+9kWKXUmXEHZtBOruaDoq
230SI2IsUqDRayWWZb9aqpVJ2k36/r6yN9gD7D12Y3htt+d7nMxlACb5+CTD+Qcba1Rsurv9kt0u
OWASnN1NdnXv7RSAcKyNd645fOlqKW8lCpbxFGqgR7qzc55tYdnegWf7mbQA8dfuO/9DoY6ft6Tp
N3TLPXFKMXYAu2UKvR3bGweB4oN1XF9v72kzvIaQvsLw08F3EyDknCokZcc+TU1nUYX+OGoWG7OM
PsXlnF7aHOTXLbOIldme2fiMsxgQevO/MU+4F5dSKZWMqMmM/cyAEB8VRSiGi2mcVpNFZ/7D653h
04KLe8SzB9bchMBkj7jNqCcTvhQfhJ87azGSdbM2xmv8eDx7h1IhFMrvYcIEktrs9SN+FgethV8J
+ZUn5rNyUJeUwDxeCrV3kNO/bYcPa1PfnLW7C2y6x1ELUCJO3FyDVedQW27GDAjuWB0u+uQPz5S7
vW51LJwO6lvYrCQVmdpR20Ywm7tC03DTgacc0mFD7h1lAsCMMF8yF9jFS862Su0FE6ugYwYKO/Zr
wZqZzu5rez5+DDeLrKLWc2OQGYOlj3FybTVLf3Oj5J+8lu3sV6gDxpTxyCL0fuDCAJAUEpvpwAuy
qXbBc9bQ/kxzJSB9iAUkR61HBFjCEJNDNT2gIl4/1f9t3qW0u+k7F61nq0NjWTaU3AgP8k7/6isc
gTDmzpPl2wWpncWaokuXmMOMxHAdyCYRnd5gPBHsCRLKZMI18GHPg/uZL3rRUgRDdltmjcldH8Al
lDlDKSidJRL3ifLireFcu5DvBHMTgy5+p3cD6VmHMCiAIoxpMdwGTkGPkbaHMSFoo5xx4cr65hHu
EpvIX6VuCsVdcpgo4rgqp50Sxs1cvNHg6HibQLOGA1g5MTWer3fkUbOT4e5+a6v02lsS8jHz1EF+
+1CSRXG0sCh9iUXl5E5GacjcggNNY1XqdVz4Te3npEDtDT1LJNaNSTIR0zq3QRkSibgUiAVQOyT7
rT9rvzQdehcKIxQm7U1wpwNYnu7S9rH0Nb42olUsuAL/Ev1eosOuW8v4FPonrzwSxFvo/ZYU4lEO
RD2NlyuJ3cIUZn/qQvi1G1hS3GdW8k1mUFjJC73DIM1uA/NmPEzvmqLWFriH08Bq5B4uIC7URu/9
JibS9bzOOdCXo9Q5TwUTwT4Z2niWsNlvIYnpwHN4YOBUEf8BrtYop4xsLQYg1Hsqp01ZYhOLW5ch
YPKODVCMvihEip26qNRCofmnRmKWwhSuA587tuY3iR7KEmyZNXuWoxJnx7k93x5Joh7uO/pkRaml
ik9bo59xYdkDf00WU9rfpGlnp08fjywfmk/SI1PYnJyXPmciXRI1t148PXAQCP+jScCWjBZmjw/t
OYTPhDW3/PElG7IblshCz1/1kP435pUtjnEIcbMNUhGm5RGcV/OwY91inY8dz5Wkbc675G3OXTFU
uZv55z9Me6m9oCAWpUsWfwW+NHCR1Z99r3vUFv3T5EuIJUoHzoJPzv0n6K0K+vTM5AEJKVCBYVhV
KC8f68dvn8Z4J63Gfw0WHUvHTPsEFqaWUkSBE2H40TlVJJO3xRHZjY4oA2wy45GRgO3XbbizIN3Y
PsI5rhtiKl/9xMPEaj+wMeEAbpigsmU/B+fXBk13lY9DXSAztiVXrn6FbSr6CEWd2Xk7YW7ti+ry
3LapTi7vFyCZBaC4iBnyTViS9mIwYQ8P+DXK3Eaq1lSTIvFTNMqOJaExwfEHCZXGABitc0AoF+xe
860LDsUCqekSN5Sb+xii12HcfCK/Qna2ah965sxTaCtFpy0+x29HqBebWi4nTLfigLL4CW91QapQ
SNPqym8785XFxE8kUlOXKa83jo45YO1iVfh1SRElKA+uE3gfZMEzNx6aNy0/usPPKyYWQyL7+3Wp
eIp/yrNZWT5BS8xhG0u8L+yKBUu4AtvnHIfVj8e9/pspXyW8j9tXesUp6A7pSBLq+Tn6T+tfhSOf
GwcOQjneTL5FaW2jzujLvlg7UaCFNyTMVvgiIc4cSzk4PjFdODnBXx40Fm9enoyvt1qjHf/CvMgZ
CqsZvpZG23u7Y5AXZeTC9rXcSgEtvyQj3jxA2qHyaZU1waWaP36MBZmi9A1HJc0nWFNGK6PY9Ofp
E3fdUcyGyAYMncnFEGmmNQCqWz0yO/PFS4LD0o7suHmf6XLVXe/nkViOW1v12b73V9m7mVqyC0nB
MBNklpNJjuj/DPg21QDX9zsYq5AR4vB9Bkq7mPlF2ZiouY8yltwy58zsJ3JoZxVf43ZOS/BAUCPx
XoWmNTQf6JKMWRdfDUCFoMRp7pCw0z5w30z8gxgSLQn+2kGQ6bAE/5UVV5tg+si4gGDeX4HRJ+d2
chs0fIwkrsMEjOXEkAFbthoRya10kyBJ3hSoBxWMmsX64FctEt8kQB2CO38aXCDjSAr5+L3rkw0f
F+l3h++cwlEdD/WYEN699S0gKDz6TFssACbPhfzqefzlYhKXvwIcusSkK39303nC5AdHlzA7ba33
b4qdwO8h0q0lUWmKDwQg+3ht+40zEdeE+Dcl7bo+v/umPM2WDJNocHSD4Vw/gVZGu1nBJQxPIYuF
tZT5crT67mj+BF9m6cFk9DiPYHzbYH/aUI/AeysO+p9ag/+/po8FmXn8nU6jvhxRJd1n9N8KLsdL
TzEgFbQrboCq2pHk2gBkKl38xKOlxMf4MdpGJbm002XDivSTPcCVIb0EEgle/OIwGmu44HMxlNkj
CtFieZg9z9NOJM4v9l7nyJn3olQrppcnh0F51ux3KK22cuzffuDJv9TFNvL45Dkpy4Jbq78rEFps
pYysJR7f7c4vA5+/4A1/LDnuYForfqk0ovRXcCj8nzNCxA4VCdxB/AcngGYRLU0jyVlqmgsKRuWb
bKi747J+FZRUcJnFFna4+PDBD5EStuMoQHHam2DRf+VR/lWkTvL3tc69gquf2FN//eT+TyabIAn0
C0pCq4ZINDz/csdf/3dipSW697lAWGP7inMUREuqK6reI2nTsiNcgrig/DW4Yzg1VxL50RyIp3Mr
WOsXQgoTcgLrX8A71P+Bz5QIh9ILxPyHpi5/I/9fG5AB6cNjzmmssJpoLX9Y+S75IBLE6CKIIVsj
cz/LjmcPLqGgnhPekQiOaULnbTQ4Q1h/fe85QIuIkwL1/A1eRXQh0xL4rYdWw7XfvImRfbh1Hced
Mz6hfemIS0wsB1wpAbS9WQTWUJLubc2UWNQUoNXUwZBNUpYpjgYPbkPc1cKW5Cjw3GlwY87+Oxpe
KsI9h9yfeNa8pCfgHLItsACYCBMoFd9VbyQAG+xnVU+ExxXyzCaIIOc6hiMp6bVEnLSL9g7Wv2f6
J1F1M8ZuHJo/J1U44qhPQHmcC8RllsKm1es0G2nJPIt7s2cESe64cOZq6ZBp89wu9nDmWeV+fiwt
H3dhus0H9J/G+eTHbPQG+E5q76p25IYPDFENl8kZe8O6oloyf3tSYzNJKVoTaRMaHWQPJyJ/p7HN
AKwvsoXyiDLHBQ1JHnRQjodptJkeH9Ecou1oXghLTzSJ1wyd8z0dY2pzs16QJH+8V+JaFt8MN1jT
mt8UnVkq/+LMJKjkyWOkrXQ/RZsbcWW1xTxHXUj+7V6lI2t3CcgWS2i6+YQCzjgGLcFc2NPohiuG
D4zGiVI12QIW3TkU6a7I4REkyj0VV3/SgkSsAC/fPfiXtsm8nyHVamLVk2J7B8MhDvfyxzBRrcQc
ftzt4fig2oQWVIBFbgjCTdszVEZZRulPprXdeVjXJ6nJB03SdnLB/NzKTkrtAq3JSppFLA+/4vPx
8Xq23c9ThW2uMP2uBwIFGufpKl+WIIJS4U9Y9oT3ea3pj43pVreGVKXfGfhRpHik5dtlno3opkNH
vTUDGgUuDxeoBT0zZ1CiIRcdhM9tR63IjfFQNhVsUcwB/grgeP37w5cGaqju1+aDzo+W3Vnvb6kb
E0EzZfQxfuj2YuzoaS44UbkmshmwKqT0rdF3AM9xYjcaQcS7n8czRT92OQqBak0AgvUWEdc3zDlW
UuFcDHgeXWIHizuwQeXCNsqdQTlxvp8hNxBa7b1mjRke16d71PmmJUhwPCijXUQ83YoptBgcwY0S
rOCHD2cc6DTg5R5xHCVbYGTqpLX6cj5JMomZ2ACFvGJ3Fi2VG1gLKu+VHm8LeAr9NH6MJoWBdIy8
egyL+1tIll1qfmtD4I2z+jloqcYXGwa/4yzmWXtW9b8UgRm0qvjQVbzTsommnsKsy2D8MlDo5MRE
1PGP5xlOBd0sv4Z08yPMpYuV0GG5DtnDlOBDSPDyvla7C1FzFcMfCuacC2DVfzaBzoJnpX+c4krZ
+p0uZqHtq0kQ+z5nHinPjkSavBN5WIa5OH4UBJjAQwrINKnNt7MggJ3c1wylgMc9LxwCCmc/c3Vp
rcWsn0WDTcFd2U99u8x5mVXRCDAYv+uLoBdt9E0rh/gEYNvP2X723o3dKt9vDAXisBHpkMuZ6j99
/YfthtguTRm5IN0nNAG4BBDcSUZulBamzjaKUKsdBFL95BGOkTJDsnO6sXsCP63jDbbGQRBs1VZb
BwsAGXZJ3E8F7cRmpvVL1vjhBGv42cV7dkfPun87nGpIlAlH1bUZSpvp7kbGntNzb3d2RSs4oi77
vz2hBossa1k5JAMfVTcpiAL/zWaE1yeMqfsEFYedb8j/kdaj2JjKJqKbR8WxN8ppU0a5vamOtVeX
OY7wCYHRfgevtN1vYQkt+9zIRRQwBs3lV59do8pvBKGrh7/tPvU5tBcboxaw2DK8Gx3sa5z5Q6oP
kD66sNRDUH/mvv8q+v14Pm6TvE4yENKRzKyt5ktEyiBij0SDk7zXFXjL9wLs7cNGF9EeUHR+6kB7
FXqGQrxzGP+ssZ/S9cElZd6HSNwzzJnyrhKt74fsA9KSKEg3NIAfPBfkbajCpq6mOn1K6aVWlrL8
AZVyst4jIjzaLOQxOHi07DjUB/Npl0GNgBr+pDEf5eK17eUtXB5ITbAMv4N2zt0TyBw56fvAgobU
uqD39BCgHthEy7jEpz+/xMkowkFpSqf4ZIXe+RgMoXZJKuY6entaizoabYdLoFoPwjB6iTr9gycz
Rd4Y3vCJ5+kRZGDDQG5Zr8iechL2/Tp6QKuQVFM4T/VYYw7FP7+Yv4lJxzahaDtHYx1C/PM1Vwat
rFbLKwoDO7q/u1DQsb4XESAzfbPDrantqq9OZTJmdxTTcIsk/YPZ7Pq2b9lsl6ovm6r/kSB512M9
iWsvIwEbLe+GIWO7rcUEItdO+DVyM++7wMUK/0Q5ro2ubKYWIPg6an7nk8s6Hc4CwxydLsYUgQGo
FVIhsWOUEw6pG5GvAAdMfOef3aYx4BFnzwrNRzzPbKk0tBnLXw02bEZ9oYDtM8TN0hBQRKdS5iZV
PrJHcf1XU/EbYTsWbkB3d1ScJuHpTcI6TBbiAsEFlZvsWG0uCnPFVgmw9QpYbu1EdQCErbNWywD+
NSpUbFX8uWpkj12CmSnN2adnu23cLDXocgGqOC5mIbgIlAWZge0a1aGtSheYCkVPYoDRrWG5ygVN
0YVqEEsm2FsfXxUNFbS59KW5H9bmfwNIJMTw/cm46V1wg3FoUnS9K7TJBsimY/XPZb//VrmlXdF/
XBhU3imS1/bYtBlNmgfEUo1XLoGehsOewHatYfsz9lY3DIH2Dmkgp3T1QYvRqrh8FXKu7ATuqrHI
K5Rw6FqeOxNe8T6C6jwOcjyxRirl9/lBYWGcDobjZ0VHnaAZw/kKgWtuOcVTO8zXlc9E/NWg99O5
SBEs/HHSJ2ZB6sXi03ZTzivX0qKkBjC65olvaoD//NNvZUHymMC8IFj1H/Tinw/49tuG8w21eb+I
mDFhq62KVRzSKKN5l/45t60gYDylT0bDkAOxZqNjfW2Z9PFiX+tcRowiMy04VqLAeDwz7BrQACm9
m6mzgc4GDYEVNkad6/3B/UBAESMBPqHtT8FpAqAGeAF4OFRyykROoWLbYR/Ctdlm53cpPBDmejue
MFquz/kPSt12mt01xLVfDdhal24/7c7COLZ6/dS3AAurcbsazXpZRYpDSq5X6/nyR4npQMZAg1HX
At1mK8bXYrJkWNrGIJ0zzhUTTYjZ6BsiIZGP7AaX4eAz7OBP6YHF1B8qFh6zE8ffhs6rS/2J0uKR
EhWGwgYBG7tHTVgnTi2j5TMWB35guZhXEZofxKOILrB560nbygBilHOw1TRbVmF97DuS7zyV+86k
UpK0/qeAV7zbgAzOjMOYobAehC7Ud2qkxGKrmpRU0OcNCuVF+aouURigftQH65+DCzMXr7axCr1T
JNQQWj1p2a8jaL8CRMx4BGEZEhwH0g3fWeeovotft3cPEnyLBDr+ggdcuaa4rwmo4IXylmtFO54O
lrYbJd04lpsxNYjDeZ0SGeGxf8Gafphh7OX5sbyKvev9edLpDbfJ6CTdARTTufiutyGs5f08xG0A
jw16IGN0B52t+NRBsNK85cNUqpC/AxVBgC+bQt0jkcb+Kxq4tPSOM/9QAh2WSE0Do13T+Sw5opSA
9driM7yWCpeYE68sJw7PmozGLudMLgym5+IKyUKRUA2zb015QZg+ngf8PPxeQwOVmsrMRYch1POl
nZ2mCE5Sn61VMvMmU4T64NnyOVRLVHXb/aAmFrKfEzFJRfPk39DRZh6EFQl2Y2RdZ2AqaJQwZOB8
CynBR8Ah+WxGFCZi29s81JytHmh6QNM4a5U+22RbLYh/XeYO8BVW6LSnWj5XPmzgTEw9hp5e7g3h
z2vU+1CMQMmYrFr/XJLKU3Up/gGkyehEKbIFgidpjGM+0yKRsA3DZEjMfDigvfuVYtnPcmC83t7A
HLqJWO45I7V8sSKlPaOy5+gNQiP06jZ1ak0ZjoNEGv9rR1Mi2uGQrhxg4ZoetPhllkguOu5Hx42S
OT9Zgs2mRIKu4hg+wvoY5VR2cVEvwKiyC+GWbKcOYttDRwjs8VRViS+Fih890HgA/tuE29LWJ9Af
pg+tAF7srTA9DhPBh1UyJl2bT8t9Q7aDvI3+DfUZ4sf+E9VQz6yAWCrpGjQ4YXBGqN6zdAE/5ym5
aVIE1Kn4Qn6IEzskT5tvlpvvCnElZ8+Aa1iaRM7H5e80xyZ6FwoERINRtKZ2sJXpE4Y2J/NOo6OQ
lXUh6s2WlCVmfc8otiUEXMbKlFQgp/uy2DoEDfWSGmlYdNr9bgrPxKFHCZpp1QIdS2DWnR0Ce6V8
4LTAxV1ewB/BuOK45qshxgXaev2saTWUJGDDLOF2OVqZfa9TABJe92qbjKcuG+dqZ0dwY9wKYujA
Pw3587P//cbm0+2MyYIZsQPoekmDT9fBMl6SCIT0r0P3pGlBipxlO7N6K/ej3u6y+G+IVzJl67ko
XDhbKkuTLO8K8jqu1TewAKnaYEwHy/ZVAuKBspClX+qUF46icf7UUKN6VV8xU0y5TsaXaMTxrg8B
cPkLNoiSRmZ+JrOojWQQlk4uxaQR98xe3DYzT72qHfXWaJYR/xW45yhw1pW4FgcK14BYm4JsrXWt
CgXiwzK+Ms2b7sYRi4Hoh1R7TUfOn0OeOTE+EvEyXVduy/G7P/q2nj5QEcX++qh/vLnIRwZcTC7H
X66nj53IxU0HFMmfhHMbS24zhnjL3IxGRiXQXaVZyFzwriiWLyPr7wwL7vkowr9SiGF3bIBhKGHe
cSysdt6sHqw1Ba9B1DI3d6Dbijk9zlaXkGVRXzlwn2YaQtSONmLUYYzk8MDEFNbGjEln9v/ondoy
TpfPRLWFDkGU3mqbeouV9IhWIYJxCWxTVqcpdHfkA0X/sdVh1Qhl0KIL75tK2ArVgE4HcokDtGbx
Eaz32Wr0wNYak5ukwI7T/1omTxyq94xVYvm7C2Hqvhf3waZcB1jQG0exbj7/PJSz37jUaJ43pEJ7
6TUiuI8+3WDa129k4J0/mzwHm2s2gYP6Ic4DE4gfeCiHQKORuKItroqwWqkCGMKVV3Z+C/aG0CpY
J0VktnEjhSv77wKL5YNwF40c5uhz8NDJpdPu2lf84TY1JrrkAWjbb8jkvqB5jv4NP9VSe8TIp3yE
KlbRHl31M6OXIvdp6UJYyca3XDbPy6TXkBx0Cmk4bLGi6kvsrfR0hSTndfW9dWU2STC19eQDTq/p
glaA42IetUseO/yhwqJGQEF2hCIsPy0mAnu2x6FibFSi1Brs5QH4JQG+vKTcfSO6/PK+RiZ9Je+Y
6y5dT6sG+g3Rk0Hphj5uEjW0qDOR6K6nbzPAIcRmJg8Zn5aj/aCPUSNLWgyvGWQ8JoYa1i9kBcaq
nLALf8e5CZA/NqLOwYlgvrRg/Trhoj1wmc49P1sa+GHQ7TsH6pReu6gQ3GZCNTtW0NqHsc0UhcvT
ElJFxP7pAUGTcoEpgxpYCjBQpd1PDP15m4UI0VCKWsayEYjwma49nV8mHrzpadLCC5tYTU1Xa6VF
xQYICM9zPBjXGItMJR0syfjPXn32agqZ8efz25If6kRfL1XSkIQeFFiIavICdHcI1JxGzA9cYa0s
LnrlIGIYb2go7JnC6pTo99wnfBs96u8+BS+um4iIf0Qx9KAJo+qK8zXAyRdEsRnDxxMnHkLor+61
3LWkf/aaFxiqb4XtB8vPKuEmTVlQ80/jkvUbxIuIlTOzGyP+NvV/k5bbtq7UpKHUySIA3HpvQWZG
prf/Iajy5KMDbftCI20yE5mSVdIZbEgrFoOiepEVi/Zid5u2vGttf9mLb9YFGurbocJ08VXA/qrM
s6UzMIaWz1XLRTg1Y++0nX7bKnY4MR+2PLLJksTbN/ng3a+bPqdGgbdaDmp8pQHSKAYg6bikALP0
npI+0HhbgnPg2s1VkQqxdbd22Ijd/kArOT8pznMqnepHfV7QM291AkYhCE09+uk0LJ4DQ8E0XgP+
bQVT+Pi+F9/z9vZa4fpZc/CUofToZ/VyYloFj7NyV3ejcpVVmnhJXK8AAtCfPhvpnVSL8ZB9Ij9U
HH/++Z6fQJ4n/h9STrtscTkB+DA0eSnqUvn28gbqrFJvJXp/8SocC/EjPgm5fLtMchXVK60fy795
NgdPUvvbINpAMJaAaKxP2o80azBX6XF6Rj5jarA0Cq9qPYMRurhsLOnBf7O2Whv3aweeKA5irCUB
2ndMO8/u0cz3K5ZJ/PET60a5CnlbaWghzOYZMNBCuBEihkJz6VkaF0YsySZS2v3ZaI9kSAGUjalR
xckZYbfV0BiVNX7KtPlzK1lJaBqQdfdUbgxbqRFQxKY/l7H3t3PKSHiSJPAQygV9L3MhzKZ9axyV
aKbTbeyd5UuakHyeQlD5EOsq35QbfsIg99gdZySqjo/bwCI0Vad2M/54jhSe9627TUT3SjzKwpKb
Fy0aexe34fGhUtnPu0maIY8DpOTxeHfMjxUU1xNfWJolStNV5jIomNLzuPU6c42AaiXU1kzKB46R
8vXVe8UuUh6a6jkYenw+6++VBa2KJZbyamoouRYjJ8+ckWhLKSxA9cX3umR4MRLuWVnYeYrNxiBv
1kezHB6dUiVVF5BcAnTk4NUBfZt+kTkXmkkA+H7POz7ntt9+nu+7ME3YLLu4SzEYnWExFo6n9VaE
CHapuWkD67m/0FqCs4F0rWMYvm3o9Rq5q4bl7Yy868CdE59984tSoL8Am1otYEWnBW/DtlkGjRXi
9CpLGEcZ7qEAnhOsp1Y/kPgQ+BjsFIgLOrHl4wT76h2O74KIFO3ZYR97xEhXwqGoDHb1IpQjnCrj
hNfXy55xA6YxuvMS43p/GvB8RW2BuypQig1X+zPrYHRhzYxrxDmD/SNGYhz0aZcch4K3QAQfuJiN
MH+QukBncSjjmBYp4iYSo9nlb4uVhOR1iJxMWtVownQNPXkgMX3ak+RD6pyzvPbxUsGXYxSZGpoB
2tYcFC9QC3ByQDIof2MSZjG9EtS8u1dOFz0Hbb4LqXNNGR3z+JojhgklF+HNNzBAzpkU++XkJnnc
j806IzDBvfcrhzH4bgW5sN0g/JzSFbwzMKzUPLwWtxv13JkDGUfNlizT9AzdemX/7xIc+JqNUNbY
IUalRZJvjvtAZMfaa0wE8I6jz0hVrRQWDad80cpRLz6gwrlTk1jqkqPW6M3UOdZEU4ZV+PEE2ztO
G6Or86ynYABdYJLp0YZLX/0YY27jy0Pn1bI6QGgj9s3v70nNycEjt47Cg5H40i5/CZfY7zEyaX5M
yr49Jm5yD6/UKJSMjUEHSkfOnj6nw47psEPqArwHXBvfTDIZ+fzWJWzEGW+vw0BLyzP76HNZzNxS
RC9sVfda8zhHiyXRtT4i73vlyMseSwUEY8DrgFySjMHo6r+Licb50qRyeVUHdy0fDUrJ4C93u++/
lRrdQG2Da6qvJHeuou9fZJilSDkSRVCFYA6zEPqpzZRqWfQCcBYA1uzx5DzonVLg4n9cNlUO1gdX
yYTy+BGBOlCXMFjco1c45wfd15OY/9ytnbNqVNJxau8oTazRbsBoVhILarLGvKUZsRb04wftomKz
ayDj/XUwYhlUH7JwtiqiKnEa9R5Se5gHFtyfAAlxp5g9+i+ALIDjwFNEg4hFPtGGRZW5SiY2jtee
bM7A6CLOCda5ikI6nCXhwJrOcJtpvlAyIHI0RvOohw0ZPz8BUqeZ7iwzaT3Q+MvvEDT3Y7GXzfVg
ASWjWn5Vu3zUEWuE0ajT/VyCggLp2DmEruEoahg6JnFR4pqwiQn2xJbzS86nHgDf1MKvk9ucsSMt
7NT5kgRPaAEbjc/xRXS/B9y+D7SBFvfZH07LhLF2lMr0hCyOxKKTwSPp1qrmjMyEpYQX0nposQuB
2aipg6cwyGua69HBMX4HscuQsI42I4QtdJz49h/XK3SUf6xfxG8wz7kR1yCX2EwbXqdObEpnFhbG
ykLSGQPR1OfsFMkH9eMYae2dad1j7GaUML0s2bxDKcOW67BOUrVwyOqdmTP3V+NHYFRE32TLH5IX
Q1X6TDip/WLq6LABN8CwCpyko5FF0W2NogClP2TNHjkI160QEo3XhwqEOHtpIXYkFDDacWoTNKwE
l2+WZcl7hUHR35M4lnTSYfeIAgEr7ikbLFuC8F4q7IGCJvQQJ05sU6bVpPLwKWkiBxtNaa3e6cOd
NLrH9ZhjOZNsjJ+0tXm8DfFD0ho6gQfRkRoH9CUr4zYJ9F27JZXWz4nPfGAoUDwE405+t05YP6c1
/NEBuKUTsHio47Fh5xMOrlvrkLJvtnabRSB+KxqXxWjotOHs8U3o2XpexhSufradwZltH8Y1OGRi
rA73iSmOjkoPwv92OXgTmrH8/d+x2rhxY1timp8LXu2wQRWqg2cz/ndLM02pT2dY5Q75+ILmeL+f
k26F7R+e04E4ldp50qhoZCZzIxKySWfQ/ceIovbME3aR7pOPhYCI0vX+n+xIdAd3yC2T6C8H/orn
S5CJ/LNttsjNyXImWFoj3U9Xyy6DzifIRcfm6iuifBSkp1+w6QbGB+wLK/zgl+IwS3EelDSecsJW
P2fDyJiT41+ILFGDCfY2lwl0xbbt7CsfwCCw4FiVHUtugICSL0T8DSlB7dCY60iJdmR+wnC2Ewrm
5SClJajfJA4IV3FhZXRHefSi8OB2NrG3cfrR9oBI3nVFZR3wmcMY+zBlnELQ0RH/NsJUvy7xtJfW
3tZ1mFak4ou6NT8G4MA6RHY+pYEggNttnAIY2rx5fZRLAqeZiHyWYHSJJ2V9mmbvJCeqwgRPUYWG
St2twTMfbi82MK11z7zMpZ0C1+jo/kxvPcY0AJbwzv6SJxpJqNO7G3jEScT9+rsHjI5nXpPL0tKk
9hh6twNBeXgCH/6/h73re0CcdjuBEIpLMfpaoOrvpAUGMnQJUHR2Bf9SO1mmHU7lYMZvrEULUW+D
+F4P8LuD76osCrTbsWk2zeygq8AOIi71fY6GueBaKOl45PgrRRsu/QIonNCCytD9iE8Td+J+wQ8R
7XU71ei0kYLZLyBb7MH/cZX/SHU3uiP+hdJoXj6EBaA1ZGb/Y+ulsDscjHpEk+Dukks4zB2duvHX
K/1B4lYm1P2y3o5vKGtBf4A804OrBhSC2AsBxzEYPonzu+rpQ/cruPO21uBKA2QNNV9xGT+8dR5S
lQKJWM4t/xB2xWb6AcBatpmmbqIfs/uN5dHD+4AO2zZz/l2tAtvgFy9ea7p4v4qP48XYt9Ql0yzu
++MAN+9BP9agzdU4AtRGCN5/pqSAQIngpBuONYvYf7/YrA5iZiozx0s4Q1mBFVtzo/rvJtExmxcK
pxgIfAFV5/WpD+Z66tzoB6+kuk7EFb0RlfvBhOXJBJ6q79bKQzX97YdzHSGTVgWOS49gkW4Y3OX+
MU0cdXsRjF2ElE67ES+8F9lGZCRKCIWlEFlP/tOo+kfqG8QnuerdnwkNFo5rKY0juNnAdiR3MR/E
b5sgPfKcqJfZC2Gy2rN2WfLXAGtEmXIzM04vRlqf1nBmpEUv/5iVCpdyxgNsT8mUZs+TEmzaOpoi
q2RtcD2a7wS6AxMP7IaZSNd7ayGuiJ/lykCkymB4fFAgNiPZ5YKpWnbSprnK37IP6/d6GwFL3iM8
+ekJZE+kbdbsZyTh95TPMSEeZqzRFaj0xl7VQsiCt+AbaAjEtqvJuHHbHmyuFfRtReySrmlqVqzX
PHZhRh5NoJE/RstrSjDqniMVyB4vKbTtarbSKFUR0djfuQG5lSyfuG2JLc1Yhf6vcBeOwLwinZLF
f7befzPSt6XeL60Cfwcsd5hza1cgiBvk9eplD7qIUZ8Os6hNyTHmkwuDmkeJT6z5szoaeP0aUznF
yGjKwkPaurFaWgou1SLhMfVLnndVxeC1OzRH80kfWWwDthrtUzrtVHEy8Wfx2n828Znm0wWvFNHr
Rypc9AuVBTMwqP24P05IEgElyzPlLMeSUlY07h3lufgYax+EOGZdHeAQ1Krjf9RrV1HEfVuxli0+
TYJpkqUs0ZYuFF1/jFoTeG/49EUeXBC4oi1JXVzh+YI4x+oZB6sMR9qtB8O13fUFGihNDHOwR3GT
gYBU7tBwaT8bJ9nSbPeRgZX8iFCGR1kf162BsVzW2k+9PMpgPeJjS1tRNoEDyYZBI8YInpN8McLy
BUWGIAIReMSYlMMeHnJDHm75tLoLy4p0D9DSjE/MXM+2MG+UVAY7eHBO4v3WDYN2LBKDK45Q1601
ouRFaHWukSuc/HlQccSjeZzFHNX8Ovdwuu4ZlagcBfSZ0jx0D9zeNzCfEHSka771Bj+ECj/dDiBB
3W+EWAUt71NX+Blf5cTSHDI6E6Lx+qrEIu/Sz9+Z8ylBRnLBPffAbyVDPHo4SjxN/mQOwlYLB0oi
qCHO8EQCbNEnpppwknyNRaDWVBwsCUosvouLpz25Eaz8C46m7sIjBclE7br7eVw1sjqqmdECkvqw
kf2MUbxxjQOzwN84jLfLRso3PJpHPMzIFSa8I/BJRLsTMTFFj/YeHJ3QZE0OtKwsm2sO8a8dgPG1
Slzv4zz/VOBH2T+Do4NjyxUb+bUqQslJGUUagnRXU5H0RmU5F5+qkk6PTVWQGatPQMeh5I5gR90l
kA99VN+u8fUqx1A0fmtPd9TDhK1/UJ/SKutHjqNK3G+5UaEkwv1m8uUQ8pjMs+a3GF2Zf1LWGmGN
GkJ79LHaVMhJIRkaIGSymHxwWBC20J4/1tIRK8ZZcaBbkamuaCGQuby9lT0VRxzt81yxBWquc1EN
12Lo6YFphhzmEjJiA6RP1p/EFJZTAHmBBhGWBJT6cmkGeEvKgrY9BoZQ9SC69k/dE5Id68cQ3FC/
FHywA+dvamSSCKjNOzAv9sLxXJpDScFq9cpfhc6xB7V+pMfEzH3sZpUBpTy9SePauBS90eT68j1S
IWRCiFh1ra3aulD1aphut4gCbQAqbz7p6Si9Q2xGUdGSiSEva6gdgMIXue9qKjnRUF0eWPtLZ8G8
KqsKFUCO2MEuU0jNrEI3PnM+m8y1dEWspk49YLJGAOPm5bD3TGo2FxG7wbXX/myn4II/nASRwO6r
pkreRLs4NpfT2/jM8gZEad7+Nfa7olo9pU9oryG87AN1we6GRWcCYvL+PfudUrslzqATlwB+sHaS
Dt8VR19Pop/c1DPswpKGXwN8GBgAj8mXMyqReo/IhXcIwSV1k4wwL7S2rl7e6OuawWsbdflgVk9j
P4ZttxqksQwJFdJqPnKAEAt+bqtUYpzphR1cmAPadlygO3FNjvtLmSlrie215Qbi8iiicJK9mQDp
auAbrykBZd53gsa3iI5lg2IwfVYcEbtEJSJ8DX2LycillB4RnullRn6oee7xZnTyrr1O8xHspQ0A
K1eS/n0hqmVYm+KIAvuO984pmeHgN7bIyU5VSgPkRSO5kKhwGGU11ysWd5Hwu4PL/entX5wNpLDb
DKtJUxEuD2gE6SQyPsO8Ofn9Y/tVOX1jjJJ+nrFUpz1Clg8jlfD1+3ZbtO6yC3MhjxJCJtrmGTLp
4EjvWgO83KOBV4yIO4DfvcpuGYctHS6zuhfOwjRP9vjGJETpXWzf1J8IQZmvLOXgYg1t5te5N7iz
GTd2CX+hZB9oE1/T6HZeTgJu9DqKStFSxPLE/QoGHiFgvjBiHiGSzrFgissoTMa2xxBksx58XWUv
/Nh7eDdveO8lpuqiuoZ26HJ9mpQnbJ7c8KB+ZdTwkPdLR92sanKJqdBVEOnX2b3MmpmfD7nccAlv
uAs8bUsZGbpM7cpyXNImwG8+HrZCwYjoejlvhUD7tswAC42qREo9o4qsysijxQwGxXHP8c5IJyzb
DR72O6nhnFROhmYCGSMWntz+L1qMlOtGIm73YGZbs5mcmwKqNEZUe6s2KsEnpJmaRvOUs3F+K9We
Wu/Qw4/fCm/+Bb1571plWn6KhfJ/8k9y1e4x71ol4rapJBD/lzSA6ARNlh1n1wuHRm/Ni5DEpHVK
lKRWqxFCGYyJR+BSI5A524Pzeib/Yo8+x1uz5m5ZijWc5CGu8sYLtv6lSWQyIPlqsPVbNhwomI8M
fzHv50TmQl8xRZzr3KJhTbH1MI/1KsNxxdwuViYYJETHHbFjKrzeKBGlx/xmbfe4CVJLFAJiD7ZD
PpL0aWYoQ5Hm/W87OXLPlqN9QyMHe9ygBcMsrdfcoM7BK9/rd84lagTYVZIazF7Ra//wo8oC3k0Y
+Gtez2hNVxC9nQabGa/unhGdB4h/90tUyc723jc7L25/hpce4WpOKRI17YjD7DcWHL1WccMYDhe3
K910uAnAaveuRXOLjICFvogWDGonH/bLTMMmG/1Z9bYYRdZvXgl7keI9I9+HslBoTDK16QkQCpGd
YXjreY9A3IXEPEtHvrRlCuzdztIQb3d21sUbbwgAXuu687R72vBoStIfCWywxkZjvzSC3us+lTi2
gmCrwIm5fs95fUL9S0tqt70A97l6f6GKqsTRQz4EMuJZsBX5WT8pvfcN5DR+DW0cQ+urJQ2Xz6DJ
x/mgp0KznIx8CKoaCFpTPMvh10SyzB3FuAFnaTzpcd5SOtIYeqXpaRuiz1pGZsVfUF5TejfWPbDX
FIbOfWcqibkk7ITQuFW3CHEWiUz7nvSm+4/RUiFlCJTiSmH0FvqdTI4H8wWYDvSqn6sfwvKcJzlx
LwVFYap1sTd1RWFjb1i/2skX3z55PIwIe2MVfCDOq02QawFnUUp8rTXYQ0M369TaKHbx5yKrkxcV
oZCA4R2/EbCk2eYtj8jQE+aZoZ+mlJV+lHSs7pl63hOwZBcNPtvc6No6fpkpJ1Y1M9AXjAVjV0qv
yT2k7neyliosVqK8h1ZnuOXk20fkmXL4jQ7v0wQUdP8ID5tep+vfzy9U4JqjcjyQfhAD3srd76o7
33nRCgh+KiNzkBPrawXY1GkS2nN3fGloqC41IBHR91OfBedAJbGu1p+h1X+CGTE7nuidz5TYIapZ
MtvAMxF3MXrg/gWhJLEN4yEvs4m6lZ1+Zuje9dMoQdZohmDwoItLeNzH1q0R1wG7JQYT2lA1xE4H
i6zBQtkx2W3PXcWZns4VFIE1xrv3REZlQ/FPa1MCe0bfRp4Wv0WhVJTcmIsX/GVVwfOJemkVogJt
nKaSBS1hLW8E84uFUOTi93BO7TMxjfh5UCwj6xKZK0EfVpH+l5HWejPRWl+dNZG19+SVKjpMBShX
FEPdWAdEy9qe/DaWcAXn/pj889N4+zUk4E/9TFbObwTz4UO1OBM4yQa33df+ftHncEuU83c8j8Qu
KOLtZ3vwpwvUo+8CGiZdtyPdILaGOR4zSjtaIUHpNuX4x1Lga3EfNOQXO9VMUP0oD1rKhO3eZokG
MLPzE4BZidNL4rVj8NhPpN4RE5+LsXWbv7OkqGnVBpmNSeCOaG80ofiBgL1ds3kH2NFhj4fX/jR+
ek+LIAaLaec8T2WJbJ8E6VmUoSgJ/d2NUrE3eT8CHfmTnKssqAo5RW+xZOzs7g8wDY/DZ+prVt6r
NLJWsq1NpZSZ4Dl/JcilgR/aMnlyqgkeNWdUlJTcnu6LQq9JwgKHpB6eqRJiEQJGFSY7VcE3i4mg
X0RXnumwMFeTeFsNVkZrzDBjZPY+/ic8BKyjbs023uta2YmmLOjW+S/IgSXwH+29ba+LG0OTLzy8
/KlrPDHjDvxUR3dlFNoaRKWWUTS7/MYYzvyzQWqOvwnT/GRDRy/W2hq6fvLrWV0OCYqLdkgqYxTU
XeJTeiOvNJEGmNVFSEn9UMG58bH/vuAm7eyeWuqSdwkup9jWSb3AOG125HdfNDyal8vfZhV6/ZJt
WwAba9YaDvb+Jl7Uc84Wlm7QBhhG9ZFMGzPl7JAvB9fso0bTgQ6V7+uAG8/Ll6JGAtDaXsbWMqyn
PrhH8hDg3oM4aul28c0pt1J9Cx6SD0iEdbe7BCBGFjJlcdo0mLAbe2vuS3iFWBvP0WQLPb48+EPE
M2vu+eVv1C6onFS2x6e4gA9EU5Z15/RqTPDiyFvMgYP+oigCHlzAsigiwcWWYO6IQy9Iao7mu18J
jS7JLl0tzVQEAPyzVCJ4EZLSgQ0d7hpr39lDeT6bPGSzxB7vy3Jw4WwaZbxRFNCBcbhJ0gkfrAYH
1EGmE3lccgAz/ccFw84XmPZSjbKNRoNwwcQdk/HHm4/jTfNLfNDT6KGwY3o69rAtw6wL0EQ3g5jB
u//1UPdQYEzNA/wkwBfbeAUAOjQ5CyQBTjtvD7udHyV5wYyPihm2CDB+CM0yYgJinp068j0AATwk
aFcxjRX5gE5SA+2pL9DRMDvFq/zritWSEO1juaSaP6nVftZ0xobvEZo8IVdJBtQG154M459Zn17A
m0HuMa8yqemC9KX4Z4rFaOlN5ZHypebuNvijgPDf8ZGpPHloyRQj61o1xe99F8+5WXiPWCFnm34n
N6OtTG1cY272/H+IVMnAUgm4LGw34n+MJixFrGfg/VwnhoMBCivnAXzREtkIrsUOdN0xF8Jw6jFo
4++XBR1B2TPMFlne3bbE5V0ILEz/Dc+tJ7Z7d8vmpmrbWWrfnFLdeM3SCfxf/X2abSLFmPTG5wVJ
ijz/T1cFJykFfbUrGgHC9o7ntPE5hkU//VYjqOTnNxkXe4GQEdqKV8XFgJbKqmeJDFwzbuP8NW4/
D51E6mRp646KJ11hgulw5x5K42/BOcs+1HZm8mc5Pd3boS8LmxjHsK8TIp1fZUdPu/8DzHjasrs8
IjZeIEmgmydkU5DC4AZCCuUbet5YQtdZnA7WyruC
`protect end_protected
