-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sHN6jC4FUvBInT5BHa4boinkqZ7j2SSe4rHmRLnShJXYQE3RL7f24mW/RbNwZBM5
AXfzrGH4fJszb80nGpma/ZXiD9LXGEjhHMzXLUOWzfXDiAsQfJEonNYm+n/c9T6h
LOU9TrPZHniQM5k7YHE9/QqLXNkLHcsGeLgdYvOfe0A=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 12000)
`protect data_block
jPm4XH3E5LyziA+pGz+LHHZds+TcIztWpgVmfYmOJf1jpdS68ejmRq69CLE7Vq63
M5Nhz1ZKPCl7XinktmB2I47vsz06h6J/dCIkzMHhelT0FnMiMFBcPHy8/XE8sxsN
9RUKUy6g96ocO9vFkLCVKEKbPX8ZqyaeQDkp2Kr+jEDz0HsJQZpSXmicK9DEWQGp
yHBEmHZZs+b91grjkfeUdjmpG9Xxz0XFfVKfDPIAnnpdXj46rH/N/IQMgEHsrpiD
v6n62efR+UEr8Q8uCGmjZAt29apNpnZFOmPJWVMdfsOoubTSe1l1Sb8pn58bJrmy
qCVEUjfy+vf5MjuZNCo8XxaGhzZWPzSJ+63WTCLC+p943C+OkNIhhj77nC5WMXXX
YeStTu1lrn66Frjw3h+Pu1JkLQ6kZPXlf2JDzpfUA3C649963S2kDUhPmUFUJ48I
eYzFyUBoh/noPiWacgml+5XUfkKfW6ig2fG55YVBZ8w+1QjNOIDBC0+RySjgV/ec
oeEicKSlPHJmOeEaqwe7vN6yVHWaDGh32I/+ZAFwrPeAHfRo4yoAagg/SDSyCsVW
xHyHuqxi7R3LRcayG4+mQb6KQOP+6a4i6edDLmG96+oxovi7uliFb8H6SQwF4f9+
as/M5wkWQbOYMu59FL9lfDxLGqZUNdodD6neeiO2158IXeUwyvgGoUCZ8AFfgInD
Owd6IOROwp4jIYK/4NlNwKSjIdJrMPPa+0tebzPunn0bTr4rVboQ4kd9vqt+Mxbn
tgiPRkNr7j6pkAD2TqhX3lUnoOMLOK9QG4+lDAI87nW5dbE1Ah3iRhnaZiG9WDc4
Cl3W5N1+NotxPhLyN+5C9pRDCbWVYTf/ogh3371rHE2HDU3jqNFfFcHoNFswQy72
1snFK2O+KBtcmqXWuoFzcb4XPakJo2FN4dX+7Ne6AEXLbe0ifgOtFNBtac6X4eNA
X8tdUItwbrgX6GRrRdoMvhi5q/ZYb69W8PYTALC8hfnjz1yhBusBa9H6gBOJT+X8
DKOF+14J0H5JS5nCdTu23Z0VWrtT5RdG7UbaORHrI8lacZLYM8UlL0VbbuFLkKE+
3BCE78mAls47HRLB72W3MpMzc28EX+5YZpPU2gcJOj6jL0ZK+2VlH5uzsdcfsuXs
Ar5xjReVqEkoYWtSTqGPwn8mzaVwLokkwfRTpLkoL0fLNkWBB05AuklFPojapAA6
UZQ0NR/s5vhN8vYqpcIB3PCgcu99TQu0QSs1R7B9h3LaOnC3mz35pk0/urmvvSLl
0V0ApasoPZzfLlqYljh2h5tiynz9O6WMnsf7uEF1xO0AdwFPa6rYRJyw4Q5SOwqw
1d1gjCwmqIGcc2JZcXcqGhkMSYesjfc1dg327Qee59osOmxScKeNYHYYY8QCvsvF
4AMQ0n2txt8HhIUjjQ5B1DwwhLrSkO5RbHqDJmSrcaG9ma3Yx8oBKwINO5lX1Ty/
o3iVEf+MvJFVv0tThuo4yWAUJH1gq677MJzTgmb00R78PSdYibl7vumoanoIqMJp
6S7nUTIUQTevcQtl0+y8vaPQfpyC4GiMa37wCk0Ob1WOYJEx08WEmQSc9yHq+dwA
i+fyygRwmppmrnkvCxZGbkBH+PJeef4yCavi9QXhpSxlnPw8WGjsMhkgDp8iu93q
h7vO73Y+oVwKx6iKgSi45tR9GRbG372zUtOHl7Ssfk6dIsuurERhMt6xkxCCLxHA
XSPdZbWqqVv45QukLSV8KYpLtq1UAaqtGSjsjyBM4KAUjsOfOExc7j9NxL2cVMUB
E409ncQDcYMVz7sW2O19da1v1ppl/3pDuS0lm5q19kikP1v+VhD64xfF2NVWMq1M
cpacb9750Gg+Ik9KVOUCJxWATubEl513h/YFsmjInTcltiBtYhTy21gh2qUoa10i
ls+owretDnBrc5mtJQz0hPzoRg4diEkhnLDEddD0oCdmu1pHQMFGhGwxDmyu/5Xa
NvEphCG1bqvgnLJ1n5j3MHA852uaSTeKr2+jCrL0lLCnfWZLpPH+xm48n5jsXIDm
gqCCUsDV82IK+AcgAstoO2w7H6UXth8fp2hsIelZiplxR97CVbRX9F8vU2GX75gU
eCCEaQws4ogBWHd1WhtkKrbyKGXjuU1H7A16ZfES13d+uMorXSGnVnD3YugAUUyn
a98aL7VGUQhKoXFTmovpXEjoAA9L+urKUp3WNAkIYJrvKbbQj8lBtac9dc7gPbHE
BwEmzUwQ30d/6vwzn0frglOAG2sClF/GMgEayCM8IPWp4B2+hOiXw0VkKYgLeix6
MYNJEvgFrYst0Z1gqRigeIodjGrwvrv57wTd3EEBAg8lnX5Dxt65QH+ju6g3Lm+N
/04R7p+TAdQatkaHrqhqJMkWod61wmNl82V4h1z9S5DK6Lvm6V1Et2r9JbHMeISP
AK4PO2IOPdpfwjDRDAN2NzOb8lZEhSUiz4A8QwSXQm8hIwY4x6NufQUcZY5nWRLn
86rZnKr9agpwquublzPjsNqzrUpOpK1MZFCroZz9zIlX8mV2LaXlgwCYAhCiSejN
GwVrXZ6m78tKiS1xhIr1RcM2c7W6SWkW8IX4WTiGPY0vLVcBhmk2fx5t0BIEGFgS
ghKEGRv4aa6M4r55810uHJZKRcasElAqQzJNd6GYbREdu96kRr32dJBixGNswn0k
+k6M+zwIy/oM2b//pEWj5M7U96U/kYK/b+A9SHBJv8FTt9uHItySkd9m6qL89jhq
nLzaJ4XI9nES04EM45U2jcOT9b/dA1GdRrOx0NhXDrjdK+k6X3USzPW3R0cPsrtO
LsLkX4nfQcM2mWwUrdMtDBKlFa0tejq2K6wcRmiEaCehJkXA6PCpQf1keyDyVcn0
xiujzJskCwGtoaNnhL7d++c0GgPwdcBUPi7xzrgT5sBxg0YGhR0yrP/uO1OCCV2U
wMVNSH33fFTs45JBefFBtvsNuVDfleRPx8u3YI6KWzMA+9VYWbjB/X9Ru7iguytx
HtlPXAHqhVPVjhUg0HSdWorMv59478JEvBceJhal4c30tEqRcXH42Heb9IBqwgA+
9zJD3N3QJ8Mxk5FW+3AiptFgrfLuldbKzxJLABbWV2G3MQysHD9JZDJFWbyDXo55
mSHnLM11jn157GRrjabncJT2uuNXhwy0y/xkTWJKIe4BTvdwVB0cgUvbMGJHCER1
f4K8Tdfc/cML2+gbZ2xFBFVP74ciUtWUB1kUXtpktsko9djx8TWJ/ccXRRCpfOEE
vjZ6g1jJHHTN6cnudK+hB3iKXYVJkc4rj3x/xsP8g/2qSKmqAW1GEalhOfBXhT1j
Ug5Bu04F+7K5+hmPJe62Hh2mzuOA0bu/SLhm2npQd4IGVVDZjNxg3S4AVlDEuFX5
NwHRLwlQJNj2LcAyPshlC8nZt2IZ1rMbaKQliN45HOW3/kG42a+4+1gdayGIxhO3
+FPiiaAZj8bx7RVgDZX6Ab9UrMWyoNDZInp2j8qCnL7r80D6u6A4dyfw7AWCLK9X
NVy8PaM7UB5e3sf1B18vfqJIKh/mgYpz6xzMpzxytXCd2LtqAMMZumOq2vcETUtp
KGopNUUITyX5hpuU8/dd13UXL35pxzKxmFMISAc3UipD5kVDVXIav491CIMRtJLL
u4HjiB/xdLE3YejPhoLBIZiNYe6QqXlZYsuMHfrTpTePlzy42GEdh0k9Nm8usVSX
IhArh4OyvubqnS6akNv0lVC5Cx33tAFVBYH9t7/B7OEQU0JmM4dk37v4Q+dNxVox
U4xTULeNTCcmFAGV9xL5tGvMMGktloiWmlTDcuG2HpFbk91ds3GYZXFVAUFqe9wu
Jcv+7V6UVTmdwgpv4lRUnAyt7x7jpzbnyAc0E2cGnBBc39aF/A/Vg9QwJ2R6snyb
dDQLXKmEMyA7RTCNlz2u/kRnq4y93Q/V1Xjq+mZ8L7llHvCYeGh+r1gDU/nTA5OY
RR//AE60J/zUgKWGnRgGR8FNOxKVrw+/ugn+/n+l52FGmZOsAzDci+3SbPfiEYhr
Vhyi0uWyQcupGU+38tJYP79q81J+hGtzlxR2v2WDML+acdNpIG7o3xsovNg8h6cx
sj57m5PiUF5fPmzlWVyDdkehiYZkYIK9SbFuGSuTbjRtTKUpvOozo6HPlE7JIhka
Jl7lioqlIo9OmRIcHAXpd9IEthBmpRMhj+USDp9UM46ko6ebv/sJxrIzNbXVzZTw
Sn0xH50pgy9xfoxifWITz0AvqypD1vluqXQGTBth/JbXdFs59haz14pSd9/KC2Gn
p7qdyAcWjw3JhZTgmZ7+cfmTVMoX0al4QrowfY1prPK0T7r9Ocll2wK5+N4xZSnd
0GWxV8MqgnkVV7sMdunB54AqjZfK2tAxwCdWlgrwCX3TTAXcP3Lz3gcAgnEIUTQw
tsQWO8lqaRBRGzRGBtmSlyLfirPLlOJgsTRPde0yCPzDYUI5HcBiroiJGUYxJTee
DLUyje2/L52Ye3nGMnel8drAGdDH4FIXVS5ogs7PhE7sYLFMFvwahRXrDtO+8QDb
gbST/NE3/V83bAhelAnRk55rE37zB6grxAyf5lmlSZ3GjxiaYSe2bahxqyNetv1W
cg/SxB/IymmmKB2pkekGQMiK6qww4Sf3GrlL232u2Tq/Fu/7uEkA+maxuy4vOvUz
5FmmVuDrWNVrsPbx3R8CK0DZnQ0CpAYlWlYWEYPpipfYjfFsVuq6KbKM8aVCIBK6
wwWTKfNq14/2/ag+7E+/KaF2GwQIgyTXDMOrHOu37Gcrc3KYj0K7l4af0QucS5oo
EGRRRh6gmTn3HZu4RumRBC4oK/YJN6vAliaJlnw5DUom6YBw82nGjjzWWfYYRw4M
uyCt+OhntfoKJgqDAe9mmR/HNjs+A6n8VsdFzUnZKG3ziqSY7IzoLQ1jHHOv1MW0
fIPyXXBYn3Vo2DNmBPOMkd5oIsNV1xl11n5Ach1FUWuYEJdT/ijYbKSbc/itFzoQ
pphDO8ITK+iYDSTv/A7OuCbz5kdDnPv/I2dcZiTuvTPSKPwsV4pc9PC+6ssaKC1C
sUEnl+ZA+bj3b5IpKleXS/3VGh9Fp3qte4MS7N0Kku6n9DHhauV3zpWmZaH2X4lV
98XRZ8apGLURdq0IIhsiiTauSWRXFx0hblbDF12IgAxhRApUNkoo6ZpMgQK81xgg
/Uksr7Mu70qpJrEH6AzQ75M7wufrBy6Iljot6ucpxQLKPaut60r4IZBluJYFmJu1
3+xFyXW7ra6dHeNJmQw727NP7DlejoPSLJ6W5OJ5DE7uQ/lVpEGgqhk1nUg4B2WP
wMyf1HiaJ/CxO259Y5RrZ5vcUs4lwjzNZJ/k3Q8JHWEAHcH5BCL6pL95e6FlQitQ
QHN9MFCXZAoVlioV3pisSrd0+KKOK3yGD3dlG+sheJBNOnSF7E5BtIMQSNoGhgxv
anWsFQ9cAOWaGBbCVThNHnvNKMoaijhVROxX3N7OeSJ9Ns+/tZpffemJSoK9Siom
bSPqHe17yLtw8Mfvg0IdtjXla4Ep/HVyIS/c5N262hqMNLTzlO89BYVuDKgSqw/U
MxTb+c3ZuEOS1wQ6NweRESAx1vT4T981v7Z2MYoxTIVJJEd7KIEXUymj6H4vouNX
AqR5usInMgQLypASh/xBnyW6BE3O8Uak0ScGnTp+0XSML0JJbQGR3M0gEWdwTLsg
N3aIGQn7M/EkM/5qh3mi2YNrD6nIiBM8iRn5F3q6phdtqOOKb9PTbL7+wK731FZc
8g0vCKWzs/jfILIQ38yvUauDmkF3KOtP6h+3iPuuzlTHwdp0NjACnF4kvUKk94Zk
KojueMqdymojpVzm/augAIagn1/rvsRHGvg3saOn5SCR1DL9MQn2pjgvePqQyU5U
Jr2OPwRhDQJUNcYbQtmPY4W3z5/EERi1tMi3sugFLpF5vpYfphi7JAJsYGhucDrr
IplD7ksC8g3ksSeUdmmRrrRKyYuX0n/X2KsyWwrkFPmxF9oMpsbxU3b5zHYhAlVc
81mTGHKiuocCNPDAUNVbv7dKliW+iTnN2koXQdkaHF+AukPZHWa3NV7yMMKwO066
tXMgk+ZalTWBWcm9Ol7o7MMXA+5odDnCmVP6tfZh+Sg+fGkdLb68BEJIb4Z2UnHG
DRYdq2F9oFRtFp+ANGBmHp44wsKmWAOTi2jjMAzdsObP+67mBaADeKeV0EVNs+j9
eLKlNtbY33f1r1w06iYBlB7blK7WjZqqyDkWIplnHoyfUWCSpN9pZWGg1khoS3c1
z/xe+wOoMW2Nn5/Hp4FOkLY52kIyL3IzuTJoIFTB2/APcpL6LBR0P7ZXLyf8ZHbQ
4t3/MJSLI59nYuEhTA+k8gvHQTxO9TUjb5aKZSDWQgypOOMf5THouyh8iga+5azy
/cZLEyT+QdRAB9gzefhWk6SMklHYYYA3lClenpEeABoLFpuGOTiV/2g/IGu4MKwM
5HCN/wcg11aw7liZIZO9glkBe1pdSd7OD7VssUwIZCTP1yyaps1Hqeqj1TBoslJy
uDpaSofv8yGUna2OBwH6Eu7wbA6WOE5S59daqX3M6J1MwwDpQ4S3mBk0KAhrIUws
IstMyjDFI6D1Ua3MiozI+y3I+p7hqy+jhdrSQYOzNJqreREwZJLlmeJwMKO9h4tl
LyPAy7GJQ/EctfgHswnxQ65SXHrmvPsAD/GiHMOKgPTAvkEfV8EEdcUrKIWYyTf/
y8+5c6zdYLeg+xxaGuB7LWeZ7hvD0Ec8TOtW/OpRCokkpnuGz6BKmxKkK3ULZF96
5+1RVkvryAac79JtqRUi9CFhfOEzYb7/dRRFuSUKGHvVxQM0NkNBWvF0tqkrZgLl
onZpKB7TzwyYLkaTSxwgkI2q6RXlFV+P8d7PE5EfxpxeYT3+hDrt8RPk/l9e12HI
D0ztgQ6+eM15AJhiiISNi4ev/4AUPHWI9riEKK9XJNcrH7JLZaMwIurHBjKa+MBX
69Inv3H+yaVvKPSIrxWsTJZaFwOQxvbvUlgevdHbZz8c1ATAqW5qDsvlz1oo4dv7
1Z23HHgclbOYnTq8Fgp5y6k2vBHsDwND4vhO4s+f5ald8FrnIEk70DOc0hvunX1/
GwpQgaU1meFvSIqJ5k2lzsxvu1TxEnZNoI4wUf7hprlpGoRwRmsE76klaV+x/uwH
6HA43T4Wg83elOvVmkIrfpTligMlO0Fl1PQYnDWopKKZg2rlTAMB/Xfi+B0WNxPi
03CknPvXxI8GJV2/HQuvP0kCFotyKYIIyQDI2EqI0H1gJZKVysvTLw2xb/Qgba2C
mJBYnI+62M59M3vuvaLo5Ecq8qj3VBTEmzi45Dg4SsH9shXfups4ly6AT90Xia54
mY39JVKLzpMkMBYkA9PnvQQUolxZpLcbjYwb8TXHuDNe9RgpZ7vrA2rwDUwMGrNI
8JylhRUqMFXSVEcaeXxxD29xQSMM/ivVorubhTcg+7mFZUQ+739o9K4HlT4ldpJH
XDl8RK7ykuwRh/fossjB3HjIbtCl0Oc0QVEikHvAj086yNzIosV1F4fn7xKXTlgJ
ZmMkfC67IvgFJJk3lmeLUZP0Kg0itZRsjcSYy6Hz2RQOzjpCoATV/bEAkwt8YgRi
7rAnQrIlccn1KWd5VhCkfWUFY0/fda1Wv/U8dLYFDnA10/48a/BItj0iu9lFT/Y2
LJGet0UAlfkL7kESCNPzjXZEGgRiJFFbbBYfoSJcc8QwVkL0NxZkIC3ggjs/Fveh
U+KshN4ZkWbLKoN1U1n+AQqyzhzNQU1qLjAD4pZjaF7hWd4EnZ5QzdNXhYMQ30AO
6TzazJ+qpMJvrCrc+vLD40SBcdDz5GquJLW3FGn/WVY09uZsvYerPIbtByk9LrAs
ksqcSqwcOBR7BdtTvPZkQWXos685hKA5MLvOfqeG97tbewMTEZwojIfO1/3U2ZIz
P7HB+jER+NYwgKf6YJU5sMv2A0L+3CCTI4wOWFW3XMiOKP4iu0xKqZpKZ+hzoglr
5f240CScILqpW6F8E+uHkHdEJ/yr+zNal1t4ArxoA6p0fjY6UzRspbZTdHNjPwTk
Gf4eth7tDyWLbebL68W9w/FONp5IYU2hyYPZEliB73wVPueJVylpFgMdUc9ALMzJ
h0wzt4fKSA4bjLXxRg/PsG6eyAgpTS+c3vMSwKj78P8S5UE/o7Ww6J2B+IdXkWGw
AMLbPN1ExM5xDTLFCV31MHMzKK8jydz7F9Uzhksy1ERuzxGSur9NzjAWw9BGwPd9
fWG+x/eS5vDSYny0TF2I3yBRn7qU+xv+g+Qm+MBDhZVR+pQe87LBdN0J15WM8gSD
oBZqrwvvYvhAfNaABwYKXzXageKt0I/ZZIzTUq6M44Kau9AbsURyXy0uE5+jXZOM
qweCddzRlcih+qOYeXrzK086GebAe1NG8XGfIyBKO+Ojq/SuPtWY+JeIui6niBnR
ALWMx67OW/1R4c/kjVchMPVp2ft3lIifP0VNj1YmEg/SWX3QxFV1G3xcWlaqJoDX
kJzuAOMoRxqyw7Ae4CTaiZ3c1aYxnPfsUfdQHt6RUiwegsl5jxBJGcUBFnzCwKj3
ERgWRCHCXW1JQ5G/dQTRV9hR/eWNA6yyfydeopRNBfzKU89h6PLA9ZFYgTvepeak
GppHGW+ll8/+UWoOKfLED9CGVUBUpNwZi+E3HsDj8QfoEJfqkGgXn6saYrsQoGW2
oXA3Y+KcQTtxvidrBk0kqKHUViIyDMsvDrXC5pFsL67CuW6/xcR7kBhQSI3mefJ5
Ja1yVa151XJ7uQL9TjOjsQ/mVdEu3BPo9Rc/5tT0raah7UIebwz/BanWr91quDt6
ftoZ05q9zbXE/anAvukqg4O9AzfW0w6c/zYkB4xLU9hNVesCHZfWMe5CB2NHU4pQ
HX6cvBAi0XajrrHVZ3t9F6rFOvEYtK+nO99eKrd5n6R6nlbsrPZjAggWoQvFAT/6
MKU7pndIp4LlNoFBIMv2c5HTOl73jpn3kgx1rhICKEYxhMRq5sBcOIfmOmYFCwfe
jG+b+8UtfBnCzyZD+r8zy4S6J8tF4S7mr+Zh63mxGkUTtP9VlH19UtvKNB+MeoK9
rtORhpB3tDDQxTqhPlJfu6qKyIt/lqE+6vmMlAcdW8aHCHzRzpKvI6VKghmll4mi
8tcqK/Gh9tAIVECxeaf3vf2sL8EtiPGuhkkwDULwyhItcJnpb9ej4bHC70J6MuZ1
UuTyWe+7OtL4ehyUl/6CMGYhztToKQYxGlPRhGcWn+8e7Mvbj4Egme48Adwm2I5d
yjN4K8uFbqUjv+9+PqY12aMN63QgYyyzjj7dF9vSXHDKYMpjCn5XVlWBZBPEcr/p
Y1Ipl6dwBuAjfe1NVyGFVRww4gYPy4yQcPABJ80fWMfC6XlRy0xWbSs3eaI2K/YV
0p6B5rvFmfb7gs36tRl89DYSzaqekQqgX2d++DHbcCky1ddNGjMv3790Ot9yuhsg
f9QDrmu3Yn+d7W7BeahuIrXYKOo0R3RB8vnJG7ot9axL77n70kmSJZtrtpLEPsE4
vwbhfdQmUC5tfoVVMFWO2H+1jYA/h6H1B65A5DXH0gbLYxc7WovU4bz170hfpeUL
8rM/bikGJD0v3sFca4d3I8k/Ilk5rrwFmdHBQ/vs0dtBlWt37AqopMt5W13slRna
GEF8vM5N+Vf+6Co2nXX81Y6fYpHELk2lWzx5psfV8lSAXYL+wrTiySyWCkJ9Fmlv
JpiLAwipuat6SvX0HNXXkZyBPODO8Y6CsG1ZjGD7YFUXOHJIT5VLj5OJwtw2Fx5N
LNouJs83hFoS8nU924BqKtBGuJAGf1xy+WphVO4I0/xQLaDjcdk9t3AJgEFghYOZ
skQ0mFiOTarLwjf6YUKo9qArzI1QRozCdDzTSgMGcv4NYvDLMkYqSIv1MO+EHN2B
FVzMtsU/1xcgCs7VlEORM75e4MIlkIMzZfpK4Zu0sUy10ZhMJDa+j+zkGe+4844M
vGdEXySQe00988Ci2xIwbQQ1TySMnwM+v9VEk6ltazIaRbPz2xm/Qr82i+BnNW31
15x++q9IXbeZSIjDBkgVAF6rBwcGuPnW+L0Q2D0opqIKFhkSoZTjU8m9yhmye0Ji
uy9cYcs0XE/qzFMGFSGsoNPhA7suxJe0lrrzV4EEbF7eKwYWg5HWEDNF6pwkrioc
zSCwLIZOrbPjwfaCA5QY+ordzO0aUWHlsdaK4Wx3M3JQOZ0IbpE+2zSiI7G3Yjx2
dFFLscluHehXvJXG05qmooxhbt89l/GGHatyoP5+qe5Az1sQRuHnbaO1Qkspuwiv
jpCvzw/hGeO9zHZUNH6J22zjEw6Qq8ITUJQg6QGZiYIef2odaq6X53IoCXApyacw
ESnL6XgKoSAs5Y8vRvKy0SYs/J2c1vSTgurakiv1iVP8eun0QmeiwGO0JDiWp8ZI
SpuSNDYeKTl6pfyi6LH3lFOWcO+7aAnpEvszhW0hn7jWN/9tEOAm2XJdcSixrlBy
1x9o3T3YMJZer/gh4oxTJ9ufLmkNYSASL2zwOJ7COLRYIBSjYNclzt3VFoB4w9eh
yWE63rivftMd+2kSoQTF7dz4FbkXPEAZqQEOJPJM6SbP6ITbp3k9mz/qHVFYpcf/
Y09tbMN0bVN+gfxlK/9ntzSZug8V3I9FpJgaSWzWbgAudFRLFj9T/21usicf5Kkk
Ks+4cRWPsAGJWNv4boQu+YtQiKnqbIWz+wfPHN43f27jucE31rthDmKF53w3pVdl
uc/WSTUcxipaKabM2yzut5iS1EPnqyqkJPmdEJqPpFxfylgygBeWKSAu9JQXh6/8
zS9q0WAh/qkEptGm2cfBJwL3oO75Fw0Qvyb1xIQ6QiAzeLnlWK1xyNvTPCiRy+Fv
Q5LcUktkCre/ZuHV6mtYEK+5NNbkEaOrNNuzTcV6HobUkTquOw6TombdswbvFCiw
W1rKdFgZAuBraCQxlkzww5g5kGjC4u65dlVd9PhrBwHn/WSLvfTouOwTTaHQPGyq
okhaopEJS87MF1KJzGW9ffaBKAIm0Rat9pSfvHlVbChR6H1jWQbIi258xnimcxMP
TI7bN1NqiMR47a/LeWC2boanOx55uVZeMuA4X2k9HRbYZaO54pT0hItFXPhLZsSs
B99lZK7P4iBFbn2V1+vGigfZWd2BVN+vnOkdc2A9DEhraNnLYXsgLcDBy+p8Ak9A
dTIxlL9v0TgZacsGnFsILotqY7zCAlXsxq3p8zgxAbMChwfKwD99MFWmE3J9iRae
AOIXVCigvTATyOXo97p/gfIcchhkQzm/41Gjm20n7E6ywVpzqodjHQkXbnH6BRj8
K2QFs3UyGbyRuMHI37VVt8DMhdHEdN3weHcpfIfprN/X+bcikMN89ExKBdK6BYoy
EvIoxyZaGF44t+EKDYWWjwpM/l0qR6x7SMwIeii3JlxHdIPl8DvTpDQSGxZvf9Sm
aomszT39KR8ngzMNv0O2lf5cGNi8wMzaPoFfsTWc7axb6hgEyy/ZHigKEkkNb1ub
XxiOWS8sNCrafry8mC4bPuzMzovziEjQMudJErr8B1wDXzMQNGLv8JsxEEx62PVp
GnQ7EauWTWJap9/YPJSW1071wZw8U8eJqN3Zzc8Htx9sxpMOfhT9whcCacdV6Ai0
aO5aNuBy4W4f0hPNMI8/IZyJzeKcMrUOPO/AlzRqdEIySShtYe4tXdh5jy9jVCsM
+X1PYTMyXzyhz9O73aX3z1uG9PzumXKd0XAB38f0IX1cYpOr+tL068x7vM1oV72j
gjC57IyfdO9k4/AbVdAzb6Asu9+lHCA/UC454CI93DP3k/TENcMnlC52VzmMovBG
FpnVuhGtzG6hbjVIuVrdN4YXY59h/Zuw6lOLKxy4K0BBne3iWiuVJECnBbqYW7az
h+SJrrZZtB7tHIyk2NrOMtIveGIcCA0/GchgWmcK//BPv7XFXAsWEnc8QYZpjgrn
EyViZg5sofFyb29qnbCOWZ8Lk5znPWttOuM7K9vAkFg+6PucCAa+5l3wCD4D/Uz+
ilCle91OMB4kAr5m0WrU1DhmYoutshohuOESZiHFD/GN/Y+8AoqAOGw8uz7FKVkm
rZP2vvQGyXcSOXUdtBdrmX06XjNmPgtABdB0MRkC419mu8/5xwE6XPOG9hHcLTg7
r25y/0XVkdh3ZCDFZCjG2D50nqsTrpfTRy4YRKP9eLPa3ewumhWwX8oVZJtRS2M3
AyWquG4uBJU8apArtNK4Ax5vSI0t1F9BNBFrTRkjKdVNrtrxrx1Dtvi0R02SLdbS
7r4UW8KxGg7T0HPZfV+hOIu8KtiPf4gwbde4sjINb3mLswUDyjpwD/Bp5Imifl1G
b3VNrtFgSl2uESm5C2JX0TVMQA0ZiT55AnihQGcpsVJ2ywFx553CZDSogy7DzPyH
e5K40mk9/E7C8R+8GSisSWp0OsKc0YiUE6kxIiqYkm7myNhLUoDR0YelB5Hwq91H
PTWz0cXYR3xhw1lbjpxv/UAoS+fYnL1BpFmTKkLk04/CDlTupajXFs6Nj/qTLbOB
0iflcaOT2BP0SDB/sCwyZt08Y32KGaor8WyacW1xf5eujj/knWV2iY5jaVmywWcL
SAYxVFwuFRCZzzvkhRNkT36vGxnLB0PHTbZTIODEUqs4dIQoLZGDC2V/LRnj0UDi
0MFFGywVfzDP4kqmHBkp6ga7y3pwB2d+hIoAirV7VQrpGGUFLIXSvgh9sDjJ7yKn
rpA9BmA7Yvnvrt0YEMASkdWAhKAvCYOTsBsG/YdpbfTGmwuNkLzRqPKOXIOeoVCv
Fb5OC1NNL4kNIREFUb9AXZ5VBSYsyG6MWJmCOJ9UG5TB9G9tICFYwI3yeuH+i+JE
o/RyzyKYSK1Ek8LYEtj0yUCXHv/2JOb32CtwOCafsE64bya1wxxyiKTNLQBapyEe
DoG0yWnWwDxcHR6/zpZCWGPZC1dJEwc4KVQYhF6+Lt99moU1SU8MPJutUNPgVIO0
Womp3/U8gdZQXjHGwrHM287xxz992C7yU1ljEMXQzRDXNOInD4fDheV30wpMDR5k
E4fokHSdj14OhgePmgwP51Icu4O6rEcqpmauEAWYyM+Y/HjjfzHl2+mdEmW3+W3/
83olMYzO2XyALzdBuZOjjR8CaShElSuiV+ziHc76QeUwo3c0mETiRTL7+ahMOaei
xpLkws93QkqY9rHeKFsYxR8KMN8GNmOYV8Q8BJqgQsi2nALD0aB89VXTSTIbBdIT
qU76O+7k0z4JO9MhH9WEEWTIiPFu7Kz3NDk7RGBByZUTWMBgcd2z+rJYEjpnAaiD
JXFJFfiDFGmXeqwkPtYOfF3QLG6kKTuIe/eYY5+WQzLH86pg2jKbMG3WPFSLmtem
Hbool37yXmlAPXteadvtyFFF+p2DMhgHB+SLr/KRGbr2GpGRjGru/f+hzV2AwRld
fCPGKV1rcs4IJ/K6v/ml6PBiWkOtBIeARbZ5tZUcbHiUbSvicj5X+cjzsbp942x6
QUyMvtzSBYlw9QLqrWq9b7aS2md7UW+PmvvRoZ5Xj1hw5mNdQcv5NIHRwKgPI0oW
EbgZWaaoUcxEoRDEfvM5FWO43PKrToxsRQSdJeOJTBYjEnKn4yo3N6blU7xEPM3a
Hc67nAhlvgV+ZksG9s863YATGaR3Ti81HA9TEpx9+SZiL6QbePp9Yh2r9bVsPoNE
tif6iQ85lkz+DNB+inrllEStBnOhJqRk8NlVWMMZGP0FiwTgMA5J+NcnrlYpzC5n
hhnzPL/krB3JD/rQ2emT4ukKcz1hvrgQgCtrmMy170+PIlPTzuaM4UnZ/T9KWUII
RtiR0euevbl9BWk+GZoJKpeogMM/TwBMHWSQY0Q4cBy8YnSrZatf4Cefz4TGqbtB
ECzJRWHI/+0c52cGx9wepazDFQwunjlzoxlyQLrredi/smJUjXgM2aVloR+2VR84
CxYxkCBPLfNbEezMgg3zlW/yxvwlEyAXMGG6I7wN+AkHv1jQxK7MBmOjsFOLC47c
0pxtUqMA1Tynttjmk10ukABinFC1UniEERW1GHVQ4/Y6f/txH/ZNu6GiCt5UcTN8
tD32wf9x/gRWe9XDa2HVvsOGLVBW7eonmcZXA4Oco1vUgpMhtbZxNNV7fD0lx7kk
vixrrAQBQz34MeKcfv3oID5B4wA7YLNzW7LrNHTJNNE4L5rm0BmbfnaV8kV6xSPa
TUXoCpoVGjwzw6Tp+R/piuC5JhGYAPXj33aX/UuPZR5RZd7AuuXJRxKbdy7qncmY
/MTCWNXkvWY2A+g7SJIz5s0ZFkTyUuVutBotXFR5pyHmPcDf7FvIM/6HnIZqfxm4
xCCpsoo6wovAiSp+hsyQtajG9YbE7fWsWxWesEzszEP2sCmDxdo9DFWpmlxBFZK0
MVWrc3Qy28BRe5KIad2CxJ46j/dg3hzG0rygmwcwuDRdKhvNRvGssxWHg8rHIiD+
2QIewEX8gKSm++djE8ufB3jH+bN8e15iWt/J4LURdjQJ7PKBld9bH5AWf4vlsejo
MvVa/q1ORzFr//lSIHlilGShpiNpH6aDdkgDulK2f7oSwiHJPgRBfJ//c5J8x/CQ
CvCy3gRrF832AdpRlKeRhwvdlT7brnclnKSBE5cbPu9YeAEbdPBnDDijI+dCZSGW
/ztC/X4WODCG7C5rcBJSyu6Eh1JSweEkTzt/07fDz6ET2sCs3k+RS3Ta/awM+QMS
rpjdSeRtLkzYVLrsZZTZuGgC8vR6PI7eqg05vVyJpNlc80jnH/wrW7tRRLWJ5WAs
56bvO83KapoKNEtUbt31xeedVsjBfYkdW/X7haiJVT4aAvzQOiD6mfcqhBWZVeWR
3/Nhg3hjh3oE/9xSReyOzMe4Q6hX+oxStEtgDEblgPGWMrp5c/xpCfLSF+RlPRWR
TUw9K/tKorNKnlVvrWMAZ42sUVKyESsrJ/0Fth50PTSIvQaHTmWEeBwZwez7gcsr
Zeke/3IuEWCm0XaJNQ8iaOheKrO95COXjG81HWrtmKEoBXRYhj4l78brx1VKFgrv
65QsHUXJQe4mJa5bKWAbowk97JHySd9yyRnEjEwBQzfcOh8S6XFvDJV3V20CH2pC
sBblsiNHtAuS19usRRiBMx+zEqwdtJbQ+fby56C3ijyHdb/ypDZ3SyR1IqXaEzLq
Y75wIHBsT8FoIhfjFnzO8CbeXakhBY6Xl1vwwbbZqQLOGGxBZ5FKWgB01Cm1DIVI
WkKlo2oAw/bZgWIAbqUjekEsya4ltrMnSkJ2z6MC7DziBBKcp+0qRg2Yoxcq7R7V
clOSyM0igTw+xGuMUWPknETsBbpTniXBVl2J70UEXx5hbSjmT3Ujn71YxHUkxqRP
bBRb/LTbUdgqQDfqoFfboyrA6EF0GB6oWufuGuEPBh0OrSefPennvArAmN2pggAR
Z1KMSKiP/+9G/EK8m4ISa0qtiFcHsmz+wKxuSfJXtB/9szKb0LrB6Pf4wiSmxRdm
m31ACx49pKWGl5uzVSN4h8+FFoOU0ZqUPQiV6X9tTarLY6rx+1NM3sa1Ng6oEoW+
gtLdcaLVTuemroqTjHSqj3o8Zq+H9+G3n/MDT4r4+UO2IV7uwytT54pbZ2AoKm4a
mENz67y3da0kJb/+Rd7g8hkIf3z7PoR/7taTQZhfUIXrqhPcBKkUCANZitpRE7+C
ij3qq796FlE8Y6YAqZqVy4ne5Ud0eNttoyK27VgXM4W17qV7PNEeIdmRgjfcqyRp
r3VSJgwxfKS7Y8nSK0NhFXAaKx1VHkcyFXgJoXtU/Qsxcvn7Fca5aXLY60JMpRIy
jE9Rcre4mvKx4lZkhdYoq+ZZb+OlPhqgoiJBSzYUmX3L/tvaxNgVg1ENazkiJiwM
heNBxTcLCjE2BTBj9QXxnb57Y8PVxweSHIzvP85vZX5DYjXrpAuKS0U7YdsKSWC7
I9L9J7OA3QF7qg4hjCpXPOUwmDlAwZPFG54bMca3ZmFFrFvsbyXXUFqai/KnJtSp
`protect end_protected
