-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
nOnxDVbPzOWqdJ6WvPooFTCUctIjNrQ2cTpor3x51kLrAU6XdaxwP3IArKCvx0TN
yzCJL0P0HbyX7S4GTG64LQSt4kYU+H27uwNisF4CXihfcILi/K165xDuC+ASorJF
SUUM7hRYWPc070t2HqQZJ4shaU9IpLMiYGF0AifTJgA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13024)
`protect data_block
LsCK6cWQ/IcWORQpMbEUt5UNhb/EEdVrz7PcprZks+YvBNmjtMQFu7hzdy2ezyqp
0r7FCL6q60uRYCpBYA2g5ZhgGOsQ4gh+eKU8Ud402kNUl/ZXg5mzdvSMpV/pLdBj
46EIfkHPd2YUWeHNAZRfa1E+q8E3XDip6UdZBDPYG53BtGbaYt62Y6dMO3SiUIBB
TIza0ek9vkpsSb7N9uuCwENNDqT5Sfb3AA+BIQ8pa5RVFN659DXV4k07CzrGX19W
mCMz9XaMmeWvJcPrH/z2SqiGQZHbHTSusS2zMtQSnEiBCjPhgj3+euBhyKB5ILfO
NBo7auU0qO+8qaJ4KlPecPWLCbw28YP84YKl0thY3czVn1Q6Dcixvwqm6ETfe1ow
bfiQy9nVCEmHCXw6gFt29A7fS4k6zYDgdfHyGVgmaWPuEBntgep1vbkfuTf3gGWC
BsSSMckzm+24cAgAcWynw3uMza1lxJgoW/l2sVT5TOZ84RdxbCeUhGHfkxHLy18G
3Zi2Ih1z/Cy96It9ZeIQAzzoF6W6SNcRDAlwg4REHKgoDnUCnA/gW2D8muPoS9a0
Hn6OJOQd8gamZFMFXsNDImcC5dTh90BT1OAtgov2qtGkjy7qspPKdaVJ5WHjpcIb
n5sQlg8MhYCwMLJMxp1a7/GpT1uubvfXtCYIjl10FztZDSaxXwFLtoTwyP16/h6b
LvruBioLHQto/v6GOYXGqq61+sc1qDGcRCVV+bdE/KxLy1T+lBI14d2cFOq/a2nz
iyoIzH1apfwY39Fw3XkF2pAPGNNQu9R4pfFfCe33HlIy6oahqUkWI9PpHFN4W9m0
Fq4a+VadsfvKeq8eTP4wnbf2/ejXqbRZg5+paOSMrjp6APot1NWPU7vL8NYYasgG
Tu6p3Rs6swDPPZc2OXNmg/5phNR15FiWm+kLUnDOAb9Th1YrboE7hnCZK1aKzrpl
R52JCkb2By+vFUrgP69RdWiqZU55fNum4Sf1Xcof8zAiDaZxUdrBPhygVM8ErceY
IGo2ibVqaewKsMghqk54ZYzdvFWjBfSBWsDp1Ef52xCJ9H/HpdQv33Mns71OT7zj
Vkbax3e3jbV39Qrxq5OCL3Hws33YegeyxBNxaJ3zx3skhZHGldAnQYVy7dkElZUC
FzoS08X5iOB97tnCb6ZyfFSzy736ot+/qmtr+vgOHBbWcbW9ES+QjNq4X6j91TCH
HQnGGx+GWvWDqAii88TjO/Uvf5a8+Kc6tWxC+j39LUqybXG1MoUnVlVfWc+jEpHI
5iRrAu4lbtGNwJDJpzaiCvUxNoIff3wnCZ8m3EXOGA9CbCzOdq3d4loTL5iALx3j
G0xwCJD869wRLvg2ZwA6cvUPQjbyoWELXGraUuvAGM9E50ejqm3qlc9UKfZzMGoG
qZKRMbL3pkIo14ve7V+DmFt5eBsRo5zxt4SiHe3xAE/QgrUe8OfRkel3h16c0KxA
ypf4WyjTBwHvkGd1n8KM8/nQtvIYW9hx56dmm7BaB6GYiQ4M9vWQR9Fs7K6xpuMF
EQ8fWKb43brR+0x41+XOGD/6c26IAasWPozKX+b6+dOohbLUiXLwtz6EBNBgAQ3D
asE/iE62PO9QCuCeJL1IkX7WLWf1bxqSNXETHKcKPs0PTzuZzIZdXCqEeDtrS1C+
46g3NtyUOjBnGFT3YNDVvZ3PwElSlH0QqfYBqSXPFOk8C7x4A0s3xnwTvpvNspDL
2L/RjlV9DqTT/SgWyXA9j/nPfQ3V2yDel0V0pS1iQNWCjlCj3sdZ4+Hm1f+ZnfWz
il9EQFzf3JEXLKzAEdiqjZfU6qhcgtgB8pcZh6PVJFZnt62sSY81FG2e4o/14rT3
2PPef2jznWlgIGcqyCr1qKjn/O3yRKXbfVe4oRC3RSEZ6LtiRH3OBB3YefRFbzBN
CWSXyBdcz2GBgawsXpA7KQfb38pxWoXoybffCy5biRTrHQ1sIAOC1B3jCQzdnGSV
zhCxvsj58vhlks/HVschjo5LHYJ8Vrp7YsHgoGW8dm0zDKTT+BfAzRw/TdiEdIZl
kpffy0Smf5Jo6I52cad7Rje9i5MTr7YOg4/GKDnhqbave8WpEAz9xds1qd2dGwr9
WPeuxsiC2t3fTzgfy+3lCM4hl1N4BnuHXHhE0/HTJ7pbgLZDOKZruaQ8A5YXEDpW
7Q6BborD0b5DqvTZAjve9SfqtkCD1FY42PewugGBkUdrDhWbXuw2h3MmOvOPa5dx
dBC8I5e7VJSnNddJy6Q5Y9yOFlkE246+BknGYFOnFUE0bSyqO2bNYgr1Tn3ectcs
z84ynYYn2RatzA9I0jppFUcAyuIqEmHPA/XqzOnKXJow3Cv8QW6Av5dPKsg6+Jhx
5gD8bbI8Slu5/T0uDXX5zmaSpSRnrnsynBOUe0SZI/8bqpk3TUexuBi3zdwYA+BF
9T6MxE7deTv8e3Z7277YF3sMdRWnFWAYoQY8RC16fQmgJoU8o4dp4OSs3ZQP5WfD
Kx9txL343aOqLBgn83/3Yf/Nb7bxLQerO+xVXhQAq3Jdfx9vB87KasjNShDuUjnn
52N9bCn8oY4+mrtti0M5MAqbtrfJuhuF+FdGmG16xLL41sAxb7pXfPi45pYGJt8Y
tmK0qUCroa/obzSLhIHosOlceiLfF7Dlpn0W0IHZX+YaaPuNHnv5UpVa4QtUY7gM
SCnl4HES+wyyNDk41SfNrgg6iYTV1K74q+wG+d19hmRjj2YPHAyO1uysYGA+oPPL
77lR0tm8qUtjjdTV/GqKWL3gSfxlvpikqjY4CJi9FpHOSr+MZVtZW61wCPvsxsLA
arTT/0QnSAlXENnFSh00cEHy/gj4+IseGYkTjQIwAmzjTIuiWAWshola3uHkHXzb
2gYiqzn1IOjopgd/dpmTSPI3rybhAFWSmphg5dALjZBZbpCqhIcs/9OgIpBW+yIm
E2CX5dSbvNeLrCLiVRte5YIGMQlVJMlMwnWGiOLTYXFSloFji62lwyOsD+y7hQ9Q
KBE0WMvVInzaA9ALC1cJ/rVfEnaWjHG+qYmQOozC3yXMsujj6nrR8gv+LwTGQxag
y3WzXhen5XtbRHuuQZegmo33KpYqvD28RHUdNfJzSptf1sbdAEsRO7PhZATEOHW9
ZHz3M99I5LifMrEJIbADE+iPhGdrmZNKBY+MgCwul0dUYlKa1Z6Mey3+H96YViyy
qaoxIHfTGlnxYCKwF8n/Roeu6cbJPo6Nx0XxJbMqTWvUY81uMVUjgdc/7O9dJB+H
jMLCGMgDTRa8zGgDu/g9/B6xGmBxt3gyaHBJw3Hd8wMo58w3jWLDf+JmDD7lo7E2
WkkSYZpYPuZkhRxt4nGdFt7mS0G7wdpIsC1k1lGO3+uivpd15bNtYEm8dKm+m25V
GK6e+nNC1lSK6BdNMiBsQltsut6oRXY3Nb2PdoerUTaw7FoYMEgiY4x4R0OsSL+5
rtz2aWoQ3h9KnAVtLf1Md21OiiO3t+ZkKoI2spaE0J2quK+wK4LDk3v6dPywptcm
gSVnv2lAngLrztMf0tA71JEOa9lrd37t8HQJ7hyAQ5hjossX6TKcE4uJsS8D2S4P
10WjXfqmsIaEduZBJokYMc52AHi4M1oGs51H+TnxcXvo1xp+4JYYNGVHAb4KtX5d
ZZ4JBUv2oZ/zdYzLc4BhroCcH+kpXArrBSjJ5Y2j2kodojQuzsgLjqu7bK4+nHCk
2IO9jqGU2QZk6Zj68PAwNKMvIfcbIJg1nKUMbOh5TKChxEBPF2uElAyjzpW6YrHp
Jpla8dQe6wXOJAjC3BVug+grXqfd0vSbgFEmxadqgycxB9NvrFYDORKQadXoR4Qk
xsh86fxfLR8lPU9xp8X/It2xNi4O67ZwfTkLKggAZk4vOK5Ygna+j0OF3UJ45t6d
JfaAHJVl8LCLQLrCWPZzoU5axXH5mwNMEJ2dFFZYUBkwLrx4FkuHUTwhmOGPkAKk
Ev5VbrL3HdfYTrBxhtgeN8ye7JlOv0eoFREK32r9R8FMG4nySvZqwIg0Ljs9J4Pu
KQ5DOXBaxfVZp6xfYezF9DS/OoGA/mY+GEtHmsU4fMJAvz+aLqcTKA31OgqccHIg
HAN7xBR8Wg3rrVzTZAJ1jPZCGCiGLkYVB0F12mMWSMt5kH8htU+zIoRewXK4Fq4b
ZHdDsQe5wew3B3zj4Joqw5yYyifSGdYiYseTbjdI7rSoWOmyZTRY60vjufnNiRNm
Xun1WB5YZp79uzW96NNLSwWqTErNvxh1s7jVGdvzwCNIuyDNSvVOFAtNj1p68ZrH
pOKp3QB0yXUhA4JMbb1r26C6dji/jB4EbohSAQTFh6hgGNi3X/8od5CPjlh1kOGN
vioDb3LV4uqrLHAo7u25Jw3OJZkdvP1e4LpXJn5lTIwP0KtyKDA42VQwfQJ1zphH
d1nsbOx9yX4/TdXR9L5QnjEGYwDqx7uoD2vZOml4Ai1HpLJcrsxH2sEPkuGwZWfY
cCHYfCUSCbMAvZr59VpKRgPyrb5ZXmBNii1FEBU+4PosseR8eIKJJAwOlEDcdIYe
mq/RJzn5YBaZ77AI3+INGT8KyU0RxGzvtgVlwK7YjW2BzA2gGRpFP1LzQYx2N2+A
v61QCO8afKUqyhaRih0LPvz/wKmvxp8ZdSexv49xZZTMhLrbr1BNWO0EhMdjTt4U
UZ5kg4D1XWyP7HyyJTHYLA7XLBqxMAmNtcn8Qn2qdVlwU9CqrQaVXQ7l1E8QvEcR
yUx7k6fNNjP+wZd4XDetu266ocvtIqlSyAdK/KhcyYTkzu9hq0HypSJh83ZIMmM2
6IkZhZXr1MOonzOIG4XUdaiKa5mfWfg441KtW5EuLp5NwTWYcaexvYy6RMVD1nJh
bS2hwRELE96AqLXzYdqzUGCK8ujQbHmTCyqmlYSd9fpGODNphpUmIpV8i15xL/L6
BSrj5wQvvVeGOjm6xwavAbhBoCwdsZR67FDc3N4JT0rbPPBaIP7PDhttkcFxlXPi
pnmt+mxaf96mzbUktJ995Hfc35sJi105PirBXZ1rhYY/tmPkCw2xqHSJPG+AYCZb
x/C3AU+SzOyMM1mJnVoXIs+p/NsNi1F6Bh4lGGtvz9Wy3ZT3bKhrjmaX/pYypsOn
QNDa0IzPkZ0ZOCU+tL8W06TuBZtTmSCL6YbManotSel3c95bmWyyickZByLmvaqd
n5+Kn1WHh6EdHUKwf3CjpcKrFilszLjXpY9gNVeUUb/P70miKHMh8zbTRcmqngFs
YxCE1nodriLMHN5uizoI6O7D38Wql+9LkELmulXWfwhEDdt9wW5bPOhpKOiraZjF
YOSnHniFPpXUC86RZshNhFno2N+t2C1+D3k553LcgX8N6gQxX90Z3pFsh7+p/8mk
ftKWgYpTymUFz0DLZmMyv9AU77beHNxS4BXtCGLB4FpcPHzDwKm97tihX3GQ0BIl
nUtRwnAVwEFdQ0PhiXq86SrUVPJ5ggcmRcEynZ77Ltoo4u/pBXVWA/mcoJXc6auK
1fKSxtGsUoBC78I6KuhbDE3CPOCYcWZgtsecqEYbkg+3OOr6BtV8i0MaSFptU+de
B+4K3C0Y0DSKJgzejdZelvB/6/X8ruzLaXZTJnW3xII8/Nk5FUj+cZirajhHs4Nr
YawiaqdLFmh2ofzVfBjYHlX/SYC9yJL8vlRLAd0EtdnCypbvSJX/J6pDjQVB5dTh
T1QkvGTYVdJr+a9CT4aEsbA+tvNn4c+JBnsslKejHXgnP6wtdfFpHiBEymKX6n8G
ruHV9CGoApwZvxnMmTsyVTXr0IMCg/sUXJcSZNzzP9au6WGw9lOOMh7TfiUEr5YW
pjHr6CN8IIaG7XKqJN/kz6mjxa2iMuro0qG2C/JdHcHkDzNICZWJ4OCVKLHEkg8q
DtkyQx85iNIDSrlMnN4DzYkYe1xQBjLNAl5Op9ryvPvPxuJFIjK0TH1uADYqHtd1
8GEI3474QDklX8zF85YBbdNKdfVBpWW6EfBmXtEhUyVNNiTGS5ht2Zae+l+9/iuQ
M0CV7hjxUl8WISSWYDYJVl+2IY/StS1caqyMNC0oxCqbnSLGdQ2pffclyqzLQjI4
h/TSDJPeyZ/rYB9aXeZEv1bvX2vfMuEsLdPZrxXoKmVv0QjGv2YFQuUhq2ZcdqQK
xcWalUI3zuQWnRsk1nlDeKn5V437N5gBi+rwFo8cGoHOBcFbpLrbO4W/sQp+wcz5
9lb7ofNmveMfFf3TmEYFxkWRZyvsctimM31YiQi58k/aD9E20CqxGwY+RVFocWMt
1kZO13pPk2eiBAnxRvHsCGXoEnknFyYL+8TGZAlKF4ATk02vJFL7hl1C3Tb8tx0B
JNuuuFcFH101enuhf0TQpmtWY5SiL7ahyjNPqDKbv/E4frottNgnt+XDky52dTGF
JBTkBTy72VkGVuALXsipfXrNh4O7KO57ASt1VH+3DL+oy55fNGMThiz1EsX+X64K
2EFVA1bUN9kEalmPJVWM/u/TkXkgtSv4ewOuHL+DN2PIxHPLN+wpQt2irJfas5lb
dDRT4mGQmsef8iVSGqG85UTWbaHrw+WYUipaR+6jlro4RuhvrKhgM28CDar2bnJz
R0mkkuYvzWUBHWx1HRtVR4free4PPNRdZQXrWa3JhXWRF53t6XCZkvU5kSB+pA+5
xKSLsABv8csPtyZ1B4kVkfsA8iFELcpoZgIbMUUd7NpPT+0uwZkGhC6pb8IoSYeY
S6KS0Byg+QeEd9+nBSOGd+831UPnHo9cwDZABifpq+D6ri+7tB1ab78MNNMvKMhA
KUCPwGfVo9c/PmGE4wq1nF3YPHgOC9CuYrvtqqmdkbCJo29+qFolHnknr1d+R+yQ
er8kyhuu0YeDPdN/DR6cjSFrHNcjO3r3O8hYWuYjZXmnNr0sOszjT6f8TnA1xtXa
gZ6t4ALpHsDBFh5YEw9Vr1G81xC+nkvpuF5cY4KjOt/+BxsYpWeNJqVbZtmEphDY
719htFYi4VXEUwTYXwym25z+Ehn5kqsj9rP0dq7Un5aNaLli+bpJ0Zww7OBE6LSj
0VhrgEto8xsehijbTnK3MTVjI5u5APG2mH9YadDI37QFYw8mfVZgWhLpiNVg++y7
Tfu7NhLd2TlU2RCZYHfFNcu0vQsxBKETb41mYLzVOi1hafEl/zaIYsk170PT90pr
+XLPyVpjdbkFzabn6K3xNQ0hh+w2ak0pNCphH5GTAUF5yupyz8z6ssTVOMLT9ech
uX+nZCcGQSkVOBGnITznbNf7swcAsgQy9CZtFiT5lbrT6arDgaRKgaEJo0L+/ck5
JI3LgHys9rJdbqXG8zRFfChbei1HhDtlALAkltwpyqops/zpUrhPdrZZJYJQZDLg
M4vrBO973uI9ymrLrafH3GsqiNtzNqGQyixsOznwYUVheZjUf1IP4+FxUtN39X0m
BaT+EBSkv3BL0xOeh97VwcU0lMe9rcTTL7mBvbJO3Y9Ynr2inzJ/I+U6I2JTc/9w
VLjeGeotEbN6ot0Ua9KAfApVFWcJDPS8BXKtK9bNTVifUqHJpXdrMWya52vIpES+
kbuC3iWwyhNkPPPYhVuU9r51uqwXzAWH1E1qaCU5nNAvn4ecMS1DGvvNiJVchTXW
+S63nc50lGgWHbb5tu9tPtv4t5pz3NNabsYGZ9ncphIPwgu6NqhXznxYE8b1xMMu
1wekgTIe4JS3mwgKCWHdRfGXElZDtAHfumLgkQAaMt/rWcb5YBwr+AHC07vNuGZC
u5/QaF7IKD2iaWktQU3pk6QqQm/THVUWmhCyuTs6APljh8onplA77sSvzTbpAqa6
2fAHEcBbVLbbc9zRMAKYQc2DJhium2vOuCsHN3N6vIvG54YBPLVD495789lgRACj
FqmpCOGikbx3+KGqsN7yC7VayzS+L92pw6gTU4Gq22cqIAwJiMeO9OrTao9X5PzJ
CeEKSFrYNlgKk9+lSRedrH5mufmQRwaOAU2zI/Eo74fyWxlKIt+R1ZFsjVIP8Edr
oXiFE5uhCFTLzOLCmsCShpJaiB5yfNYpPnF1apLjLGZR7EvEKPkHCOV0TcSMM8w4
OLwDvd1SpgGQgXh2OXl6R01OhXsZpwfPpSczVhL73aouzriYbC2VHRe9RLwvIymE
g75moKTwjlFn35+QPaWJMNwmDXpjYvV46k/V1297OgelOhiGQEwuABmjB1s003Nm
141ott2AEM7E3IdMnFg4ljnvB+3WCLOdL7Da8d5P2Ucf7EGBuo/fS7SJExS+Qdwh
KT6yPGuhWKvWjyUE6/brOW3CLmHFiB3h9NehWGw4sYgblVScK+JYGiWyGX88KRsf
mGRX1HnE6ul2mK4v23jNLuSTahzui+TosEG5JyT2QjwtNyYa+xRNTEK7xeJp3o7S
R//kS7sbmVN7dwWvorH7OqqVP4gOTJ08PUbE1GrcAI/vsdHOhl1ata1qa4t7sZar
icevSNuduTuhwwI/Hd3njCfYv27Q6rhNZG8fyetMTU9PTrvdkruNPwkwuhnT0T4Y
14bkw6+7GF25/eDWCNHNuR/RYmbuos+G3lc9UBbZGkZm/ANwfbLN9TO+j1tGSF4L
wpVMDxr3VsONsVb2MRKaZHGGtbM0TFTnUIjSL9FOcXqcmfZrlkOyBQFwiCdVSbDj
0W7Md9wJwMtQvzjTJxPaAsgs0FjHiynHxWV43Tj7Yi2Q3lOdRAmwM29QcQ/wa3U2
KpMcUmv+aVwIG3t3DIOLv9gh/236zJruHkxeiT5/qpk5weISNQrI9GGxNd5zIG4V
Ze/nWN3oIOgfZQE/PM6c7WywS9xJ49hExyD9+/RdXE9+jhjIVNFzYBysmN6evkk+
27F2wWMunkf+xHz+SHfq/Li17SLcBG6sptmeLn/DF0EKLdgvPN77F9EarlMI4K+g
k25Qq6OnuS++r7QXmBtbTekeKvhTT98N5gWCYeCafYp4vYgEf6emcP2UJu8nKJDX
HaYQKtxBnihrywIMRkrpMe4L0DI6aEW5NuCzrf07oIJK+58FAKKNcRBSV9thhAyh
UxHKTXcKjARWNgLjrM3PtbKnmoHQTmht5RLKS+AMRwCBqQwUAwnJB0fUeYUjRO26
GVv+8BIiZO1ceJDe7JkF1oaInLZdLpMsk5LTIdboddIjmzw0VXFGFUy269PHpDTW
5qf5Vl4wfuvXbIx7C8d4bJ/BqYVolk+pdJN3v39xDdikXIRkAjluKscIWUGzPUuZ
khTIFbL5uEeqxXVfGKKcBqjOtvdpX032DtL33nW3xi0WNFcqI+QnmiaHjlgf94m5
eY/HB0zMCPuo5eueCXcX1Z558erBzvGpauKUVh1M07oyJdN0+AYMBa+DTDMkFXiQ
Lm2IgDbmCL98MDMPckzQsP1SzyYDE14JvGwB0DTWPSzmxL/ho64bIBUl6TE2ukDx
lDc8p8vvY4pbHx2rCv2tN19HiQ0taDEWwsyvXRXq9zu6C34QusJyzl6OYGcuyvbS
nD3gADbaBhiCjyuZM+wCAhFVrqSamcKU0ghe2JZSErliGEBGfPQAItHizyJdzB3j
AozzNLLFYyPCMuDkwQwXaEqO/e+aG3BAGdoIUMRmNN4aCx+1VD0wIdoq7svR3g6X
NhjwiGWz7AjSCLAHENmQtnKz+yiRgXcTBum1Jkw30tLMZXmF4yfsgRYhJSq5Kabp
x+g/VEpwNTWI4lbwkJdAyOnxiq4kVFexvIY1cj+H4HNv5A5v1h1k5xpXf9V5id20
rxR8qOSLwfELamStu315sGeLM5+s7vLe/RBAGlIcSxa6yisKkMPLT432jDLXKX6y
RoLrRZ4aomo1XZSrFpdtuXFUNIaWlpNTjfsHIRQrJ587nTwmy0e/ykh5dxZ1thvM
zMjO1+8T8qar4NJMnkFb5XdNm6GVrmzj7HvcXfAhs2Xpt8tH8uWgMv5/0xeOUBSr
gx1/9xxA6RgvTZZ7yYRXGLLeZDYi4skLmXtj8yNaFO6q8FTbPDXgK0eLA1Z/BxXe
CKVyhoJndzAEvjo8BRSiKFZCU6nvtXnTbpzzZ9mBjWXYucoLJejmpMWx9n/kxo0/
rdWFvf9JGbJzAp2NBgBaI3tL1W5Uv1qqGaMigtwOGLFJSbz/YcRPNsk0SUHAD2kT
qizjn4vUWffssZmS7yaYb1lbu+OnylZjdit1R5A/wBhWXGghYFg65Iw98zg4B/O3
whnhzWZNPlSpC7jCkEQxbRTtsJEwQLkRQW/iz0y+MBfR2Z516WK3IoCn+J+MCM1a
kDRVthWTdQJBT7gVGMWtsBvEGdiOVCYTUR9KERl+aVeRZpQRv69IezMmGbcBtYrE
OycDaMqDk/Q3e0UGaK/9xZDapzlMyaZW9BRAlJeTVACN3TDSz9lpt++MlvDC1rrV
u5/JjxPlrvB2ckedoj9Tk3VebdwfXskblXLvSAxdchFXgcjYCp4d1oLC5Y+d+5bp
gV4nupGM6/9iDwk9EHlBRuWL4AyDqLVVjBKXRqKFEDYcRNe8dXpwcDKZVnnyyHgt
Ea/qf3pg/cSMDrZfJvU+wyh8eDNx/9w+tOq+UHc4Hb/V/prEk3kv9cBat57LiEl1
JtDJeuL6XWwxEQChUqigKeuWM2RchKJ4EbBPUWFiIjgiHWCKdK+Zfqq4e/atoGTT
8KGfZpVBnzHcoowIT0WVAJGXtFU1i2Qp5NMG4MoeL/K8fqkFMY/lhr/HASUUqE8E
5zZWEXnoAVZZq3qMx0pM/G+8oYfzrBcY3HarQJJIfbYOXBnssQSi9BVcQgQqUJv/
HSAqsd74dHJL0ovKRLUylK+BWCDUAsUN2VdAxtZrtNtBU6oN63lSkwdVA22iO3Aw
0zIHtGtVf0MEWIukWyTMjHffdbxjt8JYt8itAVxBrONBG5LjY+CD2ul3j6eGTf12
9JcnII2/np0iJwBBSCKpAm2ZBSQvF2Da2byWGQeVtllujBDN3WZ0NUHaLGFRkaL6
MKvXllm/xzamcp7mXTCkRcmVlQTtQkM1YGuNJDYm0SqBFgs2L/m80W+/puWkKEUi
kMvfvjcyls6wF/ZJBM0Ij0uSoA0/7vXJAaZeW4rAuKYoBEbzDiC6AMKPnxOjhGwH
qzOBU1Sh7BGQdV3ECnPS8oYGlnbDJqJHHe08rNeDUJedzFTEBb8yBxlc97Xot9sy
fSHC+evQDnKjgcroxjeVk3T0F6KHuSKdr/h1sqeCpGZ9R8p6cd2PVBCwNK/qajFO
GsZcAlUca5HUeKgOycT4DwzAXat8TjVdiJE8PQ10E4TqXwKqFirenG0/n0KUYe+t
T5ZQ4Jz+C3yAvhbWI1d047189Hdjz6OrzkgV7MYW8MmbsZDMT6Q1TA4CxOVRYCoL
kYp2em9Y8GhUUyeyvRvg3l7VPXaWtmSm0mDcJETE1ikAb0TL3x7LwrF7uN6kfW0l
n6HyDJh6TK8jsfzE3kelCsryCtx5gNyysHEL96+tLRI7CduKjodfbcDhcU6X75gI
zqqnifOsDi9WzepjW8+/whgWJxk58KWuq7/9qhPdwQka+/lxlRBCZfVQUT1AsVve
Lq8ZcaqU5Ci00f7EZfI4k8afFwAMBvnpI9XrdaXz9+ySxitx7eDdEMqr5AtfqGvM
tCndBLjFinU2Owj/Goy1hCi1S2AXNfw491YOBnOH61UtTQc/bXbYjdeVfQsw0/dy
KIseaayQ54K3WRrIoXC7aRrxqjFf6KZnND1xRIEEAyPkygi//vbBUGyQTTbudkm4
RAWTcCBAqRDPVpX2/GGFFB2HAJ/lLxUg6yk4p1FiabPKzhGxTfTiVQBNkh3XM2+e
2S06qSOfSPtCiNoq4Y101mHx4tGKr2ZArmwOL3mxqD6+f5xzG4WfvlRGpuMoS8Dt
ea19MMooa9NGFrrsIbwYzVkgUKAoWLgJij9C/BP7pxpK325tSbjaProuU+VTAobX
CP/7eShq5J4zsw+4YlGE7fCiv1zSJG7Vx8a/c0eZg/3pLMaHuwUEcB/y2n/g+eKb
RXHaTr7cMHi8TpmDrL2yq8CD3fgvxMH8O1fHRZdUdC24cCLbXqNo4I/K1+uc7qCg
T0hgfahduM/njKc2P0OqG61OM5uL/c6QW4/ghHdxQGbGGwa2mDuu9ZCLU7c46Isi
fB1rz0SDDAfbjwwInnDU7qCAQeLsdfbnhwgzxFpO4Z4MnHmh/lsayfJpTj9IAXiK
LMDRiyarGkmgdCMURluocV8nUxug6hxH/sPGRBJOlO0zE5mynY1gb0RKUbUsfjUg
xqjSFttrUys+54BasRBFOt1MCfP6o0iwJSFumU+6KaP7S+312fh0HildK5Kh+4tp
/mz/PSSp0K51iaConBo9CmMRbZ75tOm6xF5UGUD9iSOV6a2mMwPnBDOwnrUTEU1o
mBMIYG4RzFRsy7FVwSB328Aki07VmlS+t4aPNPv48Bvi9E3ELgzC0D7o1Xfs3p/w
d1m21FSYFf9+P88Sn94KJNHgkxQk0cRUUr4BIFlZRmk/TQumZQIjJiq8+eKu/Lkk
Bjfk7RinzcinDOUMBIhxFNXfy3P5Suw2sCxSYD4ZrlUNHqVvVBlrn4ArU0+A4rZy
DCEmSOc0ju1u9qsuRBFlekRlnDRzE6E1qCrKHxeIevPW0fSum6fKocFifMEg7gBg
N88CirwaMcW/b+O/jCqwq6bV7g7mZGemLCgJjwQdyYBU9NvHeTJ5C6WQ/4+LTpgM
2XO6eCBFT6wt3dyKOLQixhOJKhVPY4DpuE1N+kAoO7ClSUd0mof9pSTP71XZVhbQ
q6xTKyd3guU8ReQ0JeyzuUjdmRzYSfgkvYVGJtB84qwWKuif0c0ajIM0ExZ4Z7X8
QnifPX3eEqEUNajo3uYH2OZZdI6ipi817qtWiFMF+VIjF6CwToB1tFCz0qh5BLFy
piDRxGcFitTwDKjbG/ZkUUK5ohRroOihkmnUVO3dLz7+VayNSy0Q6AL0ktjQ8+Lc
3So0EWPcUjZ5k/ui6/NHimhih2PtvdwFPzZHJ1lLV9OcMHvei5gMeIJe3wfMh1XY
N5VyAnaoHpkn1BfhWGD/iATw1122lr4OwSOwlsyl372Yn0Gpfsvpj3HBL44hy4Yv
7OfHToXlbGPGonRjnjwWnM/GyhV3Lu9FXAQKjddGlAKBeERiNvPI2MzuCF7WUusZ
ElD4znJjFCIW8mwfctbsXmAHiJi9w4Qk17Tb7uYxRX8xRm48oFlJIpgn0bypkiJ0
+azABlmEbSGQhz4zmVplsf7GJLKCzbgueMmBnaElqXqJvYNWtGopva4nXw3bKbBr
JzstXaFSpZZ6Mn2Qutf2yuwyPABRrTaAO6vku0sFgZB7aBHjGb9iFA6LEQOITr9Q
UEw8xfptJnQ7Rj+C1DWRqzUNiVF4Zx0TVPV7RAmgKfLartXkPQXK7ZNPn6oR7rG+
F+/wvZo6CwN5e74Hz0YcWv/gDd5JlPGwMcqiirCUSejqjvcd2AsR5Er45Bf5aqrA
T6/druwEUMcFICOPzj+vcWIcQGaEcI+JPqQLTOiNAyxQxuLkXqMEk5kjUaYpkHps
l7C+ppztCwUn4UkoSR9XFiHY1/stLhHiyBj+05CeSQ/fGjMLThMQiaHlcJKxGzBR
fqKTWEh2OrGPfs20aYZN2hnTnsC+bHstOLZ3I5jiVxyH2k4pGXXwVmkDssMPSxYZ
uN4dL3gnmq3iHezIQiPfVbgnLyC7E3kz0S7MDPq6ewM4K2m7lUuxSbk6/SRADPHl
r1F1xelHlXTjYxei9DP6S17kWWmNMwxT2kOWjwKEUw+arA6sAX0ftxc5GkAdTdzE
ydpw1NBx3fl6FAF5H2NFtjKBcxws87cvbe8mnDo2dg8x3otAAoX0bbYkF5QRGijG
41DFUi4paCWmchMEcV95nFT0ia0lhZ4MEQ8sjOexm+epDlcmmkU0zjyzuFlnMSip
Gl6AG4KumvlfgGcwgNKloCwbbfYaBev8HDykT9Z/1S0EVXCPfbR9qXVOWp5QWKFp
2+wenoKQfDRyIw7U9br3p3Ubr2aM4FAb/9d+Zp5mC8fK36wn/bjLTwJhrQLgib9p
76LPLSSzZLPXzxi9fCfdALVn4KQfVQ/kWzLZi9GmGNPf5FG8tF9uax8d5o5/DnFp
LR7ffr2rSxcgkHQOAg7QHYWqTQibG9hDDzXaJk7JSCCUosY/uzSroQ5SaE8r8CMw
FnPJ2YxpIpm17ls1r+Z6DBEv98syLD75lTVHPj7k8QqH65E3Zy+BX7EueCy02kNn
AdNXRszgNDC2ah+BFuc73gC2NUN4xDRTMTze0tBvmNMQfvIUrhyid8+ytVX4VCmh
hLBxGFHRO/7Xmxu6AtQtIBYBAPqMl9JLRKur3H7L2g3nEbNGV9pbUF888vU01tHF
SzgAQOivQvL4NmKK/dZ7v61pBcUO4o2Hr+sTifCGCfnRQ/LVrPrfJ8vXxReWCLt/
0D4tktGUQ1amcjN1xs4EiRmZ0Np4PLUFLuwXICtFHPnu/kGb5heuvry34VHR3EXl
NnRX7XY/XH1UhSQc6Ag8YcIILPZcL5cjZ/ukCexu3/rveeEXhTYGjucX9ifKEiqU
AcOiElKBBarRia9VpAcheEYd7Zi8EMN2IpB30Nu2NayRKEGDDK8AXbllNvhwYljC
XEwbaNVnAHwTHQk9QvahQwsJaMdX7aFq59Du5dJrzkBaM2o6GvqkISane92FuZJ2
J4Q4rW9PRuS3FMM3F46ZB+NEkpRLvl6v0V2I7sD1uiBqxSOvcQ+yxeBHFmVck7Ix
xFV9FU63bmkH3sN3UO74SA70/W2kIOnWroln75JpRUHFyRGKUQhQO6GQpQprEsAj
cdgtmzqtDnLCMrKQqSYRf+CKdoyRdWpuj2sGA10pdZVywbRZSXYGgFjIzlf/dZGK
bdwDk39nrh0OEly4QVFRHY/XPD6g8dSWCsHiDDF7+6GWkUuI0JicD8ZZMFEO5A4J
Wdv4UQH6Gjn5KzBT9J7mMTGH4slDSDXYLnblaGLryGQNpeeJefGU/QF+Ro93j050
lqrlCx8cl9J6baFI2LT+xBJbxltGJ3JCY5Xvg+geTdr2m8HuUmLcwQPVdIXLC/nz
ZoH12mkUPWJfZY7z+ttVxJJTt7sb2CCzVuZzRQ2ZQUzcCffVIsoYQlYifadh7rqx
q4v67ECeGrkK/vUcH/5v7m5mWrfqWYNFZ7xErTzdLlnG5jfkacXJZ97/oWiceVaW
S2+99iqejiiln+tPuDTpRHH3Gpnmg2c2q+cqW8MMab6wUOixvEJgWsnw0NRt5pGZ
lpaC3yk1ES/tpgGZ18OWQish0MWh2EJI2MOsUjr/j9yaDs33gCVtsQcNcYsjpfJw
48MmDKL8IGdarAnmHEm1IHDzTlPIeIgUv1rbY7Vp4R+25cCymBFAcM7wt6ltJMfh
f2LfKtGlvVGPVMoxkAGxkW0Mq71Ph43sHUzmT6h0sKl3yVlkzSvSiDUVOLCG+DAp
56rPWXg9ReQI3Z75DIQrDVz/3FkCYHVk+/1WyaxSFGsUQgMCtNI5WM2lhBIZez9o
Xb+h4WeWi6RaJpT5yV8U71zCFkrTjAyLyY+DIP5LUy71qpW+60di64H8QS35mIml
NqVYSRhfHw+9o8KEKa+pHqLCE7sQgzZBU8BVqLgpdukoPiICS9M0qFvxgIjYY6uv
HC4YDHHBu1olR2I0PKdXeBkPeUchR5X7YeVP26If6VtoI41uvZ2K60ARGQn9YK/J
nMV9rqiua/2BSJcpaAKP2Uol//6l3skeIaSJRRo1mOf77aIL+N/poYkcD+/jNr0H
EB9LUypbF4SuCtNixlUHxGhFVTEnI1ZlW6LnpHPf2IIAmxBLdJ4UOveM3Q/r0Pd1
nkmb+xxMV20aGkxdir0aU3g7pXqGWv2lZHB9YcQrV1M4FEcHz1PshJ+tnrZtTtNP
GudittdtIcCKZL+x55yHvpgL5oOx4d2y3Nj+iHcJu0DIfbOm8b1gqwNNUGv0sHAA
1Gk9QcCoN8BfUH0D8ybcTyadiOyBEVf0WYu4wWl55fkil0UzYkZHJkkgthoY9o9Q
l5KOXBIxMp21WkpHnO0bmpMsxsA9g5ITO0tqhoP5y6d2bY13qME2JeqfGxyPOzl6
edUn31uNszwLVM26QIinnHGPcMANDcDPFCXUMLDggLtkKDQRwbtaB/+BDkPHeOoI
8o0Pa785ejt4Txiu53Mzjne8r0Gf4mjEaXkO7IramxJwK5kZgUFJtP6fIVTpfMGe
OcU3zx3cEwhoarNZdlVKRyAVPok9QYOH2Yzb7hzHbsg34fOaGYVf0EihgxG36LP4
F4h4E74jkvYo9Sr/E0N+zwdKWgSuLiWwzQt1vLwgu5ovC/wx17tt3bgHNvKJTwMO
KgARLEXjJ4uJ/03ybKpLOCm6pdWgubQy5p5mU4sYtlvPLO9x+/s4PieQPtnmtd5A
tEA91lIAFgA7I/6HnD+HRh+binKeCX/Ipewwq305n22B9VILVElFSR1tYQxpyr4u
2OXjfhyMf8Svg3sP3Vw2CA+GEjEHbS3os4otrqcqmapHqxzoMd1xoWu22ll4rlpo
ed3fpVJu85tgjTaq6s1COdUCmJYPs5vWVLxbfMCBpuk2UUDlKaxvZm32LW8fo1Ib
fGcCbBJ23FuFYXfyZNTxRZoJWy29903T+45Xdr5sBsm/hXCMAWD/LjkXMKdKTLBl
K/vF2Hk59JDh63pYsO1+fczRK08R1atZapuIuwpS9B0Ou4B5oUWESF4ls3lNlVkH
UPeHgRQKerCgiv5n+fIDxyw5Ga8SDKPsbZ/Uzf4RwgSKGEefg+oMacsOgWwf+gYn
yZpktdBmmNl2Bm1UCdO6tO1YwG6qKv1V9o7yIop0Po6nOM3Ds8Y+QbgSnjIRAZem
p8QKNg5egkP33WFA56F8kSQXx0RyT+ZrjBi0/f+puPIGT4PjXplAxWuB++pYZ6YX
R6XPAjaCJij7Zj9bw6UvczMsLGO+d8tf83CuguR7+fgHIUVLeR0uqvABsl1SHqaX
GwQg/fXcHWUSMGY3f1rSVJMKqCb/ed5/NAcmFBuZnRvPOBcgzpNHFy0YggotRwmv
OfbDg7qa8DuiFT0xZBngarTHwVAykqyPpW8meFZrmRXNNJP60WrR3nx3pjuHOg92
zrCYm9l0YELlPyo6g66F65+ZDHfP8UopCMAAaW0J89q34FEU5+Odmb9Cl/D/ZbQP
9C/YHFPHqwh9Yh9jxgaEWPVwFFhsL3VGPQjbriItmrcH+v4MQyZVgXx7piB35Cze
z9BHzjv/6TA/JRkLKgGKe0qy9Mp/sZDkYBCMFxnpIh5BzARbN0jeIu/wz0Uvhwsx
oMGRsSJHq4BaMVvL5gWldjiSUCz4OstrVNcbzKI11pW1ugE/B42m3LiTFvzpbjpX
dKMGZmPymtw19VRvT3jyRQ==
`protect end_protected
