-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
C9TqoKeJogYHguWzZiejDlUU/N55D5emT9RmhF7LFqENFRz64ejVQriM771yTPEqsFLmM+C2G4fC
0DeWVvKNaZdWXaWUnUb6V7F//8pDJ8KpE4cpfDWk8WN6xjaD1ITi/ccFjye6fIBBF0RvHuIaCrXs
U35lEB7gsh/b7/nAAoWt0A3I2J4Fd+xwz52A3Jc0qaBByN6lMK56zCmWaY0VfzkmEwu5yj+lS3dR
+bBhD+w6wNZxgs/Wzos7YQPrf4VtvJiZiyOPqofvf9ScsuFlJ6IiaMU4qWL4JkcP/Tfe4iNHxUiX
f4+/NZViYL4yUbfVUv+FYIWryfoIILyzzE1wGA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10496)
`protect data_block
gG5FoINjU5W2jIQ04/h2SH2bOLmFUNETBy8EdA+MVxPgiDtVKddwnLIkg7L0NvRwZZGdQ/AMmJlx
mBFnRlJMPArqowcYvovEQrLlYihkoELVFrVfHH4ZFV/ieRaN12I60vuC+bBO2gRlHog+FBaYtcWw
+bMdJmKTyhTnOTWZULAOlZc6d3qBe7EreF3nHio6HxatM6S8j8e3gHICb6Lsx0VVHh6PYToz3G7m
efWRXuM3ExYSMUDuxKHhsxhN7qHA05DK/GxicCx1rPaJDPgnFFXgLe9IIyavOHkLkoX4mr7lZELJ
Er1s/9LapY83CoCxrl726QkPVid1JP2YweDXu7igRzSOfpgrrElPtR8Hsshh4E0urOKjWkhbRgs0
spf0DTLLtDIUqqAjbBo1AtM2FaJvvb0VQTd1ym9gzsuRRj9GCvXY7vFlMIpEAB9i3DlZEIH3vLUj
IJA1waoKlCYbfNC+zGYBb8xmPSzPqMnwIqo5VMGmYbR/EhplSK9u0VQdPq5FhDU8Om9WWVaB0XG3
vW8o85kfdiCiLrgwPShHJjH+GRyZpTjKtK5WLCuYkAwZe/HVBgsB6Tth4frGm4GTea5l+TaH4XnJ
FD7t3dA4Nw3EQgFT7Vgd/o57WMFsal+5PQKJft3ZR1eDD5y8WpZy20ILCCipxMjLC2FfkwTZMOKl
Dp2/kCPgv1qByr6Sn5byyct/QFG7VXPt7gIcYChOsctah36rsVLRzhvI+TKDw+xY4oKYXNnhEcK7
nAL0dVxoWZT7MjWQqivBuyQDK6o5e2w0eqg9yj80Cw3Y2J+MHbKYdrQSxumqc/du36cNIpUaIH3t
ejjhtcOUyzvEfyI5tT9ny8Cxrlnq+ddA0XJyXDtZOIG+vIKpSfi+9Z3Znd19Kc1kkRtWUVWDa6CA
7VG3sj5qavRuC6ooNI4fBd8zcd964cCBgFNy6tG/LxrEn9iA+NHkspFXI8BARzrkGNGBJwInmHVM
EtxOXyFTGvOjHa0R+nM0By9M0YJiYOOolHCTXvA7tF/jFer1dUWcCsXrd7+fxNFk1TIsCR0cCLC+
Q9YWob609lon3XbFhVe3F29CR95szIbGvEVHPxxyNZanXfNx9YIUVGd1Br9vEk4bepKDa3967bRH
FB9I242WhQJAui0fgjR1xSciquqjskP3Jbrw7zu4mfgF+p09+3CA4naUoNLvZYnCPnP3Z/PGBMzl
MV4ONkszJ+asYFR75MxijnW0OlXRUixgiPkzYMWGC450ESSVh7p9uFE1wZR8K3TC5o1jmuIsoTFx
y0BmWA8Qq/ajylbMFwmucrA3n0JCUzm+ou0NNUAtoDeJQNr2blwzCxDAe69qwGdoZRvqAImpZFsA
uq8a38d+PThEYgIrUItut/lVpiVfv06dURhPjYxoA+EzIhpOgLk7xh53Iv2dyND9n/IsTl3sCjWI
mDi2l3UH3yg36wqoJjT1AcqCbmuwK+u0Lh34N/q4HwGROfQHEXPwY1z1oCemX+r6PKmBGgymtxJ0
WR3GYytXkkMGI5VgdAL6He2fdaexlrhJw/072Msyp34oiHbRdBrScWwdYuMcaK26+7isDnfBkWma
iHGuQOGtSE2EywvP+6xVTM1lImzppc9YCTgaLnfSLFvvEXauYdjWvJvpKPUl2BSwXe+Fvblp06Q2
x/MAM814fTNC1/3C/i+HXh3oKI0nY5qMIC/j6zxNB4fhiuSXIKdtvGnuSp9YQ37cJShiE+s/LQVC
Bay4VIXqXgT32GDJ8z4jpfjn+wSJCi2hoH3kzjCEqGBddt8i8xvMADU1+aDj3fb+8/7AvnuUUMQX
6FSZcqWbd7P2+504UezeLz+Vg2mObsdD3dmfcqpS5jaoVY1X0D+MefIxDIJHJmf+lVYQigOgWV3/
o3i0EMYIQPldC1V5BH/mM17JpRCPxT8J5HBDGcFPaRrItAd6JoAQwDs+lQrqkAk/LsFhGr2EkGQ5
SScoyZu+a4lIEp/0QT2f6hZSPehSGjxfVtQaUJ3LhR+u9Of2CpbvLkTOChhu6M3Qffm3u4SR1HnZ
A38YuzqTxW5P4yhahSog1+BrVsLJcaFfsx6862Z1sfy/Ul3eHBzAWMrVhpXDLApngYASV5bnTYk0
IT3GgzGsiDLxmpzKBL+7YD2hdXhQ6OFn/YJJRDGOvVSkqXkVzDMDOkMmK8FENEMTMgOdAfYXVWWb
n8YLJRgtSfVq47Nk8+mgGmtY2JcnuFL6UdbH+VW1UsFyIvh9sH3pHQVkSRAWEzU82fJuMEeQ/eEn
o0Xma1/SL8qUgg1BGYDLl4orVwtHtM1zJnfhvIwUs0wQYvK27PFV5aQnojSlNV2cLCJLvTf726rm
mGtZpv2Xdko/TwcEzAfPXDJA2rTEPsxhdDr8AdY+rxQJQFwj3Yiw3UZRpdZRTwbCnmOio1vt/xXe
rN9Aug3Iq7hb+nxbc63Da4wh+eRZkixxD3WSYki7ioHzeEYu+ZNWWnG61aKDJ5ADjE3rrr11JJH5
JY2cdIKAeesyIhjrXv5plJZeWuBZ2sOTivXkiNeQr7xOxnZi6EGX0FPCKFpYQis5GUiXimfRndXo
WzuT0bNhn/fivpVfdpcmbwRkVxPqIU0SljmDLam91ykyq5keZ/aKnw5PLV8dyvBooSRu4WBXT47/
u8rnUYxBt7asnRKeTabYnfCeD2U2UXK0TghYthVex88Sq1XdYnkQnHQ72ibftRHMNSeXT7ndZC61
/lxm9TSaAkrYHSC5aRnmytdsySa5DxfMJ/wK6bs9S0jka840l2B1S9hEAyeT02wgBi8M5LXHjdmY
1nYGEk7vqCq31DPe+Z9NdTnBMdluV+E/FihHUQZSnO0iPW9FXYGlOtImu7A2krJ1g07bSuz8g5/l
BI6W6XWQjC7B01YSz5cAwxs2pAV9o+psI9M9KBFx1ZLsmAJ9Sqzrnbd852JVT33rPT6g//EfSFbh
/76IQSXy5Fl72D1Y+qg77lzCGMbkdPEIqfxaTtvThwkfVnswX1Qu190/dYFt+YhvaJdhZQZnm3e4
C9W7BOW1nVnZmwFcigM3ngjzFTj0ZBz/+klhPGSrwX+mzJt8cP7PDDssFIBxQbzPhdUlOvxS3cj7
4pXXQbFkXrx0e/mOxZ2V9QDqUKADfVshSMJUu0z1Tf0LdUa53vLNif/SazEn5pxcoGHGZDvkmG1E
hU4iktsU1zvA32EJNcvpKb6A9dDjKY9WvPpJfr8okhBHEhMZvtcvjeXC7Uoo2Y4N6O5WqCbmDy1o
17gNwTvR37dLZlN9pZNspd5vMPsfSUEe3MNz1OnHi0gHpXngKTBqfocgSMn3ZwggK9RyNgl3ccMZ
alwSS7fceQkf8iYzPLNp/R+ayX2NqaQa9qHCgPk0BUuJI+AEMvjHf69QACCNXBEztZBnQnChZJja
PYMSbcL6se6VmfsCYExZ00/kPOEcO7xudRjANlFQR4EENjiETXAfF7zdY2G+6dkQoyo+pN5lbos8
RBxXBbshu+nXOz6UTAcBnz/c7ibWjV+/kzwYmseJp+ubnQgb34FDSA7l7UVzon23ZvU/59nnRIA7
IYY5qCI54yVdybRdoibGqhsSwcQbb/96kKNAsVaDnOCKB+qt3jMgJtZOjHsHg2fe8iuCM/6QOIdq
GUBiMKer0y2CnvzAtoJhk0lrbdqBBaoF6yNkSutpu1xD32JU3ViHqlbvaYkYgD+iFWn5zgImDJ3L
jYWtfaqfYnVl9N1tz9DDOeAbVfSENP3J3mdR3BFrWx0UBGX6TIm5i3OdXHXeVGwxAvh+uN1Yd/Kp
HZlgJx1Ht2/eNUzz2vEy/a4RtrEsC0NLdC4IcJX0y70OP1ZPIS3XVCNiMGaxWmWSYtPHwK+iuYqK
sx3DXXUCrKkhm/x2g0Ki+LRC1HTh3x+42NbPQZzC5xFDPUvIGnxZknyDcwLnfJx86pzcL5BgQNxs
yrTSvLujbRr+hEHryfnxRwIILRFmpF09z26veABS9szRbqvtq3RPw0FF/eQVo3BP3MzBNB5PF3t2
k/bF5kgsUCso0que50K/SEDN5sRtsH0U3BTVcUlGrXl7B/nJfLZpCMRLLTEci1uWv7IlolLmrla7
x+4M2rI6dQXtShiPUwUN6F307xrssYU6U6IipuXUxaf+g+hm1CCC0bz+LSVqM411R52HukGdG7KC
+AAQEgz3p0aOyD35L+CVwVNCA5/AFdxgHNA1khUagcyl4Fd6T2x1iCIkpu5qRWxdkxe8UXVnxLh/
gKXIP92ILgiWQkbxd4072nAhNXF+fj34NjLRh4m80GAPdWiLjA3VrP0uFOvq6RguQzZJ0ouqGwe8
hEDqbmvp7ExXc/JW60+7pwM6svJ8rXjDClJmRObuVP35An2Srw/hf5py13Qshl3icf8lTt+mURSk
86xLuL8BmhFwPQcrLWThaWcc7WuBQLvwDSBO+tngZTQm7svzcGcUmhryRt7DPxixh25kquw/qk8l
VKucBxUTxCL2+Wha7r76RIHmvTXP644C4vBQWaSL2Qo9MPvfHDKhrDPYiOb5O62J8lQTeyFbZoUK
85gSiNu2TRX/aLr7MpP4W7m4dCHg//LYjLFxvFLWFwZ3mrmFmcC7POiA/UOj7R2VYo0XZJgmiVpS
tlkNpGBa6JdQpM2YTV3lQ8AfjjOH86GKWoHDId83NxI5hwlxQZ9nEr31IBUoaz2+oYAmZrUtkvVF
aJXIfIk/Je9MK51QgDhmSjMXYJhfvlQVmYsIdD9OOOrd6npM293pUcbXAWw/Ldweb41IcWNUNBk6
52ssWN9K1WQxhefOpmDEmrGwbWGCVNJ64o3BAl28bQ1bOiPKJafEUWwH4v2ZeGTS6FKK654wsiBo
OP/Uu9rqVr2hCKtiazKJpCVi+ZXK9w0oMiTa4PM23zA6u5NsM4PU2k3pTR3yDgkPF5T0U8fD6bdF
FFNqH1fulfs1zmt/6Di6/2bnURgdfB1ilBk2bhsV2S6POtI2pycV8aBQb+W3B84XW6s3V/wJPTrD
dM39mVnThRdFLGlgrX93aQCUsJJ1vzpbGTUwNxrCJNI6c5walB9FgR65G4H+OYOiDbrBpSKWofyL
0YoW+OnMD6u65tP1xnPc/9xQ9YXpTGZOBsm1mLG4gN1UwzgYeuXuDXRjUMl2yU+XYC0g284Rg8Sd
4rDPiIO7MzJc3LI/UgXITvKWjxZzO64bThf5ILBR6bxZ39zFYavjnOZ2GW2p/qsqprCJsk0/DOYB
qrQ6u/2UvOcwidnn2F6KjHgydopsfhx/CXolKTv+uA5xJjOP/eNgn7Kh817zhVpEVZxQZxOnxRGY
indGASb6ec1TtpPwnAWJFi4FNg+1LzzRXSQLacrBH3qt1zO8OILN8nQbYdgMn/3qL5QP3Egv1il6
6bwbCG1ll0rnTIr7DZZp0dKT7KGsmP08xsMK5DIL6elTOrDrLYrvFdshSIfEV56BXUKL7bDtcEX8
u8efmSRow/vjZOAfoIhD8vk1OA9xhnbpGSnop7A2V5rOSharXD5FRrRZn/cg6Ybl7NpH8eG5igFN
sOk6WP37TevzJ3XimWCjDZ5aGqmkNYciYIDu7D4Ir825BMRJKjOIOri2Yz3L17O/B1MtSEgNBZ9f
1YYQx4SzuegZXFj6BjlHolr9Fyj2MQUkIr1F1FwTrPWiddt8f9QiQRCOv/kTebrSkCh/jYNwbp0+
ykjY1zvBNyx6pAls0x8qJZCxjdZtEUQ3QLsgb7O2Q7jru9/PW7EkrCUrqmn2PtnBEoAUPA69XD/k
jGCZ9ZL30m5xRpIQcPBfFpFvoIPYzJMa4UNE6fDl9ahJRFa5ZlQXcZ5nLWWcJPJnWpAOqVpQtBhB
FE+lpSgUylwvOl9S7Qy1B7UtX4q7ccMPufX/f2mSXq3OXz9HYi4uU3GOvFRCK3+nrTGw9Fu8tJsV
O2KY0DQ8TWKIoiH3/mLv9SgOAVKrmY0N2EYEXZIceQLYEp0T4sJzyE59IdKgQXFaJtDHWU6JdZd4
4PNEPUweM3EN0SPXmqHJqK2C9Z3V4yT3Yn0NttF67FnLhYi/T0iD9WE010E/busZZQemYL5riHBt
6P3MA5ETnKUDzYAC7Mk7nmoyHlxNV8PGTKwXxPUE1kjwk74jBsQhWGvuGMz8aidDtcKGzUIN7Rjd
kmp40Lp+Unu39iYvnrYh7Ddfp2Z6kH72I1NxPZCbvSTX2SmHDI2FtVEPyRTS+TF5eWELm0SSMBsA
uoqmHPHVz4RuCNJKDriGHRoZCdXnbC5h/i5JWD90gbsVvNQIfM3s+NIHIdtWQNRvocazbZXLd7Fn
sNke/faE/Xs6+raaI4tzc92WKt2FCSYmhFvITqYjbEvygPmI4dVxTQ6stxc5DdfKywT2DqR8VjIn
0Hz5iM/9YyC8mU4qpWfh+oMASXvKLAYfvwuOED0vytVtEPQJzBtAX8UDEysdO1DxaH1dkjLovvzw
YDNXNNL/UIel74+EDouctVZ3zy3cF5MOp+yh6QxjhUoXNxZHVkj3W6Lb9SiSGq6yqasg/VdCH+WO
p5rRaZ29YrcmmyZBhuKRMPzYguON3vsgIN23ZI+KVAl8x4k65wISt7KJoY1mlnOHAu/B9SO646mP
IYACaC0NiQKQ21aMJPLppXdQGEmAVb/brWZxl0hA72MOq2ea0iWzwAJOC8yeRPG4mVwLGfKZGnHn
jX/74+ijcsO4nJ6pnv1iXfBwHACbJJVwZWlVSm5fuQ08mhFPfRmaLVoBmOY2WVbrvx34Ov/fd4m5
aFRfI+ul22S0xGAX7E5R4FKj/3Zt0a9lP/QkDfV909SDQic8Nld2OxPX9nI/L5bCmPZ42uaOvckQ
FLtC4+Qa0NY9chToQ+EUkSDpqvzW3ZWznsZl8pbo9XcCi70CCJD7WxZk8KIqjGtrFp2yGXEelz3o
MDZ/8aQrfRrw8jLk43o0+PkE/XOSOAtPl34wUi6rIOe1ir1gTseZ/wdv2IcddJQpWPey01U6uaDD
mZWX7KZ1jX3XCEUrR7299ji1vPvAoDQH6gH8iMkKe718mE9FV4GHwEMYrrprUzrqhsOgKXRWh2gQ
D/wuYQfWdk/kc+Ad49o9S+BqJni6Bq6E5LRhXpdaxaS6Or3ncYJKLDjaHWRSXhv6Y52V1z92lIlm
2HTcoeXQW5GWyq9y3QSLRu1W6k9fbsaT4ZMyC61d9T/PM9pyqk78zd+16c+4ZpWf3+JQBYtPe5s7
im6bO4tDUIc95DzHXA4xvHSNbe8vnzpd934/qna5V6/UuG41oY4KHaVVuKyuk33Y3mCLgewlFdOj
Iwr8phr61T7fxA0y+RlPd41l/hlZKTJk7JHvLCoML1rFO5qDcKTXTr3Rxr73oPUpWS5SnCdmfW/7
a5igBHCc+SrQodwQzCAl4ZhD4WBtw31my7SOz1ngMtPMmQ30AtoUErvTIYQHD4iFsAw22tdQ51ml
aJZfCgoQFwQi5i5Rk6gSSUO3ig2RPqEIopGH+8NQDsp7EaCae/Go1ebIFlpLj4nvV4rOw7tPKjlT
GWClEJeOA3quHflSHyUtderMG0wle322jPWSzuhu/n+RIwcQ6yoCBP1V2MW4hCCuh7q1XjmpwYPe
b3SmFqeZtKGb7NUX8U0O3VFV8sQ37ZeKklXTlhezaFBMypPLGWY+IZKs63D+h+Ko8Nj659BUlOBz
j3cQnp4PWGuiDpVo8YrWFeKh81E9hbxzw3HQHSLb5GnC0HF3/MG/p6rCdTZ+QEIYnxvm+O4MpzKE
c+tcLQSaf6fp1uGDKKoPpX+kAZR58x7L/1yMocFqb0p/l0iJprmXSidG4+D0tVOqg5oMwMM9+CjG
ZxurVqBqdCHFM+BOtCuwbAmNXqat4BukaB2DBgVCdw8nrCwVYIDeRx5dhEOZryXBmu7/26wCFdwD
10dnQywpmjgG3D3v8A4VcXSE78GIGxuYBpDrfo0zOnNKj5RSAFU2O5EpP5j+qX4yrdEs8i8VaW0S
bksN2CSt2Dkr77oh93vEIuAxcQGuBtccmS8AdwJ+flOk1ZKVeApaZ+bcZY08pGchw1aq1rvayfFP
CJI4Sw28Pf07YmJo07U8GGzvZJTQGSfP4T99EQ/5+ydc2hyMO5xfjaW43tmoeJYCzFdlPVfTOMi0
UD2gQyAttFS3gf9Y/L/SRvLcERFIZWMuBE3vEAO/Q2bja6OJTLfZwSdAGT9BF2nrmQMvTzMQ8/U8
4kQHGd2BOmYeSAix/VJ5LI4NNeGZjsgIVQBrSKqy4kfO9PgqO61+18fJLAyYbDl3x6LRnpKuv2L9
S4Qz3SHyLEsJhCzffZSNu5VHwMbVevWLMfE2WFJFUT18otdgF96dp4E9tFVsogZ2RfvyTyPY6B6h
P8dgiyTkvr723tC14Zbl78oVt5B89Qla0SjndQAHd95uI6J6wHaGm8NZfNayoPz5ALwHlE5V1Zxk
cWjlWkGlMHqE2uChgKhJOOnFsKz3RNESn7WM4hZk0YPxe/Gz/+G60Ym1DVO8q/Gv8LfP8306L8t1
cu3kZCtEfCWpHx+SofvBqPmDSVfL1E8LNxz+pDg/YnENhAAPggLzePHEg/V5NTgy+/kSjDzm3n1U
LZN9TnhyriUE3TV8gR1E23YJxYERiosjHr0YC110kh341IurFmDPfFOb1vSZf1UaYY9l1TsBMIAq
jnL3z/+6Mpj5MLUr3IAP+pemo2vxS/fNetzTymHX8j75D7aOzB1oaBiean/gG9HQeG8NVx8ajk3j
tThkaxWoDBbQvkpd9xTNdyjPIiQn1BSd2xEi94fSzb3Q2uwG6LCm+WJJ5VxoGj09ZCEoCTyhbrUG
bEGF/Ze503IviVxYEm1rHBf+tjo7b+RT2Etle0UfT0juZvETxNZxfLe6r/HVnb4PnKJoZDzvWItQ
GLCeUHtExAUxJ4YAJDQFXNHJnFFI6R01WFGwvrBr9aCXud6xmmsnNXIKWuiWjzriI+j4eo3RaT6k
dnKy5Q+KzCmOD0dhl4p1sOF1wNY7jKLMUt7A7jNmocLoP6LTgCHftJlqXb7TPIwjcxFr5cIEAYLr
GkSI/XDSx+JMvQXBKu0djU7W5RbWVNvo0H1RlsUVIjPUSUHi/Gx6zG5WYVrGP6J2RwwhcspdFODw
dDzl9zxCMNWkzFO+w28IaVk5QornS5aLBFBD8Su1jerB372Ja9DI0Wa1B4EpdAuWGzIdkB8d25T1
uingPzFBjU10nZkcSDpRM0iHfJQh52eg0rZP46/XYOF9xpGWA+1E+feM7vkmtKg89fe/rYqYZzAw
tvaDhCu9berdMmc6G9CnZD1cwX4dTW3P5WFHj4DxgLVzr3vgzYGOjl/oS4hFZql7b1JVQlSjno+i
on++l/jrJdTCj2b5Ezwj870ARLjO5WEMdaX0sOrd24DRxwOL1E459TFHi+WgnvQBktzZ3xaKdsUv
tLDLjAQFYZk/CiId7LDuVaMJ7y2qdG7PTGlqNfbNONnrERilI/usdKkcE7P9Gz9T7fpTyoREOgYZ
Xm/hZA/e775c4+/hpBOxlxZwBfN+GfkQ3jDKadMxfBJHDD/F2kqFi7BA7+sGGACj49E5NoXXCECD
vmLjzdZRcpoG0SlVZzR7EzpU+d6s3TW8ChSgmbaiNMDE1Lb/+O49zSC2mohMHb1Tuvv4eSdYF8du
70p5uV/8Q0TqaBIUF/MT9WvLi7pGr11AMNLdf86Vtd5Kq81cG3vy7eaOQ0b0cgXiOIjeDBOHPybm
c1SFn6emJY45euDz3kovd2A4bNfMx0aQ/bmMQho3qeYxrLAPejXaIntfu6IRgMsVJEJfid/Yhsl5
Ee9AcV+rEYcGhIb0biK2c0FIaPJx9kpCFEz2xSzAAno9daC2k6XrBI0FWILkHShq5xgTgtIAZ65X
X9Gc0tdNAbn0N54hE2KNYQEIBJoO6//48kTxRDMpzPBKG6QHYdFyQzL4qvn09AFrmxzkmCxj1vDV
aejuq2p48a/Qy7WxT/S3VjWWiafJVW0WcTdSjCjGQT9p6o71PgVQYR8Noa2BC+/XxLzgQCvh67vi
e9VukqujcnK+0D8f2z5Z/1TGy8ue7HxOiguYO0Ay+ib0q9noAYzEULJrJ6Rc8x7pExE718lr0wng
9+B8f7eGbU9OQWNNdOrgjbfpJZ/tX3l2ESNuNwLvRiEH1RxhMN0bRqo3LYFZ6Ukrnts71rOC4Sxm
iTtVCmZd91GuKNuzcME7+cQer5wOrzYcmPxLVJJuzR0rDCGmOVzBYS6Nb3CPdT9Yb0B+W015Eo0i
ZFNqq6DVKNp7umeXgJWKiEd0kUXyHU/7UJhQzR3Cx56cMOD9RSd4D0LiwYeXrYgy+DSp9/s2V71L
z2rM8EFrsuSMWdFxlaaF0ZbHLIx0ElCj+XeG3dHCLR/RVxOwAthMLxhITLqQ1046NDQCR7+72Igm
TNKnyqDGay4ksI9nq2R19YWyM32Yoaz35JTMdcQzLhXY2v51w8Xhfvp8rrlUa4Bt7J9YJ/i+XZUa
XuCw8Nafkl3srlLJeBf5zA4/58Mhwvz6hpdHmgjvUvjigEi9JNh3yhKtt5MBpbr7hn3XjaaaCh3K
sgpfd/eBc9kSXQx7gGXqgFTHt7Q9FxGUUc4GKT2xF0b2/Pe8a2H2Qa6VQuYyB4bXyid2bqBt3wlR
3O2aq9loCaCPm9fc856ALzfHNaRbPj9KsVjsquifkK+M3GXXOxcZX/GIfOouM+gqSk4frvnypMPn
4rivVU20XpzCYxeCcKbuQoDU/P9xGvVYM8Hp/M5VwfsBDaW6JsCJss60EW1CGDGi2Mbv/H1zq/d2
AT4bFhKmW6a6Vag7FswxAnC73kicC4PNZ9dpjtRr97b7f+TwpoQQptzOSG+XpreEK7I2+Q0GN388
mvT9x+dvd5RlP3/8uW68sFuxIY2QNBF8c4d3EqZ+8MZd4gijW8pSrNhUuc45+4msnJbJUGK0lytV
Cy45Y0hAYkIF1AtVI+XvgL6K7A+ZrKfh6PJWiCvfZEey55TU2K1DgNWzXhKboZytN6+ILKMM4Aiu
0B+5V28R9yBE4ql17O0I94TL0F00UTnrTNJXGjDVbqwSACZSpjq/LhiGw79C64RYrujXLVmV6vDk
j69//y7fLB6Fj/kfnV4n5rudNHconYvaqOhT4Ud7UmQTaJaJV4YybG0ckAabYp16U3z9C8fOnRqz
PmeTUFbmirdq7iADXyL0nJ0nfR69kC9bGCzJLX/IhiEa1qmWRiCSGSSTZYwhbJFocIc5La+pT5/H
XKP5cg/5/5a6VMVtJpZ3dAxjfGY6qdH+GHY9PxTKSlqk1JKj0WpJYrJ3/BhxM6GhEG/VeZCD9V9G
2D4tVPxh0a/Win1DU2egrK4psKu7bJDO3wx4IeDjssO4rTv+7CipIt/dKz2RytP+dPtkxMxbkCVJ
8WA7XaDdr2Q964H3t9h8cvHJkGqAiJPE5H5lKjNEXPMEDYwocy78YzuiqWsOpfAjMIQt/5zIrglM
NVv017g5+BaUpxZjonkL3IEOwus5auJj/Su9B37n+3+WcSBmKoFMG0Jr7QTr8lf7JlQCtOdVTYZ8
I7ThJDG7Qmgi0dbaXqJSHhEkN8jpWh1GS3q/Am+OHFTDrw4iB2zEIgXEQ1cO6emX9tWTlGs2mdH+
7P+QAIgs+lrGR5OVZPLagbzFC4C0XXe8Zoxp67/yvNpEvni3Bx6b5jLKDXfCHfLx5DumnUj+v3GC
caB7Yehpwugw8kmyXC3wZGIvubsiEhYO5A5Wa2YMKZvO5Nkz/2uxSU2wb3xzq0YJRbg2g/opIIm5
fsJo+uNaKE6AyS3TRjyazZi6qg9ABL7Uk6YrjCPvTLvy6xmSYwpHVHNF5JomNPSkncqNxkOPq6Zo
T4DZjOMs285zhFpz9+Q33JHPDUJLYHMmntzDhUqopsR3kaItUBOGV5b0hpgceled21ESIAUDJFdQ
xMyK3aWNkXgtgGEGLgkpOFwoNlcwzsW6mQSG+7y3zG+09EVTM/0nF1Oosp9HpBsjRDa4srgx9QuR
/+6EvcGJIxb6glnLv7O+0aBflpQuG5aiGuX+wacg7OLcvs05Dyui+c/QifvoyipVRPHK/5jMjeh8
NgdOlleBZGQT/KM0oQd1kPU7zPLHtC+oqMeXZ7YDQ+Vn1KviGfsknk2Fu/mdwCziozl9+6xuIKg4
f2LsCogcsI+j516SkodCeyl1doXbTvQ/NTt1AV3IxxSmWrsYBQCBqvylf0DCTuquLhTtp887kmuS
wbn0PQQylLIkNAulL8lIJacSiYnMQQVUbjTtiLvEw1AW/CDnFUuMF4UD59yfVSEH4pprNI3oJ157
rR36YdqaqxF5inCMy87p74yhRhxY990rlaQptBchdJ2uUpQpVtmyzhyBT1cwHsEqyV8HFQLbWFwl
23xPMI3UhIgZ3bR9JMEfpPbioGo7SEkiAaIYWqD/hqJWyRtu4IxilTO7X+W1aPOX3QSY8+uvxFFq
X3iToBxpc1yNXxR2i1XOE4RRIqFhl4Fz9vH6gfInmm/gasUGd/EIoGKOpbmHjutIv96/5aG1YM7S
2nxBRAjak1TKVSG85UAU3g6z+62yz9bT7bhPSak7wmgANnV/6gCZjxIZFb+pQV1LQGr5KkNcKbqy
q9rRus+HObvRCLdUPXvi29xrKoo1t+wk81uFTHnMTDdsDM6+RatPtYkPPiAinWz7nkAMSJP1f2Xx
LdUbrgGE5E64ARLy83KKYXWb1qmUt97jEBKeL5MS4QYBe6EtMgHDNt6JQdFHH3uy9rbWEjoeNbnG
dHP29qhcajImpnH2DSBB1xmkMTcM6bxkkQU2aRo++0VDv+7KoqCOTbSu4rBlQgWXCC/T3Wvnc1Mq
rYYv4cCFIEYUmXo5aF4sLVUVjYrVhxb16rjfZHrbNWaEPV/2Cg8PGWsgEkZq4QrBnbPkIzbXU8y7
5HPI1QPdkItavjOM9biurkJaWNF4MeRs/amvA5uk8tvxuz55QNBI4lhrT9w9Jj6u1cl6lgUUhHzZ
eqLPnB8ZkdmKq0v4DFwty/DnX7gnFWo+etE8m4B6wBp6r6BeiOm48WEMiG6ZB2af/H05gcIGo1h2
OgdVGbYEi7rrHwrJm80MUXjm4Em4ltAvpb+aA3pFdaRjGuHBbwiW3vbWgZbb0OON17wBsYndXaoo
EnnCBjAohD1lPlArzy0B5QW1wh40AOoQnepliDwUD6bl+iWO369vUqyBjq9VQb4qAvXrmI8E1aP2
sLAjGrAzhSd27Y4q/6X+9jCHsg0I7XbelSZZ1iPfSWXUU2NudsUiXMmmS5XvXtgMfqWOF0EhVa85
38v5N3ZZU0hiPg1kal1MDgW2/cTmnQdA9mC9sKVvQwMmvNayRBBK2g+no4rE342u6O2doDNfpzfn
U4Tt+ACwm9GWWLyPFWCtre8s6u2v5T0r1+FornInkDFNS2zqDsWdb0YxcOisb9/bm5d/tVGUGRqP
06OLC8Kql8neMgrTMvnHNtLIr4Og83zHJdb7hJbP8XTzf6V8IjhPJzrVK2OorQH0EFViYIe6M/CS
zik06F8TOu6SqexS9YR1OqYnuCaIdM4BgqL9uKNL2Qg4t8UEWHrotETzqhOiYi32KhsOmKXN4csp
o8kN5cIqC7suwugUSNuE+zqIFY4xw0eLzbHLcX582OV42j93suSF4UjpJpJ+qnFgTs1ajjdc0fBl
uf6M+UbzW/qK0v6pXNRX1OgVxNs4I1XKv9IkbKdLpb2eFdEBXDcaAirtMZYsDeRXGLuytD2Ix2bJ
jWvL/1hzRludfQGeoex93YPCwfnYPn2yGiAtV5OJPfma7Sj/a+MuaS/mjQBESe95WpuYQrBqwLf8
XnFowU3FtX2oOHmb7VunePPX3S8r/BAgghNg92Ea6UZVDuUqQXmTJZnvt7cLzd6z2LzpfQJNeaKo
MqZPTmhfr/vh2uajgKN6onkWAnShfmQ1OKRh//3ixneLLn2vRSL0y2MrhjY5eGIH7EDbdHF+I6P7
3UO+C7gyTaU=
`protect end_protected
