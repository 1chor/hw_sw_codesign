-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
B1JpkASPjwDjhWuTDWGM0WWte3ZHM7vOvyeVrsvMKPvD1140PXxfCKwfxEmImgvF
LidA3VOpM02MW8k5dwZ5NJ++3jvJU/QAe14OvPY2d9Y0f9xCToNsCDb9Uh+2VAzE
Vj0e1jkDYhYb1pGdglkHWXlr2iIjV9uxQMXcFiay8I+vlexcgPsq9Q==
--pragma protect end_key_block
--pragma protect digest_block
+Q9J8xlN9or7/ZKSDLvLSnHnVoI=
--pragma protect end_digest_block
--pragma protect data_block
rPxbPh4hNE+qVhrGY+e9K5bI9akVpE1IcwTJHIleqT41eD695az6fQMRR9g2IN1o
nr39lVFEI+KTpbFKuvGWAZitBJZYz1R5vrQOU5J5b4zc0l27NVGJkuT3lddCwc/i
X/B2kSEnNXyiw791YuG93vJZwHBJdFbigP5dcwCwt3oSVlm1jT0jQBU7LbxrLzFs
iSeC78CDbeqxSwDaZzKVHeMecDKgtzfRWcWyaERubDve5u0JDNYV3mA5vGdMSEyB
h7d13DW0AbESnw7P9qQnO+aDUWzihiLOCoR9+QCM3F4R2AVuqPl91Iv2PjH/Y1Hu
Y4w8Mi6geYXuevOjqnczywAHmdbYm5xmTw9VLdHuCnrGikfOw/j/wzMDLJiapIsH
wDt+/rFPyXOxCG4omrHSB7XD3UtFCv8p+swamB5lfqyJgGOjOZSlJpzwBAhHd1Eg
uIscr0/YiWOKczMNtjv+527OVZ/NoBxC5JSxouzMBlJs4Ccxr6Gia+LxmfwhQ1qz
5Jto9kgMAIx5028AIN46bDtrdAp+hY28QB36NEQ4rY7iLnNo2u9WUxOxxBqhKZms
KKHN73Iu6/GzyySlisVHETP7SmRWuy4HXxr7DuX0HTeD2psTTzwbNd++xLb7imxo
xw5jN3asW5rlEYJUVeJPSzHmIqVUX1urzLHJLhDoGDo6/nN4w68uP2YTvnH8s2ts
BihPF8ogvxijC8H3iGB9GXbtPb5OzpU+FjeXhPB1NG47RYDuuLeM4mWsZcD+05RP
sUqnw7DmAZp2wGeov9DdoPS7nXlCWd8yyNnI/qGED0D/n/4CpgYCO/v7SoRZ0s2h
1rlxnLJtfvDnuLvqq9CtCUNdkjRD+Ctt312Sl9J2hznoq9nsIx0ugqM5ei4Ctnhm
SI4wZu2VFC93hwpky9iaqjbb0tByrllJgi2m0uf74mpHcDPqzkI4iR7uLpyqgLwp
ntbEOpfmNV2bIqF5N2WzTyHJONHuXJjb27Kd5T50RVmm6xe8nn+W4p1GvcWHPqjq
Rf8VvSK3G9iOO0FFHRVSvInPqkuUaM1OgXX3Emp5pDHQiSemOgfuY1HHHpQgg0/d
PiBUmaaF4BDEAYXD98c1UMCezQr3aoj8WiVF+5bjOaJBdwAU3LI+rzeIabLnWS3d
dnvHfSH6eROR5ivtIf/fp1S6g9MW0a5xFLRurpNlObVElXtPK5uaWyuLgv5DlRUK
sSjUiUJfkKprIhEVD5dd5Y2DYmO/WwI1v+IRgh4YIEeys69c/7chp/0LMYKU2OEP
strjGFGMxEbMVOFDBGOxuQdq9hds/+cGhdrl3t9VnAOguHaYbe2qQ5y46sR4pI+8
cW8G8dQ3YI3un1tVwYQskm/3w2vZMWiHhrYQO4iII7zomsoLrnNPZGi5vJTs/0iB
gaV4WhLK5f9+k9R812a5TJdM30Dz7+wnlw2KFl2xDobXOIp2et/JuIIXu1pzjh6e
PRDmI+hjVMwdLMfpl3j/vx49vtapPOFE7IjbrvMJKzLVkD+w8D5dQBe85rszFoES
6hYHTn/Wb3jjnlZTsKTK3NNo0G6Bol8KPix/nYjhKCk+ycwHM5s5crkPs//jedhK
80FM69MSnVuz2+QUgd9MYFAyXrFzf3QGFpYVD1wJEPIa1BUS2b8puUM6kJSQ2jYG
n2Fh+JcjJwWGshjw15rOjxkwWKnA9+VhGqyZxhyre4nMn3l0ncV2GIUixtFlt8o3
hbLznGi7VsdKgHahgD/tpQRKBA5RM1MEgm3a378MR9WszaGM1k81F3t8XbjTkr53
L6pC9wSGfc+X7RPpRZUspoUKb4nijZ0D70cf0CM9Brg2+gMV82iHikS3OLMmVpuI
ds3Jo6EeIzWOr0pbKbY4r7yEiFfwXyDmya74OQrpJzetRPZU1OULjpc6uvbzVNGo
48Jb9CUz/1oPKfSWSNQl/7o0+VHnJSUhOGbcc0oauY0V81Y/VT8oOSKgs7nXhw0w
egklD8kKYkUUzQ3aqyi+M5rx45nT2uTOI1QH2rM5siKdGgiRvLgP91NOEB9l3rSI
BH5n1eJe8xM+RMsjJFI1nj8X5zIre5CDAkRyl5rIPVNGjeRBV/fXtjI9JpYZCWbX
L4kW6NmTuGSWQiWFBvifS1rtR7tL4m5Ap+7ngXYfi/bmMUy9K0THQc51maXjE2jp
9JGjQAwcMU5soNh7scSTKZUPcSwBUjWfCNOgXgrqvK60xgkKqwZCGgVbD2UFhMA0
6UVvYxenZvjkff2OyrddulyOLfsyrXkDfHysMEgdkWEPHGdSQjCOgq5pJEMRe4wR
Tz4GviinEQ5CW4EUK70Wx3mhfiBhDYHdCx2cG6sStfXdrTAJzBDog7uTaNkgMHCJ
P75rVFNIG0IizlymhpCPzEqrviof4/sSoCCCzOCdlAG8bWusbQnFLDUs6qv1MtBI
oTskNaRE8JtmIX6wTxxhwBn4tKVQjXVYepIvJLxV56k20KI6P3vKv9KMykG+m9+B
YUs4ZE7e692shlpowrFlQeGyryLSwX52A/kLwMAakKoEpuBcwKnB1jyTWif2VVl3
Ti9QW+BZCYs6PhS8IWJiUHcH7D8C2BKkb20m4ELf3lMwYJY4mq2Z9/UxJOSPQZFN
YYbjsfj3wUajRJ6gITMD84gNxd6p+Eup7ldYwcxwjiOehfinZ+vwavSLP1ERGPnK
ZdhWUBSyQMY2S+d1/WnLDt96tfFeMXgMfK5y7XK4WJ2IuA2D+B7F2ou2UF0Qy4jL
q9Pc+ofRktlcJm1DPMNkO5hujrHBG/CYxM2lfXBdFmzqbm0G5phRhZLSqD1qxNll
kwm/aoufbyenpcov/bmkuOqkVOdqPi9teV3Jt0vkhoxZv5UHzLTi7v0a0QKi2nRd
n0Ycz3PXu/RykLxBtHg30rPffOukvsnP4gvih9VOXbl/itF4tGxHWhXyZlo2pp1Y
YBZR/U3eYVJzG9IYpb3F8rlLHUBYvqaDFMnTlDD5XX9/ayZf/gLVEvPOy8HkeXF/
/W4rN4hdMayy/kZEWwVyWbkzl+XrP4p28NAGdxLjHYDJS7mPFPFXZZvtzFtDXmaV
VlVxJi5bgtRc/VBlIh1vJFTx9jlri8wCJcGcGzZ2llSxwElwKB3sMP5UeBBv3QEL
aXEF0V2+QQr8eNXDqNSnUakTNHF+BPtlaMfjlaCgLFLYn1+OEnmmU5KDCmv4up1N
8ZOfhliJYYPRSF5UeQH08RRUyhvhTyx++Hl8kbNBbKu+4kAR0Ppa8oeCObDonR39
12ByVPz++OTW+ziR42eeBWDB6Xd2bGJS8dCR9w1aeH36peXMekWEzlZWOWC37mJR
/udHhvYGT3nzJihzubOEuGQAHDpwqZ5A3pI31Rt3Fac1xlokEqe16PTwXLrv3Z4b
LpUEA1D5+oMy+0HCEXfXxOApLAojxjTKizWcfLqzAVt3gEO8HcFi59gLfl7Gi4La
rj3JOlAEbjegLK94B3o8OAyfv6N0UPb1XBcZSa4Ile4Un5oiLHaDwPn4klC9BR0/
kHYFpY9OB5vZKw0DQIyRj80237dgIxAJsrTIRT47jShTuUTtlHNWQ4lN2UjNZQJA
knLqTWRkEbWMKIa4od+8Od0SrTvFLzGhZotDlZJcyHDgyDEIi5XubiIWfl7x38e6
LYKS+1d9N445qtwXFk3b7CnwgJECiJA4Ns2s64Bu/w78EicCgP4c+kUMvZmWFMCI
AwpyExVDVb4T/Nb7tBQLwOHe+HRJmBA0r12/2Ormq4G5rLffSmLYnNwb99tDLHtC
JXOkgEN4lccXiwan+NyGQyLiVDSDIFzNQY3i7u6q5MdDM7wcyLHWyQtOpaBXzj5i
5//u4mmV/uBFnr6WqXgGxoQdfPeRIfp56ZRW/g5SH5CSvvV9SBm6SfQKJ8dNwBgg
RpBexBimGawXHbPJth0DO6hQ00PzmTCu9C/SUcIJZPk8szngaV1JfWdROFFZ61zp
u1taxIU4MJFNF+egwNb2/rtHID65LQii0UK0J5LpxGV7YST2pUwoAZvSqSyc8uHo
KPbnfCorejucJdtAm/LOf7T1IFUUHP3ebWdCsLPNqIfmgnDO/WKKVzXZXylCnKjx
Y6nR17vCy2noElvksxFvYNYRT0VGcQhXjMXYDlsrnBBEmYF/ih3X6jfoWx+z22XZ
7VEhWqnIFH5uvhu1RuIszh9LYHe9G6ILJe5bp4DxtMq+hIbkD5UMNUomBQJ+AV7R
Mok3kqfduNADOpZH0/oltTZ/WDC9tirY+QuCcNxCHjHmMg4TVR5Gqam5Wc3h6f/A
DYNwMpMnovovJ3U2UY/C+1I+3GaFd8MTKpU7AoMMCsz8d3udhpTZQX3arPKjE1t/
rXSEOEJHcDifnw1A+E4JKqKD33OsknT64X8b99i6rzOHfCj48suxG/H/i43+/riH
nQqVf53buicoubFF3K118rk4ZEeVWEqqdPmPePzXQAzJIbWPuuUxu3XZ7lFIsnGM
dmFVsDybTwgSl95q7lEQQMa8nDxBPbX9v7CeWzNJ6xfzukwRVhWEyj8ojBo9doxp
OGM2/MtzHOSsH/L9PrJ4K+XR8IdAOsropx2lHvYwkHWf0PDRiodvgMXBAKwwim4Y
F6hDRCxQ4TM+zCQoYsLI9WgUlyWeeLRH1V3pMg8xH8BmY0yA/KnaQmcVzh5ZWw5T
T6W2yl8IVD8F+fCM5oivYg+CEpqHM+O4n73w5jAH3trwmFaDYWYT6vQHoCBc7aU/
eCumtiX1fB5uCChxyKLBkgnwo4TohwUZxJYC7JTOfiai2Wk9AbTdHDmgqabtDFT1
Bx2F+w3KApEeNbGz0puTuHuv2XJ6nG2wRruEFaTgVerix/WNxK1yTO678/EAuO2k
562S2LMnME8texVeVKiXheDVFZD2g4t5/GhGlW4DnyYX8bV8SPuVfRYxbSbskUv9
A/xq0RCLV78roQpFpl51HRacZSrSxN1C8s0CxbmUzU3o9uyHsknBspMMdmuaVQga
c/oYj6EW95K7Ju8roEX0as4bL5bSw9ZWfiCf8AZb/5opRdnuEoM8OHiVjgOt4xpg
SGREwfrN4I6iB4/Gtgfi+tOUIta+R4yqT6qwy1GsbL6bhwqRGMccRhxBZB+IhZMu
7rzr/jmADfgmGkO4QO4Nh9BzE2IyX05WLD7jZ2pmo+nPPCS8izSw8bvnmWIQdV7o
kxGoiiVvJ+uOzkeiXodoZXO2jmaTd/1FM1MmM00l8QjtZqGurlrOXk9fOuQwUYf0
MHXtnvts927yXnLOPwXauqePC7x2RA0JGKonRVg4ti6wbGvZYZ2mcc3LG6N7cgzZ
lJtMpM2SyFEinNgm0Svd8IRFraz7BmlJkXOfIa9ZwgttUU+H4NietHhc2rr/2+R6
B8CbBlSvbEPk5JH7sfTf3lThl2sDsHtZnr61+9pOQQvPWF8RMGbpgvRK8ygO2yeW
0qFbTHzHv1ejsW0SlS7KIyOmKq14Vha76xAkatD8qkWa9emcNyQdgxLiNi+D9Kfc
2nSGbeSdFTavMfqEOkOxTub52qWs5jozOU2ud1U9xb3EHltxPABFHCl8kAaSQ4CR
mG/AcYPcejc/RpBTJeu/InMuPrpWtKGJt3JALZQX6BAdkegF1xWnPV48LNosexAS
joslBaLNUPjq5OaSUsg/Z9oWu1auhZCkvSHKJl+7ZE/8tP8qDZ/Az/xqG1FWD131
gKr2OpQNuO+RHZkBdXImgpfj7AXOa9isv2FFOfarosy8JtZRmFS9GpIbs7cF+dca
p8OK407gYucY17RUgCPxI/lKwbsPQuLcsmaiz7TTUkX/RWAfVtcg1WHLHFOAbVt8
mMzdpEbSPyoZMLUt184pBh9KcqHsmcwbMb48h0LJeYUJWPQELpkcunb4koWlmmBY
uMAgDPXs7lMPfTDH6gwm/t4u3dafX20WQfWk3idW1ijDqosMAdYfCs7yAx/uJhR1
6BRoiZU29owrOofjPgoFDjFSCSJ2SxabrCDijslWTS8oa+zRyJAWE6dAypqkp0Qp
SR6bi4qNFp6CYODpm0fS2L46KNmh5S1qxv4QPnSoItjR1nsXTwcAIzIJb8+Xp7b6
toKfqGqutoHot2P5wL5a4Q3V2Wpi7BGqWCbDzDsMDFKbzjQUuZOpDf95kc51n7Un
NQp8K8SyCgypQeb5zoMWwMX9eWbwoKWsL5zQpWukFBXY9LfGQ5nlaN0bygTIJo0H
QfHSAtedpVxTY8g8dpxiRDC2SfCDZ4X3RY6gw2It5V6A3AVWFwSWIlvTDfF2yc/c
K/l8IUi13PjScnRpOtGenn82l3400SWk2d6uHg0DphffL0/lKR4JGWmauvqZhmmf
k35CitHAakxRWSTiED9aNuSyGiGYMngTpwtCaw1k8zQTbo07QCZZAwFXb+e91WV8
J66TrBHn1IPjlEYsqZjSN1dLymWGKXSQ/eWiP0TNo8beSopwwovq8XMKc2iNk7H6
icpWlUUNJ0yswO53RngHXuDXk1mCtXHek4Qwal8LVqEPMtJh95iGn9gx0pwx5y3A
K53nNzEC26VJpFz4AaTw8f00cDZUCOl1Xe1RyKKU74G/n6zuw6SxtRTqPrkAh/TV
SiRP6C6Mh963Kd7Ix3zxOlqfpevNz3iLGHWgdPkfQSKj4MTYHw6HYq+29j9a0iuB
IdeAZ2uVWa8Q8X6CiAwqPEjvEDJEu7uLRpf6e1nHpFHUQgpuz7loop/sRv7DK+qq
QHwkW9cCc5nNKMkkfLjGLy8nZYFF/OCSWjZmKjPGyGo/gvR0BUCBYdyZejnoMe3C
zgWpvfkFdI6Bh3i38Xp/MNtWyfqwJhSAEB12swTRGB7oCXZIW+2MVgTPlUCLVNl1
MwLSEWCrYt418VZuG2x8uAiU8F8dXn2u4U1fjIQ8i9M5uE1TH/NGbRcZDRYrhEgu
qeNNLhBMXNeFhM8AdWEqu1nA9Ee9ovmBTm9lojsOJ/AncI1ts2MO4IZrzKGOkt15
B0+O/bq+j8gldIaT9HzAJKSc+kXtxKZRBnMwYuF8tlriv3IiBxi9ouVdQT+E4M1W
BnwTsVzA417y7mIusaC3Vk/3x3oSHx0JwGIifXHV2mfCw0+yiFE+NTpkiElyv8f6
NR72o+UtuiOr5H/DJp73av18g9XZA0PPscbL9xkk20QyUJpKnZ6mydHVtds2ExIB
lw1vOoi5GQ0GgIesr64PjS13BV78331ncrEE4UN7+09l+4odgZ8Id3L1Hjh9c5TN
OsQ0CA40KViRtcK8M4OYEj3hA+GXiLFyZZM0f1Oe2cby2o0BUmoxLzAn14U9AGnH
wdPQSyjcjl85D05/4NZL5pxmxdi4x4HdqpIb2m5B4uG3Ypa3KtL+1ViF9kkKPS8j
pZyOaptgswJr1MJCGnDN0OQCbdA4AFfswti+9wSCsKogJ/FMqe5jum+/WJhVt22B
t5M36AYTQa+pzTOnzWHdYscSuwM4b/mTH+sC6Ko4JxsyWyJHw/V9yAUfFvS9S+uy
iBUycLBQkUWH3Mjpa7OelKsF97ER6Vo59DGnAg4KdUdUvNRcsqO77NmNk5BCoOuF
9Cn7jUUrnwa3sjVhg1XBbgz85FjOrzVGDexh+axnmZcCQhs2ufW7D4R+PcF9pxO6
MhXTvpOncTFsY0DFuHeJC0qbMZ/syq3hSkmUCp1M29FVDxpo7JXGDNweyYxI4SxA
mRZsAmpiFJvrrp+cFCVMyGiGfnOtiqsmgKim6ZNNmyB0I1QsSbCtEc7VTU2viNPH
K/YawNuMjFj39PzxsVfJL0DsOKHiZhCt7dZ5003Ml+TAIvg0poyEpqOhsAM/NYRt
NMk6fZHxBynXbVjKT+JvdQcqpb1ezqBAwFo4g7Il0yvkBkhcvrSp866Fw2HDY5Sy
b3Rn9p8g+JPhgJbUIRknxhFsAcyq19jyla/cCdMLgJg3R7+jbug7Quxbjd3E4O8w
TcWNMB6m72YXfVY1U9GaNjWzKOh5nK3VgAMbeV5XpEDmL3xPumWGvUHHb2g2UiPJ
s0eI6mfLwE+7gIukCWvL99ZjCLbExbPbTiJxNKYkTE1TvkiCZnzR4j/BD4UwnnZ8
5yf3CeScy07DhpUCwYxIEizanFyY7Y3GTDldw4asMnWoRN4RwfnL9eQilAlxxwmD
+sc+NmV27CSqwKkkNkMRTKxd0WmVOdUj1YOgosfR2ALl/frpZzPAQbUbecYSTzz3
hloPnNh3PGqGp0MgdKpTGcwC0O6Ev26hQxLkBOonV5QlJZCQtjuimmNAF3MYbY6Q
UXhKLCiROvMDyJfIKkamLzRvcwC2bRCVuUSR3BGdMmUKwGOZPkK/0qGJRMbz5gbQ
ha/54Tz80Q0zxL76GzC1WRN2YU6dGJffCAM7ht8TWVHj6CuXZiERSw74oILrzDKD
IJfzCvwRhBGJDolX9gB/713X+R4LcNTQHb6Vags1oTISf6c8DYPJpnzCkpAuZkla
+K8LoTQucp28uH2hPV7/0HiCfGL8m71VCuc0KF3mUEDCXO0EBSm6nCjTZOAykLrx
CXKdekO4Sv0N6kfpB9XANFf2zKS/jyVE7FK3JN3HLyTjfXBsHFs0wx8bLae+gcQz
fyASE120zLxxHQAPFf/+E+Fee3415QXjNVDJw3ONH6r93po7lwaOsurtLuwTkxyy
7IiAoZLXYd7ykwn+8vWvZsrvHbqoEd2vddIBSvVD+HjCUvZurLFt/glfLP81xgGu
ORZQTSkV+HHdAZxfL4I8h45kdl5QKDBAeUdUEK2kyHS6LCry18ZBxDgms6uz2Eck
HYdAVm7QgWeJCNqhmQM/67vVVnLd4qHNA3/NWpKiJNsBk3bL11BF8iRHVpEsz6Ms
PNx3AVZhUEbqiSJcV66rwaxGa0SZYJ7trOgzapu9vvY+G5DaCrxDqzxa1xSPgSjw
iAGfsq5bGYsOkw9/N+I0Ip1xGqUVkf8U4Z3tBdiq/pX0aEfI83g2Xv/PvWDXDCt3
i20/p/qlNthCf0+nL3tzXwguO9QTlt3CQs0LZkgkoSXo2JnE7rR2x0uGfMmBTuWI
4ddlCgz21LFctOKrjZoGFX9+vkDpbYrMpVvseRXMW3Q8FxCjCnT4kPKmYYnJ2cQV
NFrYR+DTznU6cqE2bQsrwZZzG2qyo4qRCjrwUc8tWftdLeMDhpeJ5JyDq4djYfXz
EOodhOKplVy9HituW04M+ycy7io5eUOECSGObqWuSpv1ch0RWx4zXVk8L4/1/ANp
YqeL+2fENEKsi3W5bylB8zwFIMpoknmQijjLntVe5Q5L7CbxktEr8GjGaDkKH5ul
mtCbR8yfLg4zUsNPY7t2mL9n4ZTZj6N7E000Im5pl3pKodl7yobof4aeqCKawHUy
WFcouk+YObVRyy4imJk6VYPswJ0w8PsDAnMS1RR7JsTpCEui5xYuQPWuHvWYoqcJ
evAk/JIF6TiVvBKtZRMbrKwJGw65vsLUOE0yA8U0g/IlP3RXhvYwnFbH1sp1CObi
wbaC/TjVznCfgA1+8IKxwMB6/XpVdBJak3tShOhTSfT6LSD3HIBOhkVZ1mfx2mAh
7tm26Jji7EnGc4xlcScXtCdB/E1gdQK1TqSLzRarNP/U0Oxx+cMkJ3rkm0DkBj1x
PlsLXOkzddZnNcB2wwoQgcbNmp8cIkVs8uUU2pmwAK4fw3yfBzx5HE7daK4uJK39
gggAhsfyTu2Vv6aiV94xdC6QI7fWHbYG1XjqUyxIQpEbrYfUCcjZygJTUxxqiinE
nzRA+Rkc5CffVYBiS7J+bxCmEO8eNS0GZCNtsHRFwhuPhG3KkcJ68lyycRPXUbcs
E0mbSGUsLZ77Iqg/SVMQS6+zcXZtk6LW9fuK8WgEcYhsuDKZwl8mTpsNufaRr3UC
N/9lAoryOVcm7mrmmZoIzwbXzFJzsVwo1kYnVo0mZIQusZcuXgA8vCHHABIelsp+
tdOaD9MGmVeJHSQC54ghiz02MXxLVxDXKjV6EBvFMpx/w5lY2Q4AxqWjjVFFjG/j
YQdcMNWv/Av1asLVlactesBUMilI6MbuGfV7QTz0FV34+ntBq+hNvxJcvX0+3NwS
sSHL+m5TEadKUrB/ICwuwa1pJRG8hqwSRP6eYUEw390j1usqE1jgjeRAaminUdWn
iALmdECYx5EsFIPkNmj1rjOWnVM4W9TMiB1INiVQHhn/1ADn7PHMlVu1IXN8QGpr
w6MjwaAWJXC/5LzJmXdKPKR27LfiiKu5JakKvk8Wnm/h2MgLDU4591q/Lb6pVacx
zEK2ZH6/2zw4DF+USmEfPzrCetpN0S42zvy8e5MgazQlMZwMfxIkb+lPYKrLxhE+
vV4YaG8FzdzMhY7jZ/FvA769tmiUC9WoNHNBl389khQxPCzbnGxn9uH7nrnIyKus
wXtSgj0mX16ACzoML3b2JQs9MXNecqiR62lX59HF5DQUHwWbef60NTsZOliU9DSf
z6g2iPid2FFwb1GTnmM+PX2A9D6X/ORaZQll/89pBMfoMcf0hFS62e5cpzZZ8Z2O
CUfnl6I82fcXdwsFtfgLTtqEr10Tmpkt9jeQAnuEA499hjjJa76pQl6UMWVXYDXd
1Ou9x2sTOw2vJHo+uEY6GNOcBHrde+kFQXWx807KQ1xasjD53+q8F2zyj3a5+vtW
KQ5elQ3gjYtFt6GxEZPCYy1wCdztyQGxmdKwWMImhgRvXSPT+ZDx05hzZirepmfg
RHeiP4PrykQaBaEGVPOpu3J5vEymSPJfy0ZFzpsfaXktrqjQcn+5giuPZrc/D9Od
2vpA6RAKwM+uDq1qQ0vBBWdOLtwEy5UrEg8J2P8YfCmN/4R5ITrXzFrbnTt2E5bl
JbISohnF4LRwbvDmhgICiqdLJKL5GA1rqY6FffaHg+uPiv4Q1RmmW1Y+cbS/XXzh
Da4e5m59Vkj7ukyMIcm7r4gnwcg8wWw1T9v72kndIqYdz7JKhV2HvZ/1EOduWp2Y
aqOvDljTffiuFfVGGq42eyVxwp/97Ut7eBxvK85mp4B1hHZfioCsouVS/droFkFT
cAoLYF6B/5KGyFJR+rI3KnYhMFhWiLailPkV0hmNUA0S6lzmUaZ0IK/twu+C1d2F
g+l/9DoIUdfl6Q8qDngPqELrWkMDh+5BUhp4/pRKrx8a7pwUSJ1Sud7XMBiTGnK0
FHKipHr7j8qy7lCdgPSkxm0o0fcblovNfrEDypi7sWigxMyp5td2AbZ5YKigX/mq
stD3LYvHZ7oqWfnP8xpNhw/yysrnG+XTwt98aCtyjQiKpW9mRn5K3LsXPDd/FWe1
XAkPTqJLkO8JYNrK5pEs6a5+pfZ+bdpFFcaMUGU7G19XL0sEdavmt7pvSUOyEZBr
0vxk98hFJDPR/9CIYZ4yP16ogBjcpksDO0LfHYShfmj9ClIPvWptyc83ZjOxJS50
8VUVl1vMmGNLZ1xEW2A4lh7iewwaJ4ZA1KJ4uuJ6yRTffxIQiET6gOeKbzPnXCWN
kpO9wERemtZDByeqgJ2WNFIA6rlQTe6lsSBBaGG3wyCOYQ74uFPu5OPO+eTK0XnE
Yom8U6XDbU1BgUX+Df/PXv+v6jXWhQuIWiuMprIUQ1p1lZPzU7xjS6F9rlb8Xgpx
f/UHk1goxO4tubAzjh543zuC4krC6FD1pLzurMjTj9LU8t/xLjNEGHrELLe99aqa
xUIq8JlHAftqmvOcplzi1MEQk6U8uW3NSXkJjTNcWfZidUGOGL8OFH8XjwHm25/T
+ibdMS/i8O2P2nL9FuGwZb4A6vrGWipwWp3l6DdAwilB91HIY5MIeUjgOtnAN21P
8WcSPwkaB6eYY876orB5U5G8XipaGEyLsjz1ywgNaBvQPFjzyXEP0YwW7jEN13hj
lbc1uVM6RgW2Mxef4Oy5C/S6NvijoeHLXpn9loAP5XFWB09TKeyhn2JW5nfyQ/u6
C8fCubEkzX1YGpabdObVZIt9ocSbCwJFoaARD3IRFlRz+D+aYyBRFXhcOfDdzPwM
Jo0a/jF1gtGG900gyeeXJn1sBxRicer7GYTL7mtE0iVZZDOkUfr6pSaVkfGP+qA/
LsosgQytbuzKAEn8B0+Ex+yYXyAJaVqAiXGNCl7JtNx5ThXKfvjrTpQWc04fPRTv
9yJTFW4bIMyoEvX83z2LK7w0pTozToBKAapXkodkUsn5TTkg3dz1tumkUo5/AcTp
MmFz+SdcQsioHmWLSEuHOOPzm0PsisnjwBMneibf2hZTwxZuQ5dFVWUJqJr7YHDc
qs0CP2UWbIBpNcsAUCuOR9MoqoWcbLasUcBbuPzlY2AMENSzga2qY0kggf3j0Apr
DIDJ1tK4Otmcj4Z8IpboFps7KkcJW29MIAq6tskb7gAa8ZgiVdJ/xJInBXOxTEHi
1lOFEF2cEDZg/fQ71Vg5NFxTppWwevEmVX9GaJxl7LjnQe5PCwmFQ0nSbpWDncfj
hf0uABd5JcTpwf8c5m8lAF7wB7ELywZKsoYbBrYbgr1+p+t3zqSJfBECLxKFdUmo
yfVfNxt9iARHA49VKd+3WZZJva9vi2VkTuYsfjZm6uFo8bhuVc7vLjbeC2ZkLrVP
i4QlFJv/YeHtBpUy9FgUQYYC7WlYBCD7ShAWOAqhwQ+jO65m1QhIsLwoAEFAynpA
NtVoXucNVpRfAZORdtRca0y9F1myYBi+ehMe2XbHxjEpl/HBu57420UW+LZ/Jy8l
PRdW1pAai7b63OPgbuK9n+exfRgiBdHo+ITQKk0PES0V1hAiFOPITB15UbHCOL4t
+uOOL+7/7OFYe4tZ87whleqYJ1aLytFgbuPi98QPkiA3ELZEkI2orArfLDX7fFIK
8L6kYVzpsaN7nuE8U5PP/aSlQ3GnuwHWxFhmsNdwe3EQ5Vrn6p818IcQZDGicEU5
s9r5Xz9RcMXZLAYkh45VTKhLYwd3jHje26vXoTgQZk5SnjqIaxBaVpwj2hYbLqY6
WGEatKvFLbMUiXCOHDO0ipe2TDAihtfgrguyjq14MDxuRzWtHDW1ttraE/JiQUx2
7UQAbPJwl13sv0MnyKpKxKCcg7EBOOJ+JaRv6ysZiycW6v3v/CoGMLliI7rbc+Ru
yN2X2Ca0xBrZXmz4VcBXpYYl2uaP2mLf7x+JWCihAcwrCSllICi2NtU09MM/JylQ
W8/42KmPeW2XCb/2hEI+6wA0MmpS4cjLyVds0GFVD7Nfa75HMiMBhnRHceINQ82l
N1wDTmzpgCEcaMNHowPy2LM0cBnkEEzF2k1YO5Adq//6rkl7G/6LnUnCY+7s8UMc
+mGCQbCJ5iQIqvt3gtZPisNn/+aabS1YoN21zaAhHvMWBT6IXfO1AyNpv7oct1/g
8/HkgxEBc/QRwcIJS3TXWNa1r5RfVe1rXiun6ZYEEGq9EvveuYAewUgDNeEJNamt
XNou0gq/nQ2O7MEK1g3Jbz+VqsomPz3pREJ93pVPzS5VCfiAE5+nPqkRWgFIzLhW
8BI5lFvZpLi4JKuWs+D8vp+Vu8c9fR5ABNlFtjVtwRsyjw1IUFeqNqkdJMdflN0e
V2qwjnaEUEnTuzRyV7xTKluoWYvwtQ4bw0wx7rB+ngMyp2oQ5NFDbvKCquFIBVLa
MEF+AED9OWLA6kdRR+g9Hlngqu3sU1XZIvztu4PvswV5Rsqu5DJOkl07fLDDdlJu
iXWwBuBT0d7jPaux4uz0JeXeI1DKKMk+18X/WRH7XQ+fmPzJHP4qcN3SWsEV1tM8
zcAWFXtt2nuuChUiUA1IYXh9FT1KQiWFhkRWsYGkrdLBdO36lkwAHQBwDkhvGyOn
rDO3dUasIcpgBF7SoJq70GZlC/eBJuTWIWEwmgx100wR7xgYOsW0yIcNuXoXR6Xh
aJSPT20c7WOYRHcSIkjznYooHYCIrWLmFQ1AUFpZXC551MQNtN5nqAGQ/lLnBLCw
uUlyjTSN1d9dFaZywb2zn6faxpB2Dx/9WXqymzj84f2ohOOAFAuKsLg5mXz24rEu
p27ilz5/WeI4JHWTrxttFFYmL1QUUK6AUJBARdKTEZ4lzwKXpV+WkBk8iyKkJ+Fd
UqwnqqyZPW2Vh34k+ZAC75OcZ3RxfY4UZE1PN35Y5JnbeS+fLOhSIxgiBVRzmYAM
8wYnxBgB/STrEcUfIpRymt5iCXpcDwWqHeCyPKyDI5pEScRCkD4GFctiWAUeB9uk
GgPmj/4M6Hjx5q7NeUgdqgNZlhrATuMFqCVdGMJu5ohDyhkzZVED3+KlbS8Bdx9l
6UdDnH3k19eiXTbYUD/sxbjOOOKGWAW2yGWXsL4OBiSd+x+HkE7Ancdzhpw8O9L3
kskeRUuCeiVvgDIycawdi5GZsWd5WqRbmH8Ds6u4MYj4JJZfSVVbdAFwzWwdVVUr
hHu4H57/uTvitF/c7E9nlfX3dyGNjDN35hVT51a5f7AatAQFvikpQEf0CE5P8SsJ
5b/emJibGc8B77gQvf17qBM3BY7I6baadaRmbN/s6mwvlhzPOuL9C/UWBGkBpVN5
PnqnHsMxb6pXpVRJko7qGJIJnxR0oKzqG3zpukJUJQaPTS4TgaIcgJdpj2H2hHuf
3zgivZfoODl9Wb5D9pq/x1RRGSir52agRYhOrr8DwVHnJmxbGM/Hd6vecP4zde6z
XOTUoo09psvGS3cZ6K9Y7EwoeYDD1kgcc8QvcpkBXJRwK0XeZkjjY1dNQ5TvI3bc
zR5gB4dCx+BhG52Uw1XJE/vgfMWHdBHyxP2An9PZtyzxPZmUUcH2SBry6DMtHrjo
BYUs9YH6irQXQO5kfYDvLp/o1yHqBhOJvSp8whnGaXJR16KrCKd0U7A9Xpc4B3Nn
t4ahnwFG0StGi0/gdt53yPBlqWkMLdTvwsJXhTMVXrWEHjd/bpKQzyE8tVW6FBSP
BrZZk8efa2JI2fM5UqXO5oYN3DdnUNTScrDVLX+oN2G1Z9aqdNT1lduF/GkJDpxy
sZlEEFblvLUZLPrJxq9Iavng1HeP3q2nTjIH1K3xQ1O7Zv4plpQaUmY9bRsVQ39E
Fb8+gmGLhuMhJvIzhqAgWxK3SG5Okd/WpFG33I2a5QbpDWqFgR4s486pkKrtLbbT
U6FGTvgOzEiHH1gM5Q8WoaZGJYyZV0FM1HLNEacrmb+oL/j+5SEPwQ4KewRnHfkf
MnUpv2M5eVTVWINoGPnOXTceRyvzHEXBZnWW+DApN9ducvWIZT6X4AE/C6APwrrM
Qv2gq/K0he8lp0Er/E8j2sq7O7Ms02J3djUIOt06xmtQ8ftRGHUkODMK86lghekY
pnP/iwP0cHM5V8T1+LxaiHXkVVSIhS69h12Zmk0ZHK2qkkvvhokU9+Sq2mbBvLMz
tSghpTkbQyvqbEls29J5Qu/w7+Fqr1FQngjnvWbWwqshjdxb3h+sP0uoTmyezF99
FJodzN7MiSGxLPdw4kPYORFsk8z8oz1YJvx5fqtmyUsBOaq+c43SXGmh24NsfwkF
MvYXP5Zy7lDg0S1yaHO6z1HUO079CaF88wWZBbp2acn6kvBtZhIlQM6hL+7BSxLr
ukA0ZGO6nfieugcXZF9AXSTxf3brC5/mdUdaiaInRmVYBJpK7Fh7Rj61szgg+CAB
WAcLH+rMTfyk24Vh3W0fUnfRTYyT77IbC+kXknlzBCE1KBOUsPo8PF9/ln5bzXYR
+x58XWMzhDRS+R/RIWrXPVGXWAyNCTwwxbfQmaLrGeYa1yAsVvT04o38/yaeq8d2
I+GyNmFY/NDB3yI6q4S6VzCkIOMqRzhMHK+T+jfCpcB/RKkGcgVhuegm8cfXEMKL
7yPBqW6NNKtWgh645CAaq8Nd2t9vq4ZHO53fq7wu1x968yxYN8jEZICH9HIUk/YR
+gA2YqXLMKMM8ZgpH6ZrUA==
--pragma protect end_data_block
--pragma protect digest_block
hO5d6/TGOVH7sLvWzxOK+n7Io18=
--pragma protect end_digest_block
--pragma protect end_protected
