-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
jspeHaUHyk0py5I2ef0+DH0h4v9R3ptglr5mXs17Yv67C8pzOPnpsEgx4IgC58jh
NrkW+88ewQXmu8DOJ1YHOJLlfyuXfraTEfG0LnStTmwONFy5bpW0SBpn2bAiyM1s
mtvt3Kl1dHenI+PxWpCW0ni8H+s6IwOq+6WgZDn23Cw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7440)
`protect data_block
jWv2Y4aCmsqrz8JoUig+llT9h2IIitPefPzoNOQ1R3acEQn4UsAqb+ksAkSonnEl
YltUMzZkESwa214+zQ7Iv5zYrIJAWBtokEsoM7GMr06vEx9QKW5MheTqZS9f9mJC
4m8II71FCT7XYRKnDtUn7da0UE8IAQEbYXrTTFdmxbfB9Pv8Crkghkqu/iqpttVm
zbC57DleALqJWfkrKDmAe92pk5nmIFfDKkVJVFTg7ZenOSmZOi5BYRGWgvcR9/tl
MpZ2W453pDuxVhfG3D2kSORLGdxhhzGmuaUaTPpbvkbyX6QH/oUgyCh5YoyDRxiL
BU9gz52x6842U/S4Vw4aRyhFa+Uqq+TME41mFUOljXYrgM/Bdp11jfr1NzYNoett
hZguzchi+IIC/4GRv5Dsx/PfhgeD2BKL8Ozp6ALajOt3AizsD5dCAuD3k1mnmAhr
TdOFuxByuZRwfaOoYIwSJ4RdfD46EGbTDMR+yEbO/hgkYUhFCRs2FW3NBFkr/oaA
4WT28dMYzxMajvEA6pnQhJJMmxqwvTTZFPG5XpMe7+m68uQ+e0cZ+223u5eO6r3a
LkVEeTXaMowrr4khWrtYHzScO4UAIqFsE+ZHzhtVPrHJlISvOLVSrKXsNRSJ6tDq
KfFwpYzKAitwCsb3ROI5JOemzwq0qTZ6W/VyT7Cf5ZS6NP5KRV70l9/I/JVhD7r1
4KyoECnft3+GkKP8DfWW3dzP52TVwdRIZp+Ko2mRwPrv2K+2AjtKkkX9zsPABWRf
2GYgWx1FM/tIPtzfcZy4LHgli9xhXm96YtZonn9hryux6FfsDcztDmdiIEbr5b/H
DORKR1qYGx1iCIPuicxztIzXUqklP9bydFtUcSq8kowWbkoLr5nQvP9OOn5SiDpG
fMuvRl2arbtXRWzumAJRIkCicxijMLqLSRKVHixP+T7qwsH5SrtIboeNu6JQxU1K
ITZ8vYYYtZo+YTTh2QzLxb0txIevxKrC/i9vf6tGLt/5ferM+Q+bDVUVnb/QmQQO
fB0zONa6PpUbrLh4mYK/cIXIhwBGdjWirCJMyd2Hgt6NFe5C6N+Ld+jF4WzwRjPy
tdQMa9Ml+jWoD8cYgQHbtLcTRU1fQC9ilVG6DWbmZ62HV08xF9WIkSqxBW+QsBw8
mCXLVk6i+NblXBEsIe6pzVg/w3ao0YEOuJuQ+fTYfTPDBWrEHQ0WlptBrUsJmYi3
A39WRrT2t2bdK7f4hgAjY7Xxtgc+HIIrgSyIw0i9kNAhDTDUNoCZN0awQbnkvfhs
FNkdTFDiWNOtXD8Y6VCAYk6imnIEr506OFkApAGQf4ijWDLl/f6hTPf+PFg0gRsC
XRWFfZUdZX1dtary0/iYKebeuPABvlGD/Y/ZLo6FgI3o0m/ZmWlRWjwjf4XqoiXL
n8SsOi7yT4DXUro4FHfmlLajPXrW2qkXnhlY6KLm/jpxtjRdMluw8Ok0vH81IQC9
PPxBmusIXed3vPR2lJXCvk6a6m6GCgtW9i37aEenJvq12kuLfTs9+P+SxK2Fllti
vYFw3QPiDQzml4QO7kTYEAu99TWZAZ2jshhwqoPLpoiZjEbhk5MpTCNiqhLI5wte
hQFmyZvWlS44A62WomQZ86bLparH1TeLFFYxFEqlMENx1AypHazzYVCTa7y7l+7A
hK3mERoz/q2Th2jLoa6CuZMLBbeS3w5KQ68bFlkaejacIe3eJx47nPS74SmgMJ+8
DSpAUy/r/eJjfb4xXf7IdOREciWVp7mVCu7Unw9MvU5p3SVrQfxxwtf8IZhyLVon
9f+eFShdZEEjkSNoLmPgUaf9UQowYXHjTZCDZHOsV6YOOGD/IBugAX0Usel1HfvA
smhjmfVZTD209HHn67iYax7xJQIZ1LVZNTDqDGnUQFD0i2TiZCxN/tIRd33r+1AK
qlWjeQMGM0sjP5F9dPawp7n7LAQwLaMch1im7WNYIXqkXGXElfIg18xycn8S45ip
eQOESRcI0uQLtxz/+tESxSkfJZtKocpvgTFEjlPYwd0VMo30hN77oP5zXq3Y0TDx
omaNW4x1BmME+LlUxkTrsWNPq3axymj6u4b39c0w3JbakoNN5dgDOOYU2tYqa4h6
zrsvF9oqTJDa/s3hMjw95F7/fjYheoPw8JmMR/QURLEYEUwDmxNNvel2DFtyZfIE
6y1nFOO3GqQe1B6oQdzffsvVUIVst2QkrH/RKLLeDyArKcmds7YREXGHyzr4BWeu
mEqx3S8XOxqlJWXGbWMWzFlta2XFMSOI9ElS/DgCiBPfsM83JRi4fHt50X/HQevZ
Nayxh1iEqAiWbaF4/mHuPhC/81IhwpDnAkELmtYGkSomeMVEU5DjOawQHGp83HXs
F8vk47wGoS57GmL20hmpzK6VYME3wmZY1iQ5h7hIrxm2aAvfVFFjN2bWVfBWAjef
iiqvyEiuwA1WT3BOdORnOyAqzqml5RP2B+VEPCEx7xQ7vaIRaPcb93Nji+AfegRU
VFxGUR+feIFj7eh/CJ5Eb1HXTMbKHMlVhCGtH4Wiho54q+oT/oNfp3YwPk8ZsrJI
ASQ3nfbIC76cp7yakF0AJZ6iqgYGmQ9UxfWuU75COzHHutuJwR7icG5ufPbEk6a7
Fq0lgcUX9wryzHcfkikJ2QF/3j1BlZeeQqMhSLoKiurlzljuaHTu4SQE0LSK5qFN
BI1wExIGx3DjyUGrTox+qgfdgmTVusjBrmKjDlaKLxJIulYwKI2T+vF4WYoVfOeo
gUfCfJpvfncSIZeL/wDo1QG1zSjM7skRp8+58GJneNAO+CCEuwmOyBuCUJdGmN4Y
3E4RKgee3XITAuQzsAxuPWFTmNNLqyfwqysbY4vVbZgza3UmO0sws3tBtL9YhKRc
WPYX9IPFoFQUnKr1uDFLq2vYNoyah/FBXwLzFP9pb+OLMxucj3SRb/R/y/87+RvS
VXcBeTHAuaGucUnO1WsL+TPXhQBI410E/GJ+K8XkIL7QqFZ4g17L8FTsHgKkezkv
xEylMAWSCgo9nuLVB4sYRSf8p6YmWKkdzaYoSIpyiD8w7Y1eG7DIGjZxfwqA01zE
YsdYmfp2PexGXir+mfuO+wtrhPktj4j1IF39PZZi3plrqCTGiWYx9vf1RYeqk/30
ujJVryQy++EZbzdkqdr9LQAq/FI/7+qJ5k17ESA1wo7mEnyZcMGDQjgdXe5TmQH4
xnW/F4U/DtneXRPgOjzwu3wrZQvj4IeNE9ej0LaLmWVCQ4UpctqOXivPD6DFI1n0
RR6M+XGjIoaxIk4qMmNSW6LgcS07xgBgDJWoaXLp99W5edo01RzNvOX9PNVjwB1z
quji7X2UpsC44jdJJ2HpyzA8W/RdQQG+OnPxnNbcPZmgpyquK+UfjwhSOOHR8ttf
LJH6l/oCdkOlBc9wMn2gK/FNrktxkq0Pwt5/y32p/s98QsZyx/vc5lBhI2g0w+ro
SITsBtZr5sv/rfcveq1EYfSJKq2Y48XMegfGpwZr73WK2yZuo/D2MGfadmn6DLfh
J6Lo2ZSAjS8touDToFj6tKY9GoqAXOkC9SSVqwmMHHB7oSaV+ph+juwzEyn8JJVK
Vqdv4zpn8SPuuh6pd/wkWT9kiv1I4mc69+JCi+bSVJ8WtZ5TerwEb6nXnJLILYfL
6JnknULg947gLjDr1mYzY8yk1b/JlfhDcQ4FRd2lnJLdjUgOTA18gqYPTMKeuK7g
AZj61iW+0g9tBhWwx20NN+RT0tNbkLw6m4O2pAXnGYucN1DRnJjWg7+43KlD+rBh
41/CE6G7GmaV4FV1IXpLB9Gu0/xemo6GZuBRKAA4qMHmoorjglYP5JwePHNoD/6T
VR3xZj8txSwTi6w5BToGDLpqn1ZwabirDCRWYgXkfnzm8EjWPsSG5UCPWlM6jv+G
TjF16S8xebwdDed8jCGCLdi9FYzPNWInWKVkpcWrn/Z1OzoTay/cyyop9VLKjUzD
5uUEGBlH4zlLPsTEYXov2A2mPLVYGuIgc4IFI+sNriM5TEUqaVYZvNP5DXY2Z9CG
V2LFxaObNQLTI1svhrxzMMutpYwi2js7bFM9S+Kw0rbEt0saEPlj/hp/9lUdSpmc
1mSFrYLy2iuxuD2t9B7Lj4JNcKeozyuS64+sgsS1+oYw5WmDP3uuq+belr/v7+cx
0iiw5PfjasTrr1i/9hU+9cou7NAIQK8eddB8ya4oMofrKezstbCcYms7zd3hHxaa
hJa5sfND97H7ojJ1T4i3ZI7hfiqG59tnhEh73viwOgW+PpEpaCAZoxzlICayc6Vn
uaQ0ZoKzMOI1XjtgM5mgNhYE5Jpc11rYlRrYcmiNe15lT3EkRT0llOSa8jMoEkRQ
7FwsoAKVoMGP+hzhbfyAFBrxjZhCI+ansBvGAZNos1k7IXkN6GLLHqsX6jCEuOgw
lNV0RNm/1N4zq2L0axeOiV+KuRsWPap51yb8nFpF5ohNi8UOlQilDkHcS3uiNtG4
ccEnk8iwv3ma9Qw7x0DIoEV4GMtfN6Nd6O1353aiGdWb/JOKm19Zhe1hVNV+UAwz
ed4c+st8uyn1WokXGF7AdAioWPIgahNyWvkur2yUYRkl8OYby7s1GT7X/ygSUuno
jyLaZh8Q4Itoz6VOetjB+Pi+cGXd3/VzR6mXxYNMWQwurX2cvZxL0Fhw/3hMhIFy
EvsFvSPQGPrmzQX2+dnElsIqmchIB5kg0HnU6ggtVNespuLrEHe5fulwUwccxLIO
9s/UxZq2XM51Ugm8hD3tR3BH6VgGqjxyZzKu2m9hxqJjsIq2XHOM1zcyA05zemiU
HqPMriON8KCT4xRW9Q2naU+YsD6b89MivyH12zJY4H4fAijCBA296Fw2LFyAP5CS
AUoY8rCxbRZ5z91Hg9Yq7l93OtrbKyJzW3/V+TNmgPX8qdycxZHM69pCCWgAPfuX
8nzGOsuh+tqqQcyaj5oBSWtUNl1OvMOZGs9zj5PBSLiQOS8wvvcBwajIK4QeHMGL
SotA6F+kh99MZF7ILHHudnLbkDVsi5DBorbszFqNpadDcvlqjOPeMbyY15BvgYgR
FuNPTUHxOnq1PPp3CmqaDDKbqe0ZsX4N+3NBchmOz1tRFyF8grDihIgjmDr+YclZ
6rwt0EIP3xfECFgv6ZnnHHRKEaEvCzusPbx/oNMk0cXrVwXF/8x8+46jYczMfdyM
2Rpv1W8nWhseWiYFHIFgfq3NsSytdguyX8l+DF3LGqjINYEarCxUzf9nFwehx8sx
J0cHo9b2eyPoiAOAOjYbiulWcbkZIxEvrs7YmmAMKEr5GiVETQKAq3qp6+9JJUqQ
6RxHK4v/MCVz0mLXhcCOX3tTI/uPhmTKqv9d4pQmBhGjiRtbYIP1bZDwL6zbGY7I
dcQIVhRs5eN3FMnkNiw+Wu1b0/YY7Tsx8AH6qB6jXc5C0fbGrOhaJInK+JZ1ui7T
tfon2R2d37D1aVTo+4gZI+/HXcdCFx8XdhToXJ800QmtWlh6sEe3cEXO3sTCMKxJ
yKZbWXSpgPa5GX4TRzUUaMv4gPWMOHyK/Pm5T9wUp8s/2Hsc51Pg0yTjiMY5ocR7
xnXwSkNW3whnGG6m8tgEQtdSOu2YS0Wb7eSVf7eqLkv9j6lIPQ2BtzRhvxFAl5/9
RpRcg2NS+4emTgNWaDZdC7FoiMIP6ecoHhXylhRGa3FNJTgw1zHeRY4VKEOnCwSR
xFXJCaO85Zg77ZtHVUshbEImqg3aGCVWbfNJW9OtTJ/5clgMdnk2UpJUtnASTXDW
krJ3PMro32oEj9fB5eMAui5OXCRQfKiRywvgotEz454zG25iKTEsgqaV9c7+R+oq
L/9RgnvNF0lJpVGGCwpKS7Hb5xEO25q5l3FjyXP8rsQmBjaW4sZ8l6C0DnctK1YU
m4DWKSrYfjLjDeVZ9aPEy8IEUCf4yG97H/TArm8fTxXU+s4f2JeBlmO0unMpNH7g
NxDqKYyPJQ2WeEx6EbiOMfjgdqZLBY4dGKUd/9LAyFocpEkfS0ON6txzjxsAQDvc
MUINk8xXGPVP0/R8bkVNEez9bcNzx42m9Qat0r/Ipl0RrG7jGLJ+vFXdF/b1Q5zd
vQhJgMUsu/WW9qgypzBjQfBdKNggSH2HyLj5hbtpanaWfgo6EzD3vO1iYtL/fRgh
bRW9FV2fdIghn8IaxPogX2v3tbV9mL5hUH5o3gakTIy1fMwaGyP0sR1hHsFLtsge
nujIVEARdg5pdV1TjS72iTxIA8SUhwnyrM23gr955Yl5OCFI4zXO7km5MEYbniXP
8vgQrlx5xGtLChJ7Wt/QUbmp2UdClNWzR4g9POYWD5o5DNzsMJAyF4XS7DEP4/o2
j0wfTu4bROfIyMriU81aqkBMzc6qheeLznQhXVaeOqOWfRcmMJ0dTE0KmVEE4iwk
qtjf6NAGR5ELPKrnxmm2IZiywVfskeupdh9No3f353NztMA7g31997DZ9J3apxg6
pWwNpxXC8PRZDtAGTLNfUOdsEt+RFwIHBtkWLi7QJ7ckuXA4oYo+L34NbwYXZjMz
MfJTDsf5i7VaVc6PReHh1bDA3fh8k5QXBMWv6QrGxHRZ05j7mkF1yLkJik9afFag
dIYi8zBOmHTFYdv/Y1ohhDhiyY2Gm9728roQf8odKapdKaX7IuPosvMYNwW1km7L
+1QhBzeaDiSU/f81u9WTZX3k5qIKsO7332pPFGqk4Eaod8hhNLDuACgsI8FTxR23
dGzwpd3oR1l/uAziEpy02/ZPxkPOxgCunFUOkRWb2d+XiogFpwYxqy/hxK3DcqV0
N7sJYQjQBCHtQkqfEppEuTbGkBW+s65dlxKKFrIj6kb2LcG+bJWdX/hvT2uEeBm8
1VuS0DP6wufm/WrpOEun2BcjeTd4zHMnM/WmOMgv0secfuAr7BvdiEaR/YYeQy0Q
BbJk+/6N4j9WpTHIdEGuW5iuVpGlfu/uqksw/Qg7pjajyKJ82ZvjlxFS1krkuYUQ
jSTrgdTaZYI8M0KRPAvKAH5krJHp/f1Dy9JMohWLtnu0J3ocsIES+dQ77oqebFJG
CUF4/Otp+u8RKrcufHHKP/AkB0VSuQeDrkboF5KNxt2xuwNeFTl+nn9D6WiFAc0v
mC6GG+JtjdyAEybIoK/2KPr8RfczTJNENMUsYbAHpqsG5Yx4gzApaf1yKNxk5ayi
RVlqwk4BeR5eIY1S2d9IFRVbhEQBiD/EXkfSSDxpYaJWqWeypyauQYzGD5lV9Qqn
LI9eUDYRwe1nYXH760OF6PjlNc2Iz6F1OwuSSo77nCgqWXKtj0zWMYdC5Xg9T/FE
P/mzxlxm5qVBdPmu9jqPej+TIRIhB5GWc4w4KpXQ9hsAdhdBIKTpJt9iLECVmWKg
BMtU2Z7JeCQDp4HNExQ2e+DeuE74j5W+YozpGAplP67GO0RBzeZFIEfmFRu5HWNg
ey72M0KXaFbgfq8RmiP/6nm3MK/dncUkVkEFO3TArf96rfOnAvmwBJfb7MDyhElA
Updzae+N5lq0+8yA7C4uofxcs6HHQBIxtddOiHjNS/ki7IcXxuh5PFFbX6J6bOzD
s/QVPBCvUKj4z6RP46MAfuBUSXz9XUMSi0qAWAAH8VA1CzxHEZOSCcgJIQBkf14/
sMV2m7pu9U+Hql9bugz+l8VEoFzcW788LPee0D7ZxE0L6WnYZjp3wRz3USweuWVY
J93A8rpXvJRZ6uQFmFSr6a6jaa3bh6AwMoGqPbX8eOQsRgwBXD/tPPnqM/0q0Cig
0SD0MOFoMcUajKy1OdU9lVkIVNI3OLLHOYYoGS5DuOTjcEKiD1LsYKLL+BCnUzFR
c7qPmjrgLpmh3Xu/7kVjaGmclWF3G7FVYdASZeWaf8fXKi29Uc6Qpzrbj+x8C634
Janl6K2n/koPnFkntJWvHfRAjZn8ZijkGsiwQ7M/ReRIlge7PQRwuqeioPcrxn+n
GGHtk0cob8BESRgln5vWnKZFSKCW46IZo7DOz2G9jSocZmRimEEc2c4nUIOtqVZm
wvgD1mpPj+ZxCOwEDtwZoHyrJn+frU3kOurYS7qp7leYrj9f+E5ftodmQN3V+/Tt
nrf2E5RIeY8qykZ/usUtCWhwaoaBw2lTM1IcVcWoRNo3ZrOURUJ8QH7qMqOPAEu0
3rLMDGfjLIPkIiofWTrLqtMHU9JF/8QBHMPntZpfplr1Dj19f11HpgUDgvr8jlPw
P3YXIUz2URu/EhStrZ5x+nACOUIM5KHr9OZYTx/8CqmcdNe3UiVpd1/HVidRggAa
k92n/gSnbflx/QvxyEKweGkx/ssVxqyhhg2paCVdExG+w841+62/43/fePTnvtzx
4WDezM/pNUqReVEfWgHh1HwlK3y7tz/xyyj5x9csMV4fatozoLmLj/psywuyeNUI
EwqlKy6QuvptUeo2m44oR/uahHa4NqeuSBfz9WfiEw1b0TVaZy4IHsyLQ1GuYZeG
x38hbdgLdGL/y7GaSJakeDV6EHNtP3juUN2KueY6LZjPMT3cKKdTgnLhC9FrarhZ
Oqzy+rlQGQBGgmdgGMH9+RNSlAoRguWDwNE4Wv5nIfmK6v7lGvt4RjJIYrRgHTZ9
L3MZsxckUNL53+emc6bSCR/1c291AuoLb2KEaLBq6ozra1ELnkptZuNCvULW86UD
kSTO/aHvBT8BOXmBk5DD8o4WhRC5otRlseAV/x/ecsWg2TDzf7s3B+XdYJlRToxp
w+cpDwm8J3ESYiWB/SLpUHXwODMR9499rkjK4EIS1/EvxXlRM0Em6KvcVJY2aEqb
vVewOd79z6aXCOBXPWsf6RbiETWBlRrFXiZI4DlrhDH9zWATmYR0B4r7pLMO4IsR
gjy2gGkr0Tjf28NUEfDvZqCpqZSvyw2RBSqDVXeHo+TkUrDvr2vLfsNdXZoN9e9H
Kgn7nsizq8tbSWVb3JCO6sGWNYKNT3ehdzZcYyfR6Zz0zD4vsTkiNjWc4v/w+uHI
oABZHgo1GKMbOs9Gq88M4qXeEGyony6EY69YZ64BtcqJ7oye1X0tKmzawe80pqkl
l/TIumqDfQRAotd7DIV4uVCubmuiekzQFMQKCs791GzE9SDChpt5UZY8o69+U0lc
oBMWPXISVdUkJmhB8daLDEFDDvS+bAVDaN71bTQeKn5ThD4wj1R7F8fFf0mpk86x
L3LCDuhdwkzbEX/ovkzFq1AM3swzBptlSjzDbSsxquuXnNwKuKEr+F3NJcPy5RdT
zZvJi34dpT8W6jmDeG0k+SnRc/YpScKSbsVGyqmhhvHo9kl+geW44U0Wx9je/tLE
Mh2REApFYuzrbHCk1wz2c7i9YyfnN9gvnl1J0AFCblIfoieXD53KwB5iEQlFQvnE
8jLoee4Bs+ftAIJ5vHU8cOYapAo82rhHct0fcwNOUWqt3EAlq6YuPWFoSKiN1ZwW
aBZ1xZobhGJsjxf8LRtdoSJFPRDiFQqBzqEyztpXOXTysimXnUBgFiFfTiznR+K8
fm/aC5tq87aoaPOSjlL409pxvs35Yldx+PfINpf80xPcYxYisHL5f16o2KbX/cR3
Vd5c+jL2nGagEnP6KewmVbbcJ+Tzns0swicglltPnwfoVj3XUAAXf+5R4pg6qCVN
vSFkWdr2hxdoMdJE3RgyXYkrzLv3A+n+QK8ZI8s8zRwDNb3sJvh6WqMmAariva2W
SmDjNiIzCwQ73gAVbiLXHse4mga7F507u1TcufN3KP8SOCB/KOESszVjUpVGt0OG
wtyUFS0q1yfEPX2ISu7eAzVBYrr3WE6iim/1AMQyc8GXNNMHne5B0iudJgQKD3xC
ZnapshBzLTT+SWXYU0+F/CftmDg8F0as6b1RPG6bUjLIymZzo/jWgZ+jCtK0gX6Y
QgdVkkD7dTl1Jda0HF6DQQ4wdwbG+OC+pMrdn0sNYAT+uiBIp31II4A83vCFFH6m
`protect end_protected
