-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Tvsohr9H/poBtwR01vYmH5rsZm23Kf6aSxga643dDgeFTBPNSBKpyIdCCknWB2Jy
ln7IlzHiAUhQ26dLZICWupSjAUYPedJO8AHKrgbKrqqU2cevGFU8AQn4rK0HCOVj
bOE8LqRrdanVLPVtFKMZSm3zaIaebgApeNeYw5y20Io=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 20256)
`protect data_block
C8/l7oi4d6msOEuwRf8fvL99fz/HYvMw5S/Qm1O1eFwxjC3jiIONfG+Ys6UyVMIH
Jz4HUdzGGZaMV07BAJ1ZgtKp8I/4APqIj/P3yh3Bf1/MV/O9/tJCBhLiYSDKtCkC
o44OhWPyCb/979gxFQPscLVTK3DX4l/i8Q8kinSo4itcBHSJwHFIij6gzGjwRpxT
2/ebGaf8nqi5V1iqvVk9F2HyocBNaF9+L9vaulCZOp8KYtMDOIu2FlGdiLrQsD4Z
lRH9h86T/oZZB5PiAz0ZVBVPYcWi9eVCfic8LppMfiXgQbZx5DBxS2h7BK6R9Wdo
8mUcP+XoxVf+/mbAJrZgh9xNVp0DsEq5saOj25Fe3F4ViOkgAbXEwutb6YLdjU9e
l0zOczirp40hSIvq2cGbIlFQORgbNAtPXQVqxTQ3GJT2YGd9th3Sx8rbLszdh7Y1
EqI0TRhQfn7Qywcrz61K5PbsqI4fvYyKX60LZQ3JThfMd2ii+10OuGeqU0TkjqzK
A2M0/mZPaYx+PAczpbCsOqCJckFeWqs0os1heiEB61Iox+S851vUOoZQ9n9e2QtR
a2fS+iLNGtSdUzxOA7SU8bNVR3/q8SNvHmgdKamjctz6fUnUe49wHCp125WeO39D
60h4jrWrp9QbVXeLiDC/5+bpmgqDns4rTEnIOl9XiK6/fiebBKKD6hxrgwJV7RNS
8PjrVRxAkIdr3wP1CIlxiy2h6rHnWtWsj4pQV98syjN58mHFxl0jU1yFY/NOp54w
QN8uSdXw+tKYEqtml8fHDiSKVA9XVMAx1Y9wM7eW0B2FZXhkFqQAsv7ymNGXIIxt
2KToAuS2f9tJfdFSF/GoUux6YACcxkm97xN1P/7Y86C+JzI/fu6tE4DC/6gUGvGY
dN/OGJgs6Lr1hn4031VzvCGv+qi5yWKp7pEmy0tstc+BVD151sZlw0KNnoAO9Dc9
WfVQkp3BRUyz/kU+feEyxrP3yeg3zmmfSmqVld4D7YJA6hF6shjSDpxwCfQHDSHw
EfemXQjYd8BYxbg7taMHHHeHHo9dL8RtEGncUoQcu0RlFw1X+tpXGITYlU1Xv1TN
G+V3GuQIzeE+n07C8lprYI5bUEVGeNuLTcP+Dp3xCpexu4wtzS2gr+1i5cpLrVkQ
CPnni2av7auU9kB/2sn8wo9nWFAx1pGRgc+00enQKMJADq2NWyaXz0rsg6GQl/sC
4j29so9nJx6UqRGMPMRpWjKEZIuBDTHL1FAh5h7ZbZzOVRyLL1EpRdAQ3+7GULep
H0cygHgz6OV67EKrB5LgVBchU8Brba0neyxcrMzhMGj4NqT0DnAejEUgDC2QDAh1
Z0GaYBhvMdNzi33FGH1xvClHY1uFZ4cK7IVKvtQJXIzrwIfYAlmPwRphSkmDWhVF
sAtuFQm0xb0fgGeVXu4c5uea6VI8YVuQoPQIU5TYVYt4eXK/rJotmVlSgK5fwsrd
8MAOUrx+ZMHHc4kYc+ONd9D0ofor+egBHvSGyKgRpGs1uns/sRT1o5DDVt4lJZUs
EQk9Ij1D8yr6xBK3mvSibEVaexji3cct3ZIg3dAKIXko11fjEIBg8K2wc5V19vww
yOu3kOlMPIqFfo3LhdcQUJCG/vI8j68nvncEE70KbCCD4lUy2aiQRiTTtIuOVwVt
OS1u3fgD6+dB4fnBMfmeqyYw3FMdXSL7A2/HwwlD56BcGph4N+WOnoBsNSIXL4/+
AmrBge/d2PWGElWjXoNxUdHg9r16y6dU9zx1xbW/LO9uusaaUY9D4YVdA4rXAzSD
pZHTzVmF7ruN4JrRDfCl99tDYamd3N5bIAV9HIcV/hrfdU1Sc3LnouVNtXR0HL9Y
eN+CI5fBMB1qZ/y9UBQ2CJsQ0el9tiRvRC/23LQ51iGoyoWbhnX6UC8OwpyNebTm
9jO8GoZo5tTJjlxp+zfh73c3kU8kr4Ll+IPTTRWSeULGGt86fDuPeL9hIBYsj6iE
VTCYY3UQ5AMHyNaevihV+lUw8hSImE/SmHXzj5DP8pFSE68bI5hU9oSHdeTth4gM
so6pU0a4cFivh/2C9FnU+1JdZ4ldZ8CZQteW40gTdXg4VCOQoxMuPRoWG5Zo4B1n
u6dcO4nvC7tN2AwFywREPuDjk0PFfSAewVupO+c8NjGhDYE1jGdQar9RsITkXUGQ
wmMv02XwPpsI09YdhpR2aIsCgl71ZJwI/wyvr2OQfGc5pb+nqsyJsOibvp34TU4z
CDNdwS86VuE3I8DgUVMrBNlpiZROcBD+l8vNTmV946fUt+qP7mZrisX6oYl+5vC/
Os39Zkx+oFEX1aBso7P+6ojyPMQNvVjf7r9D/4q//0712l+yMX/PboIjvfSKdCJD
Plsdm7vHbMthkS6d3EzobCD8Oy0mzHtzmUkQQ31CUSJ9qnXJ8/NfNryJI2BYYh4g
eu14Fnd9VlGqRQJF89e1Mci/PtuSM10X9IHKyUnl0+J4ySU9EhOGN7QFx8plRHP/
3Le+q0n7PdUA1w4CiQFaxIh7SssMA5SWrLM/1nS6PnitJh6X66VhHU6sDMByTWWi
smN21PKQJWSdjItkfrbPledeRhO6izdFcNI4yOP/ZEBtvXZahby8E7XjV8JHukGH
OMz2x27vHC13tAwp9HDL/GXEGx4o0G9erM4mAkEwXiQehsLDqPjZCZQV6X0I0FjO
Xc+pnwf63Ifxf1yIMtIHBm75FdTnE6qehnkP+kZPxAsaQREH5p2cSj8Jxuzu8q5v
mFQ30NQNpRyXhuSDXPvlRwfYWZ2O8qC6pFUculmsnAmWdYaRj2ZsIVJ3LPGUlOlp
XaTV62Rf8qYBIjh+sq2BgrcLh7bpmYok2gFnPgQupa3PpXL/vyv0uAlOowXWuN02
xcYD/f9hLGizQuTVIVA7ZmFgTmCfYIq07YWk778J0k4Mv114H4WQdx80Ct6pi09E
ib69xEjqXbA0ZIT6B6Gagp1baOVlZIHBG7D4dPPMvBOie27R5ZPM09iYeD4ghIcD
WcxGV9GB1xOBqpK6SYX0T4kzCuZL95LFy/TttF5EQa6XwnJ0IhZEYmaRgWTnE/ko
1b5pB3UWwTBS2i48xGTnuVWhNjq2tQIeoU4m6TjMjAm5pxx4k78IY0Fi70BaEhw9
5JDJ6ZwbCWYwCD8DRPERaF6k6bTv0YrMo/stnA1BeAeaZHvdNibDZ4Cmxqn14D8i
+ZI1aqnyxOsyLiYV4mHDNNgaWwfWfLDR2INGqskfCc5eWIvrMN5fw1sedXFH7JKI
MYlW+JJ3pSDNxJbnh8Ov7ieW6SICUiBhR3HUzGYB1zF7Kkg2My7MmBatnfWQaN4T
0NxxlnzA4lS7NxgMeEyFPIBnJeImSXpGRERo1Mazgr2y9fFGF9lOmcWk0AAyRECw
xihHvULflaGw4321cm5kMYhi+52cA4v2Et7f2svunhbtzkZtswgFbiLZmPK0Ju1N
I0O+quMcEpYcz/vSM1yuIJMI33GXB4zzNWW7+S+u7KXAoS3WSglsJjeY/fCVs2XG
rzexLUmcDIIkBK46HllSgLLOIcrFuhX7HIplrqJkoVCB0nVbKiQfirQFRireAJjR
1CO3Mtml3POIYZSn2y+3WX3xV0oZbv4BxRaMGtgSoW6qJEdsbSHcAGhRvK4RpAY7
ZmCtTZCcJIzWLJKFPMolmrTtd4XIDY5OO7KMKt9kDBouJ8X01x8A8LYd9Wu5+xpF
u+0D4I6nfD10Iz+CKYuRX2xu/MGhIeiZyhTgZP8HKAOeIzSO3YH3fo64590npxl4
Pd0UJFj/HsxxRnqfRzzgJau3Qhsg/DsRcAmfcUMDlrUBY6PNRdiOqlOMnRbavZpt
CGfzdOa6WmkYAiX4Ar2HJhdBoTg7loUdUuXIoXFthYYELTpGhimAhqfJsz6cT3kF
WVc6VqMIZaD9Efc38jc+CnpY1u9pmDHrmfHSVAL6JfRSq0eOyMBSDGrcSKKuzONO
2DJJgPaApd8KeyRAFE015Kjef2wEB80y9S9tIR0XcMUwXk75pCAnknliJKZvGHH4
fsZT3NwaDwLiwCeb1Mwj3R6mJioXHyQpdwYQX3vB0jK8hyAXHCybPpNz2I2XqShz
ZZsd1ilfd0jV9Eg53jYC5tcBvxT2+Ma51llJsTRwICmpYYre8tVqewifZJcJPfsM
HQYw6NPttbTAeQG6PM6tZ4Lydit7eIB5p/rbjDuKnq59LOfegvq3W5qvfbROhJ9K
2RIVi+b2S3DAVCDWjwJUqaBliamHwWrZE6/X0kBCfaHTWAoq5V9jSDs8uETRzIX5
L1SATEEMmwiOu/LcJuCCMvEGHGLAyTN1FpAoCpn2RsTcB8EFCTs3+5eskIPMbP4o
VsBWOvQUw6oSUdEFBzl/aKMseenG4uptKTGWSZ/kRCC/DyFAvupx3zjwVgc01zv2
FCEbYdc78E6JqZeMcH5c8L245MPUIhR2EtPkV6/J22wAjlnRMNACHoUEkF6nreK2
ELZSVHBosSOir3xR3ZDzGdQJ3JMduukexRUiELF65BdaV+gjxNHHk1Zx3JWZMPFB
QxyszOtarAfN/f8uXKxwfMUwXOBjmIXyXmB5Q34HoXaza6KnVm3GLX3T0LDklyvf
ZTzekib+YOgwvSwcp+Jfj3CFIlAKtuEupO8LZmfSUWqpLjBbpwMVj7E1vtVVha4i
LSAz3LLvbwPyxykFzcsVflxciDQeNopkZbsw09nP9l1INx1VAQnvQMY7cEUVP4mK
heirYuyWKOt2HTTxE+m/HjbOiMa/8747vRWmi4setnKAVdX1clFlyA6xwRXZMaap
diE1REgsgt0IIvm7gQSmxq/QWtnzK0Z48fj16CqCK4qluGg2wwH2D2CQDd7nJPoX
EpakvCPdwutZfG6/xusqboorUoGXSxQzHDjCV/G7M81ug+hpfUftnNzV3TYxYC3X
7f5XWZFqZgkB0OvTag2l2suCWygw/EBrPuoXqWHbmthHtoyQolEECif9cJVSUXT1
piogTQNi4aikfwaoNzouUpct9MOdXrAf/K+Guk4gzi9gETDSRR8s7eXhFHxsSZFR
5wdg2wnQWm5Tm3X+cp84G3wcwxF67Lggb3qYnsDlP7JGKPHMFe3eJ+n2imvLEGAv
jtoZPxIF3up0Bx8zGTNZAWSeD5PygD2dUio9fKkFeiDgkTzguokch3yVIzwIVo60
Hfy+PV5jpb89Gru4Zwx7MAV3DpQi/Al10DS643TS1fVP0MRVLxjZLROPiyiJ4vqM
FcAkOH1CZ8Fxbmg0jRbYUlzOPqt6ibjrwzmppXSRPuW3xQCTJYzsL3oTtbS03q8n
QqC5s6fMXR2c4lUPLuFF5TTZvFbbje5ekodpMhtctZffZxhAXN8i7vlhM21QsjOR
ERFL+5JsQ12Q5aNZ2hsvkSuQmiSxNDTSLEgJEf5KVi0HSbeyQXgFDt1FViWML/LO
MW+9tTnNbkurMGxu/7JCZmNYN6uy16Yp7eXMuzEZaJoviGEwFywR8/CYqvh/2XjZ
xnvH+5YOGpaaDxpDYetnFSQBLKm1gAuaHQMAdyFf2nEU8YipBMQhRLmtQsoY18MB
+XidT+5OQfdkep4c+NUakR8qDL511oQknAJcYhncHxTOwvtzPj7JgJyOL6NhS8qo
yJMHhwVPsK31wH2QX3khS0OkSl/+0tL4WBgY7wdU4tQ0b6N6yv45LrzD+JPHbP1+
ul//Dogz/KCRUP15ilMKnq9Qr22KalybQN+GCu4n5ixcxEPwv/ikoorDbktolDtu
VXzLsOD5PHELQcaY4BRmM/vua1lCEBCXgJxwZ+so5xF+xlRNQmHZ+qFNnb3k2r72
vnj8fI3ojf0laEPdCr1bsBHPqOhviKjTeoie0zMbSa6VkWP5aX75/rgrlsC4+yJ/
7KmWkoQFEzM0DQl68JvtO852UK28H+9sHHiOr/n/MWdYrRqwY/DzuPkKKJio3ESk
/La9LrFWgf0QDiDVrjHVQ9rn/R1cBe56KOjxSrNEfi/SQ6xCXqtC+oGU3/SsGPOW
KAxcnk/ToUXqEOFoq8MRK1YZbd44yuXldcLRLpS7wev0MAH1jZIJ77zKDBA0YoTX
14jdYR4sBOZmUIrFhiQW4GRT2/7xYwZmTSshHV0bylQd/Il87elIVokT6EqZRqUo
idn9wFK1NmxJyzJLr6Ph6ElPOeFnCmMmIJPqxORfRoCVFT159d//n1sheM44NX/Z
IHGv4cc3uCgo190Ve02espGYkkPtIidDYl2QiZfI9GbEBlQ57UnwS1c6sYffbr3A
7iABXvT5XSSnhBEDF+iKm6Dz6wWexDvWF4Cc257r6F0rFw/Sode3qXxtT2e0b4s9
HfV1pBaHJErcfLkbLKaxUk9p+gJb9Tzc3rGchraTH9KSpXUEnBhrh3PS6PYigmmj
gkwCMj5vUL623XK/eR1sqUFykS/ZRacIp+fFhwOjlVtYCFPIdwloC5QlLD5rnzFG
2bpNIX/XpIzNjDJefmWZB9w4q4XXV6iGO//BLX0j11RfbhiplANiS0BR8uB5afMn
XEjPNn6nKxLtwjLccLjX6nx6aaVRd5h+UdMgl0FmVrF0o88VIchG0Hj3sy43jtlq
du1NI7GXKN6yC4uL1sEjAoTmU/1ek79P8PRyS73NdBv4LRHQnE2KiLSO9gvgk9m/
E2tk1QnMIaO2QGNulzCZKLrFSfYwAu0U16TilQOAEetiM4gcu6xrkpVob71z1ChM
+i5v3vP5bs7ZJDoAK5IvNN/Cszr8jc5mUaeWgoqbE2MRqLs8oT8lB1W/2c7aUj9F
lzunokMTtwiPzBNEL+Rl8cBDQdoG+sDhU6H4bn9Qkv3yYUDDI425ZlDdNffxruUN
GTx0wAD0/7NopkQDP20G1ajIxTuNAJbg7hpx8RQ48evySCiPAPYHs+7+nqyqnGgx
1RZAjjZR668aTWBROOPthZ7J2XGuOkmVw1LqdcQktjrcwDbpviM20ZiSwmmtMM9I
dQWui3tr7wSaS2qE+vFMmMxx4rO69a4iXfunLTWRL+Erm5FCbBZQC/JNjMOqZBYZ
cAGHfrZaO66g1mVoc1p2d+OUmuWKDyLoEcbJDPVEnt6/A9D3Ey5K8B0RLRfH3LxG
VKziyvIhAY1+ZR3s6pQxTMPc9mM8xrxBrF5P0IJguNTX3zT3RGXRLj+q13RTqkLo
wuv0ZL7s1eoUc8kltsMf8wYo9pbW8Bx6ENyYG8zA3gdPgsWY0YGlu0j6ZylE0ZAU
9cT58SS2gZlGmGhLhupFm8v6RTf0hc3P/I0Ho8RhB8Jh7WXI7mhBln69qHlsu46t
o/oXVBJwHsCWtUpGzim+Qj5eYmX2dsW8+HMVi3/Lq5Bh1t/XYZKPaAB7TEEeHCo+
0rMY6HdCI+FJ9eEoEkZfnOHvWEPaG4fGE/XipxHoz0NNftkjCUU8Trk2stClkFjk
MZ3k+y/RwnGCY9mF7lqBplK00OwFH0zBzK+pPuJEJv5y2fSqHO/ddza6eSqEYzxo
cdOcm0IXHFfbic1AWChiQ+aaBgh0RArqasows+K6Y3aVOHoOZZF7Xw66afZOL7Bf
qnm8yXXIDSUgQsLeSmzQ7QZ5kC9drhEUxLCodq6g5ptBXSB74hSCraU9gCqdQWnj
2pwe2mqNNpqoZ4U1LTl+YS7pRA0WkGAGINvisVIixcxcgEyvJZMSAbeT7jNnABN8
jdd/uVWGpa6auCNsKBYxcmKt8xI3DAGCSE3lIJ+nuVBqGuX/RqdmX8R1sQJ/tvp8
tboyZQ9kDPuinMD3j9S5u/6WIkMcpwkFkzYJ4kPwEUrCk0HtxApK1KKX+SpvC0u4
Jz3PBqMgwQt8CL55zUfA7Np1uAB32Yzcb3/GFjFx+K6DRO3DdC8ZoDFjUAsLGENj
XlYKHWOzKz0wyBMi/mophHm5btv+KFcUdUkIASSnHGRrOoAq89n5jotDjjsA4ppM
/tNz761S0cd8tQU8i8vjYyUYPMtObXhsMOzxQxk7IgiHendWaCfkgXv+ye/JXqOF
d0HNmaBFRf4WL4Ij1M9BRsF3vDqLQx80KtFzVu0sKCJvIdmyLb51PB/BWf0j6JB2
P0FUwoCIV5CTHEUYq1/Szs8vNdoSi5lIn48VVjm9kShGiJtueaCRooSl8BFdGrCB
Es2RSvk/LAnD3ilSVlrxsg39h+fmjQiFKbp++CZGGmXblTI2tNvs5I0IoXsxftyi
jRF62xVXcx0P0dYvRP1VszGTiY4v7mmVo+rDzzGRe+u9SwZCISMij/L1IYPzXY/o
CQ+8PukzYELJE2Wf57YxG2rloz1NzH+01gBsNtWTdl76A7jTnP1NiZ2n97F3eN82
jcrVcb4JLKW+uGm5BBDHWXv9t+ATi56Y+oMpU3pZmYAxIJbdPOhpYotLQFV2BJqK
WmbfXm+p6GDU7zr+2zMLYZ+9oCR3t7QhuJCaepm3V/QoO12oAn9/F8gfLmUi1MV8
cFE2Df10q4oOq3SO/AsnaErsfDPe+iCgUiXeWtIzOwqJD+M5u1g2WbCmrxhMecqK
CFXTXrnBPTqoWqbhjUohC5wB8Dju3daDiChgTcoy5h3VmgrjNhTJl2xv2qIB6/6l
i6JeIiQaz7B/mF8AQ5OJ7iTRx+aH66tKQGwLaDdGod4y4OTqCjhjMz4aoCs4Y5MD
r+pi2FVfsIjX0ZDjM+0WLCPzQm/5dsIQckr0vNAOhtXI13Re0Zh908HzIljAuAyc
7Gdot+cKhNtuMUZzSCqSKrfQ9BzRQcgOhDTtHDlihwx+oFJrCgXj4SS3bWu9RYck
jZiH+D3hAVgHNhYNE8rLdPbHHXV+dTWMcSuEop8YxPv4BtgPJuBzJL397wNMJlLc
SLlkT3fBs0MTzsGP6aK7rFGLyGYDYBjqTW5G5870GzTOrJuZyhh/5a3+0ktIEjVn
OPdPgg52axXYnpJDXeHV2ojYn0Etx29ngAuNtFqY3ME/nxOpuuMJa+PDVc7FsasV
KJhx5dS9uZYL07uICAiSybl0KMD7aNVDKapOl1mvoYhLSVkhITreH31o+nSJPk3L
v653gOB8x5Ih3ID56L6CvANs4F69OCOR7Ybx7d/vrt4YStKPWm0ys/sQcrM8q/K1
qmc0GyLfUNgR6xDXcL7zXt6USZjydPWnhic8pxuw1TKTtgbVZRIm51tnPNunJMw7
xliRv2ySe2lF/DwD0tfQHITZb1eZd/qLteTLykBUxK9LSwH0wTVMF3f87+S0UOxW
GPtErFHwCDP8tX/TOrTk8TPg66KaS13G9UuvyazO45qF+HjKbNVVkoorj273kNlv
TYu3QwlQ7AoU5GtKoDy/+4tEUFx7e4c/OPXevA6BferElejv45EwAIiVbLuSJzUz
MO7put9Ox2MrpQicTaagid9faWdqMdJ68zmSYdj/v0g7OZWpmrlodGN6MQIq/zKx
xlOC+YHa8tHxJ/dMg4AFw8rHOgAfge9N5rHgqNf1Q5mcYfQVNgN5RRESJKIfgCYv
YgeZwav0ql7HlFnrplrzMEFlnLbDVqE9bf/3MfzgOnbyrmfNHP/sRKZDctgWNwnU
/knTBTB4LxaeQyIZo17ixKIVNKKcY2Sol2vGw2Inxup9jYjKSgCCASvLBDmGVJ29
pVkM2CwmcF9OXovM59nzRm9lEEKsSaUljKT82k3MOaqFO3gymp4EAHDxjXL+zr4z
dx7ALRJG/EfG6eTAxYj7AcXDUMZG9aIRxrZ5CF6zvWnNN6vfNOHfq1d58WBIWHUB
W4hjYfNr2hqhlhbwLUtcdqJY4k7cCPA4wc1IuKUsfCsr8QZzrnRAGCrZzOvJtYMT
trF2pbGq3V4MpnEopp/ZfcntUnLCLrwH0mdTTaF50zOp1nXLtNlnJ4M/qQEE3X/E
bFTKB7y50E8/Uw7mc4XRJoMdng/ZSVWAVQKvmHwQ604kl9PWWJIoPGMsiFd4gT0W
cIlGs86VEUap+2wnBp48bsAwDLBXDLHrbSspKH9J6n8cSebjwFD3XUF0A2b8LHfP
c1uViqsrfUa8OsyukuFIrKj15GOZMfDw7nzXG7cwlfyiX6rEiTQhtNSREmTxYOuG
Atzm+8PpE2xlOV5gLGL/IitegLdtZBAGhp1D8UvT6p/QvdKzLx9xu9iv6i3XQ5FA
LkPRigTPZRMWRQJcihHfZnFA2CInclu83ez/8cGoH6PM0DlDPzVLIKNNlciyiVyE
Bd5SWWa8vMS2NGvSJzGdXACb60Va2kUNgi0r5ombACEk7cIKCIgqgL1vp/x1rlwZ
OhviJvY00EBU/uKrB6Ug0+uhtKPghp8jd6ACmoQQVj2Fu8MJJMIIy3jZOQVJiDxg
FR962TDm0gMybhG2wUfa27bAlf9Fv4XN9o+5gXqh3FZQaBWc+bLy5jn389UVxj3a
wmdbeHl/AFcT0a4vBfu/w2E7gPIrfvqD98h9S2zGWNUm08hNMhKT5MhofVtYMb1B
VEcGlZvbfP4wTYMp71ZYgY4PVNaSffLPWr4UlCYpA7XW+96To7jsKC+Hs2hqNna8
/k4ZqjT8ZRufXSVMRa7811FGqIB/7jGeoH2YYn/63qlxouK/XbpengWequEyBu7C
EbpsnV6ZC7hMKDhXKCtdtrNXcGJItu2fqzAJ+7PJzYUcHO7PgIfu2olIzPQzi7Ib
jDqMGz5UqH9Dmwt3hDdjlGH0ky0QXiVxokwVkaANKtMZcW32BantCeHCTh1m9D3F
nNs7y7DvgtFpVFNJSStvFjzCc2hXYoM8RbKJcvxbjb3ROd3c9fnwnVQxhYyd1JNE
wiRgEnfFuuQNJwTL2ZKKPiBJejIU0iR5knW6IBj0kmzEBhCn29gN0+htUQwbVoqv
9+pj77ov8nd5iEWpXJOfs8kjsobs+ZZ7KEjgGPxHgQRw2EH1MzyaoMmuv/MGuJpL
5DEEsqfHdg3slNhxhoYl+hUhIqHq9ufmBEB46COxbG0BuO7/lLZeCy2/Axi2w6Bb
wqL1qAc2bmq/7FAIf+S6W1mJ9mqXH95Ivrb78R3U/DgFj0Fir+vmM8JVyTltnIpn
0KIa2bVHdx3/EAN3rc8uptBa/BxGEN1P8GTjJIbmKGGNWdtCtrkf3/mbr08wn0EP
+FnTFArxVt+GvwQr7HujyHkOeENSZUR8/bOQa9/5pSbq2ZLB7Q9ptSU9+PH03YBm
eRUmGuelnF7y3BDYr/bC2jAsz+jFgWp6zXyybSwU8mkpzXK0tYsDUfbwoZ9Q3ogo
EMIbzcBydOjNoYtvZssw9bHulSFwyJo667LoGZaThNLdBUQ/7G1rIrsVsveuaVna
NOenr+pWfb1cAI2wmMRREEqaxpMGTEA0UuS+BuwbShUXvhbnjDaZZVULSYwss4f6
IxBm7zqU8/akK2UIlIhDT93EXem5jbw7dGxhjejk+CHlSj4wR7+bvIinPgIHmnWf
8sBUjWKXglx6kwiRTx32zuHvEXW3/Vh9PuM0Gl7Zcii7LjL2Mya6xXKN7FeT2rp5
9dJOpnbkrFC8bWXKPKeMzqoKDDHkioSrt9Y+eq/HFoX58e5Vq7L6p5Nuj64WObyb
T2YhXg8GFNRHeXGXL0y7Jw8xGRsAaHVvPkfToSVcArLFUsQOYuu+v9CY5Bj6ebVE
IDlzsRWp7Dn39XbzkjIb0HibO92taB2sCfy9anovhS0/87llSOfWqh+Vyq57jHm9
HDPaZ6yh9EYWfjByNtRP5P2X6XGjCVI3g3VqbF4sMtJfObtjBwavDooJsSGLzIRV
ZVJ1LUCGMDBK+UUYuhznCN6+85Ei3FOZN43nxNH0x4AqitNqzWxV1H0rD7aaNq9E
MQyV4ul/r3ESxsJW4hxfTQVw91FbfhY04hOb9ZX2OMa3GXiUEj7l26jgeA59lQSX
I81CKjEpb+ZjI6Q9yic46DT0oNGjl0QQGoPuikATaAJ06rWnlR3gvs2w0oNKyur6
IhGbfmcQfFYQcXQz28nt4LUFui3msJNOPWxETPRnOr6awO/256hJptjYkrGHARNW
YOc/D1cixxS58fEVb1OWK35lQsEZcJ2UsKsaTFN1rRA6J+PdFVvC1LPghPXnKXOT
j1/1ZYkPsgC1LmvRGLx9SBn/rSvH/giRWnSByS00lJE7qxJg5Q1qT2/726y2PEFS
HTb7UaQ0pHFGJlfwt0ArNcGjqJeZsv9GfWDJvufoxPjcyh4RrYxR0hfloW0DwAsw
GL7A784kTzIwX7hv3DxHZBEEaqTCzr5DEHEEi/7jQJ9IS8rBPIzz2tb0szxk1ZjF
xS3RQvt0gJw4o2Xcy9xhR4LfukiiPJsMkepw2cDeHEdn+/v7OXFqDrck3FoNhDO1
1ZGADkXCU+3YXFEULgp/AI3m4p2sEv/H0UcpOR3uWguQF+LPOcsGWmrjcG9W9tYp
VwUG1913GQ1g2DDBvk+VWN1VRLtB7MFhlbmuLv/gsmThakuPs0+yoJkzzXzRf0yR
Aa+/6lbCt9z5z2YH2bEYq2BYhUgM5iPbiakoFdPdZXo3Ln4BOZgsvMHGa5G/ji0F
X49tBK1UPdUJpIMgzvM3gyUAxDxihY11J/3vfl6gAGYKx6xJaXNuszTy0OjAhPgo
UhMYvJQK6ndvAxj3Gh8E1A8FyNC6cwC1hzd/ZQTgXElI+bzZALqf9zAK8vmDWid0
vHr+fDXYCIkORUDU6IRK04bWrtb4Nxii2ltm+gvi0zY/P4Ru/e4xrSW52WPXOZgJ
0jaLCmwpAragvR3repvNYHn2n1ihx4yMalHf9iBfmDUlcXiBUkEi9vptFZuTGHGX
rG8Prn3W2VrQQEeZ8hFMXedIRLqc6exZx9/LWi4HqvNDqhNk50FABQD0UafvNC1e
YmhVv9b6nfGyeh0urardxoBoN2K6+qcHmWmTZylXPONK7cwKjlVtND7jKnPg0bEX
9XrnDeGcDx84DRUI7Qz3gxFe2gyaY3GVe6b1xSPtZzFc6Un2jukAfYtbPj9I6cXo
djftVjMFFhzPQn65slSFMlydvAVKIEwkyEwHuNOJXGmfxC2qqZtE4CQvWEchTbrh
sRsC8FcH/j3ORq0DND/7Rdnv4JaaiggdKVwUq+T/LRTKif/RU7labgLliDhDhWJg
8qOikeczpVP2wHQMJSbGD8QddVQGsIRk4BydUsm4FHCUC0cy15eBu5YYfnD2hjaN
MBcU7XmhUsh8c81SpWMsMLEpd8waOBpiCqcJZFUlhlHRBhALQ9a1aQ3LJOw6qQoY
gb9We0lShiKel5NKdv3pewwbvo4RwMk+iEcZj9ZOWXfRXGNqI0uWZjR8Qyjorf7K
n2pWgiCRmSozuGe7w6BU1Up8Hn5J63YLC/qcGdbO2E6PzHkntIQu0LjfQGtXKw9P
bhTcQ1FItClGTKlRXaqx80wBqP/mvCtjlcyoWtV1mNtYluZFMDw64ner/TuB72mr
hFD98xU8aJv5use2E7AvAaIHX/AO1bikBh7yANKsYfem3xR9dldLBqSgvNjFQSEV
WPnJO02hptnGPrns76BliXaFQji91PuVgt7XgYhyc2OvbOX5v3MXOsYnS30TsKW6
xpbQAYFEXXuQTDXKz6/mSa6zx4iWyC/vtqmlVOOYnrPG6ZMJdw4EkkYL+7GXy3TQ
RUFfrYV4fNJj96QhY+rUm6J9KGjIS56zUM29A2AG/LdZkZ5AFMruCJxm4k9X+i47
4aQMNR76hazBMQm6mQHAz2mW7OhnUlRQxxeQ3vS7fIDqi47BZ8GJqSZ77qmK2ybL
YZGb1P5z/EzRdG49unybnADF8Yo1EKpXA+TY7rGui0eNrMqiqjcU4dYRbyagVFqI
NnX6Z3EC8BD47o6i0n4bbUsLZbpwIeMOe07qlHoUmMIEtkz6ZkrPNGIypW42DeUn
5mkUEfjnKzsHzIxRmDrvW/J4lEbr98Jp4A6SKaNGyi87nWp/U8fhq8DB/j8cjuZS
ptAeTgO822mfdzDIW/j9W+w5zoXMx4vY7skZh8m0G5TFihqlQMHfyOKakCETsxTJ
oV0mzd96TAlsBPbLbmvinYxcdD5SXYFRXffOelU1iomGt+6kGwLW8IZM5iuVjjym
0LTJuov0We+rZjc1BghxyjFPJf/k2FcoTia00nKfufHq0PT1qU0iAw+QWyrFdjO/
PeXBduS2qfOg4SsSxpJUbEojsTpoXKYr/ylWogRT+CntNXxxgK+w0OcXXQxgWljq
O56VzZlb31n+fgV8vNDA+BXdebsYFHRdtCNKUNqwFe+fVWqShR+r32HuUbScUyZA
A4BtdEiDE5pwVvtSJ3CpTr0hhn41+geliKN/nAXG5ERy1MmKDp+vLNl/FQkOi89l
5Cny/eQxMu6Bw1KDeWlVpOrsdSu8gLMGWR4wrAaOyX4R+eE3Mq/fz/oKw1CFP5WK
kJvJqkr0Ll5Sy7/t97EUzuWk2eAZWrcxpPCcwSxlCS98pwCiu2kkiRUP7VP6OTdy
69P5FjuTfVQhZzE8JxLDDi6X8bTYbhdiMWPHyyMjKU0zhTEu6I69k69cjjWwnzUP
+Wob/XtHRIvkwJ2BTm7ABKDzLOIRVa3RLpqSkX0a0Jaw8CjRlj96WJRsXTqg1b9J
XrHE6Qhkwd93ysG0yLID9yi63HyUPqKoBa6XKRi1SoiEpayQl6H6kEvW5FnQ+vFA
UdPLKfw/QyCnuPv4NznLxDEKPfF3vPo1IsUkZqyi9DfijZAkVQqg5ot2AvSKL31m
nMnIiXao2/3pCXtrF1UWlwNqspXExvXQNGG0QFJK6+cEZKdwoJClcL0UDN0W19y3
4eq+b43aBpMEwa91khPsZ+FgEV9St65OW06+E0vwY2NJV9qXID6osruSmrFvFTZx
dOhOgZKiqFf83ejyPvfk0+VaB1s4FSNYsbJ65gDrwVYFJ5RgED9l2lUZJvdFwsqg
G6Teu17cRa4dvXJYpIDUQn6ibomxV3KpeyCWT52IE35bqys55uVu4M+N1w/FBLW3
2StaaYhk15pZ5ZJA976KIYxYbgYMZW+9NJV7FibKC2DyyE7qYUg0HDOxmfwDFQ12
0RefL955PnWsDTMAUw8r5hfECtoDiG3a4vGd0MDabY0H1yBiCWYiTKDY3VeiShAI
MKZ3vaQHN5o2mvtqcYvxzHeJSxypqsnF3l7cIA1LLbyH2hnJhCUkxTfCnIAQt43K
IYvxJ0FVJoapNYkZtMnoYH7OgtN6AIe/7Nc4Xl+2nA9JP+AlSIqjCNhenHaj2q0d
KNxd5Ft1T6xAfDSy6JbzqE111URYLXniy29mcLd9fee5Cc6S5/r1wdqNGkNR5Asf
Qqn8195xllaED1E9ERR6aLnnB1vdJC/AFxMcnxsBmvH5aB9jmBvDqCeMYZTdUmOt
6TvgIUcVLaRvKJSuzTRa//E97C/6562ZD4+6/CCXa/9nV1V1Wtxfo1pKzv39JECs
o56AyhkuOnexAK8PTVWdMukDc/pWAseW1jQOpLwGPiY9QVlLxIe8pFFq+2lXqRFP
3Snge+kvyTftRAbYqi7rbGgDpxIKsYw+oL34aQX0yeHJGjJ2O9fasQBWgh4Xw749
xBm/vVEFl+RQZjj6melI3g4bbmp5+3gCpSQeExm6hSMZRrp00igsM03PHaaTlT3i
/A98pe22Or+Fu1/7VP+fHHxmXC970RBZLB/T0YlNVP6EdE8HRjD4lLMFAEcbR5/I
J9HgCtBLq8JFrTQNqc6NDaFVyixVxcRNrQh7kfixN2a7y8he5iVyORMRZs8SYoHm
TVITl4fDnkg05Ovourl7KSF74OanAZr7DfCcEURanBfJHs0PMzVzSs/5UcP5p0ew
xQP8lzMaLLBup7H8irF98x40kYJlVdgTawMI4i+nHs5eeJ7Pn2hW/klgbS5Dmgab
o4tfZk3H65vJM1NtJ0yJzv9sjAL16sphA1l0CPK9WB0Wtsts9m1YAkNXwotsEu8N
H2AUAga4qaQyrxErEzjVoSJLrNW7znFD44/ntJ/akQWPnedUqpfrYVxRBP7/I75t
4v1B0wOIsqx6JVo9rHSvhu/BNFvoO+90LLZsJmapoEkdPBBdy7b5k+L3ewZEl/E/
1NJprm1YLBCDLLuf1iYVqjrrspWnfvlM/YTVc81lNsx4hhTE5qG/ea7fLn8slyya
zD6OLrrRcvZjDhOr2KpBdTt33sUd0Bp1Bxk5dYMTqmKluwmS/iHrgzERUEJrbvK0
xLj3Rj+NIeaPR4RPqkSWCj8SwW81TWddHHUthSRV8zItYDybMkCfDMasUYjNuv91
7MN3xe29nnVQR7zDMgEQRmnnajEs70rROFC7inUqbTcbT48tk8RlDHl9S1ZoEWUC
FfEWUpJ5N+mkzBkJUfT+1Q8VcWKaQAx2Aiu/G1MuiIzLIxqoAejWyioz0LT2YTp6
y4YcHZSud6boh5g4/N6IwMRf33ZdxNYV3iweeY2KdxsLT4p+yNk0zjqG4KJQOTV+
/JG5rQ+HcKLcSFGje9ImsOkDqTQxbJgmuXcdTclHtEX+vaa94hGBjRzVjXFpJbWz
nbqOUNYQKFe8wHI9pLi1VOo6yIflWX8P+NkyMtAR13bUaneYVphO3AhrzarcBhkD
Ep/Gd9FCQic9oTw/p/SuGM8S55ghhiiGqaInoO1ExG7UAn/Hiu8l+iAjaIlvwNnV
PfkSAl8+bnulsHwZiRFpVKmPjk7rXQSqNVXp21nG6+054poX/IGA8Rt+ljwv8x6r
+MmXXb3mg+Z3AeYwcGoGqeBN2LLLpRJMvljwqkgF+uuPy51pGxmauZOiuK5/rzHQ
WQjuEMvabmlQzCbBSaqoT+jde/JVmgdFSUEpLmDq0Td9VDunKf6Dhe9/v/7ZC5as
Tf+kyl6+tcx31VLCoaZT7o/c5smVJMicfLRFhocVdHQC1oi6M84k1OCzvIVAVjCT
xlrsEOavIARia1N0P2fFMDGtsC4jrVT+xn1U10FBMW0+x7cGaYsxhSGp0m9QVmmU
ZL+47YC7gS5FbgWCeiZgfxOSMxipbmPfZuJcbsnLX3UGK7OH922WvmYtfJkGLDy5
Xj4zWR9Z4kv+WyHCQKGOvo5wwIJgmmsokkQlLsbjznCgVsjrOJbCWR6AocKkDQ5n
wqsIJUk1IdnjVNqfL+ph2gtIBjJBqV/MfzjHGcgwgQ8MFWqunEDN10e7d5/Xf5R+
UzXrZvzkjOOEZvl8NIHox0kSjRbW5pzrNwsXzlmcfr/lwZ9mVTviOgb8uKvumbTZ
dVFIe3PIUM7Ml0j6rN16Z4LD/pr5/A2KvQUhV1ObGY1PPfGK6qU9BBPcjgtoE2Bc
zJcFdfSH8EwwyW6R9guHmRYyLEmSAJLdQDgnen00BvNG2R6yNjP4uKsRsiKJf/pZ
Yz1MZrRRuXaBAQNTku15C+agNLazRasVGCyO5p2/jneCngSfs3f39aQOQVBxeXmV
s9RIZ/HigSl0LbxwPzr+tKMXWKgv0OA7P9npomh3g1Gw7xZKZdU0+JV3ss/o2Y0t
7FtRLtyBMkKwG6I+L0Eu0fq4PEKIOXkDGpU01L2eaHK9sfGWBEKJgQut8PJW7U9W
VhmOlC0Id11IhJ6ndbB9rtU0AJDEtAL5LUj2OvJ9re0iRB+ZBdp6LRXV0aQ8KR+5
SuoEsr9QrjuHuvnSqitxFQkzWqzZpZSDfsbuQt/gxJBIKkeqQuorejrkd3aBb5bk
8Zj7PajOmdmt837XOc/dwpL4h+/N4AYwY9G9BzlPByOqxri3hxcs3y9foBMre5wo
olGcZdQKj+WLL4IDOj9UOHaVQKIdu69tofIvkRp7D25BvPqBNjGIlRFOpfK37PMQ
xdp7ao+O04v5esRJmNoCV1UxJLQL4xPktvU4fLymzlAid1WjFEFNNtWfi3UDQZrG
kwmDTmWbaSqZ6l6KsTRMjdGnoDxVcAWY+YUAYYuDWGcmE+IjiZqpwmgsksOpsLvn
n+UlX8ZB0+7iETt29C+YQ+HQ7zC4ph9zXWiikEt+fbe/1Avbi3fDTC5seGt9A9CU
Jx48+3xOV797WJXDOXA/dYMYrZwiZmENERCWj0jzCowyQwa2xsaZfAvHvZhoblUt
Du655MD87gfLqBCihGQfyYZVUaET7dhFZNJzkS4Wde16kNHg4phJSW5PR28QZxvf
TxWdPcgZzR0ZS1hGFM66AT6WR/iKtqFAXbR6xJb4eJa3Mfw3tpTCoFHQQ4QBOhxl
SZ6/jM1BEvQbCbdoDgiy3HWhPVnL1c18zlA74aukKEAxseGP5TMm414ZsyMpzJoC
m+beOc8A/837GFbqVH5XXb+CVKIWSChqnjhcOgAFsZmmPPc/JURQvC+VJcZbWiB2
2xhZtOYtxoGkIPECsGLhNUNrrTEIkj7sgnUGIcuHdrJzUVk6j7gBCAIzqGstKvgA
PhPjierbXW4w/rt27/dSkbkkkTbPt2rp3pbPrjsX7Emnc97Cc9Gniqh/tWmqhmdN
9siovcJWqGOOgHtQhHKEdeL5Fh+XDeK4uB/2NIm1AtWd/4y0NN+uqAkLGPyk8Nl5
uGZ8qEE6zhBg6rHWcGliv8zfrtPZ1xbdYy2dd5OAqdUy6netaw9fNnNkBFTboNn0
Pk+WLiaj8ZPGerIh3C1uEXlEK1JMleWjctyQqR/PGItZdo+DHLcSOz2taTCrEFuj
V/ylHjOZc81fXrt6XUIaYdYfn8KzRe6TORDq2I12LDOcKMENXdqbc3zgqQbjE/JD
VqMnjDUeLmc9VV6DASSgDgESdTkaojGi53Oj7oIAzE2e93Bb0EsDsfy/SwnX2pjt
F2gLEkK+ThwvVX4g1PTbl+h1LXn8FOEARavAqXJYtRGq/qjwszmQreSHI5v0oyh8
FtYIkjQANnWWfqB6SqkzGTint+QCdYrrvITe49vsJPHG3wOifadL253yz2pux2j7
n9yJlF3X1Qk0NpVxdEEyN4MtjHEjSl4pgGI/WEIt5tEtG0BxQPyTnlteN3quXlVa
Rlo3oaxdIjNK3XnkDcdt+5S3WZ+cdG41JX8Aq+/Hr4/Vv+sHSqrMVssi0Vz4JeZF
VpyF28rnNcxiruR3oxbQ35UQ8aUTPqZo+vJ+s+dG/1XzNkbCU7eUkBW21rfVTSsI
J5uBNx9s9qYfoYAyDiPvdYRYv+TOFtTf+oforRn1xLSYJtvjzLY5i2FAziACgjR5
EUIe1+uAGHlo+jOFZ0Hn6W+2uzpi4J9l+LwlgoFHJWy4SWH3KztmNSM8ZkHbSdCH
8NMWFNVvlfc/qPxWNgb4PS6TxfcDBn5/59rEA2C7RuXJfO55nkGUJmHTLssjiNOa
6l1yQgSh17EVnBJXEVIKARyHgrc50mT3mf03eGhzHy+DTb9Ih9kbch/gM0sSRVjy
7S3LCbsRnPrFKKhPKJIgwxvqqYIHASIdSJ17gj3Rzod7I7re61SBH72mssJWW3dw
av9vQeuAAcTfngMe29laa6msMk48/9NnsUUgOWGZsmJqolW5RjanpgHpAP7GDxkI
HJtcnjr/Os1vL7Lc4JoKuOwOU0wwZ12JEeXrovG/hZwPgvCUfIr/VgoXxYN7+s/B
s7ISY0eooOn3ddEc9v4LaJ3U60ps4QlVmrTQasXe0nO8kmoG4Oh1MoSHsIhLhGeI
TNL0h23DkaYNwpkUcRhc620fXy8nZLnNrvCBtgsxnJKaPHoEiM6DenuQS2sLykME
uUmxin1tRTuJjDe6g4hCxSKrJ5ayLlpMp1NNR189+ZtRQLm78GS8u8Gku3OgmSuT
hX4Rzhd1c7tkieMnJkNy7ZrOt2ZkcSWm2Iw5Q7LECrr9nvJWoJN0qFPtl+t/7VgL
3XPZ6XHfaLNdGh3dtj8cQD4D2lIyVzLjwV11G1Sno0zdFYF+0hrsATjgOPQH9VNb
8SEoGuhUWPff8zz2QZBSzhAHOq2LjzJYgWTdRGuLUxKgFvW/+xb3Cs52x4Fk5unC
EkiHLpM+VgWdJbV/b+Z8b96KrRSk3S42HbZ0ZEpBeKXL4qw2Ss4WHSs/2KkT4uNY
PdJZhIVvEcw6+JwsdCX6iusq2ZPgNfE4KhpdKfL5b1FGEiJUN+8Tffh6ELLeBXxD
KAUF9ukWQhEUF1R0wmRDPh2tHZJHU1g1N+3kM9kmTgGlD+OR/s5B+Ry1h4Bs0yiJ
Eus8k6qhObnbgOAguD8bSECTt63z4jPritJBhEz44dktJ+tNVaahwMCiUHFg4Bbm
4A4AhGfjwFcKbtlu18kMEKSywwXYzVUA5QTnSYmyb2R8gzqgQfwjrUop10A9QJav
Bc4i8A/nXY5V/FTQKwc4OQeA1HTRe92a2n3fNxIYJrqNUd+z+ap3qGxSgFImyxaG
7PV/oMOK5OC2nglJcv0YrQfCkMsBraEfF0Nqn7wgoEuTvuJUZ9cU6TTK4Z3OF8wl
dao9Yb4olUdwHRDxVwBDmbtorfVDjB+/eC/UiAEm4pXE5PvSI7gleqYM0j9816wq
ZmC63a+wPCBEgytlvHsoEfN93acp8raapX+r1Cesk7pMIEHvzRIZ4gxcTup4b89o
nj6q6VCXiqtpE3e4MRWQ15S4PFMtihfPq3H7gMsjggbiulKKrmuQt9huCBHVGh1j
6kJsiLC2EDZDOfTqBpGjxli9NIwWYjC23TU1ystKfgvf/5IIB+igvNiGwjaN6Gxi
CmdC7MQPl+HkywlcQuxoTbVCnG4ezXcVTRiutFpCCGw2imUEPgf+OwR3DwVa3JcD
SzyHuaS8e1D+JxrbdMA0vHeD7Y/Ayri4xvmQJaUPkpKDOjUDhvZZeJWu2gRA0F9A
pNPe6HbaWTSKpKrKr3GYAOb/iD3hsw2K7bL/AGaCM79eqFtsUmtvNppJAptJiIVP
yIZgRiy3h8t8pl2lwACXdYwJ5nyYnRuf1w99KBnFRoT2cQSkUhy50aCX9qrF8x3/
iw0l/owOa+DoGlU74KpA0zvP+KrA6Zlpvy15VYLGscfcmuUpVsIult2qHZScLKZ9
bXADriSPy9GCt35mFK457uj7DmP36lYv98Zghx22HF15om9Jd/1SViF+yF3LGbkT
gR0ZLJiiAnd4M5flBGNXeaFZUz8+Tdi4jjKvsyrYmxOKAXoo20seNlFjT5EANh32
aI3WU8D95dRMI0j7dJcxk983JeACMXUzzR3A3jFaQQcXC4f+NOt0LhRSMUqbop5H
qzdmLwtkI/oJdUFDcCte1fZbvyKS3kAB4Ax5XvsyyjUk1sVLFIaILN+lrWgO/zdg
TS4aKJle7Vtd03EN/izTVOpWXv770O77aKK/N317YtPBiIt/RAIEOHcH1aX6Y5xW
CnDC+VWQsvnSLEos3B+mKOFTVNiC5lU4lrswWnMfxolNfSJ1hyEOpsY8aKUKxS6D
nNDRqTWlQsjjvYUttoZwtt3932GuhuYHyQjvoM36kRlRAtPTIz9mHrlUdEyNIsjd
LI7zTpHB4kKwXjLKYxnG/GglwzQdnC5I9PONNifkFzcXkfBD8XrgNJonxjAOS3rM
FagEkpITGLE5u7lycvlIwBnGMbJgiyS+VfUNzcPuDXQP4+A2z+0k/ZjxQmffeDv6
lmVrfgkSIK1zFTWhOPAigY9vRcdJcoWJsHJ2UDoUFgj9dTU5NIbICYPoRV1uCGy3
R6pAUUoDhiiK4cZRnMLnAyYrghHrFopeItkrYg4t8flJHGs6a/LbB6gbhvRO4BLn
g96A2MdLmFprufQ20YJoywh//TIc8ddpGdXrtNatTxepx+nLQB6jAI4fb2d0eZEB
W/I75Luf9uzY2u2kt86oD7+k6/arazFRuy3tWciSAuXsJjhnOhQcoT70AQYk3O2R
7deErw0x6pfImFTGcMpnVjqLl/ipno2biPS/AqwzWwaXeJS/bI4HZ+SdfzKX0+zd
A73yXSbV9vViawhgJafHzfI2kROU05pmY5b6WNk3Ns21DDtAOvEtEHQ/m6J1j8b5
dpsuYm9FWzvTLyIyUYhRgLZ5Rg6svHOrAdLM+sT+6U60CdwA9k9Gyj8Sta2kEcVm
4MXEPx2hX9gUWnjIgRz6PN4AIYHB8OBO2vxfHqg0AkD5O+tbuGcmUcNOXbqMAkA7
pouhQubkMl2j1EdDCje/GfD8PpKtr5jFPeafZ5cr/8g/BBfevnRLS8OBA2sewIEJ
UxRadsFmD3AKpIUPPkmUumSLO5sLhFLKGo4/d15N+62SXRMD/NOW+YhoEUs0KSjP
oA9pC7ZvuyDSDeNS8HnR5UPi2e6ZbX4HFRPs8etxv4Qjkyaz0PdFIjc8KMuWTmt6
rJof9lpLp12hfstVH80iEb8UPZUY2D8DvxKfikpj2WA7AhrqMBtt5udhxfvlhzrR
OWVSPCcAJQ1DwLeUufUCTbAZSi/r5fzqHAk2aE5E5wRvdKv7+ZurUK8QzSteL6Hz
dXPXq7NsZLXjq0iUT8Wg2Zxt0nPGgA8XZD2CG0BJkU+8R9w6rDS4m0m9uNR5FAXC
g+vNhy76nw3TMTETtF85AXH62cFYDp/bLta+v3kx1sM3Mqyqw71OtXFv2DYj12R6
kTLgGsBi3JHcJ1ZE3Ebw6mfay1FoNZzglFNCKDrw29qj+V2nU2XAQXIEn/0QN8LR
0R0wUCTmsY+RSW7TdU9hbTQzDD9JU/4T1nGo0Y6n7iMKX/mz8ChiBZ9eL4pkdA2/
5vrskdTX0H0+oDhweKfz7rlshIfQvbc/XoTNPT0CDyKcMCSGk5M7fLX7vReGrjQO
+nC4e6GsFlVZRwo8P2BcA/obVKVpvy2GOPfjOCMLlk81xq8nOHkiBHtWsFepPkNz
TtTE6HAtCenuGts5lC26lgIxj9q9welMG84qYBbVkfyyWM13uuM1qzxRvs9u//oR
a/zzpQ89OTQ+jCraVxeaNFukZ9AuuHQdRLgORey3WZSldle9fz7y94gX9PdmiU2w
fQZPXaHyhPCnHuLf3xVBzdMATqFHn7XtnEwORiOg74qa67QXDAadUt50NK+vorA2
Gfwfx1JpuVa4GBhRNZ20PbD0rYbQGfE8jnCnCUNwcRPGFHOVRRvDt35aEsBOM/l+
GUcVaxgTRIWOjHYxjBr7HSJ9BU8eYJRLTNjgQ+iUvOWo1s6H8/OGwsbq0fhDzpYl
EmcovuaFRiNUbGYKExXwIT5XPPsokKVQo8dCXYLOQEk0DSwwIy7SoYKVdMaKSdTZ
PgRgsvSdOHo09UTblo3IcBhlN33ev9FreEV9WJ0z5CDJR1NpgIDyWiR8xGyvF6tp
bAAqfoFp6lnv2sto1dTAt0rtRAH+u6HVL/mx9w5VySwxjJ2wy6sagXjIRDlXXD0+
d5YQInvHK7B+JjtI4oyxq9t6NxxMuxyCbwXNZEYJlcHplFxCO1AcyPn5mz0iFqvM
groBPyqO7AWElzzWynZd4zzYlz+U5zhk0b4wEp5D0nPNlV3Agqq0yAodc/IsSUCo
cigzx7KiB7v22OeAHo41BYYyy7+weAtmf0vGa/B1UCiI0GdQCEJbUcbAZInFCC88
qGeco8QI9pbWfS4uVom0ctPQ6NV7puA9q03/xhlDgZvvfRWS7g5LRMSOPB+rphAG
BCLGYDG188eun+y81ysVE5BxeFIlD5QrEYlgn0AmJEARJkg4GgvQZYz6/C/AeGfX
b7Pk86eMfcSgyADchoJaMMsSjkkUCpvl/PyVqPR0ZYGXkBf+j5iP5FOX5b5Hq4mc
J7arfcr+ycGdOzhQUHCqxn96dU4mqMqksYT4SzgW1q3yjyqp8jZIqrNAzaknumQb
ECC+06qkrPFKr/LfNnpS43CUpLaCNR1Ogz5J+jF+Vv48jkBvqJ3QVjmXECMZveOm
jxCCAUcb691HNHC2x7k6C/HtBEOjibcs/zfxTAOftlKQemz8QVGAa15UI3cOq1j3
FZ2a9JUGVJzUtleIhIGBHKNujslUPJV6C7MfBwO+RcI3lhPlWSWYoBKG+FiOh4YU
2asUnvlmBPEJ33UWJFalLB95V86G7/kNH4UfLLZ+UtWVfpkmZZJFgjOSRYMmkFNP
QIKPf82X4l/poPQL9vWmvvdbeX8h0Bk8pJcWk7gVISpusraouEjD6h7Fp50Cn6XO
scKuRpXGvSEweUobh0xbkrG+JGJowTfSkILU+kPgUIQRFExoOoEo8oLNAsTchBko
+MZ5wVK4wrL7IXTGbBZNGkPw/LpKxl4bTocP6sQAULsllJW5y4sdo7hmcPCLMm26
0skpkxOZUqiCsWgE6xXy0/A3+KXyBiWHuqg+LQ9bOuSyzUoDwySqOZRO2DKHCTwz
ooAQQBAONz44UqmtTqFbHZmhYY3XWHeocKFcs8TImqC8Jjj83DE2fL39ccI3Zx8U
PUv7wX1isZFL1fE5ZPs8TTD1YtHlE5//amC37e1asRck+QqMtTyGcLI+m8VvD3vC
srkOeS3BOwLp2UD4T3QTrben3X4N1SeeczSexcwpMtE4d615jaaCwqflJ81TjT+B
si9lLPIjpfV/0KAbnYjfdIXPmci2O0qfyqI69bYGb6tMoW0XTYWtp37+W42MweZI
yN64Q3dCy/8+zeyYTafJAIyohy50iGl8+TSn6a1Y2/1pqEyVvG+MnBQExSZ2Fhf0
1EQFuhiW2q79320Oz4ANNjvhRZ8hdJOTARl4GEtHYTBc7WqWNAv9fadKr8ILIQYj
mUiBvMB/lkt4EYPVwWnesX1HIdTT3kDxTlOpuSOT7pbZN/4C12hJUAmB5RCC7yop
NvTj1z5TN6zph7AuxSCrND/+cvlRt9Tz7tKucpfchVsyvWaegZYyznn8TTwPBmDM
aQ3fdyUlnlF5rpjrjeFnkYqjePU3AEWiDOuQ//2Yl5lU8BZzQYSW5W+df3RmPrzH
W/TWcej+44U918IPDYRI9ljlelzq1T2zecczhHGAbyWpMccE6F3b0K2vfn7F6fCn
xYaeII+bpfY4AW3nhdJY59Nws7TcvGtNlP1Dy0lBB5jPIxA+1iEhcNeQNtYE9xXG
H5c9JrRSq7BKXYLDKjHc1sfvmbOytrFKPLGnftNFKcG3QpkzNFIfyJ/DJgxQVIKm
sBpth2Egyn3X/VDvsNfTbrw6LOSjy8PDgBAulg+RY6DRPdajSX/SyLzlUbPIqDNL
Oo+q27kYVHdyyRstTuqGLP2zm+Uaq8KEKQfJzCT8aq/dsi8LHNztlFEj94tddl8o
LMk4UAEy9qwseaylGovv3B+19EEkO2YayTc3HbCJ+G9ifttDexhTUl2FEJ+ekFUY
N3ejR5Um3t+bYDR4mvAPGZ6/K5bDHBmZpaMAScqC3Tvc+zzXRAWdJmIo68jRI5nQ
qytf9WF1XTg7zW1tioLGobwMidvDOdVDmZsv2tx9w78IfGx0sSlh+HcqUKM6W3LW
1UDxjqFNfJbOjki9kRcwf2PY7qZZYeTGqgJD2UQCRegze4Jwq/UYzWMPVePAnfH8
OYJOPjJwNwNfVw+3+p7qYLvjBcsDmGF9JT3svgQxjq0f/IG4O+/IXUqJoWVAaLSj
wLimhAQ6/qBeRxT4U/P4LZwTAyHEUna8yiAvxxgGBXiWXD6bv2cibHp9hBouQyyP
MDH+RzD1HBi/jJaq/EIwd8iXbzjFXlN7fUYCP9wvM7SHa9P4qyRZYJCoFVTZXMFu
KmMvZdJUlsG8ZWYs12vmaxQTcRIXoxWEvCDJM3dSpQj/Hl5GGaXeSaMOA5deEnRs
G8wnI+dRSHTriSdNw29oX3/QBI7DJ9MTrA+K+0vrKEI6rLyXNwQYT98ghn7ygleM
1e8LEn90W0CRQZnGu+SYaTpS5WRqteRnQUe+3gUl8rQEJPF1aLE/dN6npcp9+1dB
tnXw7TY2ZAA/tvb8mb1XuQF9LKz8M4o3RIVOaTqoVUPdxxY0XNvq2aEjVDo+Q+m0
YqkfqnYjDXJbI6KtrSueSVpR12DpQ3nEdiCVQzelYjhYEuAcBghY76GPqSKpIbC/
NX1pf+Rh7kRn2cChxIgpAZsMpzWecVu4ViWf5YPCR98D6Woirib3S2wKYe6XBWVY
imPQlN6uylYWSrhOpRzmXNNLMuX0b7LTHERYuf2IU/GAKLHHb0ZmwcOCqXLmwidi
4H2dh4kkyM+XJTcasrKHipGYFZLGtDrdqkSRs6u9agnZXCUDfvevbWzMZySBP41B
bZmScnhNJYtoa7clm6lq8K3roLQ9soQbSVt+Q2cnxqSl2fadj6LYENWlkJqGPv9X
ngkRNn3dxJ5smzXH2yoA/geIRGsrWx9nC83SIh5hZ0xmr9M88AajXkh6dBJ6ashG
untkbuf1ELTBqRnVcCQJwq2/y5Qw+00r7NL8rkLjx7o+zOo27pFjr8uqv89uhdOq
XjANdVxBoqHG+dM5wKu8gXpHzPcW71EJMI/9KDQtxb+l3v4IFdDrwLI7wq3QbbnY
cY+6XwqiPkRHx17lujmks6w7zk0H+zg16Xsj58l3wx2wYpJ5lfpE7cVeSAXcWqwu
jzBEg0A4X2fYhnirlsiUwe7F2076pWLTzXItcCLpWinTpPcJRtveElQHmwTVslGC
RYwOExjHM4xLqz4pWVM248FdOli4KRhDnbu/JhEoHFTikCWf+MJqLZ3EASkShGcp
Z4iXgQXV0eTCJUBhD84V6jNks2BJ2+O2gF/xVZIM9y8Zb1TAWVoqsR1CJytTBRq4
TOg8zKtPxwPeeTGVJUul/tUpdsjL0BmK02Z/qXNtHVnBQ1Tpx5GtgJUW+csiWGGJ
EtIvqa93SC/Nui5SqurH4Juj5RTRVaftMXYEqztTbHWddvGwYAb8r1gOtFnYGI3v
nxIBRjt4Ya4hz4m7ArbMMR3YBdLfuu2oR7ACbQfB4LwnIV8bPvyzXLukJC06lNwo
dagxnkljzuf1z4QqgHmxw9pxMTBEWfU/HPeOXYdUo0/vdA1mYvx2KJrLQM4+gt+K
I5NwnnqvlaH1C5K1dJVtNACyZeBW39/Zmt4zQjogm4FOnkC4eSyGH2O7WW4VDtlK
PkPtRJcU/nb8P/ZYSkhvOICTSUhUny0r1+0RPyiJrKA+eshrGl5SrcoUvtajDtbE
WbSw3Rxrao8PlJZWZ2nBhsZgQAbSLWqsdaGZbI+bFZbz9/pZDdNow6YsQ4ZvN4CY
6EpnEgJ+CMm5VMoMbPoiJBih6qLTuvKQVAuLtx/4Y4lBoaP6yPFEySwRQCgzM4uu
`protect end_protected
