-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Ux1ACKIOXiG924xa9aQebtwj5QUWyNAXpR2LmkbhryIbwQTwqjIVGxPuEkAvFNz/
rZokGZ+qBmOjGHI0R7FZ1y73rKLNfL+IMLDSCp4YHHITxonheDi1DHD4RazZnuVw
DgO3C9JH3s3aS2fIRi5ggGB5ZxvoUnCeZK47sORpmlg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10035)

`protect DATA_BLOCK
XR2A9G3xpUtqPuG0G0GHIsliWGj9dKJhF1pIL4fWfIxBILTDr/DH3To7ksN7Ybxi
Hjo2g+F3DeYO1F8QgHccsHSQfyMU+DnmibssZe13WZjCmQeabVKZ5RYFnEsFPMap
gnYBbuPU4sNSYENjHUdyt3U1rihenB/JnP59/7zuA15WZREWaIH8aTaaRiecJN8O
bei178aARGpTsbEJD8OyUBNMXSEyGmSg9W4LB1UuS1v5gWC7XCYfmr8mdz1QWRCp
T7Hl3orKaHPwz50B1cIPCb9ZzTjQq58YsNwALWMXQj6ykZbfOOwUv2w66GwrAUix
+zipRTHoM4vzUqX3nLyFEzxAoRNsZ3FYf+9QaikzPEed6l31oVxTD8dPKToowQeA
+yW0Eyk3NBC/GxVz0Zz9k9qBjFMUNHauFXX6Hxv7PztSIbeWTGXeIez4zqD0jdGm
28rCwDYyMgUVRYnICAIQDXk4hotYgncUrrwNx0XKnp/7E62uYQTbJnYUW4haZer5
W3FIx9Ep+HyVaFUT7cm0YzJaMfy4WZW8j0UqLUi0Ig2206lJ0EnBIvURxFyIKk22
4a0BJlwmMm6rSRVFaRE3p05USChslqVk0eDXlMtuWs8G30avZ7E2YTlPMEdpw8e7
uONS++3ko1Hw/uJRQUWe66uzkrjMeHfocUP36XJ3o5hSU8IFIPCsmcT1IxoY5w7x
ZYQ1dfRHkSvfUrVH/+qUQycbtNX1uG9h4H2/Om20ASYzYV2wiAN7LHUK3QBNoiYa
os12sf2J1TGrvkRuE+nQx5fpD7zlPxUMLXC+RREWR4hyJ6Cto4YhV0bXdDRrTx+Y
fUCXJ0XDACkm1cw3BbM7ms+s1F8obVwDoi0C/eTzCfDUGgSsey+FD1CGPNxRZZjD
qObOxG4Gfh1/gFzNhuJmnWqz5Z2qos4+Y+Veb8fN3CQctxWwR7omhPD6kndlt9Um
c4n1BEOj1z2xsc1iUdsvPS2+G2mOAFotmVp3LctkKLvcqGWZXm7vT0tzLu/W/Y7g
pU8RbLOcJCp6leEcSjRi987v7Otp9jNXpRdVbx/8PyGNHJ/s3t7jQMcyc9InAPRH
sqkC8L5nxph+1GtLc6fDfYTJGt2l2TfDz1H+zQBb5/0nyrGwU5KeuFKGhqj9GVO9
3vqldXeR4p81k6vTJWXEfAxjhRMjfgd630R2Tq7ijdzUrUvTIjRpzDNif5csOI7a
uL/POXwnsYXEHtPzyRTr/BaywyI7kZjrlBlEIxUB5P3XnmAN8WkXA6m3/QkWlbB4
LPmw6QuH0ekVVL7pefUNLh9iKRoCJ9SEhu7yT7vXXqZOL5o/X9xpxlm6AugwQ6AX
vuov5qrOjjJPurILNu/RoovPV88c/A2oAEBbQgu41rZ1Tu/J06BeUTo3ClRqhfVv
TSvFsQxbAPUP58A/DxpVWN9ZVzLmOlFPVK7HYG7clC1j1IHmRZQ2G50Iz0u9udQ2
cDdfnywP4mdyvCSML5YxQc1Y9Kkj5xYlQq58NV9ylBv/JlWx3OWnv3e+cFS9BSuV
w/MiJ2ltvtKEe/xLc3bxRVdXZRiyvJZxSwmidKrYQSRU3mbEB5vG9SX2SneRP1wC
27FCTbhalaChnBWmxBXmH3FizmSy2cMN4diTaJCdRv/gBrBDtWDwKkbXWPpRFBzD
VcZMhX70g07ZkJsTqJIdoPzO3oiT6sQ5ou2LTFl19a526CP/AEbnb/VVoZGc8uMC
Yl5ie9cxF23rj8jIs71I+KJ5ZhSlaJIopXm8BhWUmSvQfHA4Q+5ealXPxxYzmT14
ODIsEFryt2D9w/vogpgNhZhwFGl6lzrPNKfDejz1Mnav9dHAfyTcnvxFgTqujC/+
5s/gLMIcD6lDObZL3JNtSZ98bIRLCv+yf+7l6p+YvzFxm11Czea0cZmMQz44q/77
i8GLu5pmi0x5jvwuJLKUrSpFibcnqUUrj7PkQV282Njiqw9NgJ5kw0PLgsCfo0iT
Ym04RkMOCGKQ5RSB932MlBykYbFeojoZcw62W8tS7zLsw9pzZXeva2cJPlXGdjzc
e9eIBcwi9ciVVl305Nkvzh5yl/He1YYaMP+HDNWEw214JNlwAIo0+TlwNN2ToRep
0siAlJbpWVbgeADTpM4vQWp2vgnNZRic8j8cv2EcdU9eRftvs9oFtzVfesuY2GAf
urSgYFMKdGCoINMoay6MBeHE28Q2X+7gYHyEqOW2firsYBCgFpL18/LBy0uiNnls
+LIdV45J6omlFhZqA/pcp9OQOgiDKpMHMbIdOT9u4aeHaiVt4RN2KaXUMjNcdtde
dnXbVbB895dJEnaXbGu7lfMdUclDaNYMA1kaIjqIJ2Jl3sXHTLdmz96nb+xZedpo
QlKEYOXzfS6rBb2ucjYhSqwZDHqIhbWY7IUqJ/hZjCsTizaAWgg2maDs2Zhcsf2y
yP29mTLJ1JzC8vPzQ2LM0JvDHZWVZevqk9sH8Hl//xj6p7cL9CUMhyw1xoqrpbHZ
rQ8V2rr9xfQ8Iifof9d8xxRPr3oNNqDv3s+UTL8i7sAS44XsOh3ZsCzHFaVbQGAJ
Rz7YGdUT/dLgDU0I6FjPwNV88gtwiR5JbN4gGBEZi7SLAqyNkjd3Bw1hQ+dR3/BB
yf3a3Usoe/S0v7sJ52hZB1lAKgWqpUqYEcFiW9PwyXNIWZs4LTeeS5BohX5EAJk3
y2t2MQqKk7RE3TPkNltGPp8cRF2iO8PRbTrBB1T3yv3dsIsq6U9iDj5GIgQsSPSZ
LL4NYbbf8QhKHV4Q+BQUqxj98T22RYnLd4nfUPIcV5zFvH3+ELpt23yvz7xid4t1
DL5DegYsCoJlIAwjO2wacFBlHDQyWrMoLoH3FjsH5av26ebm0d/J16fZsvYaRrmW
2OkXcxGS2DZT5tGo4wVfJ39Cyr0Zt4ZPZ4bXFM/DA5AK0UE/HmG0F+2LIzyujSBu
WqzAdJkQ46RZ6Pg5K/er16hfY1EGWzWvimaFJYeUoXOimgEb9Q+IvNkN6J3E9exw
VY5NRmo9PZbZfrifBoB7kckNr7HdqMSO5eNZjMSXCMmhnhK2Vo5Zcz28S1gBFqOM
510R9LdpVIO3M78U5k0UcEAqjKRyfUfzHFm9TAxj0C2PMNb5lasZJUEr//HNPPVt
TauuB7gIMs9g4UaFuJ6nxr6Va454NraaoPj5NMxN5HGdiXZyGc3QC5Fm6sVTpy5t
DWfjDz1rPV14c6t/wVq5iZzK2uFxiY79q1RHQlheGLnbAZJLDM6ImOYYMM7svpNW
XrAJvIwlmOZEhTbR2+X3VDkw/H7m3JyLlQisw5S+dl//BsEDxX+4dNy3Da7MGmag
0Ys1JpCM5xvkSTkBlYW9LzcUsiaXvIoJatfOZ6JaSYD59k6vkI6EqEQbxB94O9JL
N5VlzTCC6bxkmqxDkR3KHuMINZu/SqhPIEOyGRdT82Sgf0LznPj5Us0XChTjznD/
4pGYUyhbICF5A0m54zCFQtb3IVStzQ78oHfOfcFx0aXU36zXjH9cC/C0HXALGR3K
ehgko/Lw9dAzbz+TJ3VvSeX8vqZ80p1nesHZPW30kz6nrA8bqv4Y5qjla/ozxyht
QWfJfoRL2ZewKo9efJBz2uXOLgr3No/Td9hm9Rn232VDBSXDnVxD+zCNHsfZOfy8
1AiEq8osoh0Nb8Z/z9M1MRzZ6H1Y71xhDH5meVm/AohNKPrekjlhVMtjO6nR9eQW
v4g0/QigV1kD3/XODwfPYUV6Ky/RJ89JEVm9pV/1BezfUh9u5tXhCJNQkvZgEdVi
faF+moQap00oYorjuqvpYC48VknS3J+Zm3SRGDE4ao9SAg9/ShGZraJg9vxKlPTE
I3wv8eGdc7UjSFiMs1j3gJp+vRn47nRvJv2uA69/xhrN6AY5NmgndJiE8WlANJ1C
uFM6zko0bLmZkFhAzSXQZDz5RDFXSJMOicJwBbHexhjYy1aSD+uifMeZ2mBam5/M
Q0/QnJZzvy2SFok5GAHQzaI/zcQ1kBSm8FB4+0eJ6HInWdYYUQCRWAREoBf7K2qf
qoz/quoq+VX28A7mcp1MhHJNjrRE3ikSyab3YuBHCPV6RyapP3EHzxOhsZC3fNBC
uiIyFIZd4v4h99d6aom8XPsXKCxSMebvmy49nYiPjWYlaVktTaHXcAH/J+mW4+wk
qYH0qEYTx0W2PLzhd7J7ucb+S5Z0PiwhjQksj31m9264VTiLjanX+SAJPFjwodQg
47GZtz3qj9zsbFMFojYfq2MNgkSkfBBsAO8VJhih4r1bPhcITDxyK7p37RAzqY4v
WTD1PzR8kKD8WAHqBan+X02bmno5lmJb0nOeuVSmlzVIQBiErWKOlVvlWfLPc4DO
0Ahip0StY2W7CuUWNeaH5kzZy5KWptUXeEsJ5suwmMdNy1CVObOl9dNgEQwWJjX6
u1C1BjsHrXSzb7IpFQqD2/G9VqlK5OOrgpJ0C8nagIwF8g7/yHQVYtO73geQ7Uyf
Jplej/bo+32YNm/uP5+jfFiRdfiOKfMZOaCBqE7DGaDwXXGE/J1Z5lkxZsZrRL+v
c+pOafGDGK/jtpECfp4iWpOOpm1ora6guSO1Mx1hvYPRDBMlK7M4vu4CSVktqFZk
DofABt8ddeaTHI0A2xXyYL1UZ1TDklIU68s24gU2pqCoORsmbJEi5LPFjmq/deDD
oY7HWDusUGoMo5/ZmHcKR5Z3uNyl3d3FT26wecXAS/pBxbGDGgBMRccNvtp1i0Hz
RkVkxWmPUtSwL56WE1aGuK28L1DDw4z9AUcKwlHqkzgEGaKJOzRM+TIn0UOlHgNd
w7tqgllFKxyFEerj7t/lE6YRQ7QsM4lWpL4SvQ/94hvJNRwZdVcrPVxnjYvlko0y
7E8w2l56ksBjG9EONwTPfFwdsQeV8q/qRjLzHh5tmaznO+KEMJSrzr5ExQdlF/zK
9u0BFKVYcB7USaEA9zDukkj12T7N8XxRPfRa/NIE04CN8iCFYojsC78Cag9KNu0F
zlsqZbhXgv3xaIWENusE5T76wWNQl3VF+B2ScTUu5s8dlq7gfltyDzZsf7cXZ1le
Y8CbEBQN0LzND10HyxpUHjfIg1anHM8/xUOCdxZrZEzoxa0+parW2AQ4qHFnpQq8
S3fJwiolUuakRMnKrDX4UOb/Kk8YF5fAQI3QgB51XDm0zpyHUyzhINODTfh08QWp
YS+FoVN2i99u08GbZHHrjF3OdvR90R0al1gS1vy8yBtdZxzW+U3hGmOx07eQinTx
VzZXCGznWOIQERqv/T6FRwIVvKRB/H8vIPfSCJvVI2KgrZ7zyZ4RYHNNLIt2jxAz
j8Vmi/ktxIQiDIi25nhLg0I7AP9SDUqip8mb6Li7QSTPpSBUzjK3kDs7+xEM5RbA
8ROTEAPDDdPL2YDwDEMGpGBjLPxr+PbO1amz4KSaDIEKTeSvVqUgr0ncvdHVJGxv
KdUDymKwHisH2xrP4O03RbAnQ2LY0Tx9u9ZsadPazNmH+x4DL5DbBUu4hszKAp3v
pSjO4JfhdKwoVeo/8924Yei9US9ardejQnrvDuFekqDagDpL+ciZRcZvJy9vY/8b
DVLy0ZoD7NRapA0LOnbkcg+LCKy1q4KCqfRfiEeOIaFtLGQ7+dq1RSUfGqC9dQYm
jyMGbf9O8IkiA/GqghWi4uaQCT5RNYlVlWgyvngGSru8VQs2sEHLZZ4D/x1fOPrF
Xz7cK2nWIShNSnkiogf2wIQrpDWff8dw6SSX9Hh0QkbWhFyrYzoB7eaDz1z3p5nl
VtdHu1kzeQ4u28BttXlyrl0Y0J4p/8k+QB+9JlWpIgnVwHd1GGrCnTZUvQTA6o34
yVPqAd2wPNZkK7RhH9EVdWt4mg2xBdLyfEqTDxsz5EonJvHtQvMYy6UUFSUCv0US
cL7w5ad0zOq8ytIa8pg7bSv44NCFwfbGzlMXTrud+KwKkZmdnhzG/sSFs7RIxx6n
wUN6qeLkaISLINVPgWbdHm+6uQAqIzIjPSwZkcyKIgKAZ3yhNS9uPWRzU2sT8qNj
N+C84F2Cnz4tS9kk7PxV4MBH7VDHlg1ZpX6BAHzDn4jtAFFCR1Dmwqqz71igYX60
xX1BqbUmIG87vA4OA+Q1AVPZNL8owmyk3/gjEJ8DdrVKXQJ3bXvUAvcuR94RKQcY
5ghJzWZc3XVom6+UD48zg/qBmTzmzo7Fvy/m3Hf749PV56MJqIqOiE2pCEJs3haS
Qf46qb5x3lV6e67xal1qOXlACpMNVg4CcokYcmxs1y/SEansbnpBfP/KdmPkilbh
aaSpoYiP3j1ARdOaQcE6V83KPkEVddMHN3LUCIBIbC2tfrLbV3rBzJJWVYgEXyTN
VH3zXSsCEHaR/RX/085aPKIiMsRogTsl4IEfzq2eFXmAgITq5IgrJ0hK1Ot3Baym
kvIgTmMHv+9vFo6A52v21WaCtrlXa35IigHUuBGJsuI4IYuwTBY/c/da5oLONU8c
nKtNrhk8325eRQngfh55vaPlLHvpvn01HNS7M3ueNvCOM8gjNu4oE5q7uYPJsfqD
khir3wpy2W8gYha9/PvKwsGhF/6Hp3LrwC+uZ4zH8YNsD74jNCZ08q4IXDm+aNTU
nnmARoW6e411F/MFYb/3cL0tG48pvQFd60AoMSsiouSSPbmoCTe07Ri+s7z3+CNi
63SzYTK7nX+g0HtbDocYyrQ3BQhd8zx6PKQD1Sx4hInAX0KIDjHMcbpupgseC0QT
7yZYdTzq1Hwh7AJ3+1yPuhdurxnRyHvnymGGLvast0wXhZvQtR3s2DTdlitj56qB
L4RJ29Sfs66ans4R3XvaulQTegh2sNGfBfc5KG6OhdvugoUBtKksoItD9339CaxA
fP0r8ifD2eySmIEOVfHQ7NNZ4NuTKYU7d3loc4uikrjP23U6eCkU7evTAzOuAx3P
DdaaeNBxvdXX+HKTF9Tt5nhya3y+UCovPdwjXRYVWtefwjwmYX9RasdCL9USSBbU
SutqX+aEKRaRQHvUBXAptQYoTWhw3g9XrMgDiz2kEemvuNZUeICBkIlQlLCdKhJf
I4lyUmIoA7Mh8YqErW9V9IKd6O6Uemn+qG+bGa/S1uOyO3L6o2hovad4tcdr7K3C
BB8mouWmhav4zdkIRFThz8PY5u+pUNbCj8gUaf1XnmI8NxBz/7f41NN/c9Cy0nK0
C9pf5emOXU+xCP+ls4nVvh7barDTb4f8V+J3JAwr2im+mK6tNpS21OAv/ktDs9MC
3bUlRHJ5wc39jkXHN8VYNUX5G/mXeJopKcKibsnOJIj0Rjg5qIX1oW8CgZ/5CR1w
zhmcYrlDTOLWOiaxvcmDu6M26b4AvLOqBVSp5E2yICwXxJAG9E/PyVlTouHmZbSM
PQaExxJeNMNtOL8YsLPPltUnx0+gag+9xpHcLfg5DuYqZfoyUQ3WEs8vSezpKDKA
SQ3Tnfidvv/v4GsYRSo+pg7YDyCmecfmXuPChKjBo6G/EKJMvZoVYgFjHSdVYRsE
3tMv/dONwdwEPxK683rCwNPIKL26tSeJRLqFdOzZVWJQTP9DxZ2Awvix6M/e8hyO
lKNjVjl6NaKlCsD17e/FOap6InOEqzBuLEkS786esODQV8PpAMRmlGmuca9G7+G7
y92LzEm8vNRo81pkoaGQtwwaeJI4O/2XpIgY4b/m3/9LqZrzz58UDnHoO3BhNKOX
sf3gwnqCx0slYG4iZYvncKdXf/yvs427jXll7urQQZT5uyo7JjakWsbnfDq93pLk
5bzrnmYDXcyolM3PpTQd5+SNOMzR37PfPMqemr2icAux5mNOwwYFBFr3oycillZW
KPhEXVZJ043fmxZcSDBfELFMc4O9RHS1aIWCBgpf11Pdi4Ese4ewXSgsdXU580UN
D2+Buy7S9OEPtnwLVslCvk5J0PeKQDwcf5FWaT4kVrJTyrAqX1pML7wes/LQF92u
yla6DZLELjrjcRtZEqpzm6l/FbqAqhljgUf6WRaYO9Y8FahBQuqreKTURvL0Jdnd
oQIveNIkvQgO4jHqKXw4WSBEe+NiRdQDh+oONexWPazON4UK+7LnfauwWkeynKg2
V5ZNkz9MpuBdo0B68Cnohd4nh5VBCSnfenEj2miOdcbcyKyYqVY7Z7/94aNLQnMr
RlqNXWth1S8PolzfydmxmgcRtaj05tJtboyDB5L4deg0xxb/X77HW5tIWKnYrFMg
dNTbXzSpHGSDC4KE4pW7lXIWjeUJ/D5st/uyfe2Hr2mA4GDF7jvEKdx0b4UaOKRn
XgvfvJiaKYWnqooKfhRxserc9nmNvptQF8Qm7gEfv+TgvQFEk1cJNrEoafJ9NQWl
4qKUlWtezwEX6qNILFpNd6718m4Oxw5aevtBGKPyPLvUavAKz2fysw9fR7p30Umw
K9HB1pscfQsj4Y7nKnbSqMLHNIsUzgwzx9yIJY8PYuvgiJu3Afg8Ja843em0w3S+
uvQ7g0IxaLJ/3lNvru/+Ag6oUHtzPzRzz1IFKQfltKoLLfOKfRCN4ctHrGsqdvED
bzRQqKtD/NrEZwEZcHKz8k6g3oZv8bMKuTttxwKh54h7PGIiTA4GLvjTzbTmu10u
jm9qhlbyz3DxEzAxQR48Y3kA2l8N/txQebi8j6QCZ+Nqca6MbPEYFcC0pM2QRt2G
MPNhoykOjAZILT3F9ZndYoXPdYfDgnMWOPCAqiggequB7L+WeENRn/wO+zBF6xRe
qIPCQugGJ059NAKox0v9ur8/N/wQeLJDwzSvWBUdGEtuIR/7EGmQEQqvqcRoB3sF
UoEH0CCFazNWaIosunuuPvI8PocV7Yzf9CdOKnP4DntQss4xrk102jKY/qfOamye
ZRcZvqx1TD11+lEO53juxO9FJ1e7cigBGgR+Ldcpi8Dpoa3TKO3YaeNAwfs1fcT8
w6v+ZFLdEnW4dl+BzeY06oF/FG+ZCiMAnN2fa+Z8x1LccBqYVcdGq1H8jPtFluVI
Fnx9B5jS+ReWthO1eC88D20NAUMqHFWxF1MZBK/ShR/Qf9er3rE2halxQxHk2uc+
GyLAmwW8yHtOsPQ9gAhe9nS8fLOW5aIHmgRvskBcYuMDuqc4oj56+oOZZMN8ps3w
IFkoduCtDKP22mr6JzTEUZ7WTxBrtUqjuSzVZ6pS4UApJDWzpXM6hrytBbT43JFP
BieUGT4LkNzqYADbnsYbExiv5q23VlSzuOHbKpuy/k4pFJzckabXkUPfUIcXcWAL
VDUqlSiOEPIyrGKdiiE8mr2g9OIp7LSlOm2scQwS8knPQ9m+oX6dZDwmvZhv8D/2
9Y962a3kFfPGLzTDJIkFoYGsgdsnZeIvt/G5pfKANxITYvbmngjjd1WXfVMe1W6y
6M45/Y3wyC59igDfz2wAyDY0fN/CUOquzPfVaU765DOG4ma204UfkWd/qd0nLdaI
TcqXxYYIQZmHlo6RTw962MifgVCqP3ziJ6Gb0D0cTL7Hr4O66bH79hBDLobkjrJU
vi/+l/bw8m/eUWCwYW0d9rK3CTXofRzcmOvrz3yp97+mZDUFil/GZHL4I1U0gyL9
6H9YrRGT0ON0lw66M135WvWwnqI0FAhxPK8Rbz8/Sl1OuH3ewPMl2e1OtDSjOlZh
azHN/4ecr5MF0eM17oh5vZlFMj7jQ9gdcVvRK2kP7K2AG2n4UE3bKaA9r+fha/0Q
rOurcqqno8LGuCGAdRAMhtAjjUKNT5bPLoy/NW/s0e0nhIwn6MVzO+6scZ7M6FUp
N7DZldCsYVfgWt5Ehoc0q6QyOM7Prt9+DNQ9XodWGmStPWWtN5Z2vS+W52F2nSZ6
/marPBa8FZZ7qL5tRIiDoFvxNqHmt6bFIMxJcPri6OV7M6bCbo8YmdCXSYLZJ2KA
KF37BM2dMuf9Rw2SavQXNMA5f0RW8BqODK9jwv2DAFLTXeKLGnHntnhaRGbM0yGn
QdhExwJ+CPCho5d4pQEZRA4tHyDvBoaYTnahhjlcIg3BjOe1YIMwDbaqVRf+x7gq
EaMc5r8cSoWDkPssa0n8cZmJ8/r8qU1Z1CMFGHfpXPQ7v8EVp7fEJZk9jjCkUyyU
0R7WO4ooz+XYPfhN2DL1eo2gRC6926Qla/fU/tYwGg2N+F/35BjrxpdCvGXypv2X
Jv8GLLlsIsfdgGLBGb0z/smjgUMLV8mW/NDWEtJx5TZreZoxaL3Wxa5L095QZy4P
k/9Gi4nszm1oNhO9kdAFm5PFfbvHETG0kVMe5dxA2THPk4d0fhiAmRgkJVyAaW8C
WxzaRHBW+Qq61xFaNe6xgrkAI4WfKpk1gG/f64Vyg5aVpSlP8BoQPcEtsC9SukhG
+KOgl/tzXysHqthb6vQbq6e4NNCiL6ATy1EtM3NNyxbuLPhqZLUf9/S7CrMaOjLB
uDXSH8b3FTYCv4qwHFuo70B3LDyGygJ3zK/ChOzIfRvhVV9EbqB5awbUSiUhNIO0
fnX8umCf22JWTJeUd+brFNbXoqDaJUwri1lKEU1zzsEhXi/eGoiZS5V8uhMMRKq8
RU9ML9vWyvwQwPolc8xnhkK/Qi2flnmTi6ls3MFtMn7qlDqGdJHcZ0aRb1CZ4M1V
ozxLz7eaPa+Fvwd5h7/zU+njqWTvm6ldT2mF0+7y8ba8FzPhS5/MyLWEDovbpq7S
qKZje1TVNaEFvm6KemKq4Zh+i0Rnn09jQBo+Fuo0okSPmHVmdi+ycChUjeSgLU2L
7ZbiIfLAc7bWcvm1U2PoxAbztFzT1PG/452FoGNb+UoEGqnzY4iCRYWsa6n69mwn
wE7qn/diLy6d4PIJaZI6oYl5aWe/QQJhwQEySpp1HU8hx3qyVrcjN8mbis9UEHRe
eu8epXgjKrf7XC3CaOTFtwLU+luLvVCzpqaFe0LdQvtfBmkY1H9iCo3VN6pdTEK/
zLEjppCLv+FMmkIJV8qDb+m67Ae64WitIRZrNFV3woz2/PEtZ9q9jNxNZOPrZ2PJ
1ym+w3EJzAEkF67ZiPvCKXeHwaqcnEJY5vGkTo0++JP/UcNtISxNeHoHhybYmHSu
AFvVAwdZkfo1AZr4tYZuPLzbhIbW8eyhX1oblPR798VfBK2j93/hvnPyxKj1tbGw
3Y+dVhHqDj0OI+noXpMyOAhwXyBGF/FYd/uYej/nDSnfzq9WfBVA1iOjl4IrIt3S
Kbels+XUbvwNcNo4JhtwwM4ZaSEUKBa9G28vjHXrnYAiSIH2kAUsHbU7maoBPXoz
AuGuN59KYRVh1NkUwuJhwxrTQvbizQmQ90OPaY7JGi4px2av+yKkQak+bvLsVjaA
bqNMoOjr8B8D8EbppXFnFw2al0F4NUdYXakiX3Mq0eiCKlfG2L6p36m9EOhry0eV
yLbMSWRSmuPehuy9MRUU8/tz43hgrGDMv6BpyoOfATfgXxHZLwANx0vxE1oqm4yP
tv8TDMrtdiBqOOxu6C3Yho1glzFcdTtGQstgecCWJEDEPTW1NjRUc93NoFtvrz3L
5OlzFjL5ITZj2cxdA6/3B4Z15rVW2IHvbmrtvLLfs+tg7YP86JaFs56tiN50mExA
zDWvWlGr1uay1F9HM88XsA5WvUep4ldJkmpKmzqtoC23DmPN5qV6H246vDT7zh/f
1qspkFuRHKNfoAYB8NcmXqG/NlLGqqMPEBMsdRdX8u6N9biWy2YbTkKMInrQWZpx
iQXvsfGoV5jW/v8wAPuCdoCMtXEQMBVXrJoZhEAr8gEmxH3iYVATQwOEZceEqQlg
ibMDVE8ZzSceHleOaTsl4cUxWrId5Ghntnn2BHrgKd8a7OINIV+jLL0UbYEj5okg
CWnXPrVFZqqrxqxb/xmZlPrtVM650FQHjwuGDyjBG2bmtSfCCLFQaJiWc/mnR3Ow
79AeToua9pDpGFZllqtNeDhYegehIbvxOIbkB05wuWWIvWtmKzT5hwXgKH6CQvaI
bsMr9IN5EDNzJrDCvxTMJbzEPdu6kuxm62OyrEriJP9m3SiQ4ZdyS51iRtA+jkNb
rtBNR9TXDWq5krLfu+stJ5N1pwC7aTF2+ZFU1vkWG67kfkdHLWiZ1b3NBCbvgqzz
cd196EbpHFEqBvO4/tgdGJY5E3ANmJyyVlWLlMAmCnkAe9V1vGhhO1/s1lod+cYB
8OIZlG9kknKTTN5zN/PRWAdnWgc8127HicbGWQsvlm9zowfQO0AKwVSbMC8LqsGo
0RtSO3RwMIZFcqehQJm2NGd+6rV2Br/+1P0B40tAw7Wz+sbfJfbJEPhomG8XM818
z8xJh93wLLBm45YzscbRZaDGHZw25+hEYprdxpsm6NQwqEvzvfQyXyb8zSt7Xapu
CMwr0+JBdi7Z58YWqNISBaeWHMDFmC4aTKGkdpSDK6SWmTjwzYLng02AEb7r2q3l
BYZ7fJq0P4YH5NUMaDEAxC1PPS2uS+NoW8wdEqhZUjItfUiEC/+DYVj4s0kdrKCY
NVXUaolsX7iLyvdbKAFKE/if8/82t5NJYBLAUBODQOvlGH0hMq08+A5JFd/xEU2k
My35g+5frYteL6S08eIIeMQMjcMC5cWiaiKqPrCoC2U3JqExINDX/csg3ULrHCZy
/lIBa7BxnJWC5gtveI1hVTRjZG9w7LnEMxqPzv9KEYPm8LwtEHtAZ3wm33sbyG1G
BAtmyR4GViPhlT4W0eMTbLNGahvCKYSl3cp07AUlAJpHVGXzoOvejxzfdKRi/2gZ
r3PaeDcZn6LYBBR4dkr5cuYDtBvzRlVL5E22QTfQnWEsLlJ5TvB0tV4FaDCGJ2pt
gD5tVejLxrUlufeHXpLesfWrjAKRmsTKzh2ehmPm/vnnL7A5aag3JrY05NdZcc3i
hQG4RFs+21SuzSLJF4yx2df9xt+dCQx3C8P4t/QkuTgTW6IU007JBe59mwgaddyb
lHbqc+vBt1Z7gu+zHiljSDWJm1co+xI9FiQZVxvHCfFVY5+LGTVgmmx/rhsU8nMz
/X8pM/MydEp7Pg6lU+YwlPC/gz47Q89oEqomtD0yKa/GyBaLqYGmQ6e4OZ9Qj4vJ
0hMMfukvr+VNOOqsV5oWj6xKrYHbm/FpTLsJyUZ4IFBGuWTMoHH4xGw85VUoH59G
B5sD6LAvYI1JjkPtBHU1SoWRYbWA/gc9/xNiYITTBPZDrXZI3LE7HEQ5u2CGI7ml
qu42q7BTjO0slkL1lcw+VrBwEHo2HYP1Oi09+TkRzqbZmlLHszGzsbj4iMVQzOSl
N1q+MjJi7mU0yWu6cSh0eyfnoYP9pCYYhNAClNGl3Ud8katO2hOViYbWyrO/HaOQ
rifx3+5k03MGtAjJJovTOeum3CeZSIubFPYv716Y4cGrjbobVQT9EITIIuMnotPM
qy0iII0g5eBtqQEEGAvB+ytt3oHTmwY1hGMTJyP5foEo1ssmmUkjL4ZtA3Q/U0fV
J//ZLoEdsp3D9K7/TyANtuIKHzjiYYaOPLvNv+O5WhM=
`protect END_PROTECTED