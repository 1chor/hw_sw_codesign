-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xzqyJ+0C8iygetvnHx92YYXbodrl7i1eEup4zh1y3NglKY6v6hVHIJkdE1hHyhfbESGcjyTc6q4j
81vtbUAMVMx36WD11JLIl/RPDrJm6BsGPk38uOZzX4ElhP/k763XH9GOt1FdNrXRQuFfqpaDMxZu
UovNOiahboIE7fNrqCv3ktqqPR4uAZxr/TpxzPrljx7pK51yAEcbH5RvThj3sp+cccjvm9um4k6M
bOj6C//10GqfIsu9GmPpNJytg47fSw2hfMkzminYLtsQuMusObLrfkSCvGkM2fglimDysxKW+XUh
u9+ycmF05HsMj5ThjW2Hg9IDO4PHGl42SOfPaw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 89280)
`protect data_block
wbzrf5oWyHc0EjnbrOYfc5fa8RNHJ+tsOXBHpNvbocy14imYI5hPBLTYnVFYL0xm8J2xSdzGrG/X
l4q3hx4DeEdVG19Nberfgpwji5nD/Gc5Ti9GS3W/K41oHEoGTLFaHND7TClnS3Jb/dHdfCSvBT8a
80h0qlynzHnSw4DtU1HozuhBZvgDtH/cSlzvXIdWXZuVnTGHgyZsh0esGeqo8CPEfjVB4yIHzxCZ
d7u/kGWEL8aZ6M9QBSyoEqGyyQq6SR8C95rzMyVEt6ViRdcnpD+ZGqd05WQu+GaMXC76Et9wJVF/
EnUPLNvlCaAhKIhEe3hpNf6HJT6Ukg2daaWTPLHI+VehgGIZ/BMkiFl5Cy68pH+FlY5G15wv9a/0
4xN2JxclRII7ZRd3JYw536+lqEiBAed7Pg+NKID23OWXaiJI4T0FtD8woqi3kiaqVpLW/gia3L9v
a15cu7Ufxk2QJsyB18N1DceGhOibQAF3iTEWg3IcA8alJzBovGK8hwuIMm3xJEUXDjzWI3aC0H11
5rWck8mmZF8DJJk6ZmZpNrNHOlWt+xcLmYGEA9TyEhCy97t1MTcyA942qbO/+etVXr/EkOjXRQcd
UOaFRCMF/Li1Za9rq1ZCpAXV7hzA4nE8bnmkT2klDFSaIPLA5uM8s5swWP2DfLhDgTIoqQ4+84e9
Ng8aOQugGyrJ+2yxiXMgc+P8bJKkhVlpAy/G7IamY9ndHd6na1pR2HyzOUx7m0mrzoQii/iYJRkz
6p4q2/wlpeCwgJePwb0PzyKaNBUjjVKkL2gcujcqvefF5sYILhlYuXAgCesVdZoom2f6vTSykZQU
1dmDyA3Rqg0At3FZSm6qGFxniNMT0a2tlRRxZRsAcdWHC/MFXkiwZ8Pl5fDhabV63qgOtAnX4wXG
KxGBCi8XiLZIZt9mKqyarEYxTPJ39nyKwtdMME65RXA/WHEUEUTLV2XncjSvCfD4THxe5L9Nn9XC
FxFpSpT+gwafhJXdCvCKJFvNe85C4pC537/OpLevOBDx4Dn8AcM5sCO3DfvEhg2R3nPYTvQThrdf
wsfxjJTZOlDw4mgKNgzVWwlPBAKJy+dRats+XkE5NdSxWDevqkhOXnZUGl3VR/yKc73e6u5ESpuE
d/s5c4f5ASoKBBUpIjJLyTnhP9HiYohkiP+BZLiLqR0g6+LR8w0p00HSaUZ4oAlK9y11yUMiKgmx
jzir4TqxHXH6QbwXBBFkPOEaqDRAckcIRohAwFL+Lkxxmk7/hxG8Lb+GdqSZ3AYWnj8C+dfFZUdq
RkJsttk2wXQKuD/u8qOwsfgy50AmfKSX5J6tqCOkSIdscZI1h7bL2E+T+yWvwYUUEErBeb1a9TyZ
7HJvCOYVGUT6YbGW4lC3LL3IBz1Uj5i1cse2E1IwAAYyS9uBtBe1vrfCrB7pswvfE5takphxGJKU
RznrpKIHgmUUwmwhnJJVsr08LNei5AFbgNdG7mkNAxITwNb8aX/E3nXeQIy1NSg+6rlDF1gtZRHR
RZX1cYibwCqwPLRzlpFnWJ5c6WnJhzSS7paFPQurMh1TF21PLeNNO9eye0kZDKc0IoV+H4eqNw0o
aiWh+k9a7T/XANfpnULu2Z5yTix/CxVVCmV4ivTNWWWP8gEvxutl34Frl5QcsyBOtup6GrrgBIze
EdZ89zJgXeQalw5eli1cjeB4BOK7plsBzFBqwM31vUoOg70YL6Z4dkaj+2yMAdDIEVlCeXH/uQ6Q
CL5imZMNiO6ukwbuKhWNXVJwwHYxYTwBVI7tEBV4mGyr7su29iO6xLTYxrymbfamKgjAvJ2/WWsn
5iCtFeuCFlAtGxBwYLUicaR7IMJhLI7+GpcOdnrNhcY4FM06DcmyM4dt8xMJluFHlW1NOj14hhCn
kZS7gAPODmK/dpLqrgxx5tlAMgYWX0vqIBwTXe7p1vvxAm9mkdJ0Rf0NFSVwmjXOwrBpfqrHZnZT
mnuyKEBn4bbCPNb5Cps5qbLXUCjdvZuxeqwqWXUycfB2AmrbaAQUHdzkZj2ray6MrLI4Le8clueE
ouVjTENmeFPNGD6jrnYLFPke0hJ3rFA1UIhlvkQYshVI4IivIy0Dk2EeWL4KXk5IyhQUMw80nFnr
gY8CL1Xk+kbh2K2vGiZtiwsFFbqyymfODEjaxipUQgWme7D8t210FOqWJ14RnHe2DH//KnF7+J+7
ULQ/PkjZ+1S2tnhFfv4txLA2nLv0GKkyo+gAmDszzDED5XCKvMULbDWbdV/1VZu0SGHxf4FOR+s2
SZ0G+iBT9xizoQ8WNzR9pt6kYO2TlM8Lpf9JV/PVTlDnKsr5hc/XKMllJLwwxKrlosOqVGG9dv4A
Bc92s2zSx19yiz4Y6MtPwMDs/TJa0eXeziz5+S70PHxJvu2hJ6Ir3XN5x3BttCh9eMevb5J6Xa0Y
9lCdQTXqS4s0IKkQ6qVLGRd4zmRi8weRoeCQO8X+9IFRH/yEw8DUTc3/8IU9a27irsx342eTOOEu
hkN+k9/1B+AyqcKzgqXmaVnhAguz7kn1cbqHauznctf9EAGNw4Wid5uyhyoDFZo98HW4g9iyBuO+
Ib61yZciPAaFDqDjbOPt7Iswky3vuADTHmbebhk/atVKXCi3E2ENvPHwCKMqb8wsJ8lEGunBamIa
JqgHqYi2LlqSniVgANQpsUnzvwzmkoKGOCS+t5KjsKrLIdgX2ertoL4UXZFU+Kyoi0cij/2RobMH
Hkt0PkXl3xhVpdYYUgODeCsmYtWreR4HiWSsFxg4GPBpp9G/8zSK2wIZ0lrBr/eF/T7U+XpOjNte
8ZtHSbPajA6zeQohUzU9CvC3Llku7feGH6DSTmZmcbSkZziJMH8LM5PRmiK0P2+hQ6ohdP/d6Oq3
+mIW72xD8xaui65JskoxEORmKlj9AKAiIidIHebE1rDYV+yOV8eUsiIvUpNP5C19KrbLq9qo7nsk
8qfQJHh9HCMV6b+l9LDqv9i4e7vH1lzTxtHYptq9QzfoGlSr2CRfVzGg3rOLxcllsEJBVjDSjsa2
+hy/rC6EE4/JFCxAhaO+oX6Qe/j5rvpqjaG+aucD5BuqVu7LRzdTYgRTkgrnjTiQZBzAF0tO2r2w
+Xe+tSjCjz3Ja9Gr2Bi0nB5Qv/8v9UKbMm+SlT6BDDN1hzZTBdomDw51UE2dqNynEAI6EWxJfaVz
2FAj/x8JqoUCKCJ+H00ZLlsx6VDC1g3mD1VB6qlMro5U8YVTUZW5iXl8yT/7cM/4GyLLKuWlfuo2
cc19uUfQjvbqz2GibJCcmBBtE7al0NpTD+iOnNz+ZFDOBA0oVV19uKYBbLG5KyFv6a44RhmMmbbp
8mv9R78b7cfwpneftaMm3lhcEJhKvw9X/LXf9l5Pip2JUXbyJN99ccPp4LsY8ckITj9s2FFydMNH
7T/N0iiMSCkt9NQPM9AQvIL4XXYPoxzPFuLAUQtsrhXUjJ2u5N5xGujLy5dEcbv9FMiVhLYEpGMx
SZdq69DsxCt5Dqkg4Kt+DrjMi2jr8GrNwSzHz+lSJH6HWCnC/X9KcWY5A/njVMnkuaVkNofqCPxW
Qo9gkat94gPAQApJxJ13Y8W6eouxhYjIgZRZr0fZFEB2RNc57wHR8GXDgEPRAM1qWaV5xIede0Uh
lboQQb/5ZR/oqEX+h+fW8TmFPmr+M8un5wtyRYq84K+IyUkMjP2EfMRSzYntu4hpyUJ+y5TNj7ox
hhu2QeELqj0IPbqGAs60IcTKbdrXsqcCZa7twzQTOekP0fNgQV2cfjh1DckOEGhcKgYH+0jnUYKK
I7/RPdcyZYe3YWCzJZJxQRnNW+dO16uHx/zHYKg80jkZyIyPkg37L7XN/6TnskucLmH0CKD6B/GM
pNp8NwwxLY14xfcFmrQ3IrmPdZ38Ejz5qxkdGjNK/ot7dAtcEkAaAkwao1Q+HmLeeBU+HkGVcV/a
R0Vk+FS75XUg1HJVmgDFXQfxH26Dh5QfouBenDR+oS5/zmRkIz4jqzo6FaykNo7C71n7RHPvjpqF
Xwy5enrvZ5RK7D8Zz0GYBwiHSoUSBrhqc7IGS/KuBNNEdcG4i1VCkiKKoBoEMPzGB6vCzsxkZhso
bclMmtU21j5R0WMGasey3alEZzlR5llZO73SfmAJFGGNeB8hxHiE1uqgs7MTHZ0Nxv/fYW1FwJY8
cbGVg+EBSSWsclwzQmZeWze+zIPndWPRTxCJWVogdTMIfJZ2fLSAR6ivzKTnhK9ysgcPsNdXRW56
NQ4qHm8PG20yfpYU+E8d/Ov7sNl/AN2LkozbhMWYQ23bxIW6eH6HX/7TO474XMGt5GUd2KxN5akw
NkExCbaqWmyMjmY+zKEfFhQm4TzEzCuol8ks65Ay+PvoXx7KMpscWXlSyN2b2+w/UbuiZ1KzVyHd
ciVoCx8hw2L4lBcqBcRt9v8AAvmPUNMjquVAfh4RNnTjbNHi2iv5w7FHgevJ1BH1v04a771hZNdS
zDcn/ZUHyHi2MHYBGBNNsvGzfNWvUaMKw0dQJy5k159NPW7YJZTy/8iDpLdhNfwz/s/xzl/UE1DU
rtLVmqDCuvwIq3g0kIxTqe5SKfMDX4lsMHcjkRDLNyfjXSOFO0punATbIQiKFmMgZ2DAbVLDQ3XH
rC7PUUqYE1xRwvHEy5v5YK3iGMtpyElTzCXm9VSeMz4KydR3Nsvm0oZdIux4NTM0RnBBXe3WfjAa
YutS+TEN57Bc1bj8TusY2FuiQPUhrnYHNsR29z4uAHcttJAR8kvb2t0wSEmgssmym7DsDcgOoaR6
3GWZzaU3NYCzcXaLRAkEYo7h7qDD3VwQWiuWSlO2vnOBvYDqN+gwcHB+SKEC4oe63FfalHFudMYb
Bq6hMVI6XK/BNk3pf2Be8vOZLdTjydjy3GBXW5CyJ6JE6JuKr9s6MJjshqWMASGxBmQnomWLO1Xo
lyX6XHxbHK0zzskNseyFoRdFNNg7R3nLah3fDvZ9W2fB28IZJuxFwrZkOAflK9lsG89TF+idpsMB
tk0uy0Krl13SPFMjIaZ0l4OCui5dD8jBwySGaZbbW4jZvwHhHf6qjq0/WdRy1XMHXj43+ZIAqBCY
Mfvbwtz2kCCgVopMOsVUolR0Dq7YkBTVPtTJhH7U0ul84huV3gh4gofdFwhBWgOBSAYk79ov+UQb
VFn8zKQ4WOZLeM/YYkE31DLobFRDHbj3zFeIxv3M0f5SKIHCSepR8xlbOK2hptGeXoSJ5bJfA0HM
PwmkJZZZEujdZBBxKbJLG/RMU192NTQYHaD1Vqr0pE2BJjRmCgWq1SULm8NR3NcDfDa1OvxkuNhm
WFC8CpflEyLk4q2Ic45OMYUDsZffmQLAkitRazE7/HkBrBgf4Z49SfE8sQDUwM0GSzeA1EjLL8Gt
dvY8fD6Q6j/rm8KI9bDI5Sw1a/tOOrVFLXdKZs+by4T44/CzwWys9Cu8dyqP+D7RN7gcOJy8pTra
X5v1xyP6E6NTryC+BZ5NSxsdz4G7l0jKZrLu/18ETh970U6i8EwcvIbljdUkSyzXBXEAqURK3L7C
2hU710uSnKuePuzLsA1FpyxUYU2UcT+Pizj5+vwyzdh4llN2HX9kDAJypkPnvSGn3DPUPYfUHohB
1SlhszT3bgf8puLll+zFzBHAZhLwk5ZInW8Jxv0jmfAMK1Ugmga61BAUiMvnuvdvj0D4ebBFj//a
zNLF8HdTumxitTH+Y3vUmUMchml+ZcPDq+N0Ni1PpW1GycuQKDHRqFQtNJsc/IKbMf9rpYSfkNf1
OCmqDxszTUvFeNNxBPw+YszIZhxPWHPFuxYGTr/48VbQ8bXPmtWqJplav3rp3gu4XBVcRfp0HSpg
pmO1BnKafbkIp2vFog8HSeoAM+peA7tM+0Z8rkXNYo4C1C1puPB6d9EkUULpFH7fw2MmNcOOAQaT
E7NTSqN918gWCAIubFACMQrZPHAyoHkKa/+Me8hO5ISTWRfa1Q2gF26cW6cp3Pf/6IwAXuFrfSS2
+gdDY+gw2YiEvWTPxSc4GO/95VAffTYHv595wPbm3DlfJanFlzAObHio3VMCkDyU0IfirzVWq253
kA8rqsNbTqNRUEKqCyCcm39YmiDaJAHKwZgdZ2OcQf0HPfa3G4hr29Yf+btjF/uPKJTNCvjtxIHV
ZR55G58lTrYT8k3z3fvvNG4BhsWnD8cO0tQNlIYBzv/U+kr2QNFGF4D6sIGrtELvdymylsib149b
2zrQ1Jc82aeL+2hIFzgrZxjXaHU0Ylps52xLVsrkI2DhFEf0GCmXOOIlmVnK3bvl75k4iMI2LEhR
CosoRMYIbsgWNih/ED7pTreNdRAa9/dYINqiDAYf1KfDxHjtWli77qKHF65kv8wW/IWJbLiE621z
J9Yc+0a0ssteoyluFdIo+0Zotv7jOmbe9WiG0gtfmYIYi/ZaiQJQtCx9Pk0F6ZFrycBmCYDc6Uit
/msuX/P85cqMafHKcDc1RzuHFv2fadWc2K2VrtV8Cv+mQIj3tFYRwRFBZsWlG5tP2qHw/vXBBEWN
gcnL1b1FayghiGbuV8EQ0yzUFRIkcybw7QoLb8NhE7G+3V5iZYyjH3/pqWvUul4vzBdYpHHmP1LL
GOFn7lgwDvEDnO562+/0IQktolVTGIABqTmSAmrhMJwuThetpaMnPElyshOE1X8aaPcJA+2cVMUO
pdLhpvx5O5uOknlH3zZD7x1NOATsq+j3x3W4F4UfcWOvphayv0p1HIPYKOgJTyNDN3RtKb+3O87f
U5RsO1VrQRzBDT6h6VCvYB08WQWJSLbaf7xVdGtv7AV0MNNxpLsLBO9mfA9k8yrfqh++gwRASM8T
PWJT6mi0fzz5TZ/oGWueyRmFqhH4fBrL/jjH6YYAI5l1yYU9aPnBXGtpkc/NsqK62n0/KFUAmIqZ
lhbs95V1iGJhCTqrrSF2G3JouquHcP0DeXfX9V0DVQCLklx/mwLi/wrP9T5vAOp+3kuxq5l183cW
qPduFeskiNcs/1bS8Nw0MLWwR+ZhPFI+tnd66ib3mchQFT+pNNGxB9huswTNvoM9YnKykwvErKpG
78h7BBbWXlTE2kFM5Pem7+pn11wHIE9EuvBaw081l/et9KD0Q0eF9wDk1/5ttdzxCbFtReLzOdqr
T1Z0RCHAkcosj1iaQQNUKXBdSc1MBN4JScZj9oN3FmG0XT/hsq4TPX6jC3mqZxQoCYbuWaRxx75m
XCGwc3TpLYrIBgnv0oNpKeYsAtM+UU3rHWz5gDNFfm9haYgnVMJGZddpClaPF7CjyvmV0FgHQ33/
cX1u0gipk+zl7tVRn1p4nx84IuyUHsD94vEdOT1l7JqRLrqE/FbDzZhSOxntXiA3k9F01bs6Qs3D
FxgoXXawYP/ts5YsMfEq6jU+okrfzHUiv0ndB/bPFzc1EW2jkO9FcDzpC4mD1UKS2MXLVWYK6+O3
T/6PAVRnzV37hBCYGan3rltJO9yFz/D+pbjU67fMHVcM42EO9AIke1hf8vrv695gT4exQTciGilJ
tvaOBOdmi/Ffl+SRFxeOWQGmQEIDNsatoXzgTq6CkfrYIHTGHMux1fi8g67z9+p4MAj2VFsaXFVQ
pnj43ndoFBTOS+JbwuhibpM/su7aRvCvaJN6FziOn+t4q8sa41HDdbNgpixl9PKsxA2oz1ehEWJN
tbP41s1tMj+C91aax1Tf9l8EZxm/C8d2SPEhlg+9llYzviev032YTNlNqGFPnZ1ZSqNlYTC+fz5i
KUYMbxCCCV0wH7zl7TH8r5B8ftxiMWX56ku2GxGpJgwxqCqNokZ1FALo2cnkC5UIwZbJElNxs1+d
UWkm8jUmbkn3ZHYU3VcSufTZLVBouIcfeVjdjjtD2hTgMkhbt5uDet9BR+rJr49FSqm0Mr7QCx7p
JtU7DlG6wAyYSBRAtanFqFTJLT70ZTD4BQeEIS9w6mU50E8qGX/fKEHEZAE2Gpzz4Ua/6OqAtARd
IMX9J/0/1XUwILGsbFoX5zVDTn+pY1fFPJOLz/uMqcMGhcIIPS0Z9Lo/yH4c82fmlnalhgLdvxrV
dKtgYM9HER7ygqUL7wplnNWw7ZpaZw0iBgku5r4wA1tY1Mlb7xDOIWRGHvidsnAhsd8huXwZlttd
RY5tzTqhC1sRLwPsx2UEBaSbdtbOZFJoFWVOVKhjEcXfNqMwB+o+lzjiSQsYeDVu9TdyTzJu/JFL
KCgWt6iyuYc67dAtnNEhJoQUjcVHEJjiAGBSf11Uy0CKmxOM1JPeKLwSVVh3x6ULI64GlXxn/XnX
qwIY/75UrlE94/is47v6JWMjfVzfeu4MYLWA27lYt9wJfJV9g+2cNuwKfs3sxwp6AaYysIknLG2R
f1pS7bwTJd3O/iIk+oULku0VBtdGvmIWNFoXVGet9ep8zAm5UpvyF2O2UFQEO11tji8kimYoijvs
W5hw4fX/2HqD4mYxbDy7U74hdpvD4bJLRAAuEjAvjzV/Na40Rf/qykNbO7aGFgWutbvI65NMUG++
8iBLhB9Squdw+/9/6tA3VDS7b7pmHx65+DO5SWRlEY4VuvUzh36xx0oeSXP02BSuhLLkFD7ovFaI
PwiNsDnhDTE7QjmGWn1TDqWRl6mmZQrwzc+ahYor+V73PBnUPZz/jfjy2NuWELvCwGdCmcTGoRfo
Iv6YWggsqoLCyTl2QBzwJZdAjkZYSCxjb+6ZjfwBWYBRI8O+PmWG6YtpNmx4YBg7E4wY5nCmbIz/
KtJECek8PyztD4We/N/ExZjkHbRW2viVFjn83GRExbEbAsO28fNeaKEsVGbmWbKdn4vQpMTNRdZv
5ytyFFsfQ8OaGeDTa387kFYW6mZTXzk25Grb2LJ4jGHZKBBkmS+Wxv6lknOPBPW9qYpk2NchB3kA
ibUdawdPDaitkL86Q2zxA2vaKbnuq/wkmb+qBZg3pg9tlzCwPwWX9dTlnCHY5UG0HkO/7BGfB/Rj
NJXjBQwWtoqKMlS4z7AlSRljzetaT2vtnaHm3p5tFZUrXwXWOG2ZU72DtCDn1S7AJvWmzpH6dpHC
w5JznXE80PwmH4TAssV+RuUvBrwIYg3Sxs81D3gmvmeTMvAPlCg5GQYOGPNAnLDSloZdHaHBD9Xy
CIMLBlC+yRnMjOlFR1jTKnw3GIaHy4HwGp7AT+xP3ezrc58XdqFtkQW+Horgf/dAbAROR1l0s6sE
k19VS3Lea4u6lxxD8tgaiCTAgOs07rMGi39K/qOmxsUxu3LN8zHGz/kL7DQngAFbWd+eJr3ZNaui
tlnLetYf3IjPtTsBTIfhUs+bcg0RWxfIutsJ3Fgek1QTWJCFNCoqjz0VocR6wTODe5gPztYfUVfW
UEWUEevzycC43krJhRuRJWgaeEZGHGpYXZVk2jQEJ3KF822QJY//+kBHb1421CopuhZAYd4IWKEk
/Y3SKiRzXvri34AvIKqVh6L8NdHoipPE0+/VfTekdpaOrfkACk+znnlkxjKg0/+qKyLw8HHJmDgO
iE5PGfaEbCgJHkdX6sSkf3JMt746Dy+by+M7SLbRXt6lDnpfM69kVOaMg++67vTl9A8mi14em4XH
5bdvyr+y0/9A9/dFEZO/4pIGZMv/j+GMLDACra9Fngbo1ljikZFHiOvhesZc3spT5gZ7TNxAg0v8
Pv4wEBRcVM4bkKiohu+yYTZcShQsUaf/J7spjLjtzvKsYiYZErefyO+XGFg47icKOg6R7BYRYut6
e7nFZOz5iuly9SU9DwBLiYGssHVwADyruD/O3Bd/7gSFlz0lbGiteeZ17OyJEKjClLEvWEJ3cQen
2Amgj1lfC+Vua4NVx9bqSJx++jC/g8g8NOAoQCU3Dcu7DImMDZm5vHY+/ZyktPSgDTj572ZO/2B+
Zt89M0rb+GE+1qj4ZXIlXFdS9cmNa6ztb/6iqnDMQFGjWqw0ypVKk/5tzgKUuMWbFvu8F3WOzTGA
rV8d0f5iTFQvcWs1J6p3HJG+4RbxwGrnvCarjRMZ175Y4Y6fB3iC+ykpHg82mr1qHKHqCgt7I1zU
RMD8ojiijjSVH5ZgbS/+pavrytIuQWiyUuyXFt3bmvqMxbHd7XbZZlV1WpWX7eNGedtLo/0Nr3CF
1oVGsWnY6zsnTs+AzTzP2xdFNNnKE67t2O2GUgrgyYzxJaVj0P5+DWgS+nm02gcVnybFM7C2+VFQ
I5K+w7/DBW7igRtLW0tSXQFDV95KtZV+ux6CvwcJqpRLjZ+GOPhoffjiNXFXKJffuVfDI+M0a0qf
piKi/qOn1j0Kri3fVwapybtXYC4X/Tywix8gJAa6iiq0ruiCxzIj4zcVAjgBIMrqrUxOuxIi5eQV
t1Br2KahI/YeyOcPhndkXS/Ws65gslzaRYNtAlQFmhS84RgvjAoF6CSi85BVDFP7OU449N7chQFV
3+bvjap4tHEKsBgFle8Ui45IOYDKTWlK3IwFVTQxsQaDcBLhl4gLzLurYXFeZnngrvAUqKpUGesn
XwcaRBrcrjIqdqm3mNrVCo7P4XxukprrC600SaF+zQHnWvb0uw5TkL6R6ch2K/JOEebeZswLt2rL
0hgJBePa+2+LOepchEs/QGafBkdNB8Audg+bZGOQHVd7Koj4NnboY26+UvJJDiJ08vm7/RG3XJk5
pWlulP7HITLTK+gL6nvXTipFWoi1SYsdKt73Uzx7TQ6gRaYZh0i4E8CqYbnf2nBc+6b89YUMuIp3
bJDd6XadutIyu3WWswKYkbiWh/vwU7TP/OcV662jrlvsOm1ORbY0N50QZuo7bVwZMo6E5j46anz1
H4K3L2rMFW8K3LU+Z/YL7Hz2qdEm1Okg+Ds2QBEh74gPpuKoMC/oCHkjVMJQ6PhZSP0aqObgiiVE
0fuyNeEuszyVAAtpSqZxnAqykxw78m//iMNr7He4I4FM86VBT1uQQyF3nNhoTW4HOqDPDiX8QEB1
Nze6xWkdi5TlicldIgCf4G6/6Ln5SKgZVvUPmcrLM1P3mxLfJk0kCTptgz/KHk2W4VnckKu925uO
vmn8RkBSvoC+UGABs0Xlkp715NNDbe588y4dDxd9++rOJ+kcaaSh6jyzUpMi7vQg2q1FDmeRFaiL
ledyUrldW8CAde5oIWBUzGfuGjYcQ5JwuX6tLPqIGwg6wrpO3L+F4fm2fEUYFjtJB8Q0OnBUsqU8
Ccjl3yYNf18re8se+7QI8EwARPW6yNZI6HIVkXHPhx60X5srZBeKJKdQTG72JBBOwWX5AcqVeDJo
vI0ZAkHsk7y3MmtZ0DRiYIfLh7AABLVBuSMKmBVaePy5cRpQP5eGD7f4DRWJR0UGBldM9HH3ZXCr
nW91ztnUUXqc9gUIyOny4vB9J2RLoZWxA9MQLv9cnnfD3o18VzkQq5gLHdNO50h0bSb7MAECgTiX
Bznb043zRvYn2sZnox0DWelTq4q57zvMPLMusRNAoJkqd08ATjWFM7jALcMQ9O1MFAAUkViejXcn
lZ6+Us3c3fELTuwCRpMM3U6e1fZjgP1IdZ0KDMxiq2n0KpzRfsWdgmxVA23wdnR3cKrv+21PHxZA
q7VGYNkf6WddSbHcq3EFAQh3IhZ8tvC9RbAcOpQoCiLjh8i3sx+MgfU3jXTImn6/7n8Kmo3Ls/f5
2TMAo7o8NGo+XOPEZXsau3gNLsyqFLIK/2wCgcZTOE3WEzBI0MpQni1S8gbeUA0tmd8Sae1Rmt4r
rAEs1/p91jmBpAHtHZH3jdjfyG8Vsy8rCH53o6LlyDU551RhYOS3F0ld139TcLa4SDio5zFO64b1
CsEGlKoQGnGyKl/6RMUN48wBjg2Ych+2OX6LhKzewoUr0XrJts7F8BhvbaIJHlzNXPcufkSUQ5VS
0CFyNAN9Pq7s3scZaqLvBvCZN9Sk+iw1KMJxNNYG81o/0hf38p+ak4xl1K1p9heaHeTIu9nEwuNg
imvCVyM2dhGkMWcNS2nFsB2nrQGv9IbPbzLNYm7MFwV28CPKkCOvJPiiXWNUYMsmKPZsuM68dkFR
V1CuSNv1P2GI6JhUfCDOUAN6YrXiSLqISSxloXf0X9gCJAMzkuU+sAnJUfs8u248guA57dtVZlVk
iXl0oOwD4U2i/8960qY+NJdmU9e5gvAK+NFaPooWNnFblhO98uq4UIuJyBlJqMuQP6khZ1//T+Li
yX9Yp2M5fJoiDJ79hYV4UC2mU7ITvPK7b/vMq7L39YKF90fd9D/BSuBIGo2bh304fHN0b5dgFXNi
S658/RRJtaR2PFGddwo2AcpBtRzcqNTzEhxSythP61oXj8w4L+J9jI+xnwF3PlNUsdOe3LsfwHGz
MeP4WpKTNUr+asVMaKHW4C5WJ7UZ8f5VPhz53i6R6upbwHU+SGvjhGn4JavFNtQ1ZtSN5l+HeMX7
BXxxple8H58SqV3EDY3h4MA4E21quPulMrpcL0pqOCFqyC9BerJ+S5RseI5TpDI+kzMw0QiQSdyN
RuEiGXGu239F71RAnH6iM91/3JenfIsXFJEB4W23dV2ZXYfDBqqDIH7H0GrDgUonTdiUVStz+uok
j5rnM104lziBboJI823QL2PzBmaN27+B2asnHb/F5YxonlK8rJmp9agqCm0/aq1Z870g1Hi8tA8c
4TojZMCq8Si20RFjBfq229Ggp7vlWfoOsz+cQFnc4ab5gT+2ttxmFh0RkIaA7zVR7a2VoFgnlk5C
O+uPam1nHcS5RLDTnoYz3w3ozppoKK7JqvhEN1C46kH4oc4D9a17+j5dzlojzN3N4iZTeqd93Fq6
felVxOd2S/1TfqN1VHV36ASLya4fUKxIMFn/d8sMnlIKihn/Hy5Sf36xSc08AV5OAqAXqlGcOO1o
2s8Ux1Bv0sp/0o/hrFiFmH4mUJJ7c1NHqLBLx6HAiBJT1PQK6CYh3D/lpPNDsP+D6yaLLZVae/8j
SghQ8hyJBDfYrSRL33Px9gt8B3utdjbq9iJwkBMJmBuPp5i8Frc+mBxclA3SI1mGfNZ3FJBM/Ixl
Sg8+pfXxr/4B9F41AxpGNVfTabK0C1gITGylt5ahcAcN29U4biUrFH5S7XaDXn3iEz8bUrhImx/Z
y2q7jRwlu7dWrGoihvNdwrjwuY9n/TM3iB3lua7AOJBm52inO61jDKX+T7M7pvp9MTq6wbwyLoRP
sz25Tsym4+qadhgB9EL+4lG2RlnkGDRlCrTMPlocxuagRVqzAkRLfQRH123lQRnrYrprbQxFImJ6
h7cajvcEYaqHVy5XXndcLwDnRGcsU3JFfbK7NuH/EhYjpJjK804VU9SCMSrPdsjS+WPWZoK6pT3e
0+xjAOmhjT0YMy3apUNxwQTo5t9rw4YDvDDhEXm//zLzVWz0GDV0bj42Sxhtq6Pv7v1YqAlHqFvY
75nYH25sVyG9vWhxZIUcNxm8aRverY1RPBzNnZugiSenv2bB3CzbVU/4qAaF5rlxtkMNMQhxNU87
bmEqwpr/1vdf5RK8gaG+ykbaFsDGWey5IrZ0LCiXw7iIR6BurOMmFQunR5KFN7cdFdSV2mPPSMOD
PLWDngdbuA994OVxuWeV2Mkf/NGGczOa30vskUr28j1gqKHsA/3rBd8Rv4I9tjFrBKKCM8+nXjjo
3gNezxpveyY5OC8FGVj3+maPJo9XBsO9bln36EaPNLRh/VGZMlhQay/sRoCgnaaCBcWvPqAyLTla
hM8Pyg6kmCP9TR4womtNG5VOALzvDmD/ifljZPmR+OMmAVfSIiUQtwPJiGwhc10d6Cpnzi7GdOug
S4Y3gpwYAHlWC+O8iPXnHmkkEpQU98NmMxDhpf5Y+Fttc8HDxoYhhRcRqITEB5uuoowsirgU3cwd
tcDSvtIS6N1xYvOe8Omw7EaMYSU1nU5fxMIvYj0P7UQ1N7g4b3iRxsSQa9oYI5dhTpWrIF7TidRb
a/9zUN1lqjbqJtQzFfP5JTAFpt0rsuj1etDQp/Xbo3cXnQU6cYxgHdzalkpUsH26rKqKaZhHMRc2
xJ+BP+5STX6WgrSsRKT9iyR0o/JaQYLmel1ymSPBOuZ6PmuyKr+JXBjLIFGnsZCSv4wuWGNT7jbW
3w0LRnqXU7OPTC7q5YXgNn8VOtfHNks6APAytTHnWqzaMNqp6G91uQRKhj6deqOmJwOaPJRSYjdI
p5jEgRUCaMgSHpeE7g2POm38P6U7R1o5dgNlIq2PAC6T/WDZzpT3EgfqAuOsBeIReKl5KeFi6rHk
GqPQb5t2u59z4LkscL+CIaFlu1ZX+8J87PwDJO9ZAI6ILQz44NZp40GYwaBYz0MdFbe6Qz8xXsaV
UOQnSYrz5ymEEWQtNQN8JbCEiY0b4rYCholemyNcNjL54RZAnSD8BCFFxo41Ph3NgOdVsGqd38XZ
qqG1Hba9fQsBfxYlnhobrTSJF40Tl1kWHw+3WFO6hAYLSauuNABtkp+TD48CiUkmEII22+19lJ9K
oVvTXkdQSEGUhh/ziX/sWVeOoNJItI6S6pbY09fHHpFlg14cHNb5FdQdO8BA/+yUVyK3we6vWUcH
ZmTIUdBQo3XHXWSpYEw+NPNPdSpp61B/px95gSOlvEIRcE2me49dH3EwoiVpabayu2mWt4PE7K1R
eMzBh5S3GqEpviUmFgCyf6lQ15rVNSChHJT2OWNIeHujY7hgdzXzzdg3jWfYIQKsozLWSpvPVBz6
bmlYWjut4snEDlQ9LSD7lvK1Qm1fyAj6XViwLzY6eSCNLutmNB4f8SNlPFdgDyTKsIM+/IpgIfgf
BOTiI9W8jpKu4pmONjUIWQGaT2s4InkuVevSXCNnDDm7sn4ky4Y+b6c2XKik2C2ZlMlQF+IHlzXH
bGgiArCqamY4CmzH+VsRC+09ew5hSwA03nm7mpfUtoClknxLLEZo3xoixjjLBqU3OKyikB6YyEi3
DgIQSmOwhHCJNt7eQzNvg1vj9vyjym/n5MIsilhmpNoaBOfRG1mQYb1kURESIG0dosJrJBE+S8Op
ymrzHA9PEZBkEF5CN/45BLd+hTphX8gAQDKBzoFW+gT42naWMoS90AoxYb5qQD1tDqd/2PjPy2GU
ED/HvSM7RYcJH9MBNVNYZQUtDxdGzMHdhUh95nelCMbNT7geJk9RZEq5QeRftHzwe7ihBnvpNRYa
8LXz4cpne7JL1EiU6zLWeLMpl3or6YKNl2vRSxd28TrvPgJtGAeAeBLctRzaRE3pc2P3Ud+e2CIb
HadQJj5FJNYZw38hjaHZfTMWnG1YJWQquDcs4ysdeDRIDWLPkdhu79r6L+TnAStybyiz9H0npNqR
vncvlk9onliHqOtGs71iG1q0MNTqPyGtHDegJl97e50HavjXiDeraZbJByKkwSSXKJIrv+aQzpQF
sh9mhytWoveNhBPGxw6uKae92Ez/8Oo3o3PFtrYEApN8buMB2cU0EWZJp87YBxfC0U9+a2qDu3TU
uTKZr1E5IOgjZKwOza7PN+5I4bb5zPVylerwyvFmZL7k4JmRHcrEO/SACvnOFTCrxa9sX7H6pitr
FSHWy58ADSOYN00L8dtZ2KhUeaeqXHvbgzVy5V60qN4uVVoadw74jVGMwKUq6dYk8Y/7mPE+H7Or
GMoFR0sIMMP6djnMQWbRLowWY6OTCtRYhpJMO+rjfXJNMMZ/bn2FM9mf4ezQI2NfG7ToWrIsVJZi
kK7mRCLRPTBnQWuQNlk2YnBSp7S2kqEjWu3eTUuz7Z0/RV+cn4nDKItHNJDJMiyUyX1jq+mtjc8v
v5dBiCp/dZtlMUngvf97UV+JKL5Nj6msfZxmwFfnI+DXtbvpG8QPgcNXM3ExZPrSpUxN8dkdaRKO
vnEWRodJXSwbfaCr6oprjZbj0gWLPemzS1VuxpEBpATXVYeg0lVdJB9GczLoObuWv1mt/xeBSuB8
YHM59IEZcVQaz693L04Ql9cbv6+Ii99+28dv0H0JaicwE10LCcODwo4cuFqFb7lrNHPM5DZ1TvhA
5f/f4Klhl1AsWnuCyjjjrsjE+5OniPj47lpHkiSUCVlO361MJpPHKxwyoJ+FXkJod410orTAPnGB
Hf5e4ejNGqGKawf0LG72rP1+73N1cg0lS5rfJQTGcA0GN9abCLP9x1zwn4HtsmIlS572H3v3VluC
lmJx0VJF4NYGC1DjmSRWHi3FG/dgiP2kQPtd4NhpU7kh4O+9tKTYqrrkGLYfwfWSFK9Gqy+yPqRG
QHU8y6AkGx2p9rJ75xGU99xLHaBOEsmJTif46a4RsztOQFs3fmeL/yS6+N3QcMP7NyU4JPUShg/L
TyFQIVOswKglPwXt3ksEaFktc10GZV8LOwe2LaVE/qRfofBxWsDnXFFVUSBs8x9aJ6mrCp89MoMF
iDXYBovnH8NBAPl0l5bfpwgvFqWphrfnPwWu6+X5lflYwicsgZtVr+P5ekLKRLqLLjMvb3hxVpGA
00x5bmYX5oL9XjkHmLSIImlduSrJP4GQxj/KU8Zms9+RAubzHKTwObeuHN0HhwCfdOHLbDDhjNjf
Qi11hl59dXLuh7WkaVk+LATcN0/Ashr/qLOaYeHJS1S+wJzVW1qH+jBSioOTM2Ot9bIHV4E/tcWJ
uGRtyt25QVIGjme0Wpat8Pu0/3o4NJtm4oURj2JjuvMCOEM1Rq8eNioxv07c4nRYFa7RHG/hjWOM
cjA2GpBNMxSEJLV6OMn8o1PorXT9b42X/vIIUtniYn38kRAKBjlQQG5qFro14XOYHfHf3qSBunvH
9r4BLTn4MUsmk4BXg/8GJeF4fUyUK4KAclVczG9x8ReegxAeGFJxnB1MoGowHuSN5+rbc5rDNGDr
1HzsNiYF2VJFPZgP9a6gXtP0HcyCFKHqdGJsuxeWqXmWOsCVVXlus9qaDJ5LG68RxFRwUaJVOnWn
hLUyyHjKK5GKwXVW5RzOg58a4fQgvpEeusdNXsjHDoiZOSde5bgUaGidaXzC3M5XSzIxNs21O03F
YT+HloAsYfxRI7PVr7spG6xbV98Hnxxc7KXZPsGfl4Z9cn0pxUNCcPkk4f/49EdL4WITQwwJ0KFW
kmOEGoUXe38735Jpf3a8cODZwTJ8t869WMc/ocDLY+9hagLm9bWijen5DMiQSAX5Bkbu6sApOWrW
9m604N0EStCtCuE4Q3CNJtMjnPodmuD8zBKX7VdEa5Tutl65FPrV+jik09HvRQDfdYxc0SRK5e4m
A8w2ZZVS/e1p4JB6s3SMVrG4a929quKy1xBN0ZtHzPgStm4hMUulDJ6suPZilV+NdwfQV4UC+F1I
wEUcT4S09LhYWSoHgPRwJ3fg7S50V4jPo5VdGt9dTF1zaHz9/jHLZgrJsJ4jxq7V8FHZ4uH7LhWH
tChIgrnBaL7nuXhmLooBiPT3X9P6+7Iqu4WkF+4uXYcsuJo31xeuym54bGBK76Uuxz/KiOWfhkPD
XBJWlgf+UdOIH+Y8Utc5rTapYFPxmLo7ntYTKb0N/eGsvx4677uzAtYxOSZrUBh14LcFm0ToiGT/
HGUMg020zUkND0kTrweODmEz/w+yYlV1hVm/GdSywhtokbLTw/i+fGcSBV5aPejBg08jmLfvShMK
NdHWwILywLg7yDrLAcD3hrzcPMALgMcGWmIKKa7mU+U6UQUC8PkzsOSyhU2yQ/UmD6RAQIOKA9Tk
uCAzsmGrSl6tdg/vnjg8RUBeLlArTPqqNMOpO6YEF8OATAu4DT4w4gfjqbWUTWRVEbMyUj5qKxa9
HkimVgNWrByxcJt5YlzaPs6+jdplTB/DUgUGviPqZjASn8vsg1KtMspDFk+/eww4c7mfbWlQEPaX
nSslDHGfpgdidfyUkLnfr1XoLuk0JbvjPnXc293od1OqOp6/kDAqavp1HMLiC6EcNySqPFkdXli7
TMgxV6VtMvljDs1Nt4gly9dBUyhUftbkfXQj9KkQrNRLk59uerH58sZP012Xls90lBinr16BLuMF
BQplLxa0DPUG4R7SEcL3ToOqQ4wX4pACpjzXM+pfKNr+hTOHvNNpsNASY5+juzQlmgq0lF//N4pt
rqKTFYa1sxjkPKzXAZ13gOwKRf+1c6Si1g+x0jYyykQo5CiI4zMWkb2II6Tu+xyICVfBxcuZeSpX
tTi69qFZ097B5obcOzJ6TV3hLSJYOr/pQIRjyGEqWVUwUlO2aFUboRQa8FRUmfyOIzXCO+U9O+qN
ZVfCT91A0fYL8gtnkt/hPGsXI4cDZKe2yfqwocenNEnkONRaNHNB+88cFCTHDPP9hF7v4FnzumLy
FKnplXp87yiINUBlVwbaGCvhORaIcw5oV03P8JHgvDyQk6AkeuVVh4/XoDTOpmPwBg1SsP2Kg4qi
GACf+/Gkpy1/5VNn4UPuZG2H47RO6Gtx/Pq0jNjuHITfNOz7aQrPnYuuyHdqlS0hcWY9yNJtBYcV
RnGgPWZycztAaZfMealDJjlk2RpJ6OP+q8C1mngoqzZtFBcnxc1OrRWBbY6kVC6kT7mulz//0aCd
BNo3ubLNad+gDpjH3Ct4aRsTsi0JFwjRIucCdb2i7eT6MXHnzd/0Dclf+iysT8Yd28hDiSrq5JZ6
Adm9JT8HC1D3OvFcZdf23nhthDUV9FBe4zpeqwrDgmBi1oJGIQmxEeaE1zVMU4P+HPQQyO7lWsam
j6SmAO7ZuQKK8DpJeny+bJ7wDkHuRgkjaizzmdMQAZ11keyUs+Z7RtKZ1eRuFW9/X8XsazAIcE3k
A+a6C6mjSPM1r3DlAxFXbnROqD4o8PA1K5HwhyYR+t/HaFqX2s7NC5iY1BaeysiKcreOHV1JLpdu
t5gvOSIlfsVJTedjtobsiuVVlAiGV3lR8RcTaiacAmTeL63g4qGoE/gor7MhDzig+5iDcxiCH33I
YUJwt0/c+zeacRyXc9qUYz76wHbPo3ijLwQ7g/ypkyLGOP1+SXHIDl313fpUX3ZVzqHs6DqBXL0j
FON27LnXVq/OQpIr5kkgIPdeHYZsT9wEO4bR6TMccUosE0CZe+X4lUArZM6VPWqiW+fSVvrz1pGL
YdW5RVmo2k8soQ4vDCLu9N26JchqI/DloYrY4c9a2bQpYWyLt0714ocuVjsllQPOH+yNR0wAzTbr
k4Flp5aqP7fSdBhYpqoe5BUN6kj273JpaL9UifFa4OYcc/bRlfy4EE4/AognpynRD3yCxk5CieXx
Hp4IjiqX1grPLBigEk9ZDY4f91ac2jGgAUFgC3/EK2DCUhRA1/U2F+aMtNAl23IPMhRYMmIXjjoS
7x4cBS5QkJ2n/BnHt0PgdPrLNf160KY+HaABuoUM4MZqlrTi3A1+5Hs6J9t39LeAyDK8vLhFlVaI
mAZGm2yHgEkCRXvKqnxdCXIPVxB0e87fFzWDfqXKCtPCnwP+DeXReNusAOwVcYgbvg0pY47jb8an
uQcAEVoshMHYeshOtHnl8uR5X+yKFPrvAxR/wJWm7FRfh77PFq05kzKbIEo3Bm3vagjoXr5EfExn
kM19f8OXkvnIZMhNuGR6WMD7rCOcMvlFhGR8GOUONhvLVinLkTLmv8XhhNYYLM/i7r+GSyuf3rLE
0gUznnPd3PkH1kLrE2G9Rpu2InUFLyqeR++4X7iFqcAYICAghJyQ775AamVQFiOEa2ae+gs9c9cO
JoTi+RniCipRWUKTsZn/GPbsb1GJoYmL/l9yxjDGUliEP8n82++WSuakKQAAT/0kyeHb3AUGXJ28
/1G++vxs1J2uGA1GWjrwdM5BFi0gWYTM8sEW+nPTqw8VCoy/JEfoeCsK6QfPziJ3b0S0pfZJGmCX
qoiLGyw/puIFZOZ/0I8RRVy8Ik0Zjf175ZzfOduDz40JE5zSw2tpFWoi5Jz9s3l+Fjc5TIZ/ROq1
v6x5oEcH6OD57TC5CwM8XaCyip5JZodudtwrIpxYPJ4Cl3OE67FBeDF+2MkNgIPVM3StY1Be3Voq
tS1yxY6i6AqAjChyTtXVyN04OoEaMNZkU++Y0AVqklbtbzVgKMvmpTveVuOTv6OsWZadQaCgN+wx
f33UuPbUpv+1Z3nXLllL4KPQgZmONmIY7+LfO0Hl6+R6ImL0PUYoqBn/7V4GyzldKXMljG7gyuJb
eud84teAhW1eJhbilVST2EdJtDgnFDu8F3v6PxuWl76uzx8fFRB4VWxj/nZXE1Te6LlnflUINbhV
Sin+Etn1g4VfvHfkfELxE0g75N+UKIN1vm8vtJdkAiTPY9jpYxSKgvKWmMlrOdAuk7RxTcEw34vy
UMsY0ZnhohuJiSw+u+DuTFPjWbsLANGbiLut8hNoKT4DIzPD6K5UU37a4KAsD9RgKHX3/gIYDrh+
iea8DM2fQHCTnk+sw+4FxaIcADUf8zdguPw5YYjm8uORjB2CCI2I+8tm7Kf8PWIYe2m8UyIV/Zwq
f53NigbJv7fTt2H3QYMrPDE+W4gPH5mGJVeA6BkYjpjxUvhos7asOpkIEJdL9Kp3izQvFwCryXZE
ExwFvgvrmQfgRpTQ/vIqkBkVE+wJdKIjhgTfIdFMwGs2df+jkbqvdP9MgQlfDx/jnDptJp1H2cCK
zSV8uE/Cs5worMuJ174RzkYmbsQ4uAPjKRSA38Va3q5qWWnfMPMA6LnMfu1jMmmBxdpRUA9lnDqH
uvr/91YD1gHgUzoEf69aVE3RJe3oUcJKj8FlkuKfxI41KHqokpvydlIy1cpElAYgmEdiys3g4jof
NyBR8+k/dcqus3CagZKeoSkhYs3L9itOABF5qbyUTjN3WguDG+jDjw3DWR45/kQIWHNAOZmxIrOx
iB3zO9qIrZyQIAqEPIkybEqlAso4wRbzeLYjZXDSyqXIMiB1HUhojCiGy3fQ/868MsX+qc6DZACY
0/2tH4V0q2XKG2qgTjszwwJirTPk7gXDrXU9E0NzS2tITS+fNQc6KCoqsL0O3YS1tDrMzMsHKIrx
AhuW2pRi9w0+0uicqpfVlqgj7mBujekurG1Z/B2+h/kr0BgM4/r+njftgR/KJDMQuLfCbCRu7qhc
D8R7lQt/2hcqrdNpEtgijqWQExCWXGO/XdYFSFBn4yJGfPMCg266dtPAzxuiV5ovAvpBMxQSsG9Z
jx7jqRjGguYa/iSLaHH6liZpqiM6LZxPuWPJLt5L5VeVjdoMgbBqntIEv5YDgNX9f08cmjTQFyir
8oPDOWiCKO68aNcjBtS/QFQhJktcVkier657hVVwZ9E0N8OUueEraKj+/V4t2i6TqcsCd3luM+of
805k6dE7lIl41QQMJeVO+IfOB9etWU1MaEcAg/iJlauY7rvoFsVxOvluBR1p+PcCn/7l8+MxxRE6
wF3ZVahM+clpDsnMrJ44D0anOO6ZCSP+C6B1NdMSc1nsQf8yHVAkYOgB9TKuIT6FWrCOudQzG+Zt
1Xmylu/54C0CDhAD0f+2OfAkab1pYsxeXJpSPWPKEvJ1wVi7K4m6plf1E4Pfxgpiz+RUfbo0O1i+
JkBNffRi/Y33TaqaD4GLtm5Uj9IG7o0KhAZd+mb/gdJLiGWjDPyFEAh+3bbKsYpbUumLlrQ1ZQsZ
WgeK0Tz0qp9HbX4JRKHuw3pvVRpnhcOdRv2rPVG7OOP50WSXYftydWLM9NSyJVddbPl3wIEGuVUD
z8t/PUMyRsm+uI3RNR5E0fY3kzlDy+zUa1B74hrAFtqLKtcjv7zFZlRJOTpkn3A0KRmuplfbY5hG
qm5vD1ZZt2PnYLmtMng38Mf3s/b2L8tLohwxodM0sYfK3/FtGP9nKaMxjKK52YmJ1WGN8PZe1q4G
ITVB1xmzM4yGqxXQDo01hTKAxxz48X7rZBoOr0V3yKd315o3Jlw6yRcN2y8hygFHGnOE41GKQ3Er
XCn15m9tG+vHQarZxuFqEF0HjDy6q6+NaaIW5Qkaj22+nKlpWUEl2zWMWDo6K/n44lSmzn2JQTRk
AQeQA6Ki/GZ5vc3bRkctvE3fSWsjRkpaw1FeH4MgQ6eI0cbxi728UVldpM9pMlvcqX2IdalPvfTc
bfAsxFb7CrRf8hntLqMBTS+JtZCPsc1H9h/iQUj/pCNEzGddkwT3fnTOZPo9969QQPQ4qKk6ndel
hZjA1EVFQZQQGeo5y1c4ZQvi1yEmGwZMzxZcGhijdC/fmuzTn6B3zJnnjyklTTQebnp/fp1bhkyg
GhjUX6DoL3utsquB4vA613abe0j5Ozw4FQW488zIUDzZtA4jJ/N+egRvO0J9980i0Occ4JhABADz
0VEdpSrnq9GI5C03FktiDQqQflyse/CkDPsFYTYxWNdK/yV/PEMMxnHi+Xa6d46itlMxsl/PSNC1
9QFHw78M6EyfVXLruPY8QO5f8zUBg3VnE95s0XhtbgVSobR7svF2l3l2FA2rruhoKFVui9ofODio
wBxDHGJNJp17lAUoJdpY3N2w9Ot+HELZR0F3LwZq8DM7BUNNVE63YazK5U4yQigNnYR63SYd3Dn0
Cl3ey3j+a26sDFi7nAOoJH66ws7doOL6wiBK7YuPTnJi6CdajWwGigEZy7+HgKCJbwzJfunZxEYg
X334u6kPa7/ISd9NVk+aA+NqbTsHVVPDXEI2+bQdJTMQsKTSQaKalQvBMtV7JEGgutBF9k66xh8A
L38E0LqGYmwxmUW0UuscOTe5PtD9e9QAoNsB7VY7gtoMKTSZTo0nxh/k7/FqVF9xskXHbI+pZLoB
XFGkU3JAj70lgDUHOMyxPhz3d1XuvADYIr6XGoAQHaMMwq9AC6JtJNv8JEThB8o4+Jvi7XcYWPgq
yQtIkH1zQHi1CInvtdeDnfBcE6see73RVwnKODba93Ceg/+PtemCjrXFouh6ClDVA4Hu868SMfNq
g1OndFjLSxpKShlQuvtKOoSDC8VMRoyi4gwVbN/gSUxLD5gQVwUihtMNhh54B6UgCSbmvF4gFkHg
xt5YOl3CpA30guT9sxS6ybSpNj522bU9OnrPBfHIs0jxBB9R6IRuRNsW4a/0WJ6WLTznRjjBMglo
bxX1fiT+9xvXE0xNRRzVnRdEI86pR/mqT9f+pn8M1wAONAPjoPO07oQbYuFZY6wImd+LsyH1TTxS
E5CJW4LuorvDTBBJECRszJDBnHWQUiTG1Pyb+SHh6lavayXqEPccd8XMIW62GHwBDuYbu2M4Ul9K
MkPmbuPVd9BYdnSRe2GuE/M703glY6P8v84T3+TEZVLQaTrm0h3lGM/N4iaZYKUjcFoAKARuxKC6
+x0w+Qg3ifP7QLBsyUE+Mo7rlgyiByqVF1QJ76NOwbJiyyLkQ31G2DxyoGvVzDDTKKcXErkIr1De
5NxzjNiOC1gt0GtvZvsIObvspbpujfIj80G79b3jqB9C+zoS7pvORhzaaBX5u0LW1/I3ZK7cxvPv
ha3MjKXIra/msR1aymEUSxMhJjoEckByJiu3BijIAurC/Q6Sd01sWb7HIGRXl2ERMhcDsoaMF6ec
Y6I4rNf/o6ip06MOW4d9vYBJrP8ixEQB5ku9oSQZm6c8RBH6EjI2qwYX9UY/YHEhxwFq2h8OXNQN
TMTrqL//Ts2jO63FlZD30S33rCxmyhcNsYEfZfSbVJ9Iw9+QI9txQ5XbWqYD4rjc6MMWjRFXRBNC
e3gNMObKGZkOOb8OhLKrG0gk9WUiYdHt+Am1KJmjABUtAKvaf7bo7dEx6KBMHLSPIyvI1eFkPGhg
RB3tfhMOPMw/+viZ3x4Xub/VLZq9ln2GBI2XRz7zWsr4P0rLCEb5vC26EyxPPfE+05zdrSO3AlJX
Btq42XdlvT9+EbucHvWWhf1bloFHkIW6zzXKIT3vmwAi5bs3uKnfWkPcMhXSQbjBkEgkYWrqsCaM
OTR1wZTPKER4egjwkzziKhtKb76RtKoXG935j18uxUZe/FV1W9baWaHZAlXjCKV0Kmt5zsWUOxhw
huhfqPPIJ29qk7sLrWnLZhR3VHIqxg1KnEofKFTsMSyTBpOXscmt9iLjntmuQev7VnMts4wNt6xg
hOY4uW+hITQ7ZaiAQqLuqi9tlm224M39HmowWKFvT+jm0YC+7NY8+tZflvr3YQ3lWsc2EEg69zP7
2SWEoJYkgk39n6A6kRUlHjXW7m/LKXwcjjzP7h77vJTsIIGeuj+af1qPBnUmhyUNiP8IqorXGClM
d3XHIwFJf8ePljmJa1/BRU0EdQuQr7Z4cNODPxHxEPDJMveZtYfB9ti5+6mmhQyV2wVJzdxCeD82
n44l1M+fZHTH9dzqoeE39+FPmAgiagBBniumetjAGtxzF4dQaXwZRSV4W7UOLXyxTxVUQBpitlR5
boZ8AWxqkMP8aEGEDKQt7zO3ULdpYosNndpPEKiTmwn1rh5kO62ObQwf6ovfopwcZi20UysqpxDE
zGm6z7b2sn7HFLvPEMJ882lJKOZccR6TVABZcGsfCfjB9xZdOqIdI4abxfdnCAKcBihf1W+XE9OX
FHl4hN68+acDEG6px5VuA/GAuyPULyjcjJZA91nKsVJDiOVXV1OYKE6ynsZaBM/Ow/uEICtM+R1M
ay2vpUghqtihBBSR+Ktb2J265Oj8V4lpEnssy7TWn+IvNfctCL3foqHOIc8716GJ8L0dLBVpG0BV
Mkj9Dx4CxSktzhz+/sJ7a7DuK39yg+Z+VAdD3p3M+ETr22fRM7WhZvwPXQIT0VNc3nthSl5/JH+D
oNCvit5E7cLEPrUJ6K4E6YEbRGAuSSabkORBShtTw4UOHDGIS8tXxjHFFudOVVdyiJMQKp/HMoRT
VBLmmAfy8Z5wLRmxfTxgGaiiQFvDLmLDb6dlvXf9luVByrP1GGVJ2FQ/9bVqFE4nAq43X/zCTPF7
FJqgqcM+kyvH70VAnREd+c82hcnVrsnxrSdPHPnkyQd6MX+FpKPfTHYOLbGOAcRTyp098eVKzxyj
A9RLZ9pqzIdd1zWs5+8q8D5fmsk8oQF3DrWmuI4Vb4Qv+KiRWpQdem+pkj+WOcE+gt/NAgUdHYXD
lkfxWWqedM5MN9N4JCsp1cKdMsDZrFjCK2B9HqA/gChaqSZjjR0rr5hZAurtEW5dBNz7EWy2SDnS
67XDvf8cdZ08E/amvu2kpXQsJrMxsTGCJ6xckbmwNmYpY3+ojFz+h6EMryL1xDW2xKfKO8WIRfWe
YZ4Xfrtg0wyvVBH1N8gxUWxMgFhlZNuXmdHMHQ4kr3PR6Yu7V0AdlPqjmG7F3phDiIzZ/ApMiO8m
k5o5L76kp+CS0b/yuf3S1RBV7MCmhryzjwriqkmdiMR+3f9RhVtjJGdqyqYCValriUKZzJ9JyjyB
YhT7m79R4kozySX1YF8RMRQrjLfN5zcPO43HmxGM+wHP7PJyf4KriK+HBI8j7Rkg+cIVrFSPFSLz
K1Gc6Y0njjOkMaB4A5UJJqUPZ8ij0C/gakxvWJlP6OFMTgk8xH6et2zWuHEYQAcw6hLMKQox4C+w
oUjFLcCZICkdcjjDORi6Twqs0m18JQuFt+MsX86CrdNw5ciptTCnbDlRmz+1g7aCvreAGyH5agoM
LQXCd+cTorsiKQuu7Rz1DFbcgFl/jSnNUp/d1jXCc3PGF/Fj/QcMdvlZffZJ1Kzf2o/R0wiRAGQM
CeoYCE3v33B7+xUJus12CNq8PXBR8mR3gQ7rJZ2h4R5XuoQI+nEWe8hdBS0gEYPtQ2tZVJljYdl/
iHePm8RLpNHk+9Xngwyo8Ur4XR9Za2YDz5kWVnrkquQhkTZxcVKzcbA6+G2jL/GCkWYdCd6hvJ3s
zvwPhnTDt2KXAJg5OC9e60MNcfhS0hRn+151E0NbfZGaiybkpeeNrdtNkdoj/sQcJykyuhN0bVSu
nyA02B2eLOaoCS/IiMYf/ogj3CyoPVNge4MA1aDAL9WWk9ScwEma8y2KLOCgy9VgptoGhzNjiD8S
kO+b7gIBNsnHPJ/sl6vTf8Ch3Wa/Dp2Zl7kIJihiFZluBxUibU/vcRBGlHAuPRQNa4UPkXylL0ol
5PckUsdGgxnn2mZBwM94841UAhSbWRIUdEiatvVIMa+6IeSowpyn5Ib29L/piR/AkLbpoQW+SCgn
hZ+YnrYxtKfmlw86JVMuBrjqtEhh5ltpbGYXaC1IWw3Jp8cBiHce73OpGtuPZ58SoCU+65xfaaJ5
W6T8NnmNhqIdBvQXLF2ap6Ccw35m4F/y+R9N+3IvVZlVywqzblWB5ydt5P3CxdC/5irFdNdW5GHC
yjcIc6CYs14wDrlY51ueDXLATbzAp9gakLNmvI1znbV6/wOPoPeUIzh5FHcZ+yo8eu5vuZDIuWzb
vMaFmJhyg1u9vcYMnkBdD/6c9TYp2i51PnFnD7FwONS5S4eAOK0KkuWegKZ4USxaHf7tJ24FamLh
XcXBx5urrrbqfawxU+JCgsdfq4s/u8Xhx5+n8SBoAyUhJDH1rvYe1Ss2b5pjS/ZRKOqCwG+MksxU
YbxYm3qIc/L8+bRhWWqiBZmeCx079ysyxrKvDveNdJwAkl2X70rg2NJK7E3pWhJyofJ8W2wfROXT
5ZkLniMWL1hPVgFX4pgseb/GX5QvwPHX7T3Cfk/DPBXvyEBBLZrX7WyzzwDfHati+kMJ1P34YxCk
M5ngBwgCAoQkdpeJsBLLETsh+Z8gtgTyfxmGZXvK2xLl9ObrybPXhZe5TzUxXWSnzuvNqhU+2PMu
aqbaOFwFZBvHaSO7ZMv8LJrTcxAmqsBpwV9MjUKqLki+WXMx44El9dTzRtlb17c6zhvVjPdFoNBu
Ff0nAVMMdp7gOBp2NDFbOmPRAbEwCIrkxKLI3OUE3U+kFr9vFOhlphxvhRriLwaot/C0m2D/rW1q
Tc7YLBXAecH5AeLCdU+Avrubh2moXhaSoL1TWO8z/E76wDg7svuTjcpvKN2K00Vo8OyMw/hx0SWK
qND/zxGWPUZP270j+ch3G5nmxkGRx0BXZabhJoGWkxWWnu1WSUj5R0MwWtkR1PFGSNLcKFWdYGND
jx7zXwnEX5oBgWavgDG21MdMyKrVcw3iEhRcvOH7U6+5L98qV2yZIAi6z7I/p3Eq0JhiqLuPnrxc
sT6iqfSQKf0frQy0H5J9SfmSSBgHkjEcPiCn7hjBquzczWXp0d6DsrG4DD1r+RImGjb5sOwO2d7+
7oXyIqHcJ5grSP0M+l58rP7BDZbUWqg3XfI6U5xsrkV/N8gRk/7hy3L/gIXNVKIHUfXd4Uju3SO7
qLGyF/WVKODQS3DX2noPao0hgPYh0Dd48PVIe3OQhoyr25V0OkXykYn91Rt5k9wMPf8t9mIq+GOY
cCEz2vIWlIQBJYW8x8mZnqRwRu3nkF3A1XDD88kTKLL69anKiq4U2ry7ZGVJxicp+2OTHbsJGeXv
NN3JkamrxxkLv+qc2lzZmC9KmGvjm6ICgSVPJYRfmG8orNX950spX9RuvuDFGPm+A4R8lP4Nifhu
Hi4SUJgBmcSbrY+rX57w1+QnPO/Ex17wycgsV+DT5832P71krdqNGJEpGmrSph2Dpl9CQqJKT2Ur
w5FFSqG6Oz9dApBVWK5n1iIYowB2YzSKaHwDDzVEcuGp7xN5OgQ+Pl6vdTZCZOCtQje04DvUEaqf
d5YGoAMp8FjSBw5CfvBCCmNrJgdkX4JEcSV+Lu2YBW5loelWG6+luzMOHM7qi4Sy4bjJAjh1LxG8
7IYwwTq9HKgokel/LM17+DNEIf/puqo0R/rFn6Q5BrddaXRdovvvXeiAZdkV1LM+x2PiIrK5F3BG
aWDuE6CpaYGISg0s+KG5HJ2saMDQ70UCp6bjzaC6SmxrzJH9n5uiUzWFGI2fCV9gp7ta1ZLGrkSd
3sPsMX3KYL74PlRA1QiJ6qFaKYX/fSfJDK+QX4oP1tz4WaP9GUTVOVVjOVcJijcXKFK2cZmncaiZ
/LkRQJ26XjlwlfEN1VU1lfUHnxmmItfWAEMddrA2VN/if1p7V5Buk7eaykgnPVoXSB1FbHA2gARc
LhMthJKrDUUqQK32U+4ASFJT8PbneXKfCA7ffIVq05UdwqVRHO6Vep4BhuvmxMLxZFH5mDB0x8ki
F27VWiBDyC9230L6KHhNxivXkQy/S9vtM09ogFjx7ZNLZp6/K5mCbUvhrkXqELum/yOIBVhm0IMe
B8rkFn6OdiYvNT3J/NCaJmCtULC+6brkyJ0MSdw2m321pWyH5BS1elsLQzQcYkwbfUbrfaAVwsUS
4Cs9QoD70G9YfFSNSnYAXJn4kVtfwBx25PdFwmr6JTTM5mLy1QVsaiVAsGFDfU0KgiBO+3a3pLPm
YAi1cgWjrB0AUVkl5iQE2Gh0JAgE9UmQPAWeg7Qbc+Unx/NB9RlwE9aPjhvFcuuP1Qz9CcNOATG7
pWe9Jna/1RYa7M4855OD/nWivk58ltNBy+oZZpcw0wAvA+yDycDxAT5wPmMnSuZBdajWhM9G+jj9
4EFioLTikzRTrkeK4N7tWPbNR3WpE4+px/PnadwdMqQUP/PpDZr9TEzrqnLFwUCzYS/USbZVcBTs
c3ilsXkglYb8A0t7oEzoktxd4OFhK+4nJeVvpEz/JEKpIGJSd2AdW0XFMBSPI83YrgiKdDQsA8Nn
E090Kf0TUSOsQUhpoPJc4UwX6NL8DUNRXr06tadXLXY8WNyYMVE4Q/z9NqvBel39jVBNJ6e2bO/d
tyby5A2cHL2Vfqy9Upyyosm0B391SAGT4YwHu0PFTtYb7DGJ79hYaCTl+2iRn7qD8fhXCpk747yN
Ykh41orz8NiExztxeZ568xyKsu8gRW+Z6TeQrmHmaJeDsXHDiwUquemTRIEliANu2aeRUCS09F6z
+UL8DwE3lcCgLyFUqeE5OW6DdePlezXxTr4mcb1pPcB3/cyBUkglSpfI+l5ib1MmFEh9kTRea/KT
xGkHosjmlNFs26T/ZKLIlgx+6ukcjjt3V91Hg1crfCryfXxJfjr4OBMaoPurpoNQncHyqNjV8GBZ
bCHsHgizclCm6JBXLbYGqZ58tYux55YE8YoHrXw0PVPdfMt8Wo7CEUPIzjcDNTipswRHn2e+n+sO
zBAemWVOlpGIXiXkqqapoV2j6CXVELZ5qT/yMbSZ4EfnMOBEICac8c0foHt6e+UfpROeCa75fXq+
ar1ttiWr9Zv9ru74P+vULqrt0ErGEzllVASXhrWX9O244OtA9iXAUjuKCW4cKngkY26P8NnTgvT7
U5+hgUetBbrjlHSsodSppHx86SSs/sSMcgQdymbiQqBbZzFQ+mCaO0soWh4Yy6gcFB0n0po44gUV
/Mba5LvKXAYICeQXJwAm51IOR9Zugmy6NRBg3T1pzW6wimPtfsAMcVszCAVfMu+I9RxblzE5p4nh
xY5+fg0truwz1mlibG90U2Q+j9H0FHDnV1zk4Tk8jvNqdvw+/+yTaZ1+y/sP6PWe0er0Yud5Bts8
A/vZHlm+FQ37aHeiDfic8dyM2RfGTuj939YRZN2CVoOjuzCfziW6+MmS6/tAZWGrK/iMORVN0YNr
avT5tmwJ2WF2QkmHavf/ZEcbZAXjs4jXZGJ831CkFjloHcJjxzpWHgdeOFqHtYZVTpqLMDvKM7Nq
pdw/lsINZilVwwoEe9naB0uertlWKIgHLpTk9KG1shH0flYo63iBAgAoaQU/AQ9Nyc36RN2MjgpP
TDRbl6lzU6yOKJQWaugmJGq6V2HpG2utIWNuf2Jeod6cjLfZBJfuMfCXDfBG3gDwN5mdqG2x3eK1
BLnjpUqsoEXPsy+ENdnHS2EVnnPxjUChH+7/GyZ5Ek0vSiQq8B2uXrKrtHzYDCgqmXA/j/un8z9w
hbLXQ7EtJJD+DENxyIITAAq008Q4sfF9IQU71glCnj6YzmeihZC/pElhUNLYPjGIVtwND6Z5YQtw
W/wBSEuaNzb8r9ljeTCYhJgEV9qAaBFP2MxVcjMKM2vQwGAzJusP4eqDISUQYm8yWweKouxH4p4I
axuX5b0PgF838/CKYEyH4sVEJmKrcRrxvNYo2R3F9toKBaMXqe6FPyIzKa+BCRfKXMRnEsdeWzwH
PivIEqYZ0cOU+79TCxcqXOTx+VViUjz6hwFAxqBCy/vCsGbYCiTBn637uMOLjc5fHI5yKd0m0rM0
a0eYHZ/7plQxYiMt1aUy8EdcJ5gPa4QG5ecarJcu5aIe0nYXPUQo/GCfqifv7OSzodxgJDF2nvcL
l5FLcRfcsh6IEjT2Ug9PZUYeF6Riey/6AlYpX5cYybtsJlzuQ+qus1QKeH/SslcEg4Wzua/TFvVN
R31FqYeyzEvmKPYCDC6h3RmKX+2n5/L9v0yixcDY+VCjKVBpTbczoXW5MMZIDZDCuEIR/WbU5za3
BNhnXybHD328c3couHzxZVTwIoJU9yaUreyVpZ3vA8q6jwlJmqRom+DEaBx+UYdRir17WFqY48Iw
qo74KYbOJ5xGM05ntpRWL3YknLs8oUV+fBtwGoeWYnUUDQB2pLItmvbDs7rKpTV7Zd/5LX7PU+H2
5B1hK8V+mvkHnGfAwCZXWp61e5GoIxpIWJWdJz1zb+ijf6gv8r4+lS4+p2+bgbib59xnedzHef+4
dqUWbz6XV2caL1vKsMy5bKZb1+RCgDZzfcNfmqqrLrMoA+ourY/BueLa8HFL08RLyQjEGM8u3qZj
mmPtlICUYltIFtEefL7uN3cmUAWzxba6wf9490LJYj9bnYBfJ+UkFXTbbzHcEoTbfEozvcTHo9M8
Mz4GPCSZvDmIMQOlYpjc/bX7Hpz+eTuJWmtDpfUZk176HQKJMzUQL6mtdHiBUTrzFdw6YtmBoYvo
lEuokmBDf5A/so3XI2N5RUgsBIv+kP8hZ9fcXjAY82X3mtESWLoAJnLEP/cAo1XZGzp/2x/0+rIe
VA7NgkJQj0Ed9+wjniM3mZ/0Qn1yJB1/Uv3Vmn3w4HRAMJCeUjkvkpS+TP+NsIsXNDUuiIoPzjk3
mJrxIPrL1UpxY50QFYbuIr1wDTsS5z6Cl1G78MUYbZZ80fPfHrt3mZQNDK1Y6ODU/lowsEOsAaqf
+0FHLohnPdH5x9ZngF8+lWEUPS678tjXxqULXs2WLE9cdXdIdTAnaqYjv+f7RWEC3mgNfLEYO7DU
O5YlzvRnPygNT/EcOaLF/UbIM0UEZHgEdacon6iZJD3Ywgx9fMUYITKBYIPjSDI6Bme33rkttZqe
xzJh3kktvpXTmMrybvgES4sELX9CAZMKsVN68TiXkuiaQ5jIh9wfb8SFfEq7qNHesAH0FaeS9HB0
tvxOVFANcgeCKgDrz4ic7MV15KdVgXqmcqXf7iUOerOrgTjCCTSRf+BaDF6YnmaR3NY9afuf5Jmg
cPIGZo6PFiJU/+NcKiEoOxXvvu59WCjPq0biQV6WLHoFGqxgGASTzANTgo+kDXONLr1bZqoXyS/y
OaZLaD5SiBhfjtGzqev0GZLppPriWypvdkV88okCWPeuxshVVEGMZmoXQUFlG20PBKmySFVxR3cg
Lzv6/FNSrBJH4iB4VuP4Z9s/UVO+8LTvFMqKPedmihis+ozcnR1KV9huy1wY+/EWrhzREBGOz6MP
FUp/NpKgLT5kwe/l+L5yz9GBqEzwZZXZiugE6TXUgj0PklvUv7rEKmnJVLM5fApzdP1v8pyS9RKZ
uJXTKW67T+CAKKFCySd4xOdHrC9mbeBGu9mXaJ8QjaceAkNG/18KZXDQ/u3LLWm7ZIxmfeQYPN9A
8ROGYTZrzFIb/W8InPwOCqNkz6IA2LxIZKAAMWPAQNFdQocveyHdloxnEUKUFlFvjGho8Yd7Jwb4
2S0mLGy9TqJi4DZtlfW1jb/7NtZdlHZX4E7IK9Esq9G5ktYCnx4GhRMGdEAjk1R9ELFtByKpa+tM
WcRUQZRZ1f0L1KmzYFED9Iw3fgksNzxcMilO1cofcryOTDzy7VBMUXAEyp2GiJxqFpJHRnS34X9c
y6VDSfj88gTBkWUfHnQiFOscwqWvKG3WstRJvHp+aQBMOAvhD2dgeipLgBXhYWzKLCNgBe+Xs48W
9A7xR89flJpL1uHv+tVDyhxfwW/+PBC4ZYGLoUKTc6n1xI/ByTlCPU6fNL6Pj+vta9/LNae8kWnC
OXf1lWxwxYsvJ9keUDeNZbPZm9BoBYoKwIMVYlAP6Me52cTG3sGStEi5r6/3fseO3NG5syddBnej
yC8vjJmMrdtPfefeQqyXzqTjhs1uVCQWq4qRFs5H/Z7NYRZlwRhjqmdLUCH+l47YnhHiIafYwm0P
wG5BXwo2Cxwst9Le0llCkFkrnup6mfiFJ/la9UaeLPc3+cImih48GcYEl7vyoIlNzhYVsQKcjZES
D+IDeBV9IV2NSHxCBx07FTTqLzS56Fu1aSuRAlbMvIsFUrsEWYqxkpryxjjRSew08xIrIKiMXPwK
3sy1ReGexoP9ujTmUtmDKpMmK3mQ9Pb7MeKdh+tGuJ/JImi3I9RhFJ1bR05ootNywZ9F4JWDtowi
vEzW61LusL10Pl5iQGwA+NyRa+pIXMY4FPcLodRj1LZfWVABzA/cgcbmkvETr6FCbZyDs3Lh4igk
8/P7WRAMMkb+qKNUJoiNJlPRLBcC0heid5Jg+E4yK0dhkEomKuh7G6EktLecBvuKM/vaWGn71uG+
l4U46yvsrxQjxGhy4uJ5Ziz6+sGDCf11cUcZeuHlHeaTdE6LF/xIMJuy0U8oLhDjUEEL8XaKF63U
4hVAnXdyKvinfaYjJzWv5pWJAmBV8qj81mOUN+FiWsz7zb3ZgVRlhLkLhEWCKzIpiZQ8l1J80JEp
Tbb7FLJs2G7m5z39q7vOdJjSIWK58nlukrJ5MtrS6t2FeixRYuSpZ2SB9co2eNStk0LrchvXLI7J
wuzKfymk/T6eBQHJxFoySoWAKlSkS9bXzThlalgaGjj5h+aghST2GtTwyveaYGgtz0br3NOix2eG
UH7WmlmX8AiN7du5Z5Mkjkx4y583NfHGJ8etkQ2LQFE4LzW9SjeH2wn4Kbq6z7RrqkJRALNwp4++
gAkr+sGQacYh2eif+CxGEKMvxThF5PDIxynDEatvVQnlOFKyYKcAoG5HDw/1NDTxSQIUhvPC7DFB
US7KwW+gmBfiix6fQvoaM2S0oTGUCmVDG018ssnyXtZvgF6DCEyvFWHFUWz37DJTgr6kgA/abZNU
RU+IBfrshxYNwGzUPAN2aQRnGMYOTU3x/Vqv35X1uVAuVNH9eDpRsGBUgm1yYsDF3tHnu9eClTu8
yb9LlG/rXfcqtc4SXP/1qVMljHe5u4zKx/mbxYt7sAyPPJckc+BtAZxm8/0z3/SY1YNLpJjNfz4D
vntrPbn22vWt8SvYwu60K4eMbWfBDiJrDrrHwSp6qRRnoH2Jj6bTMsD1Iba+sE9lll95TPP6TsMe
Os0ViXrLemyoIeOjpz5NSzp+N/397lcjicEZIU6gxNRhwkCxUUesVOEZanjwbkeDQz3SMrGDTOna
nk4rViQZLC8A2K3QLvGCzXtNlAEt2g+0J+b26Xw+PeQLX1KDsnFoQxigX5AxIUKDjqfqq0IRyW2g
YoyOLiHU7Dhfud8sHp5QPw2XWsUdSfvBdf4LnNsWk5eeuzqOv5OiR5+yWCgZPLnsYs0Ey3T2xcrF
rl5O00yha6onlees1Rno+DV1oOxtwGHhJUXJ/CtqGWQwyI32GHDq31fL0lKr+fJSqbEGglGCCzmh
IJsReLtmxYnvHgGj1h3lBKeq79qighkVnWQFY82wrmfHe1FOllOwwl0eVq0uuMypnrFSROs9vHwc
kwAGFzTJL1+M5ZikkuCZDOOW8xN2DkjCi8NKLQb1tlgYqdKBREMpfri8E/LJcPHYTdar0EzFFf3N
i9ZVjVg1XXOMXWyoJkw1tygxwobIBNpN4bWEoDabF7AbL4zqsrwnufU4IkI9Id1wFVXsfKvxeHd5
G719cdyTtj948bddXgSXt7RiXSBcg2IuhngSxO7InReyVR4jmRDFCSKtG5bDbglvXC7wTkNPqXSP
g6QK8BGNCqL0+yH5G5KdfS+bozsJohObuKXXoyVVtb+SW0CD75XZbDKNnmIM9x6U5BAzdHoZDAik
5+VpDivpZ7RLVVQQgIvyktOmkgfP2/mVDvosUuHAlSmk9cBrFMtI9QTDLc0l1iiLs2RqDL8JEqrA
wDm/Cs9EBX9FaQRYNftpZEPqFvYVCnF6u8zDS4uw3d6cMabHccxYe9Xj9n8DvmTvbGOnG36wuPw4
vg1eIkrqAvmmLNcRKhJnRsrFL/9hgtti2Kj7AxX5K4ok2kVUGY2cGOJypyUBC5gS34HRHsvOgRF1
6vKiMfj/JlwI9O+SXqdXXhaI8P7xAkicuP+AzoJc6WOrPKd8o5QraqAEXaYfKCVTtY9nLPmQEwnD
hkDgFnN9ZKD6t8sTU16VUWug6aAYZKSQBbNQxxpmKb9ib/0/qRPnyStluLZIQpNK7ZXJT0D0idMD
dzd/xShmT54A4AwvhF9IFowHo7gUviSU6Y/+dnPSmA7UMqYmU0miCLoFaeuC9yTSfmJBFD28op1w
GSBQY3JWbMpOfVm5mbdaS78DXoMfcVVDodVbmSTsvUXd2NVGz8vIN5q6tI34/itRVSgFwGIZrjco
0PP09HJzqCXudFf5ZPbczyGaB3LCZLTM+fW8te32qrIfi4F5gKeXzXc0hMaVnpOzjgK50ev+1ih3
I/IGrQdsSckdeGcPVxk4EeKsWuXZH4HGprAXWttI9CtWVNQE5Er8scCuGV+GW0CpWxHwoBpBkHaI
hARfvv027syZjvNECqEGel0HrZ7kvxdh14xd2UpPoFFFTGtzrsMaxy6pdkAcsSKC5JVSeHOBjKc/
xmI4vw8fayswVqdQpCi17qhkeLs4wCPUbaj7+Y+BOFZKNJEVlvIAEDeyPnfe9Bx38Bt0Mg+fzkx9
iK7w+hYeN4beRaCVA5HSKTAIzh1Y2sBlSl0PVIq1FnXm4WbMDCNu82a/5Y11rwZtpEVHpQNLCz9j
1mzdPv1lrc8fneR34Y6m3+wWJX6ofM9R92VaPB/1T00gEHd42R1oeoxdbB1ApTN3AOkddWJBQ3PI
due3YbYP4++nz7w/cuVk5iZCu2uMtpTjJHxKko8d43RJNnob8v7+CTDM38GMmK9+9zt+dW8Q/wzt
RRRJtjxAtbHhyGItrWLUgTwXfHj4lazhDOVYMfdSmKvy8euNA94yoDvzfdJZHR7FPzswP2o11kJw
z2Czw5P52+SimYsruGPkm8PXAOO3XNA5rFjemuq8TdscVAhJ6fE+w6eruJiKsxMH3IXeEps+J+jb
RZMGEcLM/ndCVp1qRN7mywIW2gcq0ggO5pYUT1zdY5sw8aYAc8E0SXtt1SnEeLs8mEwnx4a05clv
AqbmAKwjl/CPiAxgcCeNIiZ9/NcbegLzpsD1mkYUupatkUUkRxtqpd7t6Z+/VwHteMNdMxoF8O8q
oe1xaSKVq+JJoD4sOwDj8+M6p8t/Qm+Fl6yYpaHwJt6yS2oQEsMo/8yx3T1PzExKSlUvpnTo6MAt
aSjV7Syf5hFXxw7g2WkyhaaB48YkhM04J/kxxu/6SXRHzys5RNf0mW5lJKmm48mQQ0XE0EdrnNYw
dJOIo9xn2wBh26vUidnHqtJdGu8TLzNeJ5DsWIFXANYc1WaJ6GmlI/zuaG0jqDiGArvZoLPxSQtk
fmuoDS5KZtqtyqo+tBeEP9Iw6wOMzOhXaH4jbi9NJ0afElxW4D69q0+mkk8nOhx/+HwXC5C3i7th
E4bVmzaWU2AklBQew88e8Selyt1/QvPfIps1XknPd2yLOgnbIA+3dzM49zXAfiibmbLZdFHfyviL
grQvX9x7mqdTT8ycRxvvrb9hjedshAWSbnu4MotIwNvWACHU6EohiOvpQgxhIK7BFjWAtdy5agXa
qMZ/xC6JTUtGrc6w1DnWiFkkYsSYZd7kuOTmeiPpV8KVZTDJA0aBdtGKNQigL3VCZQh24CynAvaV
m2kcxY0eidOncOw7f8VSWVV9Nrj2UtEryvSBz64dZuoSibXGhwxinMW+dXyyBKTV3j5RpK/H1mJC
pANnF3jrg5DI/P+z2q2rGMqhOYKZqKlV2WbALMNJwQi7yunh+fmxWPMc9B0WPPUQm63E8EoNe/ei
ab04G736XBNIAcqH7bGB3w1NL6+8Bg0yV24eN8flH1K+tfNMLnZDq1MCBAIZinYMcctxOt4rAt8a
mDcLB3HntMhGKeEJkE+QYkFHKilnJYpZ50F66OMGn/4YRwQ3ap4F44Xi15xWjG9TKshbGOQumBey
CQvJPZzBfZ/ZiTYUn2h6aSlktXWtjMH9JGHXpghaqjSf14kkE9ZMnfEOCseXFCOpXR+nRu7hgsvx
7z8h61+F4a6lwNTJTgKxqms4vXVOd9skwcnfmTk8adHoBr4YzI/5GZTj1o6jUIMX6AsVaYcT0qRw
L4nQGItrIPvy5AdLgJzhJIRN9eg5uP2yrROTQHCvRZLNKTMIktMORvgYsIy6CV4hUpWNb6uRIj+p
+ysO6Sx0iui9L+gGJFfuJd0N9mtBigxNhCTRCB7CsBAfdP4fpddzSE1XfR9C/goggviIV7z7rMd5
L2W7y6B7AtxFJbBdNXYSWilCPGOtQbDQWrxEamwvtm5+16hiP+6u5lsnwpVOXAntDBx2HlyFtami
zHhUp2MHHqatTws0TXDAqZbdxFhv9pgz14YF+yO/tuprbfNILEjsmuWfk9994afOcyy6o6pwED5N
hj+yyE6YFjdPUWgo9CPnub4udOKfCGmtu+qSb36lDS7k8N1IUp5iVui/3fw37+zuIM0lEhRayPfj
T+B4k5Q1rtGkhG0BHqdYEZG7RDSqouJJZiH1JqcXqXS2EcrFaKRiiGR8FFT5KRvybvovq3zttOYD
V9hjJlfx4wmm3KwjBI9imfuxsTHYqgrwJvtUICKZjfrFLc7S8H7cU+FZAuQ4LVkaWV35puk+OaOc
Coc9MNJ+8/ufCtxOkNyvDzkHxAxxQhXXlJ7uwt1wypjIjjhBG1OlC77vwbBIh/K5Ys7O925SGBNm
YXyj/lWCC1Eoug2VEPy+R0PM3hHCPQHqDH22oDteYZeAhFjSw9C8DtkAsAvWYHyIyW93ij5kQrCF
ZfwOt4fgE2I9f6dbor5YR7v8lMIpfmssiVoSDHiBQ94GNONV9nF1qtcu0FqTxoQZGA6x60qraVQi
Th+5VcqlFurRm49rKDSI7bz55Qgo3uqEm0UsIm135EnwcpYVnpgULsi9TY2tL/HcsQIrmtGATCA7
tAixR/ocGCoDYmuSefGdyxEh7vy4RMyTN2ZDq9yxp9JNM4i+OeK4UU3ipgG7hGbMCtxp4zFggTRY
hnzqmu5iAIOqxmzD5JUsgjBRKKP95Rv9jvyfxc1bvNhQFJsmSpJuxvQLVjERlONiKbSP9NXtEYLL
hTpUThwo1Sy5grbveDNdWgCrIUVluE3zT5L7OoLBdLCOnCkruLTZr9MOF2AKjwrkmI5bBzkPJ5nj
J39xtIdILxQX6GKJ7TZtPzoZWWYBbNLJmOFjwMSXcDLjVLhQAb902G+Zg72RHKkDW8xh8i/E/kGR
44n5/5GelP0W28/uon13NKJVOImPOHE57c03Sy8OtPeYfihzN8oDfu/FHaUJl7OTUaMuHeL+jYMz
O87lqZEFowPugjtR7CYlbm47ujLelbNzz4SevRpoeiDTK1KZUg9b7Swqe6R8cL3MW/8KV86JkM1/
DqqPEFIN9UkI8ynGAO9X2pUpW1bBDlxb1b8lcNtUCGnp1vCqh5dnWkBc+SuP/ibXfEX2zCRWRA9c
zRpKIf+0hD2ZDBj99lGIZvymoyAXliM3bgIgK/1jnLKacvApsFN+ZM6UTjc9/ODqptedw0uglKVN
/LWvhTe00ckcxCJhyvcKq0ou4AsPiGZ7bOd9hp9l14c/ygjQI7Gpv/dJD+H/ZdUJiUpLhdXSOsL0
RABpLjQzoZ5hZgfGBclUghNn7JiwEftFwPVDwCbyr976gFQA6JPQkLlxSsnoNtIBpMEWgQfqELpr
U8czjivqIaBR1jzLpCM4cH40pXYpSu54oHdWHJ1Wo9GjXHv+ZpmTU2sXW57Amw2O36VE9TVuW4w4
bY43Rgc6qLxEDv5xZ3QT9iHihBvLdidEGvi3Olg1h7W8l9EQpCXBAhVmb3IsDYwOw92ReoaXTisF
1c1MK6ltVFV1gaRbHp8yccCeU/LGZwevIz+V46JQhbj4jrOujcQpsV7+ShBwCozDPwxItMxCOomL
ngdx6BG+FwEUmOU57DtxQeXdPfpHD9+JJzc9sdOjSKyhfzpxOjD5zobpv1qVqNVOAzr4bcKn5q4d
eM3Q1iHuXnODXYBlZdHRe4GVVhWFzDHDhJ7KFklA/3Oevfvap7Uv7D7IMn5RxJ/udBO5T+hRIMUz
lbeYZ0mHh1Ed/dKkXltnfElq5ebEm3EDCesVWKywCyzUQ688Ikr+xfJoNb1ru4fHr77KN6HkCRhS
vQEFe7noV5qpKq3O5WjC6lnkNX17G0Co/apA8+vNKRt4AeSnzA+cquSDCuo179aYcpztKoBPUXJs
U3XVCSIGX0j00t+JoFOQlusYta9CZyde/WOnP1x6CAHMTu5BNWuTpwm10KrNtQe8jHCzC6Xs8lNi
hoFGRvZR5zborbloVo8qhngyyVN1TfFozGJE6tw2v7Mfb351lEA46mpSOXq6g224HqCyzSHgzwVH
K9GnBsK/QRhBhsWARKAfdLxB+eDs5JwB9CLRD+j3lPNO7hXe/OeolRG/TD+5WV20LdvysYcmKNAi
CmxILJH3Y1PYZ3D19oWSHTk0Om+NV3M977MiN2ZlitMNDM+nsSVjM8iumslIqVOcaTYSDXi8hTx+
Jrwm9OxBKIOsUSBN5eAXZbPkgBbYm8AwVsULPQe54PTNc5ldmEw5HOmLyVqrjMXqNZSadQP5Nvnn
logMVCZgvhOdLg8BRKECovQsnnWIEKgPf6wXCOfF22FT7fr1W2ebz1nqWTk9o69oXX+2XThtPAg2
mLTVcQB09drn1FJPdQsMZD3P/QWGWnG1E/tTy6TvqG3eEUM4DitdCyMVCvTywOm153ShQWTXCXOS
tXdiM8qSg93SBQuz/Ewa3YglwpvQUWHuOuQCUM07A+YSmyeZs5MfenA0WbuqN7/ol5dY7dF9W/2U
qX/f3oorhmTugDBAoLH2agrYUkGkIZT8zY60zsI4pvwAGP40GQA/jCu6/54vaXL5q1cG413TTY1B
eHyu99f3Is4s18czT7+EasONfgX331BKqlUimD0jxXLpLYQqEC3kWlOUCsk2Y9C4JA+rqzqTTp6N
75i7TnCQaWvH9b3CdO1dCnyKFGYkHleyD309XMIbhT2RVCsFsOtILbR/RE2J1qO77JzYZfRlOwVV
B1zcAQYZeB1rcJy10N3SSsEDTs8Nh+prLI1yj61Pt1osaE8tBdE7Wg4ji5hHoP/oObI5cZuvDm2g
mdDdVsH1Ib5e8aRpGnjZvrJOYJaRTEjI1zSnvN3qcF/UTVbIJStcedZUU8bCCQwA7bUTPtdnz7b0
q3yoNXotGj4sqt5KMg1+FcxX3NjN3x1y2i6piBTXBTMIrgEX/rwEzz1PjHGs0y3gsF/uh9C6GS/E
dKKY+giGhtOUxeiT8psg1Px8PAMQhQ945Zgat0q5IOwZoHbNtQkC80kntxJsU9J+oa7VHNh3VKYS
+LA4J6JmKaZJPV12B8aXHa2N2XDBvceejwSo/6JaGyyDdpgEcHzOBhjelccrhsJZxF8e+Ts9ydF9
OjMnAfBbUMIF+dYug5egPtjR8NhMs9AHj1ozYFsU2Of01jE7TY96XiJen8+brVdlqBNZzJxOKIxJ
3Isx/52UOOGrYCrXCySN/3TZYj4ppNJYxDS4Yrj04FcPRiMPhHjatJ1Ab/doQlZHEYc8xBFCYcPo
Ueh5WQ2cM2rw6ivVHOqYhcJB5Bw3T8Ql3amvRHa0fWKHgXIEKvJgR1j2CBkBlqHi1VjnWBK0JkAq
HCQ6I6EwI3dThx2ntCDY9g75NnV03ctDu7L5PtWHtZT+DyLb3UWiYO0elH8sdDMubDNRLBEdbo14
IZQ5k8GdvJhYH1Tp99ET4E6DJnMKkSDpGdY1xBSSrKZbMAJJCN3HXY+GZPARhoPrp5c1bIOgil9U
rSI104GePdSsVEOSQdO52ra0gMO0Kshcx6DeIzNEgVP/7Jnw1VBc2EHNnjTvU9F+An+rx/cnBZCj
EvVLtnHCHrHnXqe3CeVtMODhyobjT7vrPglsKMarKFQCqkvSyxsT9O1O1ZFYk+QtX0W7TSLK89aR
LfSHxIU+206JLMvT/7dWr7CMrgOBW31RcNLGvJrxYzTuCTcWPbQ7CSa1dbjysQGNBUEr/2tDtM5G
ZadhQ4VfrBAey4L9CGSgYNGjey0/g1J5PDAqAtrEyxSYyQs7STx+J4/U+v872osbRvVt/XysXw/x
hYuVDjPDgbrw8rY3X7LymAwQoyoKZcDmK6G7MpsVcQeTsRY4RWzGKdyGBDS/1Tkbtj/L45Zk9O4Q
K3lbnbxCoaN9xkjkX0HwlIofKaAv+Xxe7K/MWjJcrDMdezWBsHbvqgsthRj+Vh5iBfavslI8p/LM
OW64VpZtLKK/fyGlrSK/2YGAIFRY1vDZwzalqSNhGpDnC//4Jz2W9LmgoEdmX2cRzoaVETwMckHm
gL9QF0qwfgfVKSNWvTUXuqonwGOrRlCOEtyWd0DU2UYbCuTQCykuA7MZ2hYOmX77i/5wJ4eWz1e9
AWK1KBZfNlaerYmaTNE8+syETuSHuaKkv7LaoTION+qpIC9UCI99tJjv+IkhfhF2Izm7vJAqI3eg
UtExutzkagV8an35sJmjGmhBcrKyxngFrZsLkgb4zkCKYzvCkXAsO3f2l5Xgua+TbzDyJLyLo+0e
Q2ptfAVi4gxIcHqXFqVO5E1GvvQB9DzrvI08vsCubbnAgZcXX3kglg5Fp6b4TkMYs0EnmlOeANSu
ZxdEDiMkp47qcb2dXRPrdOJppSsutqxGMM9ToNpEYJSKAAiRzRjJ9F6UOrFjqqLPpUlbzzVcXqiB
1DpZr/9nuQLxSKb6wsaWLhtJg1eulRQ3+PPWrb8vs4hHKunwyPsz1CENt5Zee/QZBaCFt/b19Zv1
HAMdES43nMtH0rukmrG385zuzZKUXJ5/silEu/Ryo8ZH9kvbeMY+Tdrq3sR5Vmr6Un5T3VnLbFPv
0nNaIpvrVDfOhYVQoU+PoYE3AIKLlrEwOVkjIaI1C2tWAohzKf5f8ZUzqT7xW/O6pJNV+3rTUTWq
WgEeeIzVPUf+3ZHicDumhdEjzPFix23yJAK0rJnAsPbWxkWTMLOvJd5T3un3dVc97pF57MXSMgrb
2v9iY3nVp84rCoais6PCy2MO+Bt/rm3yLMr/WPTvBwMG7uiUF4dwxuA1yFrUhfAQlINqf0sfLeQr
ejinlgaHStnVV/xatWmI53P6UE0fex94qfzmG1wyxmbszVVkY/ri3zRbBhP1jylllQqBgr6DY1aq
PKL27kvlUBI28JLDE7FI9B/5ksU7CrU165ghXBQ+GFOdmEI5vmc57jRL22Ge9Z3fu0OagyEUj7Y3
29xZspgUp1ZQe11+V08fbmicvJvwcD3gbrpo1ZJNQ5W24puuSsFBjNCwpwxAQ3+JZ/GrMOxTFr+q
bn1TyxiMLtScM3rhhD2N6V26l8WUr6NAdjBXxo/aoQAc4wnS9ZjTLRW6fToGfvYoT9rk1VkFc9O4
iJj3gx5wz8fjfxoV8QMlAtHsCnbG+AWX89pEJVyM8LvnkaQ69y4QFhkVymrTnSsxlG3liSeFwcis
3LVzmqerZ6PSnN3EN1+Sz5kOjXjKU/hXxJLNqLWjbPHvwMECM0NKUB6jHd/eG49tGU1SomtCu25A
+68C7JmO7zJ3V3YEnfXiyonT9yZ+8T22JbE9+GjF5N8+ns1++L7arJJfV+724DclZNBhIksTpcgu
2RiEuTjXQp1Tr6uJ3CKljO03Igvp4VJ7i7KbQpgbmY9Mvfdx+jKMp8YKZPPPQmx0UWCOsbkUgJMY
h8ZAK1jTeMMCZdOL0DjzPjW86q5xa0zWQCTjL0bzN6S6R2yKozo39xbf8E9jWBhdFxXCOoq0RbGp
pR8O5HcBnhYXfaDSeB2k9kmr+Oln3TFIA+rFaq4LNfwfFMIJHtMyzM7/y4N/cdRoUwHU5VtfqEWh
o16XUZ/BiFIW10mANE3wBrxkX1bxOcXCTdeJJ2cZMQKQTRU7ZT/l2rkOdk4q3jYyi3p/nnBrk6D7
ZawMekUjz9lVO58vMW45ZPnr11WJWgKaVDJczOU4VydNq6FbKR0zZ/nKEfNpoCBtyVPfyzeh5Uj6
36QWwWFdNARYUVa3BZXW8sqGGTGJv86r/kVHd2paPOqNlY1r9HCnFwLw0RBSCkvAi0MGqh4pVt+5
Rwk7j0rdmKHtJknB62JxdXZWxeoUKHH5Mmn4FFhX6L+4EZZnoITwvEuTyLoFBzc2SunlZEyRtNz4
wZxMLM43C4R+YScaEB+G7J98Vw+5UMd5eNREN9BrCpPyL9EBmyQTBi2QRY/uzWtDBD0jkvnDydF8
ksGnekE1Y7SHkIRmMR4B9JKE+OUCLAMw+4zpNykwnlr8ESqp7BIldOLud3wi3gFkpLVLg1KJ4Qf+
OpR42aa9wsOaV/c821cfxdOKUhK/PvFH+sznTDI+1QcrAhcQ6vuO/M/h/nupyxZqCSWsmWq+Uk9X
i6ZN02+cKLaqYhV8Xg7YB7lzyj1/I1Yq/VsRk21/enSANUPvtSxA9vcInIwRj8+TicSSKkkd1vVa
QhW3ZtKrll1kE3iZZnKju+F+tVY5mdsfd/j1GVEqSxw5yriIdkXCntFst3pEE1xLUXaog7gL49oj
2jZ0IR/JHbqnoEl1OL9WlEKxmW01hzf1xCEAt1mBQN9Jikh5zJ7A0u2AjvH9c+XrWyGVoVaaOhPp
x8r7F9Wv65Y6c9BUNWZLMsC/EhHur6VYA6zp/fgbT9lUUXCTbvqgd6Ge17Tv7r0B555rhQ+Xh3u5
12fhfe5gYnHik1a5E6MGmfhVSDLtVJL25jSoBE6/31Ji1cSTI8MulG1r5DrVpOdolMLD5rdOuIqZ
5bES674VJy3WfWZO4RAulMaD6e7ykeT6NVqT5jTPAVk+a80TCf33oxeM/w7czsH0kHoYmoI0lXqv
qe+ZsebzTMe937EADwQJujcCkFXCjAVBr9OyZBsgA3TB4rEW2IsvRsZHiUkO1ap1+xrHSS1uu3Ig
L+3ymVFNf9NvO0R3l0Y6k+qFkt8oP51yA3Bgx26f1kA6D1N2OHloOPaS3y5AE8DkHDQsuCKrUvFq
Z2SugH6Zwuum3tI8c6gwDv3eHv27uFpprsVWBe0OqUcxfrXnMTSC7yt32CORZSVhmI/r/BUKqP5P
77T83fvhUNjoi1KOPGxdtNt9wv32NYDJ5CNcGCeyBKluu9Z2r8paigItgx2FEVIi5woa0tI7VqpQ
PAyKsku5mgRtZP6CFCQyNOTutoB117DWvoIFRPuw41YAim1gUNkHDyGDgMmeiHhoMAZ5Ul5uIZ+G
eY+InAPTD+rQb65wy4SXBLhlkzNzHdIuIgL1qbt82+sfB7o8vvJ7b2NRa37vYr2PhQ7SVOHIV1wJ
RFI+jrnh18YlpbA3y74zOrkLqxIjFYZyApWICYtzzwNsPPIQ0HFEvomKuWJjqKu2v6/gLhIBqDFd
d+clPw99UJ55hR2EfeAbJ/tIVfkpipQ3XmnitQN3eHD+ZfNXT5Wwdk942wSv+5owX19WUYavEy8n
yPVB6SAjpK4aXkYd5mR5Z3hQEZWT1byLiI1jLNTJ7Hnz/lzLbgb9PO4Bqdu4XPwf8bA3bF+c9CiT
L4h0gAywGrMmHuGf8ARE2wuCP8LYEINk+G27tVqTeJBBEZF+wtaSM58/rYxgJ1OTLm/IVzkuek7C
1y8Dsvy5v7N9aAM0zSUoWZaPrmwIo1PoKslCH7qPp9SI0EOOXPMu7ksam6fIvVnn1rbcvox1TE03
0VwK68ObJksOxtpIWA9Y5/yLyYjSXK9/xhNO0cLVKnkvp/p9oQKhmMLEAQH0U8yYTYAnGx28XzKu
sBq/zBDNFdfSy1XrmxSYUVKgPAeyzJWuqKoU9tMkmXaBnaPEsFfVjvJkoOkuiNcu1khpHZrZoYFI
zaQYBz+z0qfcQVeoElrS14eyGMNm9eeZ4VlDwWJUkTl9X+bpXN/7VVMU7/zguABdQeWUgm6iT1cy
/2z6Ia1oeGVys1pPJSjim/9VTokYPF52DHCElgFS5yd8bp+bzWBKYZFMczYpojXTOGV3EO66HVwm
9Z0Tp2Cf8585cKE3I5MWPJ+lV3nx1Rt/J2ikNiNRKzz7Hceh4N/TV87e6Ftohf5uZqGYN0qd7TQi
43TBf5Ij8ipEK3CEzzfejwi+yKSm5RL9u/kaI1X9r5rsk0LqbxVjkAgPs4g+wlctrOcJLth23Pmc
IuCmHC7VIsj5feqjdMqivLCAzLkFvdDig4Pc+f5A/Bog8iaYXNCc+T/8WWb0IFeB65AV3FCRtx9X
TPkD3LFhh7wj00ASHjjiBLfJp1sWAZTVvyOPT8jPWjpR8eyB8Bz/iujeCwaJFbh8nisw0oU2HS9/
SUDlgm4s+Cgwl26p6HvEBB7XU9WVMJUKiNY9KYUjWozFsYHcKd7av42au7WvpVv5zejwJWhSxD85
oigEsIidx/DdSFGhXOSGc55M644SD5nWZjadYtHfqz+wXwqY9OdChyWueMUmH/wT3wnF2gZjFdja
lJduQUSUBWEBMeTDNJOflTMN5C27b3ll/+xlFOcxQ8VcYDEeMxenVojx+ymssCi5ZDo4DWFaPHhJ
n6bIN5xPnjR/VY887T8G4N4N+aRDqVdYlP7rw1/IuJrO+WV8NJ0a4FT5fUVga3uQ0GbCRvwA64bF
DHOHWjuRXJcRpudG4Qt0s6z9CZe3aEr/6YNM4i2GnwIvZR92xevRofhO3jIHiq4sM1CqX42DyTd9
mYL9B6EcSqgh5fjh/h30aWCzXuFXbldYAZwFBnXq9Iw+pavDcad+Ph7frcjl0kxAU5fIGqiSmkV2
gYuyP0EtRJN4q+e2u6pw28KMxQIfxIaL6Ll0sCt5YEXaiRpY3FdHum/cKOTK9hPnFLByw+Pgh74J
grofd8YskrqPXtd7mOGcIAWoWrDzbi8XjHA+YgmvEerkVRVw5sEOaifuUXZlFUxzEzaGl1t7V7aK
Ag8El9KeRIUrmBIH7XSWEvc8/Pakg0iTV3XHR056S7RPS4rR9DpoeRnCskfMHPqIaXKofakO2o7Y
/KHhKLLNaFy1RB8tMGt/kZZw0mqBjxN6FPUKgMJLIEWv+kwJPdwGSB8ybgt1LnfC/Oc71nMQdTmL
diSD+U6+S/1Bm8RGaZnUrd6CwJAUMoMZaEjjAO382NgLJvbR1pR7VljW8Doc390OzCks/WQ2U5He
pKzfHZ/BZS5T1VM9XvOKbhlBdqFcZYYjkXlaFv9+bSzKgZ2Zq21WMJFkHt5LfFXGuMqwIbWUXCmg
MWnbsXKMTaf8IAdx2/HofIQVNcYViRc3OuMfIUtLkkI3yJrpt3H2V8UjCpup37wGs6LG2MUzxkuk
B1WUh0gjjLhEpzN4XIy6RiQwNqJfE1w4KKHdd+G/lNXn8XVutKorM+RrxuAX1jG7DQ6iaOyQIE/R
NlLL+IsYHgkDqMHCGxt5vnmqXf3xbgNt82tQi5o1vTiQeUpkOxfbn7PuvPmgoXCa2FaxQlnEIqCn
iit88rZSDFQWHHspuC3snoBNTBSeIHizMoqANVj4kGME3wZcp2yvYk1HvgewUlGZvjhM6EM508k5
SD8Wdci3K/N3tmBaoYHwrNzjsg6MGtlrK5i8NxoIiUJu4LvlQ9awLzwRXIKtN16yDMUDMw+2mPoB
nIJ1QjZPtUXDTJxkgTebbrqnFK8l+7aaXUGg6QvMspMvPmzIC4JN0jKZhC1jCQyVTL9LzQAgInJp
hp+8HCK6Du7Mminqb/QOIyQz6HJWtoTuKKB3qh7ZoOSCSNspP9u7bJDUbfxzKjrffw8h+f0tsZLl
j3SxpZCI+jQN7/5m7FmmxM9KL1TdA2LbWeglL5S0at8mKlSEQqcqQZOufRq8S+hqspoWr/EDAfzv
0dK/rPO1gUBJbtNLr91EaW4zse+5i1VnU+EqKJCqSvFNp4hjNc3Lq82qtapKNJnMMxuEV0Rot1jg
tAcXSeXvGwXgZi2sJDi4IXgphhnXaAvQcKB09vZ61SgoOBGUeGpy/EzGv7e4SZbieH5MIaUDJQCd
R5uOL4bHGvZ+ryHDp07jmCe6H0fRL5mSj9gljSnDY5AP1PdQYAaFv6YKqHg+mYTmpCaeV7jKCPoL
3dO637hjGZaatTGm8uohTA1Y32pxBwGrJzePwtOsDuVu47siwqUhfj7EmHMoKeSSoJeo8gWEBD3Q
YQyDB9xbqjkbC3uVUHFc+ZcOaT921jVen1WPBR+9Bvk2yLsNpVwzRyzrbuMcUSiBJ9RKbwKXrOWz
MxCXUAJx1aKVm1LA4xnRnaYgAW0xLWhbGokp52nuPPjc2zA1Ws9yWD/nGO+faSYhIuNQebpiEYjm
lQpj0Z9/QyrQi5/lRPrhNUnPpe0efs/K/I6DPeAnYS/zTcb1+UnsiLjuLY55oEIQsWjQRotsoYGW
YtpIClSjfP1zC1GLIsCvG8N65NApzphh/datHLCGe2Fhut7hNlT1GouEZA90+QCLMpM3Bf+GfYSc
C28/wxYlWN1liAJvGB52I2J8wn15rvHX1BynIFvb9MDph6bKVFj3G3m2KV8rjH2kJpYg9Qvp2j1g
khY+ZXbNEsoLaSV8V5LvumlAYelLt8wi0v6ZU9pKX9mLBGjV7PbT80FskMEdlZFE7ivcAqmTJmMU
Sag0ZozHeaXX4fEzYZ/UXV1uDRNAcyNApAdmJEf5hhC9WluZ+8WND8qsvoIoXYqeQoFrF6oDx0kD
k84UqYhwoLRofB8yxKninTxPRBlY4JFBFdfFbqPBA7+yALGd1Q1ufimDVKoSaqCYrwYf0cKWuPjf
m+fVlkG2WBnY7vmhOJ0W4ox27BQAuKWApjYyL/pkwq0IIuz2SX1hytj/7cpiVSbhL5MD2e6Dynrv
w8At2cKwJYbCozvP5s46f5g2u2LkOyR3VCye1PIfOb5ZbyS9PUDGcW4v7YcLX/fCOHDO5PvzxXjU
5e3R0tZIxFQXQ6dffltNtbvgCm5ZTMNJY67HvwYFMPrmv3Yi5pGqa4HZPUg2X6TWUTSmmQLxivRv
mnSjSVtiF+hVmQLBoMTZRxMHVRDv7ilkvThabzThNe2j/fqnksho4woIe7KEkHZ0tNBNhFa9JTYi
iTU2JGAvvvWdmtWzyY2kEwL/yD0a11sQHyGZzgUO9rE3+7lkpuEbPp0ugj4BKCew6848LJXozkez
juq/LMchaHruCVfGUsfPZIQFm+9y58jkwoJ45kMJXmPd6nBiJYGFMoV690DYD0OkjdQObwKW0dLb
PF/LPSE/cRw27dXg7mNMva0Ct3C3LVp04oDpql5/bpD346GmWzUQ90ZZjUZQxB9R8KTsALsfNkWN
x1h5gZIqxZAYspKFqBZjO0dt0JkFyF41yisZB7GyOxX3wANud0SkPYvuOWL/E+HZrA3cbGj71FSK
R99MOGse91tEnbyDCfhcXhjQkASPBnPHsg0pfz53li6Xd5L+fM+1rcLwihmKyG6CYoPALitJkjF2
ymq1mNOZMNXA/PC5PXMa1DFJjVAvMnQlYnqf4uLCVtGvL6Q0Jiel9SPpygtbNK3ubBGZza5hrtch
41z2ZtSUPRhNE2EUca1FSWHotWkBIhzfPeE78ChdSbSUS6n/wHrqQyzDZkSf0gSEkGhJfoiL5v5x
U/2AWGbGEd3Z0c0psG6r500Kalsyy6PkONo3MK8cXTpzfPojMGqskn92qFFvu3NH5RlALi4OxOtJ
7eepxleOy9dmjBoD9KyketoVanN6m08bqOXoK/k3g3UCnkX90rsdQyxrflxSg/5U1JvcUemivf1Y
tY6OelsIJ4m1iS5zQHPMQhs3aEqlgrQwxPiaBVzg6zzMLkHGnXk1uzZG7ICkE8stWSr7wsd3Uzum
RakOvtzr6Zicrj6kXqhEsViT3+kTOQO9fnVF8RDVojy9wLWP77SNFCsGy5cC5diQVrhKGt/1yrRV
CLDMDmMRPEB7p6CSESUuAtGhDZ+o+xDPTRiMmgPRy7QpCsBEZeLKn0v/9vB1A+vV04580Br5Iktt
9BEg7JLQGJ+vTN1spQcYvcGoFOUfL4FciTcXbmIXlERJDbkJCEOMHtKxmDCTWi71CnA3nAKv4Sbw
xnkoDkQxXD6caNTa6WAxoVyy6kVn1y4VpwsIcq8MBXqs7y4RDeU0YDuvs422qNztdwSn6p9Fy+Le
S4OV4aYkKA0NUcmMo/Fph/yX9irdC4Dj9Pc7famdvV1mqSA274QeTLV7pT6/DwW+XLkq0BY/vsUP
wKWdfYSz3N5KC597r9mNo7B8kySrhrse8ZTGHdPbE77O7hmrFBhInzplqB5+puE8YQiVcT4IF8Y1
NMdmu0xfm6OXc0GA4ia0v6LE6JOcCUCL761YjKqKdfwmYS6AiURkKxU6rV00izJxu/geQ5+Qyflp
+yfBy1S2U/gus5ERlfHQi2z1/r9lOBcxkWIugM0GSeGcmFYVcR0T4nufeyaOyQqik4QRpw17JFLt
FnNhGCX8UUUPSZH1oKZjB1wjVYOwl7IKNeG+6ZnSM+YvFGQiosTdX58B1orw1A1PjN0tq7/Q7shV
c3ESm42zAvLaASqdmKSOs9oF2R1HvjihQO13uwfwwjZt/9KdQvACO3zN54pCI6ldFWJiRpjMuKNI
McnDM9X/R/xVcME65CqYH9+lxzR3EzXrREoVO+8Yfx0eqR9rOn+K8GIh2gWOZfhBCxI/NNCqRivl
6zEvDqlWCuogavhyoC16AWIOulRaYE1x5veYOSlBpoZ2tyK84ikeBpZ3p/9SuUdFavO2XNyxFSUd
YeFA1UBvnItUJzCenk/86dgcBe3ojE6fWczx1tT68Cyhobo9qkLsGnplAgvGNpbgL8c20iYL8bsI
GEM5ieo+RPcUq+vpgL7cUZPOnaiRkfoOjiKFsCP8nwYwqHXXCX6I4kRXgxn2wmnsZ5yQF8uDpXET
7HYzRxOBR50YhPs09xx8cC3jEeA8NQaTjdq/Tk/T8umfDg44G1rRaw6YmYOl9XaXSKQxZi9gHcHu
MIDP9+1e6wWrHb+d3zSXocmZlj5z0fT6sQJrDY1bXkedUTkbjWBPs73GUwANYvzys9Acd4a1UydC
ixaIrHAZv3TGwocWVTCFkIpUDCoykSOhXBW0h+9do30cNxzrxVep8+gfoZVRYr3Y/qqT4k8gzoES
eFeXOkqugpBa7Ljc3ZUltWc1nKdufjjHhB2qfmH1fzvr1HUni66PhBMamIsFV/lJGo9WILNEqtGs
CtXp7EginnXnTJg6FGfIIT78t5OEzlVz+c5hBj2ifefOUJkxPSfmDi+Jhse/WHuv1iKFZ77prTp1
7mqoNso0VuHSjOmBSYGuWCpJo35BN/LSpwDVvI4zxGR/oopLw/t/8WIMIdYk23KEQN4e2jjN+CGG
OPtzzt+K7fCNdFfF8cDi2m4bjMKFHPHIK9mGhBbVBfEZmZ34AG2Xk5yGn4aDCU9BfLyscCAOWYYI
12vXfJZLIxIZmnZlDXIpDT63FWp4RHXG1naQPZyurvbDMbo1k1YmgOYNXc9mH45LvzqGzfkJ0B5m
BT4gW6v2s6u4wy4nxCVqj5Klbd3DUdaLAbX2K2Lac9q4qW0KbkguEKktqC+U9bXagtkVUXfYl7xC
dIlws9VQ+ywEMZrjayrMjMstlnIhpNa3H07l6sx2Co3xKWcoVJjowXALmJRjP4Ov+acDG/soJGKa
Hp6KZTjHe78dpPe0D0ukB/vvH+ki8FftBK5aF/2/xMFRVdkWp9H/ro58seoK7jHmP0wNIDFK3qHD
kUUhwgBHL01gVzKqMUmGKX/5yFz2GXSwdvmSRggXZS/Uvcy5fm7Kmv7YZOA/wPA6YfLlp4C9jYQX
unt0OpfNCHTFNqMmeBEzjKkdfPrOCMfEbUgw7Vs1w7GM66RrV8NRWLtps9M0JlZMXMtN/Oa3LTXx
J3+9+dx41hWEYqyKt635Ha7jFbRWI8aH/sA4GP8u+jBetDaz6MAxrVPz23/WNIDKbWHk92BxqL2e
2Or8WOE5jAANPRMtGxVz8aa6Syg1x0UkVCJJIwl5pzXlc5wd7/11mL5tdfFnK6oRGLL9G/eQsRQL
qNeCI2xNwzwd/ZJ37UDXOg685HgKj5DTFaMXUtd2lSXIv7E/Wc4eMv9AqluEw+rKFvezB/pv5Dpp
tEKaGNnvCico+v+mLqqpVfmAcWBLvs+T3nfG04ExB3PtK5g+lA6iOvdpLMGO0NVTKzrRCFSGI/kH
4aKD4aIzEYglfsRyK88ZGE8VCutyT0R4uIu4GVNIBDakbhIAtHAO9pdVodTvPIS74j5sfFpk7W4T
1R7jPUysFMBz368DBQlVBzH1B4CntUqkuEYB8+lMnhc1ZjDuiGXerBDFJf4EulHt/iQu2LKEtxtP
DTeX8NbZNz0srQio2o6Vn8enl2lJTeDHBumMr0PIdp0Tqjw4a8kOYLbJlY1X6GHdueUTCttycjXq
V1rXuzVNePDD1yaeOPewivrgv+WF4KO6KFDfhkpggvfQ8AOL5YZaXYF69wzuriCotlfbqzx5NrBf
DaWqiS5C/XoGcJ76ogZn0audatdoYWD/zlI4ipEwjQQJyB3GayHtjfJX4Q+5zm/sFfoX1zLVCpQL
xxQOVSH0uWGCrN5bOurAndoAsIZVQnDpbpkdxcgbK7ZTafqLsiCJQ9QAwhYXeZia0WP8eaALYeAm
q0teauPP8nk7O3HYe2A/TLnwn6X3/Wq14al4JTTWiC5mCLBB4AB6ozpnxg5zB5Qt/oNcb05PEnjE
Ho1H8S07AQZ1RnKyprgcqWVRKx+a2Nu8b2jRjIkOwz0/pzlaqT1os4hcQsUHvj7NjU+g9Lm9I+Y6
eOM6ubeO8dEKC+NPu5S9mh+Ep3U57tmkQRsPOtWfvCoYWhPA8CYoDL1orKBFd9dPNkOgqMmjpLNa
xDxJuAHDqCAb7aiC04slhPJG43vEiT2MK66u/XFkQc9W/7TJap5H8EZpBQwlDzEB/GzIVYMJCWsK
FC4oIV0X7+6Eqbnap6zD1XMu5KeIGgwOLVkPYX9TFGs/sBasYIsTgIQV3LbDoTH4uuoYEbXqmmla
B9UWbiINPR4wJoJjLup5VVgm/DT73MOdMnl/vnVuOYuf8IokNJgYQnJqTc6CJwvpooAcR6VxYv4P
g3Difgbgj/aLe4tQSBw1fM053y6AyAWwnSazhPrKDiHsipomO3dbTs42I9x6g4KacY8Gg2+ASkjZ
byWQa0g0kQ1R0VSwEU8Nk5Y7uxqwlSiQfvUOV0h1JEoHdNLm2KkvoKEOki2T6lw3XDBSNayDPaeY
5hDKRkCgmq2KkQD2o2LZ7yVU/YTXEzsK+FJseLZ/x3YMc1/6RDTjc5CZ613aNd5b9icVuziF3Avq
lEklQGVPx7MwNzn6TncQyiy67Vfj23tK/OeDtKMzZ56tdEdyRi9XmH2MMpj9qam0UXcY+UGhyTb3
m32f0ZgGMHmtfO0+blsuZBEh1MOfi/K/Ssk3l1NvwbO+AeonS3GndHfge4nkOyH21JUb6hqi2NzK
5ySpH5TH75oKXYnp4Ca2x8Yp3pa4iFBe5jJz6otz4xI0ojcqVSwFEwIYLt3rrfxwUMQJCvusQvhw
3+JMSN8VjIMQqpGiX+tyKevAA5Gbx/IUH4h4o1vWDQi7eDAZnjI8efoJgcmyXD8fnmO/xebKyAAM
2ecOdgqZss/88XIMfAPeHMvexc/MNmA0NyZSXUfQpmt1F6xlLsWTPy3Dv7yxw2Ohp89VBMO8yQKy
1gjXuLjqPM8dfFvKn8/SdWCTfkya26OVWQt6DcqJ0ZHKTuNF+RsWQ/m0oVImoEX/QAzRyBgkEczi
Re2sYUPYTx8wKSNii0wnooET/l01mYIHbRQD5hw4Td5zdqAOnMKAFIhV1BfX7nTbA0zTKPWoQO/U
U/i3cY7CcPruClv884TaGZuFdGuHLY2E7aPQ9jCw1zjEw4+IxjTmeuo8A8NTCjNnVsUMZ6C30R5h
mYDesK3Tbufl/uIGLjUA750H0tTLAQCHQtLu8XHmoyb+T9AydwLQZM3UbDVyqWZyC+n3DXOKnAMV
HaQ49fEJxx58gHRMwg+i2vfm/y3Ho7hnuAdLzEFxmXSnEHOTkpXBMwxvMquDmWalbGySOYolmOj7
kc/nnrRsAuCdRDz/g50MLkayNfGu92hwSGDzmQyFN0Cp2E8XjSRfRu+khxOpO7xNgsMTcnartSk0
lOJXEznm7/H5P7xNbYZ7EPyU0m1WdYnqPPfd2da+5Gyey0ZY1Ka/rTNvd4kQWLPFzL3VhDzcb0un
0s77XvQvMsgUJxkcuaf7f3KvdvJinupTNX+G8bes/3YVgO8MGGEMwLohx5gOFsqqVw1NGEON0pVP
53BYXHDfi4IWz0sk7bpE8JMSx8iBaF7A2e3dOJR6cw/0VzO5dNerD0L2SwyFsXkVwFwtSYrRKjyQ
EBHLLDt/jm/RHEF4MrswIhXGaiq55sjfihxr28n2U8XoHfZ+N7+M5bepgcU2B83dmasRhqEslaMG
l+HLwKcpivSwvTXn8ryq9EsR3cNy9fzaUzBB1BgefNZyI1Bwwe04C18tBhCkpHwj74a1PMLiz8Ab
WI4gYIg5qVN0eFzcamM/NvFAdqUEUdWjCBSN9JRFrGdNAFZUATlIUvUtoKvSDApaobO3v0jvm2iU
66FS02WIAVmuKw3TmQB6+CCxITPwlbxmlw9BZge+NXkRPtYeb6mvd/034J91+zh3M+i7BZzS8vfP
g63kn6jDw4HYiD6kl5oeLW3475WtXDFzwthpOMXuk+AEU0qjn2Ti8sV9HdpasIHbMPiIOUpyiUrm
AdQdZdGdBtanQvDmH+R5Ng1MJB4RPvqJzMQInDwpMojHze9a4wbhgojaEcaVXA/KqcNosaEZmjWs
FSNDreQQv/9jdSn/WbdTaQ0VyzUXYa3mok0eafy4jxCeKGD75pmX02Erci3KKWordBnGQJFlc0qv
8Rf6qXIchmoiv4K2Zcu47YCvB9BltbJXfHeqAe6QyqIVTzAOJM0hbvzGSzE2lWWObkQpi/xxgGHG
gz9Ipvys+Kx1883dW1Zsqa1tJHFFqIdLOBaQpODYBmarG9tLr2pCWT1wNRWAMzLViXZcVPyymlsu
Yv7Yxo7y1iBSqNzaPJWUJ795OBnqalGfz4fEUGLurbL75zAa+Hkp6rhfVmGtlE+mTHdQPJhnfMRW
JxEei1445oUrIe2Spdzqlxy7RhHc9xnXwxKkaU4W2AxIQmEHlj5YsdDFqeBbfgtQJ+9ovzTLvp4C
6lR2PrT6HKNmMZ/BN9cuQf81ox2bQsKM+dz4nkftyXocW6f/cG6mU2GKCrZTekhweplp4SXWSPrp
NnLzmojXNCJZO2KV3PMCFpDlPdPxvp59H4W2kB2bKYHeqfW2ZK5yYFucHePcrg8xMjqPHYHL3qFh
zaf8imtFruakN2Pf2Un2q1zfkTOOCNk9RvJeTvWXeET7BElOgsV216PhvmVsAJUmmgchM7Bem2sk
phz/pizwSxKYTVQAuX5Ij1uzzTMYYT3cmK02tshivogk7VgL27e37KDGOz18cbmtuQ4/ww6p5nTb
28G7PfYo1Tj2rHv0F3d2N5xppf3Dk/zeK8WUuDLp6nzRMSM6T9rCV3qxIOEmws0aPx3DRDbsyASB
KFOQEzJiV2U6ulvnBqY+eUI0mK7z4BOc2dS0xYatjZ2t+dlAXdyuu0pjxOeT+MiUyNnlSpQfaSxu
e8+kmxXt1VoNY/lUu1swZ3Gz9Lu+ZJ5cFk2ExZKkBSgppLqoCjuES9aWLD8t766wwQcxei2UDuJ2
Wr7XG7rgazdVWedJtdlFYJQKrEYm5IK2+J4duuWk38JnjH5XBQFz4fdEvsTQBAUy025cW8KlnZjB
FMHaqaY03zfg0jO6l1RBOqtqGr6arPSit+fAs9dloIR71sMDGxHiQUacZtLZPLUSMhzySuQzXemg
N6Rr8/kB3HZf2mLMRzgdTpPBolKjGr/FoI8bkBxuo7Jdy8PM7+Ysts6LQBgO/evM1pemJOSLSPtM
jTRxzxfC0O3KibjdZ7L5pmxx3Tf9BiNY/Cw3KKA2ckl9KW6mpyTGzFAPd3uMFtlwSjAIj4MGTI7F
m0N86uY/hYsdGhtGuslCdHNCaaOseP++sEoFeA5DhYatelPAQ+pC3VcuVd3GViWJZ4go8prDXYQ7
Emy47FMdc/v3XkyQZfUyO+rL4TbwpGC8t1+N5tALIW/p+Hm5FtHiyOgzkTjlciYKbeISIp+omLws
864NvgbiXmIaTPiatco5iT9uvWEZofI2Oltqy0rgFE0abLiRMiNtx5A6/rvCMD1K+bW6ZwPdXpQ2
vcKVYZb8edQpxb3hs/DrNj1xOq/nxfFmDLTcXRjCHP++7CpbHY7Ul9zrZLJNkxG+Cr7fXwZHMyV8
38h7rSuGJBTRwCduyJetHS63Hb4pO7UpxnFY9d4Iyx1fv1VCEeD4HbRNSZDVgQWkaycXHoCc3c5x
ekW2Y1T8K7DvQGxvWjxGkpASjiBRBXF+pdoza2nVtU08k09u4/AeIJz2M7ukXSbhvlr6sJgYqVfg
f0AeGvGo4FUn7ZAcYRppuodZTxoFw8zhTzl9YBd5QtVfnAjF6J7am8oTyfW/BFBe1xePRA5Oxyf5
zGFOwdOt25sbujePUUGkaOVPCbhbRl3NRdNnSvX75NMZ/I4I2y/nF/wNu+nA+yLajB98GlhKRxZD
FestHsYoKG3S0REdgSQbXICKjEZpc2V5rq0n0ALeAwfTQBFV9GhyUVGn08jrZNkVwSuBiHpPKuda
iXg3vhAuh/CJgQpnp37xX0aZaAGa/l1ilqEvwmvNyUVlyjb0D1adVfz5N/7Cx9TKqzWXrn81Qk3t
WG91lIrH9uPmYgAcOO7VybUhhv91nSzwJ+smwnsobji2FOHqXMMfaxQ2V+YSs6AHBCTKHvMwmIwK
DbS2Bfl56cr/UWOopagrbWEAXDVuVSGOcO3cITA08K6BxgwYupY7M8R2fSl21ND9seNtoj2v6FWq
wiqSNWKEylM7Lo16x3k6BGsR07vXu/1kGjQqefIJWpl55No49qivSFu23eqmZDJpWMigHg6PueKj
gZ/cyZoMkFVIah+hC6uU1ANE22ikXzCAEQLv98kdAoyA7TMMDGQ70yfVoAfntZ3mKrCRLtSVknef
xEIX8k+eY/iPs2jYdABOHzsTDJ7uN0XB5Z9OPR/fKfM2jqD8zdOi31/CcjvGRCtTsX4cS2v8WWqL
3JBFASt6DZbOQuBMP5TOr0SvfGEJwJcFmnWvPBH9ti5Dxj7lzh6l7aVSA/jWKTm4P9BAs1I/Hr8v
cPWr7rq6PMPdeDLszCrMooNbIj0TQeq6EL2ooZxemZQKJdq3WOzE9HKc5H/oizYF9FjEy7NYQsPn
wUv2dVu4A7PJ+gTR5wAINgfawGTyePlhdd6nmjdVELiB09YBhaYlXUyS0R6v/fiv370rg0pq2zbH
Sva13WWyExN8Laa21WO1eBwZ8MNV2vlX8C+5FVbjvy0PZWxNhfEos9AmXh6x/XojT7BTXo090+SB
5lnF1dbaB+Dqq2JBqHHfguJc8iMYQ94We+Z2VfApIsTYjKuyd5X2+B24JrfwGXMiqYr6F5LS8QGp
KeV0Xn70dwV/Grl+nb5BtrLDxNAz+1wI3FRC+4qNP6ublbKSjPhhTyVE2NsCw4SImY3777fCHJBV
GWQcrN8BZXJMvvtDsH9te/b1zH8knZOfLtT3b4615Pu97sXc2L4P0+6plop/ry+2e/Gan1FT1X7c
adFkrXcj23AXs1ls5qfwS8Wvoa2zGnaEL/G+eT38qom2OmbnlrYY/2UE2Aj1HcF8nBv9jN9sxpJo
1tb5AzkwUMpq5A8XiCTcBewxYkJ+2r++mn2jbNatLVg2wrfS+8vCX6LDyVe1+hXosh67r93gPOxn
78nY892qxX55NgrPGqCBVIQicEyPFs7eHa0RCCYoBbxNJ27nYWHlokjWNCZGVKS+Xt+FTXFpqB7H
Za7RQyBhKu0qLiU34d7APG/GWtsxy30i7zFQufmGZg0qOPdLB1fC119l3fLsyQzOFuxcAIqkakfj
h9Fr+tYtnOk63moi5jctAvpZ4XAkZ4RTaUOA+SNxzVkW42n3asjmUuDUKkUxCrL0HdZ7YHeDKI+u
1T3DTE/scnU6rKSRUKor/4JXrMaDJAzsNvqCZ1nEGIxqFU/DdMhZdMdi+4MPvAOPpkANGiy3yLfn
DYhF759hzF1+QyxiX6RyYMnAXYS7UGpPfyagd4JTSIOBgSHZk2AKaoxnYnloMavHgN55RxwYyXho
vjVqGHyV14o8PyAMwoGeEISbA0tKKhzl1YVi38C/Y/71QTRGf6fMYVcnTn1vmxmgEFWVdpyzDDNX
AFqvyxZ/GpummEMImPtfFpsGGN9GDyjNLDrbVICiRQj9yu383lq/8mnp48VdORBV616ZV6u0XqzS
mDyHBtZv47AY5JGgD/11sgMphTgWhP2d3SAnkIaIdDzNZ/DvUeepQUE4UiOTcwF79ZJw2mXCaa8O
YjTM6Y+/z2tntys7vRNgHv9hLjbEsvuNKRLOAZxk9TBkQyInxNwSdCRdb4zQIhSccb2sq4q0oLcU
82TRJclZAxTIn+plzuswjvBGlh7bdU0AIDLdE/LqrlP264FiTcNK4jgUsUwhxT6tXDbbb65PCN9i
OFX3T3CM4tMNQUhI6nqehtR6HpKoFr26hVrK1yCNAQ5TIFrQ9uek7qM9R06nyBnRedl4A7N19t2D
xnfXvYFuUDLlAzS21eWx+JDZgyk1n17fUSQ2qCSXJsmQ3V/hQ/DKLnijzSRsW8Fbp3bRUrA4LrdG
eI7Ujj7JPrL4FK92Lkgp65TdKApWWdRau8xHJD9gwKlV3fCC3HAQL5eXIPPenJRhSkUt1ptUHFje
FmljJ+NsyZVHx0WIBxGia3eUZNRao79lTsqH4kT5NuDkmkepFVLMYgkxHfcM5zFkkyEpxCLeQgwF
rKV8giyyzhTVLtlGAbcKCfvvPCrlPIaWcTD9+cwGU+cm5SEmvLWthxWPCn7hW5VdtlkDP1JhZP1N
rfHzRSYsy/uXWWLzSnAK1LchFZbBDUv7gEdCM5i8flwJtKltHoqfqT8QyJbWubDIEq0RPGqZ0Cjn
0yHjX2pD4Q8JREhlqxmRpF49AgxcwoTh0WAPQiwwPAdiDB9DGxlYiMK2jN4Q5/TMcVMcrlMyTuzX
Y+2OJAvaPXS9FAqK3MpZ6TZM6ZJN/2yjz65V0rM93tED01h/5BzjNok/R7kwilwaIWtnNzfhlyuO
0EkD/3KpB2KtkRJqrmny/nSIrGOV1GVvwszBgVvl57ZUYyA21Ge196+DsWW8kVZrUkvwo+nEg3x9
4IaQ+ZSeUXiYGOcRPLyOhbQMECNAdgd9jyQrLDzepfrA05fIYom3cImsFv30wtzc8tpCooO0E4gp
A62lOk7b99GieKaIeocfIc4ug9lwQ7yH1iW6VYQD7LmGiEwPeeKrx1Gs4bQ29B+NsS4spOyBy8Ic
cE/Zr2A0XZDBWn8uomx+PDRadQhtP+jH03jJQcUH916T1BJDWXDi9NJT1pk3Mnp54XjzYjFpSNgo
RLT/ZexV/v8xD+kHwOCkMEppE0hKX8JpO4O03caYnM3zy0513FnIVDtTCSmtxEap/o3adkxYi0W2
37DxdCCxDvHCeMDBWAdNEe9e2cMbMAaF50e7xjgp37VAOxm4M1OyylQY0bv+gKBsIQJtlpPjCIHs
aqH4mi02XWq3uel+yku6kSn6hnzfIv+kNnOjWYsDiuAlAiaFEvPHqG2Dk2/qZsiLvef4ZrE7cGGa
R4izFa5I063YdDsWRnWWsjNkI7SP3BPLIg/7+oDIo/B9ydAOiRBcWjCAc23t7QmU8nW6mIlAZagK
Qex+3svwm90JyOvohQsL8mmGIQt7yfJWME1qVEQkj6LvAvrKIyHfsmXfDo6FgkGfuFlqMvInwAfq
DhBtOaBZVqj1mOQbYyxN7EMoCIvj2Ddfi1kjR6JQFG0l/INLJVV0uZ6GAqeQMdSELoGqwdFNINSu
qAXCSVXjg+AEWknu7JYzQ7XHv4aW1V8SAguOUSaaac77p8gV7Yg09rk3rY/Qe131dzVZu96RgTc2
TKw3D8Z2MnMYjBpopxx657bVAZ7OzL2QGKzWUnf0ZaqAfFwoAb2ayXuqaPzliIwasgxdLYEwYA19
GuNT3i4QUn2YCTbKtx0H1psMuVagxX5wpU8+jOv+Y25HilFDYXADBkROsR3b4WHDRjynJLDXvWJD
/YtKz3DG/+QdZf07xXvk9AXK0lQN2kZa5tIQnkA1gHdf2UXD+Z9ygxlylkJmlpdsS4eWCEazQjSb
QmWgdooVcJBQqIG9lUk865Bc01Q9LUmd/RXat/b7zMhw65jP1N5wXA3szQFh5+6VeiD/li/f6Au0
4UgXJGRezGkYRphppGR6TfJlE6vjhscJnm7tZFtmVdUEzQj3Dm02gU6kEjR0UbcTYzw3kJ8dI4ca
NZZSjRyFuj7/jhWMFEVTixWI3oNNrcqW5NmPBbSeZdulC2t/OgRJYL5NwijymVEQvCDBZiYalOHG
SRHp0zDJsOYSau9GwqhJ2ZzhjA0rva9SfY89jbdh6Je2G7teiM1wUg1R/R454zNRRHVkMNUmL5DD
qtbNd+MeGE7VqYvYBoO32hJdX4B2uWH7Tiw25hqxpGKKTDVv3wjrtqFxGQxQCQeFmoQ3Egv+3ZEG
aa9oNx6kJFBGCF4p3naZpQTh7fDy0cfAj+vsSQUG3uV7VUjoVqeGHxK4QobkCXzXqMX5AvOblAeT
j8cFI83X3KO0A6O6owSZzcx8gcDiurAY00BtAjWqKrem66zYxV0J+vOX44r0Ix6yrLAvOopT6qN/
Z9V1YF1+MCpd5n4jAELsTMZlcttI0evDnPx4bsWC20F2YLrOFJKx3CrHAMXANIshJZIVoo8VpQNk
+OpTZSRy9kyk4sedFgrPbRPkEJ7CCXnSTTRbhvPGxBIsnOd54E6SOZ2SvSvLcbT+WVHungp6wG2T
SFWaxBbvTfHwU3S2UQm0PZN8lqSNH4qUG68H+1KNjSk0CepkJH+XDWDUc6fgEj1xpJsSr44Vy/Mx
K4510KQtOaNnL9mCODMespvAEHy16jILrqNNhrbUi3qkKVp+uin19+8zkA0SCIzWY3g1SD1KFshE
VkqS6XdaRRyjlt45t+Y7XjDfPvH0CvbtFEZBbB3soUHTicyX07IueE4MFbMQ00dKW8YIoavAZjfN
A78aAb9xhpW6KDZsADdMFm22OuudQosklXWE4L88h/vdHdm0ja1pdHIE+Z7fFpW92zjLdjE6PW3b
/mpNWbF1M8e5IlDaZP5Dz9RLQ92Pvwit4C5iuQ5iAG3ot1xRr1bi3sGyhFSKrbMk1UDpX68sC8UF
9Bm5R0oE4aH6T9aMddF5Co0eXF5Wzx82VEnZlnUdINHxfw84E7W6FFInAi1DnB3jdTpQmbvU4pfM
CdowLTDHVwfELZ+i+DccKnLR9kkJmYtgrfg7/D4uSQJVV5i4cd2zOvuVIupnvnFlAVzwN8uMJy0F
baD7DW6/TSAiO+bgaZ7j0LHGPkAsE7pLCsEur/tZFpDxXcjDPQ6w9qRzW2oYzo0OTNG+dYr5S0Yk
/b0SrVLLCqAGdDTEvgkwqUt3s0T/XbX9nB56VZEQsH7Wata72XSOQxiAQREL60hFXGLYA+G5+Atg
BLzz8CupFIGI9WoTYiCO692YHs6kULIASDy8xEbv/iM+aFTK3hSkgS2FWTBzzGPtMTGp6dS4cfsb
VJGHUgdviozmif/FY4m62UYJMoFYKoL6wUAWRJyi5qoUe27UYioAD/fw0Z9fRRnkxE6+tcnMV7MJ
JdSx8v8PSm9Is0LqcBsuW5BzCnLygSIZz5WsE8dUGbAFQpOXSndpT2KWfUvGL+IzfUpCRc/DOT5g
wOjaokxcxT05By9VA277QfkxOasLI1hJH+VUrzi4oQqvmSqQh58L8TEylqvfJchi+oYs1S4MNA7V
vpSI+MDX0q098l4ksWcKMpMpSSkME0YXKnY5+nmtIlon3UHvWQb7NcOU/GUUZ2WTL5c+IJru7gD1
vM03xD3uGhw7VYfyHpJPlacv0Hx/xGrh9BdKZ3ltwDAsyrc6BG/BXiHF0cpl6W1Ju0IhryVfxig5
JWsEMabjjAmy9uoj7+8HEHehkfcTtO7TAMiRHAqhzTNEyPGQn/zv758paUuVY2yLkQssbViyhly/
LDER0ymt6H/OvYhSrphZK+ZaxwVBWQA+WckXnwKmqe6xD10BVrMLr3EuXkIwMsxV78XgsmogPPTL
dzszBmu30ssZmAYNmzQwKLgnds9BwMvH2vFr0Onb4XIkhaHWahD5dqLkmaM3Fan/sWiTjF7Yh5mw
KeyMmx3VeEy4TIVgtTmdtKgZsp3dNzew4OVfphyc3rN50J7Mry3+t9vEksGe/NlX/iCdaJuMn2gc
NKdEDFngWG4/omZaPvIKuVLwRBlV18Ustq3h09REVoR3IqTn7+h5tBvnFLAnllhlGtuueB+X/1wz
f9DQyiBtd9wGgcBtghekBPKjXZxHw9kLOvcwRd24pKb+8Fy6wposamZ/7H27DltMlP3mgD99hh2b
V6HN+RL4+BuAo7/TZRm9sfXHOrZC4m5l+LBq/RGhdBQssweyYI/15IxWnXXAClWivdZF7ozbeyRk
GlNpU//GvPkyuNG1CFKrvhQpY5v93AZ3JdFh27TzqLPwT8gRJxPY16ppqN9+HP8EOZN1hUupvG9S
LM2JhX2RlWFl5Ny2+bVyRs20c5F3OmVw/rxKJa7FsbQc58mHHPkTieUQ75sRpdhNdneI7drH8axX
ikHQfW8Sb3C02kvxE7koDCYzuo+8yxdlD5PYMVMN7W8XFZNtISucVSBcbQCm9NhJN8WNtS10daoF
+1MFEfaaHwRLXshILkQwVtv45ShRsYf4vgdUoT+NBlkBS6rYmyCJ2auHBMaUeDYUr+vkSSVBzU3J
/DF+QPOdz29IKlLloe3hODSiwQPpt7ztduyRRDXVKk6rJwUmyPpZWhdVI14q/DfvwKCtNe3Cof/4
uM3DBDzyD4oYoodpj6wXLwepgy0ovnRunn23PZpGLZ9Itxw3f1U+QqOPbMjnEiVtqdFA2n0WLHB6
OdeOcuv5lSmHTyV8qU+/GaVq/Z44R2OlsMEWSMJkHEpSpOG4se7h5ZAWgF69x2cL/SWlLi2o8ilp
D9xp+aHB8k9thvQ7TiodsnOHcwlIiPKRSmDklz/EiWmSsSCpOMlEANCBxYg7ofFTMM7+Q2um3ce9
GsMx3OMcg48Twu5nHKShaMjQrgCSEQXdp/dSQGLceyVqR7r/YKWnYfLJ72D1QjXBztC48SqtfznS
gOBMUjNnsprQe+vKCEtHd1MKPXv0ndYrw4YSCtUV+/MNaWYokzNfFcqDMdqXhq0hOSXgF7BSIpoW
hjmoncJ1sE4GUEtGQHiSpMBYckdHO+qcqNAQN2iqzoQNYBlg2YJChd2ymXM71iwu/zctVJPL6n+w
WmXQHrHHxELjphm3xUEiFKfiSuLS7sxiy/dvo3r1wxHIwUYBCmsAkURoPegiylyVaurCDEI8u4A/
ad2FH02nmavfwh57QOhNqlyPp4vhUIbsYubpvU3aMKdqpOcGv1S+N17InZUnBTzarn69WUWyFaLq
Nom0L0L5xoFiT+KmRNMpiXO47thzF45sdWQsAUJ0gblPXgLz77kIRsLhwAJ8Q2JlXVYGPXpt6MV+
qrFQjRoe//lksGlpuTDVQ/NvqUhUVTns5qPGG9JExJwRfzNT8TRZqkC4OL4NEJL4ZH1X+nRu+6qf
tH3Vww2xpYPcGd4o1SG+Hd24kER1US/bU40G7UDz0D8DIgo7eLtUn6WHdwqUIBWK9hv5rief+Vbt
IdKCZr6njDfGk2K0jHPew4511/ZWajYnb7xA/gkCrTXbCb3IpqxZJWtmsATYPruUZVF2hZpoQloz
4vrTL0Mk8hQiOEfhs38B4DLNsqOt31WqDaxKXVkEKK6QGNsJBs2ZgAtymyOsyKwUzFL0hkRPDyH2
xLjMeAqxB9illTr8VRCe1ePb4CCHtX0H7en1Bem5n3hYYv2/Qxla0aG/pV99UROdIIZuLKSotclt
bQseYvh1uuuxUSQpth8hzKdkQ3dU/LL6KOYaMBmVBo4Fsf+/g0HpnGq4Ck95JZbeJsWYH3c0rRsP
5ujbPDQdfxV7J9iCFpYvY7nmrwGlchgMwk4uYuRQOXB1wfE8eAhNX5UfUlLz3pza9qQR6BEdyHq6
vVnZthyvJQioZa1QhK1Zs3eVH7uqLzmSo3pwlTkiWWq6J2J7VG+06X8mjHeiyDEipuReNFNsrq/z
NnWfIngdpEDpxmDjn0IK+BgvPNtwS5y3CejmUHQ95Cl+u/R/c+tZDiUBUwKhYKMvOdVsEB+m+4x1
G0WDnMc3UG7aQBfkYdKj0mmi1SlPpNWcbyVBnosNHtm3NBOsBreL/1KtUH383JiU4PwR/eyUggFV
NEq6WWsdHulr1BeProYKH92lGikuGT4zQ+NEbeFZHGt1CK0dLNJ0dP+hVMjaz42KfeRAalw6YO/N
qOEjiRkSVOuW85ZBqC0/GkKNCqXCwiTgF6U1NHEjmSPf/ebXQFr4Ss1cABMz1LoPeCkgCjt7DRCi
pxLizE/vlmDqfaHqhXJvLaSxNv3jYB+CkvzfMjw8HOjcJ0FLqo6grCIJepsdASAjGrJ3qqgzfXVI
upZi0nk9EeI71LN+YhtPV8kSKr866rdQvpRw90zQjWSCMGpbuimZ9AXpM9IBpOdpaR8UmfdIW3hL
NTp00xF5crnh5ZuqC5qx+xjKp8tniIUYye3sr4q0rj+5Ypehs+Xm5Ts2mi15GbgfGUUtrslB+v/U
8AxFdv0OooGZQhf17tOeRzasqS2aEt3q3LtFcxzdxGOxdsCV3QA/rt/t9ODKGcyRem16gJlRoKt7
+niEaRlDJpG+vLnI5raoe3Ab+dj4e+kmN7LQSXlLmugB00nueNQmgcmZKbpSDiVMSM8ZIIYUrwVY
tpTGa35qDb00c000pKgVqu09AQPTjgTKkBt7KF0fnc/G13lvKpPj0tbgjpBZJ6u1pcTL6f+dlWUf
GHQUkVPPFEpsb+LWb3NKbukUN2aipjLkBMRySd007u5IGdEVxXpcZoMNVh80+ScjIe4CxU4gipji
T6Y+MxYVZ+Ka50wJg6RtH+7O4GptYjZ7Ad93m1CJDR6tHdpHt+Ec8nv/PcuY8N087lv27GoQ3Ot7
Zuzvxt8hoyfVZTyCoFhn5X/1E1TzB6EMLglVLbWGzgnhgXgC1OwvrEAASYSdwVx7GLPy2m03zGzI
GOoRrtiUP5pm7HjhajGZM2IDnmWVCfduk4+/NzMXkZxs5ZV9ivgaljbZjfwT2O0aNidVEu5V+QxX
tlAXU4RUDAi6hxJa4zJcKLu3NLFh+cyIi4a/wIuZZKmYxcYJFf+4mmSNvxYs4d5JVKmiKzEbWSmv
q/Sds8Yhvbez/10SVFjnmINqI0hrHG4qtyWHSG4+A4OckFYOza65PMPKhe7g03syogXpsflt6hES
3UaQA0biUmTRaDce5WVbTp/igpH8h8hjsuqGIVQvYh8COunCaWne5Ssc7641nJlwM99cHg2RRA+y
SyDiotUjzi1yKKhUcjhO53diINmTYiGQKn4d/MsPjFEkZU+DU5GPBr8s0bT8/EguL63yZKvOG0CT
Pq3o5i+pY7mMNHl3IMEPWrgmla+965hgtuv4jzxBp56VMpfK7VXDmAt9C2As6RPyGY1CkkqCRHqa
J9pTMyPMM1Ky+j1VX4yWUTUJF4i2z1fhU4G81BRenhMmsulr88+veMtT1oYHPyTZapWuxDRUSOam
7BHeaw4tjKYqjEz8QYNZW0E4VB+PG9A3enB6quv+UMmIL57QLZU7wieGlPhS7TfalaoTTy6LI3G7
vYqbCYGDOoKdEZu66Zl7/D/8ukbewW62pK532mdnvrdoJLCCV+lEJjwJhMMG9aTWL0B/8hiDKdk9
QHHvqy2uJuqDJYLTwCD2qx+gVU6QmkPz9Tbd/shM5Ddn4zW9od8z/gMRUNUGfOqvzBtzqTOQi9lc
HA26/tn4VRxL5gxy7imEDc7sdFsGgZJ1aAR8eRE43z0m+W6+Fgu+wYgb0sJwduMS9zj9AbizsYn0
ziTtEJY3HeTSXFsX9ktWuaJjpWQEPPUlgDu95d6PUfhLqUw5tAdjY3de7dPhwTI9+UrwA6AL2RHB
MVbDFTkwz24Bga6iAbV31UOepIjp1rYp3wO58VNJ3oWLN0PRFd2IlylfwmjPhloOsaHttDwYcGIK
tIQ9y/+GGan/tXCa0QsImpC8HvpAo1fJ04lOdL31iUSM5TdVcVF1InxBUzNQgEEY+jo09+gk55iM
L/oOWJC5PWZ62UmcmE6+Ez7h1GtZvopjg/Jp+usl6C90BaQJqGT7DwPM52BX8kQ0riTMgwu3dKFF
NMK9ZItXmuKT8AJ8WGIHkk7iWC691XI/PE15WB9FzvFKukLffAN6N/TL8oi9DTHkFJVd6SqkQhlg
gNFkZmEgMzZcjeDo6CMIrqIonvE4iUqEgP6tuKukBGZJbhNGLDb03iDhqBOGi2VqR0W6o0Rpj05z
ikZFIC68nsPvdsJAe8tKg9qEa2Kf/k139OludaAaTJUSeLEsd1nF9Rz+MpTy8U/sgB+cLaLs4LyW
7rQRme+QWixs3nRTbgBKb1xZjmij4Xe24J6JTylg2nhQyqvM5u9oefQImlVH3iuxQE5mwrCuEIRI
CjUjlyaQqL4oNzoDrXi1uw6Ooq52Le38NNiStxZeRrmpi5ZYOQeRNqGmzpMGHfSB8NxHIJZvv5Hp
SJfKZp37UVtbRzvSyEZYdh+6ICDgxEv1eGa7aCD7b6YHdX2UJTYgIXXm63GlzYj5y6x0mVn5P7Bb
+xjyd2NdDc+GeLFzTu5mjox48q4r4BeFjl7HgadmBHRD0IAyyzCBnPRrgwakpFlFe4sUpbcpKfN7
kauYvs3OH+1hQ0IOL4327sQ4R+JGjoFBG6s8N1XwtpcVuFfVLkvuBprTDXpg2Mxq1ingxup8puAm
tbBI0ZybIQaCudiMnOp2468ILidohWxBCNOmHrrAkziQPz+Y/57RR6lIwlTlYTZeBOvvVZeguwZ2
pBTMD5+Bo6VIpbCWorUnDbFa84tzqeJEYW8YM1mze3P+qb370Fgke7wNBvvBx9LcgIihYPQK2BqI
fzkER8IF+1z/ncu93UxjMJegNe53+PQe4crgFJkD8JQXBInn5NRgzOe/hNf31HJJzW5Sz7rn/eIv
1d2qcUw3LSjAK4aTarVo68uYPnNWKha2ak8XLEW4Fag7OWyVS0v3U0yeI/laIw7GUTKGFBXFfLL2
xyAwM5YrqVlBZ9V2DDidk8+RI36TSoew4XOx1jLDZXNRL5fRULNIJSyMmxtR1cEOKRSwkF/L0Db4
tn033XJpdre+u6XeMmOPkHw2rFpViYlvcW+lJAwPcrNKy9vf1vHYknlUhs3neYZ+koHbgS8PkPcK
vwDBaXjJpt73c35a/VpPItTIPYO0Yamnb3fjO6wf3W7zi0sAEYgd/X7JilLE0+omUE/OiAQ1elLl
C3yvG8a980rcVmBQgQ6VNVtaqmtHZDYnDl6V4OMv2a2xtAhwNlZmQeP53MkI7TxC1IQ8G8FUKKp1
S1f7GwwANP7/OJwPu3ZII8LjY8kvmz0omP3wE1y74/0UD/SOd8xMY+y8jhSeKnXT/3zuYQqQHzPb
Vwvi+tX8QDgoU28CBf+lqvxzeemJOOWdBH7x0wLr1EP9ZCJokqNfwqrwY/zHcvWqpWGtPE2G8QcV
CEb9e7oGi5n1BWEQw4OLFXIr8jE6qpVAqEZkYBtpL0OPODci0Rl3fkJ81gyMWZUU5I57ZVlpduER
6AwvHlsoBV3e9nOGK0TyapGlyx9O68r5znp8HnJydh8ZRz0dmiDtPWYldTV+FXTCfMKVitKCnvPA
a6QluydNVmF+WcpBtxDsH5zly3i4sz3+QiRzZlS4ll90y7/1hbwG8hXCB03cf20jevg1v+t01Rd8
gzz34Cy/ZP0DdHqUW9MPPcCxzGvzXuWlwZOrOCgwwXlZqRMX/YOscbrjZssSzfbWhxrEWFlm4sey
95kYq1BXRJ3pjmOK+yDaYX+08Vj9DLAW0tdh/oRWwCw8JesCQ6ORlSy/uC0soL6AcK8H9bqKFnT5
VBLBY/59I2SwTsCn6Xq3uCWNVLIv2+CRCu6eNgHLyvJormXlzEDdL2qchaT6UUzuAfbuizKaJ8v7
+cCIv4P1KRk3v7voTfdl7WdaMoXcPokLPE7BdcvgxeNuHG5R0/mfgFDjVi9gf4SjNNJ+NceGJGza
xxyfL9q6W7Lb0XIQJr730rfGVUO64VsL0dwiSJrdCaDvAqUkQQ9hyce7uqjMcHzBmmXTsy2h7KVN
JZLBfeFedN91NI1vPnEurHGHiF5TSxI368tC95z0KNdmFbZV+izP1eTNzI/bqp6s7i7sgjZ/k1im
eotJQnn4tk5+Q2ppyaprcxSgM2KuCgu+tuYkgxKuKHPbLPS8/sUULyG4jFpnY2qNsI8SUOxR4Va0
zF2EhLGeqIqzqzanmeeVSizLAkACI7iKLMq7EDakuywHKwzLiPXvqbjsA7KcgGC8uRE+WiQBz7Qu
Mw23M5Hig6veK7afoTSmtHfFIW9t0Z7bsKigfIK8RSjd3w5wCOHAMJtQFqEZVhNksSuUmJN/nGmj
9ETe14t9HYnKQv4Kr0vTnyXBvapisehhALxxBipeyWYvXuL4WGUOhTTCdYmenf9U5UIJ/V1GKgWm
MeJTwmJptru/ivKcUUKzrbkULEMKeMwfUyWGIaSklJ/BFOd0bmqKqX6la8yysqND56KK9dU++Fpc
JqeKHqJvAMlQ/qmzLdBR5sLBrJUfnBl7duVJLSQ7Rxxnhhnw9VQEewVKH8wTobqpY465C3fhdQwO
sQSDA7zqfvQyplKWZlrzoaLSbvO1NzZExHt6r2CKTq8HQx8pWYAkJJ4HUedDj/shHUMtYH7amjpF
raA7ZLuaF36cj85GDYuXEZaUZ7NOCN+tii5oTfMyn1DTv5UsXVIMevdauPdm9i9tUB+sy8Cxf9XQ
w4CO50+hrml1HBuOo0uJSnf1KrpsEJKDVbN9Yt7EFWxOq8QVkIFHluGhjottDZMggDZF+87nGdq3
ptJcXV4CqKaY9uaEjk3pJFR+Wmwgzy3L3AouzjIzvg3Y5En0lJ5nySBTSs5zuF/4f46j/vzEd8oo
uzvlC3gttYoAkfnzaODdZnmcGuhjA/dM0QkklQ7d149c/HVmF8mMP+XZngkzHyyZR0UPgPcphYeS
cuvgcWzv5ebduhmMb5M2mT/26xx5XTp5u9PQrKscn3bn5hEp0Fj024AkkyJChORubaegirDvRTBa
nm+JpiWqbn/0zhe6/M802X9VGhPfTCAPmfBNAS0G+y9nx5mJ/N/1erl1RF12x61/9dlnP6GwvjDb
kjHjEvwQ4fBUk9qT8NkCngPHOJ1OGXiigZucIw5ol/rQVE6L5DGu5i3TRcS6i13PoqfgP+XJLNlh
VGzgZScjQE+3LC3TXmDCMOz6rBAWW5YsugB7RoVAGyUznfBVHLMMcx/rJ6WChFrut2TH4wZE1BnT
IQNYsP6OzU7kI78a/rc+TC+DbWLP0t8E6pvKg27G9uYbp1mTUZHzsc61yp0hKUwdtAFPze7mJJ1B
VrSPZdesXW5MPNsaAnSWMB++nJy7V+BSgDFlMLa/k7kOmgHKaDisjUc1vBwu8TtzpXRGV6hVL1cO
cYwdU3zsuw2odYJ+345+uHpa9BcUMSvpiRAza01mgaGGdRxI3sr2WLu0skO3DvIqdnx49DEyAId0
kreOxObuaxzyJcXVnlEZ8F6Yr4Kyr7I/u7WUqjs4z0FYEDTO4tUYvx/NGeUlBqU90ctJglhy2ytQ
9HhJ/LF7Tif5ySjoPQIjJCq7NTg7fPqEgnFpcZoFqpcMR0OYoy4Wsu/1K3Zb3gaOHtxZ8Tb0mFDT
eJKTyba52J9lYZA83qOP61bDQag0XEUiKY0dEWsfehAmYCUIIfNLkacJ01wO8qngUPbiyPVsqZrw
H2NA6DAnVewgt9lu8ROhcVcPvqjQmu/d+b82LgwKs7Bx8fLgxLGDaz8G2kcJiZr2Q4mQDaRI26k7
PyfDz49e6Jpi6S4rszrfXkmpLc6jyBcZ25Q0IrgjON+N5L9efttiBCCpqjCTeJF48yfumNV0tERg
W46dI+aZ/clhHLO7pTU591yeIE+bmcqGDZ8Qb0+qQWjSajlU1dz2x2lPUf5kwGlyuOSpy9HCyvDB
HzPE0v5jmZq27hqVv5JMPd6EvtTD5DOG8+WGdFvXV6z8zovyd83m+TDafE/pxk9ST/ooWq33o8ex
xqnNFUOyBBQca7j2lPOEsOE0HkwiyLDy5e6ZimMGN3oF48eWTYTcU60S9av896tNb7kS/YZA7nlp
Xa4aeCqju77voKkQ5PBnsuGPEGcIwxqIL0On0i+SwBxql7ZWHUmQl/ikTIb7ROAdIh0fw/9zIfhW
r7hzOL956EzrWsIVxGAJwvllxDQtI3Lw3Btx/FoGOru/zzDodp05PEB2i8Lap6tLW/4/FTnaZzP/
HT7pe1TCnU8zXwLB5Yso8JdIyRZXeVCpcw/dPXiwJVG4ASyVWIJ470CQnmD87MdHwf3UriAsfaw4
ZWmL7knT1ssAA3eMjni6STcexPBaDMdJ+e8vxbnT4leRzz3FW2aptes8yOqzvTeUww+YyHBM8uUy
SWOjw5HF7aEiiUhk7k3Ep+mjneHp4N/sV3ix7JEii0igPSh33hWMyd4B3UlQWtpQyIy0noZUuZQD
D0912LqegzSxDcSVxeXxWg0+qAtOWVUc1433pstc5+a49G+DIllQN5EgoWv/m0XEKSALRPOncauV
ZGWw6fiyLwCC9cFn2EWNKD8nnA5sPle+kdyyvW2wvH/it4KCKJZAvdiAhAQWd6I5cO8lK5hiC2PG
sxp8+z+oRzOeOmCG1kBi5LaAL7VPB4OMl9l0Dj6JaYvuClSI8csWNeKvUcHr2wkkSnkVODzqGLkg
tjjpBcfVd9kdu57c5dXVYVBx8/1HHsCy/rUvmI1LEVjxXPYKzB6QIZ2s1vMWgkp3EYsxmwsSQcSG
sf+sLyuP+TWHSvDllSNVTm25NdaRlbhaXI3gGya2Hnks18ApRfwi7ib4Y7qm4cGCbS6mSVisZNWh
+EbtSS7cTgoS8AMDgtetYf1ekkD1q24ToKX/lx7tQV/uZ4dpzSAaISHwGEUsP7wN4qNApwl7LTsJ
AzaKAGj2QSLken55eBWDfaoxAPwt/xldp2Q47IJLi6Q+cSdcdHa5YWmVfmFnUhQytgS+5sAQEa0I
Jf9laWs4fr/nNXN3unZFptuN+65Ao2OhyU7vVRL1wxDSErAC8drS11PIs2YR3RfBE5Md9hal0CE7
FdQyqhSw9LWldAYgDP6LngDMEV8mmjkXYPiEIJmtoOm4r2jBnTAPz0Vk7yk+qiyToro1bbrS37g2
kWv9Px7cXIzJ4O3ZMDiiyMWzf4T1xD955ivoRdlrJkHG+uZeoelmieG95M0N9/mddLbXWfPmyGnG
BZ0ZR7P+Grg/wRdSL7dX7tw5EHF+FSJ0TlaeRtp3BqUmG2aW2zqsdOYT47f1AATPqbFpsk/3ysmP
1CWqlb3ditlHQSfoMLJQNvej+8tIHnK6rBP+vREcWiOGJicjZqPSc4qS5kzJ7guYoUkw7CnQqNq9
JN1pp4M4V6Jt32WMAjlby0e/j0ehfRq6DY2BKlmfk0FZCpe2phCgGQiNeO030IzL05jBjYDBT9fe
DPfQGm4Xy9OwNwM2KWUHptCEzMEBq4zz/RlqqJfrjJ9JO6i2ayJSkaOo7TMD/+7WfSlB1so+nJkt
kGU5NoaCRKUZaWG6wTjsC4CmKL8Z1uSH/AVD83rLAsRDquEBUrM71aAzxZKsJy0Y9PluyD3LJpi7
oKiT2wDQjLZxCr94JwtDVn9ycu0nUioLUWb4SiNdKInXkqYrqp/qsG7OMb4tx4Sb+xfG8/BdIafZ
hZMm751XNK8LK0d2VXrYCnHBrfsVIi4jLscUuca4m5600X2XJANSaLP4L/PORm8vNWSOGb6e8nYi
zlBuVl801j4BBbz+tk5l7St0gpDK3HXd8P2QpBRS1P4k1dNAm42td210FMFya/70wxUG621yNlUp
Kd5kBWwhVPXNVh3S6yBkicW5VOYvSP4ADqmWVgFOPXylc6HnrB0+h9gIT8X+SmmDL/kKDHvdJqZJ
268vgWF26AvF1hHDjHgW7O6/bAsSDAB1KIginWlGdKjC7DuM2RmrNLLD3TsA9qlQ+fl02tqUFSwI
UGbjuUybCaFLL5JTorXJEnrZWCYnJVT0azjzrGtcqB1K8Q8w6jUV6B7iR0LP9V1Ae4ITutSoLpic
dLdqqW2yCS2e4Zl9OSYSimvV72+aVaObHZdbtqWJPwYn8/DCivYpfE8LVMSmJOdy4GSLkNZMViDp
OpZR56ztk7eCJTKAppH6hPPUn6kjNPsH8wduaQCFTZ8UOs7oK3GLB8ibOr8mihHel5DaYpRZEXlF
PccXrX2BcIKNKgAsAxJGtmbHiVzjDX8sjrKy6qzlMglEhNOksWHHLUJ5+Xsvk0KgK4jtqinWIwtI
cqMGVxcbLfbdlKKSdfPkwoWfD9j9o+0lTD3HC1JmFENVo/PXACqde7wro3DDViC58KPaiim3xZEP
BDuZ6k3QQbd777BgH16t2T2MNf+J9poyvVgFLkImuL4x5Lg3IZ8WJftsOfxt5I5zotnmWnJGMP2o
XfOjeqWuPfkdgrxwBgY5Dj4LSo1p+2jiWWRmW+PPFNVPvpC+7wx7VzTh/2w9c2xUSnfHAeRZcFLm
ag7Nbcwe/wBUi4s3i2H90NCHGPThMR7CnSEH9ha39mEVoPhM31qbpHAAg5kdNpNEuIR1qk+0igVb
jtkQHGqd9Sw+/sRWNMCxrWnETFUBAyddaFjO2E1Svje1UtSO1pnB9jEA8q30ZiAawRPre6WXkxxl
qbTxAwAmgGnDEFDZVLHSXAwd96hXIIFlJPtnZvjDXcR4KvtQKSZb8k8UKogOWnVqG+2PU1+Py2t6
HJ8WwvNMZ+xD5baGn8KLssH7yGGhkeqL4cmztiV9UP0xFYCFJNAsfqfYqRPexibxPmjOgyywvuWs
r1fhiMXn2N1aYVUEDbExxcybceT9x/tUXq2oM+XGE7FIX9Nv2+DQgMYCVTAozaHFmShL+cHN43gY
MSqjLgrysHlXHUShY1DsqTGgxjUSOEeMn5vJbzsPVGtNN7HJ7GRAI4HcW3hh7VF1OXGnnd7N/qVx
seCDpW/AlPL3rYs06Y+cIqX3tYoFBnNTKmrup9ggrV3nN/8198DDIpBbxzCIz0XFv+GGxR9S7Bc0
El5lP+MypK4Qad5trijVPcVih7P0qndEyZyRUCBdt9OduN3G+11g7TuwwlmgIGdBrhh4KlV+xHD8
IHPs8u4GY9KhFRU46RC0rdtwWNWup7B+wDIYSuJJ1xXEEPBuddJCjoWR9F3R12FDXMJVlHtX6LhW
N0jO+npo3lJKX5DODpk3nnbXZxgeuYF2jGYPo+i7zHcguZHNA9chz1Q6RjRjLW3ZVMkUr/139j89
X8fyfU0KLsmdZvZM/cIAx/OSs3Px8cXnxMmKDVuB1woYY4DodhLx+sONDHMI/MOZXw9fCc6xEbvR
fOMOlbrRIORdu2csVTTkYSxYuBskhKJDG6wDtYMBOGLjdoYw55KZpLBvzFUiIGtv7M1cjA6g1d6W
3SlVmJkSPq90hN2D5U/7edIaqHjh7Tops81yRlEmnCtVfBJgAVOFfWdmeGxY7iwMZTx6Adj7xnk1
URtcYkwpQ3UzZ5KeITNcS/qO6ZNWlljHJfgpnT9Jm+4bNjETJ6vWIgFUJpajboEd7B25AiFYHr4h
k2unVHR8MFP/d316e9q5kdxFFsRQdqhaLHSB7ASVYl5bUFs7KBBrRkqnbvqitpDTN2UQSsGpfVh+
aG4G62wTauRU/6Ev9qBijEBfVtYNeYiHdSPIq++h9fJFXp22dP523bHrBqKGR8GXAtyp3pyIWKBh
VBeNclqwSDweKotXHkcVADzjfQKR0uBANbDFIs5ONsZdVcfIloWP6gjtyMSXU9f7w2IRm2tLxor5
QRnZixHcTjfTWboEYrilIZvzArHJ23fq/8Q6KDq4ff/CScNFKQhM2VrZzLU1f/CsBWtrknDqcgSg
68K9QAjGdEuKTaww+YYEbuv2XJPzk7iZB4sqmODaPR0+NaGFz3tzXMNLP6hgfVluu8GqzsnhReWq
l9WYrObwpW598btwy5vACvHRnOCwxuNCpzSkZOBy1NBp0vbkUYewxe6/kJqEkSuj4DPKJYXamUEm
e3axjIdOQQHooYYwHiTLTCrgCJ9xb3qk/o1lStBUwme4BJ9w/EMsuZcTv1IUE3JA21tzErLNaKSj
d8Kth7okD8ChbmrmOd0/pWrb5wWfYpCtPGYh9AAbMJCF62JuDoMGnyNj6fiqgsy2Qk1cDvcamLw+
Y+RjPDes4Znc876X/fzgzwUW9hi4exujca7g9A+vXcoB7aBCPfE1znfkD8gCbjLnVjD3JvJ6+KIm
icKaGDES38/k8OEloBTZC9Vl3VN7jAVBLqL6qq1IPotvTKkHoWdXQfIq/LWBLNUFR+FRTkGQKph0
EVm9PKkC1oQnRl16iCYrzznBaHHldSkpS0+F6nX/8PgrpiS+4E/QdpFAVYHioliasPfbObe8Hugz
9KrTg+i/DwheSUlHxPYQNjsKUVIvdUCeu7z8aIvYN6SbzcoUDhb7NcZK6PXy3wobBu/A1oxYXzwo
wIL4Lb6cKSUmPLE8Jm/oSO1OIp1NkuDPu0Ch71fJy/wpmI0nHSicDQoG5npaXxPHPp1QuUoq+ElI
S3kU81niN+liWhKgRyF7SGzN7rfDi5xHnfcT2WJh0AwTOQeGiblsryzS271O/eO95dViGdUcygIl
0hAhWYNJRLIw4hiBtk0DNExz+qtIW6XGG4Hf1N6sJt6yFB1LmqHgZHxkGXAVRurI23pC3+I3jIlr
bodtdkNtlQEfZApT3bwkLUavBRBp6Tq676/MGLyt4Zo1YzEW3+el3gOBMqo7/FcJYhkH9BLklkrV
hQNlj/dvSaFVtMrVg2z9TyGWKrlNCk8s0x8CiUt6jMG1xHWeNvbPQ23W7fGY4bboKMoWDTXgt3Jn
QdpCrMAL9+KRc2Usy5vG/Mmjz+oMBXsB46gLWh3JOGtWojfE52NpTOIOKKvK5eeQZm1DvXeKUQXp
oIrfp78dWqUml6UCOf3sOiH3Qx1Jn8iYz3V1Uxd6V0dcRx7eRtSBw8auHEb+Pjqx7qLiFf0b/q8Z
22kqQHFGM/SJ9n70JseTNuaUfbom8mejiPteHUVYU4SF7i0FRW1xxwg9kENd90/qJfiutnbEiBuH
6SpBfeV4qzp2zgBGk0a6f9DP+49jdNTflc4w31LnyD/0HZs3xUyfpRIvgjViisdU6n/Bz6coamW4
75KsA730NJIVQGvMo4UUBdppOFYdP8P4bEz0DEJHK8vu0nou1TgAro/1FHF4wHhDtSjEAnuR5g48
gD2TZrWwpt9RpDkOD0SJxWtTPUYe11NbI1GtcJ5EwdiXunTywMHUCCuHGt1TWtSJO+CfxH3M31I/
O3GBoPKm7KnJUtzUce80iRS0tig3svt3gilRdMvVitS1seAg+q51hPZ1eJYdNWtODRzvwWM+MM58
mDHr63V1pQiH1kgYzpLNamDoO1mrsVO8AICjqISEaNFtAe7g68VG+Bl/X74k05Wq+fdjG8Z6ZJEc
rM9i0BwB5b6PLEkB5/oKwxnxm7rMbg9yjYtrGmYJgrXvxiN6/bASaGiEMfuzl0SthPvI5xNwKxc/
LFSRyTUHL96f7K5rwyUsXffEQowzZXFT7nYZcKqhk5XI8w9j9g1LWFqlwlDZpsIMflgxj7xm4tnF
q7PHGTelz9lVmZJUsGCbSO0E3y+TEmCo281tCIpmrhHeeUwMdWTbHemugam3UKDIfahObHbWuI/N
sFhvc3b2XbgSM2DpK9852GrORu9Dx1VVe29GbOaOdygU7Vsnucn5ZJ9e09xbD5en8ucix8lQYXTM
0ps6+R8KXubib4K+5H1cWrYQoW65WzpsdgULofaEwWJXEthGSAavnUeM8DpMOCKAGoEkT5gwZe/Y
Hc3C/LHgksEXzu+j0w8WACCFcCaz1son/hjhcFs+AEsXlrzji/UmzK2s4L3EjyRPx+ZjIkJyZhat
F6l4Z2VGwVRplmivL0+oxasvoEePr4cci/zMOkX1DUUPVjgsCqV2hK2pAHc8ny1+vOvK3EwJ0ogH
ocGe0bm7vSllMGzDiKAfjZjHxrEx6jE+Z/wD3RtNUKEFwBhOivcC3vG4XztgP8wxkgfpkim4jb8Q
fESAIBwedW/cQYkKvD1IK9C7RJytIkPEz/+ctPz7NwWYGTZUOkR3b0B1KPhnD9fP+AHhmFTyUPo1
3PLJ5oUX5LNB2tYKMPYyp1YhVbLyt8TC8XRZEYS/RKyX6FOrbRYAbrVufmR65O2t5L8W567XX86L
0gTG53jr09NJQVf0T/kdS5xCcUsfly3ek2P2QbHdRTJBEM/MOYykPbbHSRXeLCKoSp3m3SpbM4Sd
2suNsiRrDJm0A6UvClLNz4R24UwPTQnQQ2Zflf/aiW9CHkBwQa+21ApUyvOZlDmQF5B/cI70DneQ
NSiebfvaaJdFaWSKiI1fT5JXrjLWu/a5soVe6zW9s9fqCUOvr5kLo3e4gtTIsCTNuBN0qwY6j2Wt
hQRhgTQC+d2TU4TZPVhg0XEjQ0Dxx1F7yYdiPGVL+Kdw58hmocNwHN0ZrBQ1VpfuOOoCGpaq5OGU
B0/+apU3RQre8GPLJb7I8GIUY43eYvWDzvWwKPVz+f0+5w7V+dJqOZ3/k1j9p8KpFBeqJ9Xd6XdL
OcOnrRKn3xD8ollvbnERFTabAEST4LwfnEqT2/nP24tQ6cj+UzqbWEfy0B9U1MrKeJ+MEA7gQK4Y
APG6FPb9V/UBdh8KDdd5roOLlfF47MAHDBRq+irpcjk/AhaOiYcr1CUP9vijCtWTIpPR/7zRNyXf
qd5S5/EEuYtsmeGOYxxEryTal3tFubp86oYKsB2zSfHapZKnSENpUlvYnr+Qy8aFuAj5kKvGPziB
TjrVHAs7YC4FbSsPw1KAvK/MOyc2B6ojvUUdt0z41gL4UaZxhfpkQolZQKOr6cEajSTnEQpcdaSO
LOUK7MwLheV+d5MpHCkaQXOOoMua2/nE/YpztAMKnBVcNhP5ReONyiXaOCB0iFNfY0R2gsvLr/Tn
nfpxSQCWXZEoU39uKo34SgsnJtAFVoMgGjoKpJsnAbkkrYs4TJfCEX8tPVqSblpvDAWNs63RYfAt
u08+rHIel9XFCvh/3yeBvH8ceA9ApOcVXj0Q+8hghY0PE9tB3l3oXYu+j8azEMJRucZSIsdzi3Oq
nfAj1mGQ9KgGo4sJN4ky29aq3BATdV1izRjUrr3tRhQfQv3RTcuqjsH9gQ4nY9kye5sFX7ao4lzA
6SyKBnib/n8hiQp144yisds02+IvLDzhFom/r7QiyXe8AubW6HXpE455Oyg5Wyn0NIORbzCO55+u
NYAzZDQro6l4CdwmXDwFmc8s3tBEHKoUDJfXrNcAYGWBf9UOd2IPwPzISKfVfxIbjVhzAGN/fiK/
sGVbDBpokPIGQkGWyD2ZkNagkFU5+WMVStkJL4m4RheMWRq70doS/jcvawvOnfzpjQBrh3hNVLq7
+LSSd5lsMbuMnpXuajYraf4Duek9inDYIkYa9+Q9EbvTcZg5IdX/MDDmziCsAqaXGUwrH2wj0Hpn
+8tsbw6NtPyLJJ2UiLp1c9Edc7BImEH14xUqTAyNxaN8+sshSR8BvcsWilGWoXO0BfV/X0N9eitr
V0Hk43npbSzYx24d9lkHhJjCbDEJGpkPqRtSgItLEzKbEBYcn625q9h7EaP3A2ERTcaKt0JI9SzM
8TUv/RRI8Z7bFE71qIcTyaHC6bfHTtzkU3YT4UhZFnzAOUvYryToWB0sLIDCaO2CYTLj8+NXA71o
YddXum6uNyYrIGPnTWRhDrfb6J/dhcZHP9SLw9q98JKwc2YE3F5cFtgnwI6oDhKFyE2+4uz+QGJy
G5ahyvSjV2tlHce6DrBLqujtEwc/rF6LrQoI9WdhzO/3lF5UGutM13J96XhwJVQuVbslpRZPCdJx
Z0ZEjeZ47tjfGkzQOE/+Q+lqS6u3nhsHHAIyQJHF9e3EWTaEEJvNtQrNQtPBeG90uXWkED1GdwyX
EX8C6u1mrMNRCJzSyBuKiBmnskTHicwyYHBHI5tTGN20lkWMP7UBWiZyUFBjVfDkZ5gYtqURUHFb
Fg4UHisPMescoFj+axaf7D8b3Tocm0+fqKFu8rkkRl62Mv2H4WD+Bvpo/j4GOur1/ZJXtQliSDt4
zMR8e2+Ss0qKW3MIgEMc4nIx50CFF6JiwdNG87Hk8AXF4i5Uq8rqgUXmTOIUqu8FFzKTxUr1+ID2
iusR84465iUOpdYX5mgb3y2TyKvhDYeZJ3iMN+SaMAYz/VzuewNp1JlAi2CsSiVn1F13j+k7HwpP
QRRSadzaieJcqWEG3jK86m88iYZ+/jimldcAz8/HnETImphfb63LPhLemz/V+gDyu5eqGEVFkGbh
YveO84XEbnxSB9Kv69WosZMAnTerF0Hwvk9HwaefJdmVuboZKlvrdWWo+U5mSf670EC2VF/5yiEO
Ydo+K2nMNAXXerDHkmmgfU2exH3YERc41GOClJeewEhlO3xyhQ/ezJAdAxV6tehhLVx67/lFB6yI
gwvb1PCAF5Ad6ilE42RWlugMouJmOiJbsLtrTy4RTeBx4X6HtB+md3bq9eDVFEfzgVZUUheAp84e
4G2m2fbCQKDCagZy4L9fuUUOt5fRbgznhF0wX3vgApwDCpCd90/COA+gCh5uLJ8rMrKT9qiOPsM/
CPqarKoVZXf0chjeMB+UbMKFlLgMLjJQawOlzaAKR7zY105EPYHo8AfB4lx2BopkQyKo0rQ4KNiq
BsuoEnZJ4XnnS1RPTk/0qdGZelNvdhC2+Y/ziQrPb73/LZngDnEGFcbd3M9OTWRDxAiyeFhHf+IG
ROKrPBK0cIpLf9TW8zQhi/2pZFZ/evWOObGcJbZLcrI4Lg+PjdYOHGVi7JQACSdbMW20ze2Itwdj
m6uiI/YDKfm2A92fhKkEcyjwP2KdusSSYx20YVfnLNIWmtKOhSO8Nda1bbnac4SCFv6sTBfwjNeD
yro8U1wkZQpx6Z3NPZQgm8bm91DADnNjzLexaStBlLUzy07GxbgWSVrYAIrPJXtfyNEhzzbE8/qQ
A9Q37LAPPmQburUw4/9417crxd4EMk6BhQ5QKSmVnZfAKWjPqxQFrfFOA3HgQLpvmRh58lKusX9K
z2Xa9hi5LCnkJkGAukOViHHOPBpoUi6E7pyyq6Pg8D7RNdJtXmfCgO0fsX/VPMSy4VX82AYxPDxB
e845MvBIB/F4GX8/NCt3G+Sjy9Pw/r+rvO4Jmgf9TwkTvq7g4wdHxeAjnIybs9VyrooazICCpjHS
VSM5p5aC1XQIstMikvNO0Ov6gpZGAiojfuyVI7ExEm5kFTWFfLakjGiAiwFu91NZT6SsTsXN7zb4
SfNGKZmJVMpV6g4b02zPWujZooiveL+HByD/1O5oVu3xzVMgknfQsS1V3RKcnDSX+/a4GCLJ6Z6p
5A1ZBTxfhUjxKIhGzBPZNFbSgHdehYuT5vEc1chN/X+U85XUgNCIuqnJZoqj38hXVI9mijSkHQuc
8bJkLQUIwsapZLAJL+SvEMKj8NAJRIb+5iQmM7JhBs+8P00y/bW07V8ZHWcsSnW1TGWCjNUpxdiK
RWYRK9vjL7d91RNkmUjdM5F8qHkI8WLrxDnsEbRtzTDay0F3Eo92TpHgTd7Q5vct2ev6OfVtMG+f
NOqUu+Sv9rmudt8RwqpKL6LrEM3tTdRj7C4aZiDN9i+x8Uz7uVNFYYGUGYNKMivVdLuwvN6jBlpc
NKDISBwrPgDqfmfnvR/8OOxTKMPhqNEfDGPbObQtg3VkZ5UnJpk/KeRzn6x2JnFF80hWw6BcJyrM
AEzpqChxs4IDT8h6y63rdAsUvTRv6SvBNCxsPvr8LmGJScKunyAgo0xp8d5uie0RXj5L4/AOEiCR
X3SRdHbYg5Y3Hoxs/YllHHbg94YL5w8mAnNGw27/Bib+/tqKhIXMyFqsSNul11MFsFGzNwO+03Oj
zRpL8YF9w61XzP08Ydx3jVaXkPqfZqFVx7hpXeZ+ndvzjiT9BWx71mNedvuTFWB6b8c8Co2jHyt6
8OqGLo+XED3gsQoY8HphmQUKuvacciEHqHSY40RBpTaQCCGgmOyA8TToWq2i76ufXxvIrSjtFB5Z
kNhvFV//t63i5MBPa8APRLVHpNrQszN4uqBROal0nAKCN7nwsBk+mtMh+5OhFvrGQuRGDd32IThh
J+Wob4P8eV91PTb8/uxf4F/lUz2ZFmrE80xrYwJ2b3ILnA590X0N77Tdgqi9NgZVl7T5QWKW17Iz
qX0HEZ9CIFJbTzJZ5yRsHhz5fyKQS5R8mRSNheZb8rGE3peMLowWXsYXdSYzZdUVwDOGB0uCNkIo
UKzPBZ/sSo1X+JEUHVVlfkPp2/Uqq9HGrxvckExLgXR68+NiRh/ImMWiugUYyabArS4uqbCZi/8a
N52SLA/1OxLJJWSnm4CHkMYV09QMrxfjetGjHsev7FHzJDG3nAMiS3RJpKN2B+eb4vQvbod63D3C
ijF+LZR3Gz4uVWA9ZcDIAQjsKfVshCgBXZq+wSsnsylPqH1+xyTfMxbRGhMzW2azeJfFr0ym37Td
WIciyMmNJHQP2nMTJoBmd9CSZPCslukR4+JXGwgxAGij8PNP+6E+mk6dXTGoBI8ix6e5Mrvl+Fy0
B4+KVZPGulgdceGaRQkOium72ic/RJJWtFCeAPqmIPyoGtNy/hhMW4dGPU/oGkiyIBEM/UZIdSBJ
wU68imI/VVXnfGq3x4Y0B3vW2k2Malml9+g7yqv/SzyGgbg4Mx1QcgGG5TV8nFGw0XCzkvpfp+ht
B8J0ta9DrW1s4giPIYE3ZIiIV2RudD8dNtgjyBo4TLXWVNRmi1ZkVGJPteCQ5I4mhXpwYD3sCHnY
Uts21LPRSFowdpbCWpDAp6SAfhc9TbbSNvt0rA4lSQaAIPfSwNttSUfgdaAwgznz2yviinUFvQh0
vaSsgJGHBVM1gFEjeqwGvtelTZHV59+YqdAkZJZZPKxnZL472yP+0tKWUEW4EvVvRa2wzSh0ZcBW
vApOCQy3vQZTpZI8fJn50ocrEI1b5Ze1+zs2Zpb+rt6JcKIz2aK47YvIcE1GkofOxDnw5bjZsyhW
Kjq1HT6i9i55zXRAoX9yCRBS19TSd5XhQ9ExOhL2yMqYeSOdag4vaxNNq6gAzzznzl0kW+XQ/8BS
dU9JEDP3iwOOGbqAbwA6Y46JO0i9tLMtu/0vydgqBpJcFS4fFrqr8qSbcwViZTW3rrNGeO2BPQjL
3/jXrbOndFH8nUcwRmeMQVhWDeRRvP3fl1tfJWupYzs5Rp4vQiLJn2TnVIClx6mEbcI3JkW1deU0
LXx+TYUrWTtk5s9TNPn+CDoAsn7bBy2Rff5WDO3ZcNEE9+FrtlLGCkqs0l94aSQUMHKJR30Y/pge
xqk/Yp8PhteC0n5DxgbqhTBUzPYj4qmgJx0F4Kfrl8dduvd5uddfVaHa0eEZSCv05Xys5KPXUqXG
7trKTuDK5lkqyN9sa1KW6w9UBj9Ynl+q/U/dO6woXC18dOWKGhj12o/IiD/2N9fB4ntPhGBoagND
02GHcozAqsgid3WIkONN8gyGesrpsgkfEGVEyX0dDdXF0uO4bYnHqANNGbHK83CAGLwhMUHrngpx
YVvI/IxkSq9DnsnwVZLyrocB34ai5Da+HVEH/WAL0o7evyMuLbhcNSMXGTi5VTntWr/G9fEkMHjp
DKE2drPJxaMofTLfL8Wrbl913Gc9iUOza7yIP0KMAYfMSM8ATDPRiR4DZ9O6XQxCStAoFk6o/ORB
XSsXYqifQqup1xLWUgtXiNwQQMfY3LzuNk5UhfDw8IDEr1zA/Q+n6+gzoB5yCY4k2c7apFhlWfzk
9UqwpFkRcTDzKg00CytT45ww4B7Alkl5WI1jUU6EPjydcd6mba6vGhlrr59eWlOjyGc1QIMYqEoN
IT9X+cYXWBi2IRW9uOSftWImAw6AUU+glKJ0m31trAxQQcP4bT0hpcIRXoBzUuuPpiXPmJzcRkm7
mOODrLhes5z0/DG1mynX8y5kWmA2HcjWc4kMxq7xXuZ+9lO7IpG2NjRHAzRmUYh0c6NdgQbB1VnI
/WFncDEj3Ny9ltyYErJBldR4X/GgkJFlAQfSSJE3j0BQXea97f3DePtyGBXGQf7h2hcqcwYOmZYS
rJ4ESltCwamtFnElFrXg+6ow7+wBS7AGYog6uKJx3CARVbbqhH7tkwvJuzd1c87h6Ko7wuLfqVQ7
P6sXCnTXIKKkQa3VxVtS8n1BhpcMuMBt7TH4dEfOT+06AhetVOxmwGNK99QXweG7IBQAGRhj+pgh
Me0McKVBye/a1jKyY8gPiUmvs+9JTKr8KLFAJvfYMxS0/vRcj/p0qE2/B2LEhDS4hLe9Fg+XttNI
ODyB+tp05t1lN6GayWGseJ9mgeQtzik0hUPpIHtzrq9xv1HXNGqkFwDgCWrr85IfcMLX0wv66Sez
3jdSQDj1nmhhXMlLEgCmZIknwXRqSVtvR9YyXI9mTUDO3GFRLfbG3KdlRTb06vZm1Zphy/oeyuKb
PZlr9lpdOnjeSJjHcNiLptiUgMsIUhrkcDgitWb4RqFOzidgfSIhJjYK1MOmQC6UsUAfvZyPbIqz
6N33n4FTWAlBVQVED47DM7h1ubGAw60Hsc3N8KLVgMGo9aS4AhBbL+Jk+zx9oLtMHRlG+psofvnP
Tx3w8GRenOTfJWqbnPEr0b6lvnPNBZREupUZbGCpO5sxh4xwCZOkts0tPl9FZLQIrLFqAGNlhJLg
mu7gnaLv6wN+fEkP+04z0c4KTLJkCces6FmI6cDNYpNvly0SCEzFRd1Vaqz+tFPoJUg9X+VgtQn6
tmjXc8qqHSd1r45CbLtbcuYhlTMEBflmI9hY7NxWGQkUsP4SBmI2MJ2kvgD0jVt3exqIdVrJhPyc
pC7j3o66Af8/yrWU03YfAxe8pR621rX25hfvzRcBfSXQ+tAJUAwsWnSmBEAWeL5XWDJDrvxyXECE
22WJFAxxkm9WF7fV3zZ0fwKQFq+diG2N7u6QZUb2DnED+3IdZ7lCa5O9C5LYUwkHzIK88uVJkHas
lj2l4HiLcUUmUnI0Tc4HTBhnJXDTOIKuHfMS85E31HZbvRTogeYQPb6krMqlapD72/UU3nGDKznz
jZz5T+LcKrPJnHNJQCi1qYO7dtu6EggV+QHYyIgSD6MehGU2QMEsNahLFSmNJwBN3pZUkhNPRbNE
p7NLRTzxi+XHBwpa0LHrJudMki4c+eXPUf6hg00WikJgwvPEYmsXsxCejy7VkUNPzMVAEb5+/ZEW
wR3yJA2rfZfmBy3WXRDXC53GYOEDZlgL6g3nwP0vIgtUfpL+WrfdreIRVU9mJmisW+CN49cSp1qh
OYwLtnBDXkFRcYEetCXL6vN62BhO9RVwOQB7dpgT/vAAfJ/OvDPBVYz4EyOy1N+DA+V9Mfa4344A
RdCrTmLrlpHg8WS6HtVxmNgZf7CBdmh59Bur6+Qfq6gYt8VyVkh+XgXogDUHlzd9FPyv3CEPzco9
f6pZggEjnxhYvia3oQK5Uh1YPuSiopakYeC8tg9jfwhnJCksEQmn/MKb754Fe/qV7Luiwni9cD4c
fORQ9QxlB2zxqcV4iNG/jrV+5cSQEEnXENTQg8reINGOce6Msk6iF74J8jzxoEZRwZouAiaje5xn
mvo3BBQVXUWuJ9jJzcUXCI7qaxTFVmOVe61sKBCkUoYsOd56CejRr7JajHexTOr+SIl9exApXvqn
wMS2QM5GVPKeLJjwG44K23M85SusJmS6tdFEJP+qgsutBMocG9QejZeSuvy9uCeNuHYkLUtyTisQ
WHFm3B/3HZUizjOnA+LxCsyQXRCjLFixuBmc4kHl+oqkS1mSr4kvGprxG8Q4SMV0mhCWndnIkXdt
arPbZIBD1c4spg8MF6DCjlfJu7rA2f94vkslUiqndIRdRDnvHHBDpq9Fi/3Y9KPrXzqNSXOHAamY
JTMkOat2k7fUvnngxT/XKd9xlDrYkXEFykBTzNrhYxqOTr4MLYPlRYdvgym+XgXL8dB8ZJlKUJym
qlPOlo7jBx0aa4n3YT8WX9Of76eAFfS37YyneFCfrBr1b6/KBoeASaCs2R9u2bOuwtmvjVvl0KXb
7lo8uI/PQ2pNunfQWmrdRQFADvP10ZOOhNsFKn425dyqcMSoR1p0hGvRCuL43MFWKfkC+aUjJUQc
zkeFR+WNfZ0Bw23s2Cf1WsnDzy8/sf50LWqQY/qWGe3mtOzJCQbtpWCPAp7rfh7iAhIieId3/RgN
fZHTR0Jas2FzvTc5QR+5ZkOPW8bcoJmYyiLd8fSkVMfZm+3hc3DVOcol+T8Qx08T4lgRAtwnlQAH
xWTfKUvDGdfJuyR/YsMNqej7vyAvNypPO/VnpIXP55sMnrWms1oxSqH7DQnGrO7Jj/CmB13pPWrf
mWCELuf9QlDYqc90s2X7fgLw3jeUPetuE/tMzSkspyJdwAu4ShsYXz/IdgFixbfXf1L+79tZCR6y
3bFeeKAp6ssVMNB4ELK3WdKxmqbAZiYyVLXn/ZO7xRtj72I2YnwAku0cOSkabweM1KTw3VCVj/rk
NNFu0L/But3W1Ymvb5PGWfW0Y/nae/fHiXZ+9Y0anUrW5/l8FWzAIn/lEy/bi5UUKE4TKLFr3x8N
d3c318XXm0lJiDG1tUk0E+O9HbjdCUsCLndZ1OXJeOrrBu/ZnypXsUiCLuwREXWGO1ZAKV5YabZ3
vu95sp4SbVUbs0jOPefwYE7eyH4xNz3b0vrK7QjpFXTCSmRB02Yh2pkuPMzwQvemNwLg0rqtB9Yx
jOPb5Qrn372MKX05J/OWUmgi/M/cJTj1S8R1hBQu+9is24njdhTSZ3c19H/9zH7Am3wRVWe3gSmK
wwEeKWBt0HsdnPKWHetvkTisuxHkUidVEbP4p8IAqZCITAauvc4QBXfGdIc/aD973ZXyJY1YJdOm
fgkdJT5x7wnq7pfRFDTkyNKMbFUfM8GU+dPoOswSXPZsXQvQU6y5MRoSTz+hjN87mygpaHuVXmyc
9LtjVLKX6NDmaZNo8L78gJgarndLeQxDMgnyDIJMTRhRjtLOJmBU6nG6UyifDIV4vIrzFiwJt4W+
sP3niVFb53kGuFbanTr8T/NX3VWAHe6hwk4kLRZ1ymgTstXK+cSrl6dupQC/SJEm8O9+Nn5CDTIf
/2k5j2vwh7osV29MyML0Wbi652vh6Rh73aJWJsE0yp0pxZM7nZ8SursKjUH66QfJ7lDH2W+kV4cO
EXvs78pe6c5pNOW5MO4CBd3oq+kmzPlrSY8qK9n2McbIoXAtb+vg6wNjBPGdIgtyVIS4Ph1wwMV8
w6L54i4a1VG+agCr4Q7u+oA/he/zUzATUZE9zs13NarWsToHBbAgJr7I4LmpiaKqxQQrHHLtUhnY
Z/nAQzbAD+qFL5gjftCH0P/VIb9c/DF4iD67QUB57rWuDreql0PfjVs0OY8jeZJsB9iQLD4Hf5E9
ZtWllJecLqLv4tQZ2eY8ZHdkPqyxdLr/xPLXYZMJ8Ydpw2SURV5ROYEHrMxUPSZMG+em5XK8HnVf
F37upqCrlF8NcMYNrFzzTiFgf7X+mKIXk05zKd8uyCJ8h0boGRn7wlirOnxrB03I4UDQz4/dw9aO
GJD+JdKRvZ4vew/TZk6/zhaNQpbf/Aan7gV2hBeEUT2RQDjXCuoQ1hRjALeTMlnwb1AalXdOGX5x
FrwASUhRFpDP9Bm9v//VwqL0HI24SAVW7Mxh46vc+DP4ffbKe+82ucupeSv3FNouXulXgL8/kbfb
o+MGi2RGGf0feyoUqvw/PFI0VNq4fg4b4lWqHFhxg4tozT5+5gIPudAVmGWGR/kT3IYAVaVrMmhK
oiOcLMYLpQAgBfVQ0NyGd6NK0Gu5YMnJG0YuYsiDFIxk/avc+8i5X8NRXZqOZ7/HPzPfqPrVicXs
byxsyZyIpCLpHFOxCrWSfBsSmszavplB1txQ4ZF4nNxopzifcNP0pm/WAZb04Vcn8/naUHk16kHV
OASyNKU1do7YufXLgkUERQDiNudYe2ba2YMemCcH3yQ7OVwkp40mj9H8Ifpqh4saMvqvugIg5YDH
Hslc/wM0BmIv30wNIpCY54Y/7ovbIJSXQSvbQrcv5vKYnIBD9t5JYKNah3xKXXAwNeA/x6Q45kQN
lv+h4eDW5vxobXO5CwasdUd572b4YI/kjUfwv/uHL2EHc23SHTbVVrwwHQm894MdgLl3Dv8LAQoZ
Wl7oSE4GRl9aN1WAPZcmf3PM9TLFNzXnzYDOnLqqORXxO956IRYTJCm1Pv1YzsLgvSHbKcEkWNb7
VrqREeE5Y40Cj5gEXmqQ5dl0IaZimW/+2h1EKTlhjC5jIMzQTYXJk3/iZa9GnWe16DpFTkOWFq4Y
a5ZcVR+kd4ykeVQ0Nn5iApnEmj4Lc380mmes0H85uIYocHgGHvOWBm3mIiJcRs/ZWYghLuaTHZ/l
Gj0zL6X5wWd2nhK3n+441R2hFuKi5aGKpTVrSv9O9HLpKv6pHnd6NtcQQrOu2fOH5TraFAanN3uC
/3vSlcPQhcQa21RlA2EbvM+9BJEqCbe0Rx69DW808no1mPI+lbyHJe3QIuit7jXGRuyy8Zqv1wEm
BgIXwopV86ptFdfN3o6FFUh4ZspLpMOv6wwS9qUY/fg+kE4P1wQzu2lmBgFYmV9JJIgvp8Z1khWR
ca/ZnlHO5eUbNAtz7h05dH/xS14dh7zuHk6FaMx+SPFjdiRlmj3q3DHZnpCTqOOommraa+40zwE4
9FyA/K0wvarxy5SL/wP22T7Wcoq3p5WY3beXy645aMBf0clrlHfeX6l74NyvNx64sRY/14dzBhv3
lmZqWVDPRXENbxUUf4bmQMB66gDHzX1YSpI57cVGsj2mb7zK8yrsHmre5U7KBz8M+yFNAnLNOgky
Gtqs60k38tDCAe2GWqTpPRvs9ndHG2qki6kfkSY4Wskfy72fj0v6WaH9M+x3o8WN89T96YoP/ikh
5Qnks++2M2BHxI2YxSKkuWkOFSN8UCH2rGHhXD7aJhyjzMJ+kaY6u6uXVbT/kaxAREhtuXkQ9bQh
QrM4lCefP2Wn0DdiUEGY8LWx7VxbozpeF46IioJ7HsJUlmqtm9H82ksxgH0JF72cUc0YGPOsrvC4
bPY3t754gDn21qcKzYG0VQqhuGAoc1t+Oh3V9yjQAZbheADi2s9Ov8IVOZ02U6Qmt3jHZ6GYLEIY
md5Jfe3rgHbagpoNHtACHaCrerRbBc+xbPfv8eRjz56pH2qrIZeRNoJJYXEX5n7cCCoYUtTafesg
FMHqxh12csuR+1o2E0SbuOp8w9fa5JMAPrsUbLqWjtlKbKC+vu8kUsGhnzAG0kKRBiinJSyOxDwF
S2LkJ1G1a7b9yyAn1B03C2uFNCGen01PbcE/s6Y8ns7p4E0HHm1Osi4bUuCN/omwAS0ZomMIDQqK
DmROjKliCUzrXVnPgg3omrw9OjpZHo91nHYMHvZHsHBB4A+IWDR2fAxBIZtpRg3QNB/+rilpOxUi
G3E49k5nNlO+M3E5kpIZs+Z3DgSOCPTldKtjDI+Se5jhulBbCMQYFIEyG0QpiFBO2E0rhds9Lr6t
r3+pdheBmFdJdVOZxdClJ3M9xEJ3WjNCKZMWFmeHe8w72G5sF4zkeJHTjUYGqf8DsBTjzviSKLuN
QpUcuTSIaQPDVRJmaJIYnKsIAHJcImpCpXsrrlviZ7nYwYuFmlcS7CySwB6xmpc+JQvxE/qDSpSh
h0qr/bAVYASvXbyhhqhbOwiV+vgB1sByEaRU4IHAMRRBHQXO6fwomg172r/mLDWPnCqLGURw4Pp2
OSuEC6NcKrqppVf1bTaxXUqsdeZqy0iP1H69VDA9ysnoe7ISZlnmf8bSCT/nK3Gv6uqWXeh78lck
Wo+q7exqCUMjj6PLdu759F2Qtacm1IXOT46v/FaAifwOyk0OKxYk0hZx+2dn/erO6jDx1+eHyZtF
bA2LmFsl+NUBcaloVASwYO8/OQ83suPK8M8x2vJ9JPLgUGZHAnO/fQQYVTH6V0JQeNEcuyvKt+3Y
pnRqRtdYPsL+6kdsdcK9WTAH/fhBoRM94MLfz4aX6AAdBDijGi6DUMb6LcsjvQHkNP3KaNR5wIwO
EvHge0kBTVPwcWWU1RvrffT9MSGSFx4w2AVrj1kkWTNG5l7jz7NhevlXBlczQYHmeVUcdHH/RUAr
/FTRzon+uH5n6ioVHWTC10ACLVc7X7rw9AcqDz0eBg2lG8c/I7gwMQgY1TF1zmt/W1/W61bvHVtF
heVCrEUfGN772o6BmMMVWzUSjsKbyzq+Wv3ATenCDB4ckNfjqlBoD7GKGfEm5yDHT4MYfISQ8MEi
FhGH+FRioXJ0dNtOz6gyFUYvbVpsK4TsgyfY8q5DGPOLR7IciIMLQuJOQV20rR8Lkz1XZ++cHKgY
TGkiwNFVUAa5/pxyozBougQZzfcuLluEVvFSLcxZpyam5HMkKiuMTFz+Y7ffMdZU+k6VsPkalSmC
jAcozVqE2ZEdIwX4iRHtITYkwDWTYAwLn/Ze/zQZ//4TOvB5K+yj49jAJ2Od1PvymqX91COPh+sc
PZNUe0Nh7EU6Uk2yF0ABrzjrzO38oJO4ICU4d2AxM897/jDr3pPaKWObFQz9mCBnRllo1FDZJePc
vQnZpYlV1YxaQo9qcamGdzKINHWRAmabnbx8IN5emKFB4QXpJJsOBcmpgSTdD608ppm7Z2LXvwLk
gjsvVlZdLPlslmCzGt6/gv/AqxLhtVBjLqHpOvAAK+EnQitfC+/4LQZATb/AbKt5Kf3QigkvO3X5
xVZHk3azxd2/5NPJUIoAhrPHQe3L5emZMRJDCgutqyrX58l10si7gNx73lijaAgIbrqZ5TGBITID
SURB5tOsrKQ3FEnMYPl8DTX+NntOcQWBqhhmYrVaNuFv0cCKDOOap58AjuLSlkgVxBzZX1s3Hrh7
iPc/OB5lLhkoahG2grvolxt1uOzXHH659y1cdpSLHMLwXpAOkQuabuZZXOzSQhQLvNA0qDuFKXBX
k82YAva25iZ0IF7KkNZkyot9F7JEuQoU5qai9Jam31QjkFeQc0p/C4yFSabO7OxWMsXi1ae2WVIj
0ZRX0YndVR1iUq0ILfJqmOruhpzVKdNi2d8CUP2+hWXZuJeVuKMasMwnBkOXTzBHf6REd2gR85tN
bJ4km39EYRqkF5lM4yQBN730r8R4G47MHO0rsIshbM9OdgJeNS7QUFmXRVN3lw1MByAHRzDZ86Kt
MZM2iiYc3vOiwelSVbo0Quo8g3N2Ygimw+S11KBrmD24rldVMkANZdzJeekfrtX+mbEbEZD42QOF
gqbkngLFb1AoaTXXYKBWbynf0a2w85r5LdzTqyeMp1kZKtAZk8Osa/XrfIXNXDlzXs2m3jOkq9Us
gKAaqke3viEVfFM+IpMtrLNNkhGsmpYltnv/dPAIavrSouUCcXx0pQRv9lH5gbyNlnChGrVp3Gey
6pgKzM2zUEvQyqQ4UfP3ezU5L0d5AIQEz9CiGd/8YcgNpNXB3ogmcR2BSbWrkG/EX7JI+tuKI9BM
f8yP7S4M/BoBuRk3x+Q/t3YpgtAhp2ePucZmiBjgIMR2s7KNlAiHnvt0oUwVD81xFc+byCoz/OY8
inhiKdWRdDQp0O0TRq6RbgvsdypHhSFgd5KgIWog/xC2ByUPTkXzYKQEfTlPJEr5il28ZZfZumTn
9kmxDV6GiI8ZFZP0ApOVrpnezXcfsEBMSzejXXtGYbG+sIDIFFt8qL2mYicA11OpQAeiw7WVus0t
Suzx4fq5mwn9pFsJ0S4LBCeZpdgvUVjIZhzJfT8paOJYNiiko4eFAIBfwkPP6DvfPwT1c8bfYXqg
WWL+1n4LCp82BTkCe5uyIZF9nGmTO/vDsTo50C3OTndz/4AM5P/yNyw9fj8ZrCPulgJykhODeMGU
1WwRfn0hycPZj9cfHQ4rSF+eHrlWZ3JigjFQikzRC6kRztku9NZzD4WW1tdN49HAoRnbHnxPkWDr
tVEm622mA0Xzbs1FiHyyTjgAqpkJpfUeAXTomhsYbp1GSQTMnXziy13Q+SAeK2OJ4MeFbIy0Er8R
yicrFTQcWACIHGaOFa46AaPRCNrYrgX2asLun225esDXst0bzNRLD/MbOFtA67uyA6OGtt3Hxoya
iefXVkeClz20Kx2zo/jsUFjQ4jrj5MXwLFA6dYgoB5eaKHLttnPl/e70FK6Oqq/m8QYCzxDI7t5N
+uvRIxKILrzFfKC9yUBUxVL37dncF1RxwhW054ztHpa6kCVpLopYsfSdtWoH46PaeVKZdaW3SKbO
lylM2qsqRirN0L2L1AwzSUzuymHNMUaKbFME+JXHEWc80fYqExwMjHcYP3QXGzICSyveGFim0hZp
fDOS0J1k8gz8qn145wUkeQN3MSqp42iBQ1niAeUj4IBebZZGr0y3BWZL338DDV50CeS0BbosKqGK
unWUmVjOk7ahReT4QQEONeTxp5u+Zdz4Huj/+sWIbypRaLOnNHu7nS+LvOvO6l8q5mNz/Qra7/YW
wLjcRs9JJ7Vvmw00gmQKP5bmBswEDewPDL5WX11aMzaQzWXvV0z8OCZmmINOuJMuDBEU97vsztpC
rosbHMS73JmjrCE242PAaJqzIcwD5zJ+AEHUCaCaGYONaxZCEFUHVhHdiW+U7dAnqLpujO752p0O
w12Db0ZZrncP5QV/lBfsXZ2yLk1B12DqaY/qY2ZHcTnB0yOWaCThT66WdMf04t/g2bDkx8071ANy
cVm4kxBL3CjFNWvyg8wrDSBcZOvHmwd4zx7YGQIrDcxX/y+ey0rt1I5vdbTxpS0+CdZPMo/i+Mpy
NGR5npY4/Yi209xqoxTaelq743r/TQ7RoQcnVvJYL62Kivo1xvvoRySb90CWjSnHJhco2a7ZzKae
ZzCl6jjaGr8oN1lE79aJjT/qEdDtgtBSVbDK1gweiuUL6+noV9unrq93sc6BtF/73QXx71vt5CQn
Ux1F1+xsVm6k27YnYdhH8dU8QJFkE6Bvmrx4I7CAmzgD47kQbl5eD0/EnvBPJhPjUhQ3fZLUMdNN
sWExe8Hi3/IcaGy/ut4T8DLfXaZ1qLUkfZXIaJeZ1reVj17USk8G6WyiqvZ1Ku59Gzd1SwfR274d
9suxED2Tmrv/IYNRuxBLZq4hMC5hFYJbFfTqT/hyA7bgk+ipz1hGrDb9DdMLtFePKMgL779dRCmI
xNwqxYDRoJyc32DbIQUDZoHZ1QQaHZ3toq1IxczbsIA7hA5LjO7aih8shBavtqt3TrPz1IHlrg2q
kSN3mQvNN8Lim+UE5YNflKfCv/Ou80ZLsJC1e+Lxfi10GQIXRUNqK5i6FOfHrpF2aoxC0FhFVnYE
mp8wat2RHo1fcONG+bBRQcsz2CDCFIvDVlOx0DfEROIMOwhtuZclWvqv+dPX44YLKFsoY216JEfi
CyoNbGFekQSET31gnoNgjAzmgmuZGiHy7sp5woCIdMGNVJYX3AABuNIrEvu1uad8y9+t5Q+unRx3
fUtVj+de3pUJObUOydvugp6S6oJHB++2u1XqIEf918748FNhBnEYA4NfwqpmYc965NWCblxpdSgP
cHELHoBmEf44zclE8krTVSJgKu91TndD8LY5J6UPcI0SSpyhidkPFF63qr8GmMvdVdlYcb7YbA3n
hEEaJ1cbvTvWgCr09VfJ93MK71BnegtAw6lk/sz7jBVRADuOOBTCXNg+pomZoyV27mJsm7ePpjCg
M/g4v4jYWaoShb7PYJalMikw0EHCi6TJPsuRv5GmHrGk6S7cgUGyiPSfs9F4caPD4QbKutg1v60I
x9t55QnHd5L2944pRBuc2SiMvW4toMzsWrKnEfMqsrHg0d1aWoI9VLiS2Ih/vOKGLD3vBDYMXzUU
BzO3RZZgVPpe8fbCcaiLQwaSsroV05DfZBi1vpC4HfEEoE/7rIOexqmPP5gwYDkD2QcBIAo2FnWA
exY0licqtBpZgckupoA+88QwkzG8OBQnzw147oT3hmeOsrlASTIjpprqSSTDr7XZPNBL7/gE/BN4
OYR156rFX5OT74BJ0fa0Fa8XBX5zWXlxBCWYkCT1bONQXx4JYGlVI1oJK+cjHbYv01Xbj/WJp0Ns
iQArjHJN6nOJBQ998tjNrs/bPiOukNe5s5K/h7dOy25Yz1/z9FhdXBUYym6/aeGiVID2pJa7l1CK
9S5+/chIx085iOQHryTKLo96mXIPvICxzq9nILQhJU2y2JrLwFStyvUx0K/ClJxmxpsU1JIQ469M
qYi7oVUiO9qt033LAMOFRDgar+qVEkUEzarrFFDYmJ3/ZpuBfG13tqbbMt8a8WUHAPBCpYMB35LJ
3wqiwPGWYmMH3137a7Bd8FEYXGNJn+Fc48lsVo080uPxDEAyET0vjboakBmTWQAGo9EHqgo5PU5p
QXnVkeAPY6BIn0l/nTFOnnJcWqRHs4EzBwFUhyHvmsQc8MkGHAp7di/Y2sfu+WU1d6cHwp4+cIDn
pTnnVMC180x1xz6KEDGvzlKraWmzzyzQC52PTZdtMY42R2nNMyRbxFdGp8Ys5e8IqfYQKAW4AgTG
R4eUASP1ZWbggC1OzbYL60gpBFcocibZrzhOzHPbKwZqxak+gThcqUgtNQJuY4SG+ZjpM7i1zgqg
HebRRdsBikLcmeOCwcS27pWfiV/au7SGR63i8v9Nwp+WQMJ6JcoBfTj9xo8yp0FlaWRfVZBMZLll
VfUEnUBlO6LYIuL6ZbnAXF3e+V5aOazER/A26VQZp/5i3tGM25HFDbu7nSRvrFP18MWRxnmpGkqa
uwXg3egg/xCFNS2+w1uD7feEYSC09wL74Mj6BOZK7kXeJvo2Y/SZlOslJnRqHW9JikhtmPth31In
7rl1hrqSPRUcH8F/XY0KA9/7ENNt2OwkPKyAx9Wz+dDUCCm3TyRkEvS19TV8xsawd2AIFJDPTkhw
4MRM6Zb60oL7NqTt4oeUPQteQbxffBfcs6kOPOOVoWzLsABrzbMlUzztnYiu1u9UaKxeKiYGK2v1
3OFw/Lbta6A1vmAAHBo4dTiuQg+OZRd0gVNHMiUhnFmXN73o6I2qLX1YGlEyZ3pC3CH+eCNcL5cH
FJq2ElnTZ970Ts0Eb7TgwB4/zMJzDNYEMYvq0xsmRfP6Y1a4nm0VSW6xAI9jp+N+COMs/T6p+G/u
iMmqaWdrxewZLPxyLgwDdFxIw+zW12ILGoAh+c++EUqZGcvnGlM64p2qxsURBg1rDZSUIT6ImLD+
ZtV8wcn8MylsTYn1bxBiZygVQazST7Kbk8os1fmsuavpWne8o5nipLTWLfkhy1jfexK5DXmzxH/j
D+KpFuK4lsl7tXD8R+6ViLuqPweunGsFPTnKeDaSk3Fc8pNmucbToez8Z1TujlihLmbRJA5oosQE
qW+IRP0SJ9FZHu+yUCFsvrbFSIEE9wWMpcyoZK596hOOSXUbHjlbHhpvfTVBufkyHj0nSKWzZekl
+bybJRCg9beFeWmmK8p5N6UuMi1pHP/GbQKs9VEppyhG+cSlChT0h5qXeCZY+7qPpUgcK47+aQSr
PfeZmrBke8+pQpFZ817ZiL7Y6OL/UWU+MVGYMBG1uA3HfvfRKnotO3klcm0SN1o7ngSS1ittbfUJ
GxfcPcfe+1WsaBsNyP1LcNzS8c/L4kvt7g2FKSoQsZBa5kUtF6pBf+HTn+d1ZnW8dg7odcBxn6Dn
gJgfW/pLmcytYhZN+q/us4oQQ3Uz3YPIB+Gk34O4znROtf8fHv8EBxWJDg71i1bkkaIN8ZLbrwpe
xrhOCOYvFO7hjU944SQLZMB7yXmj6SgogGddohXF06CHC/w0XZNy22i9+uW/fxgZ9E59khsNzn3F
2HRTpsGK3USOCXyoAuxhxfPFa2SDHtaagV5nhFoYWz2aF4YwXrp9KAphYewFma1EfZnX/+TUkU03
Og8npfGlcYiGuDg5Nq64jRBbN3uS4hpvaOlF4DW5sgLg/6EyoE074OtH/rZ7x9Wwv7EszjQst984
CS4OHa2r9a37nYAF+MkoqsWmm4tKZ0le38T5XVtifsJ6U23+0qQZwV4bR/XhY7ruIAsNa/64/HpN
Fz4V0kILUpjzad0rBhHasdwe+qLjG59ZA+0Bdy2/hR5uPuIRvO0xw4GC7fy1iUWiRIsD8dm/OKU8
VeZOOY82b4C71neomJWR8K6YPYBZagWC/1Y2rH4uxoffh4YQ32Z0Ws+nF/rlgoEUPLnDr93539bI
fDui0CvEbfeWZ8B0SbDhNiH3UaBbruEGyyQlKggWItEnOgIY6ztgOd1/bURNP2blv+2iFzKQ6k6R
jHrGJDT1ichZAUTowkqQVQKq9L6euRzNxgou0qAIdByYAXxZqsQjAiO5ZigkGNc3w7JATeURBTjD
KN2KmS/gC77rMkYuNNtc1CrwzY57lMfLH0iA+Iwe7+Ev6YEbZkvaB9GuYeCxnPK55MPCjq+cq8+P
N/zdJ/lQyEAydrIUqGPyxebbGtXrUufsG1qvWEJWbhjhUG5jYhEJeTlmFYSIUv43BXifkkHE7gky
7hya4xbevD0n6ySRoyS94QveRFQa6YW3Calx5IYawQLazbliKRsaA3tnL5V4eWg2029uqMpRizwm
Mr3K94zmLTMy1sBJzVVqS2g+q6dvSan0w7o2or3wh7M+hZ8CFtgDkjMKL+UDnUHxSn36CcWcIdwW
S37HpVJUOgkw+aXIMpcnEigQ8wGwoyWA1JNt1dtzn7DHzdxG1o9a6LZ8CXYRbqfWMPvz10ew45us
pd8czac95C2fox4JopJrcv+JJHM4KEDeWyoOVTzuBKvV/db0jbWGfZLCJchdQq0G0BFOOEOXGvS5
lRSLSdH6jFyWAclhvoCzi0kcbJTBwAgOfbdERJ8Jx7alBDSyfyOURUP3shImAKOtPcfEq1IUOfwK
Fa7nAX0RrdNPCKxMYv00yu20Ru+PhjEcoyvZeYkwPaWcNyPLA8L7fnw+lsSr0F5oMde+HQFCz8Tz
I3E4GIwVJ5Jk4sj7z7jtXKhkFBJL0icMceI73L6iBg95n71EnWh2/GoK0nPoOe6o3e3gV0TC67Kv
HpLAsAazrRzLtsDxd3EZCjmOE0zy9MygmHscnmXErCnbbu1t3gb7Qu709oeyafuUyPYQUPxFvJHQ
yz9Qe7bpa0zyKSGuo3OtD2uUerygUIEIrDxmPbG9qtIPD/g/heqIRbI208o8J0pqmAaEyR29XHVh
SgUR26xD9JuOL1ZDp4l7RKC0rgVMq+Jm+syIt4vsBEJGLqyfAmS3Iim9IgShlZMATGvNbqsge1vW
dDvAZePxcj2ZnGHBv84HsbA9vuqy1J/9vHq4sZBkAXFGNPIMyYvjInu0e5BkU3Gyv4tXSIAzyzSk
MOQpjw4721jrP/Kb4jG9afFFgrnu9xJ6IXB3HQfYbyrEfx5LLGZMpAYnWkLz1xih8l901PqBuftT
MswtAZAeKIMGYzk0z9PtwlwvuLK3Esk8xdMu9evBxpx7Bo1u4J1CN+bY3CwuEk/qAcOj//l+yJfb
vyfazxBu9OPvKtH+w8MpdUkTR2vASxllX5cJ55NGsD8ZoRMQtl7ho+ul5wM61tIjnlNIqwI4dWlC
GNIxpcekUNaBUzryP/PG1vWunKyleFoDElOJrySdLaL4CuJWwf9Zg2d3H0JGzgId3AjwBkE5WnTl
rSy+plHkj6jZXgpHGyINsAjD9F1Ll2CC7yEcrv9zBMhJyKbkznUBm39jpR/H75GdnSM8akB5IjMX
yKEd8/Psq+GwZuP5WArTHtTgg17rKrhGdlsNNVe/vrZBiJs+vtdPyinLCbsqilHeIt5+l2tgRGTV
hevy78wkw8XaK2EznKU7Cjlog4w9EtU7md7TJLXBPtBz1CCpMCv8nMmAooPnRBh9VYxPeqaVCBLv
pweadZIeUCzmSYMnNfOLUMAT53nAUBroNmCMCnm+/hN83gfUhzu0CEvb7i491d/Dzs8G3pd21sUu
rfRmSwhiSiS+gBmi3aQnbkwEY0A/djOB1rd+O0EY4TfpxwczjHDElRvYHSYD69GQwpPszWOrI+wS
xlbGeyG3o+T3+CmDjNF0nOJLzlwntZFUvJSZgFVuIjzc9qgh5XfyHWm/seZ+T5gHtZSO/h6cxwo0
3TqMx43QA9EppoEr9bOgE9ma+kn1n61t00+JF/ebbWKuxQxd+OzVCagaWB5wYmrOFAdInVQgLBqW
X2lwkV7WEM2RBKc6h0GyzhbC7EDLIn2quVwxkJexQ9pA5WLJuvkdI9BT8seu2VdvwuOHDp4PTsaK
I5+nttuHSYJJ1op4lxlzTJsgWOj8unmU8wrIciCFhuvmsXNmtAVoLZrc60hrOHaEQgYzvGhPU/HM
1/vLq+cTfVtSYtDHENc1v9ICH1E8dMDNlVOq6wgS6DwKH1TX3EI6Diqr6C0En+g4XFwmLVZIUWxM
r/GjiPV4OFd1x5/3AM0t9S+uT2FWTFuha5K3IYJ2ExnKRnTDk6fLF0WaLNofbBwELa/tOS1rEz/A
WjZ97Xmyc3Wf9k+jaK4a0mwj3s/4kjSZjVG4w2IedYwk5O1VpIPNPvYcybojtYHghNOnVzE3YlS9
IiS5PmAImXovni36/XZbpr6CUMq1GihqXDJKhHdsPzCLKXXRfccyYI64AwRMoEeNCdKEkxFH/tdp
qBIzUxWNZXnox4RfceWHlyFr8ykqnYYboiVQ6bbgoZrDzS4hnBUafth9pj8dr/9lFaVHfvJv3sr/
BpS2a9fbeYsg3oRXD1sXi3fYx9AYF6GrSTX7TPi27QjWqniE/vSptslvHddfYyC7orqQvoT7D+Ra
CPI8Wa78kobH4DttS5afG8sw6b82L69BNEJDxVR1uq1vUMRMYF5jTzq1tXG1HKER6z4b4afDm9rP
5vVMyOFndiHOoJGRf4eVUA9Mg2q4f4H8U0w/Om1u/cF0mkvNCN/DxD78PQGi6v46BSgUNHq1vSIF
eE858mMGrh72FOPICfjcfF1wEM8v5TI6eLWqEqwRySEnHqYjfjOP6FX5gSWXKH35SokuyUR8S4is
PU9deJ79y22vRKxDuRnNKZ39FuOSbdSVyT7o9YJsbhnJiBD5QXsKXCLdkN8lFFm8ws485X/TPrEp
Cwq7dqzweAucbX03SLRcpTr9n+6GX68lEdMl4cngIvDLpGYwE1bAhI0KtOplwh5cqKL747fiWHup
uOYeXeBX5sMWR/ffM4k7z3alcf2ud3W8tE0nAhGc1Af+kCMPDvXN/Hp+cgbvHA62DrqINm4SGfQ2
o2oAwgMpY5ZPui7s5aGZrmTUFCL+9naPfunogX1ARLDPRcLU5kBcT3+q4MGBwpPfj175QInxw3Aw
0Gbe/1IIgrqfVCpdc48u1FSf9Z5LWORYFZg6hvfp7OOe9GrxUyVsl/JPcNETuyyhJJ2tvQtoTR/B
hHbFckGhiWCQZcay7L9gPg0XiBDtzogjB4Cr4FmI8RKKqLSRhe7orpFzskfiiVMeJNsSqOgqT3t+
+0iaMF3KX2yclhjMfqpZxM0WwqO/YhAQjFe8Pd9KJmS8JmCj7hgOxLIgAD3K1bE+2pIu92r5Nexd
RYKV/JJwr9xm+ylm6rjsvvB2Npva/tIsW/cu/otXpxIgIPlo3SOSUIfzpBKmbgU8knjE60D+LyUm
SFeF5hOzim2aqzVUA54qZfQ3yktAEkEi9gAbYZxoxZGmE9dUoT7hFTvbTkde5zLK+ewMhk3LeumD
mTWOT1KKbh861FsUJX1GHXAtTpo4GAdfgIRDuVVWAhefG9yDD/4Qp30I2Kj2AGWKD5qZiCCtRf3B
XCN98TpYMcnRqTCkkoLsrIOFLpsNq2+SsJe8v4lIAsUHBQePNhL2jWlOVzEFMO8AnwXhApCpJhhv
Tim1HwoIUZFsIQyyMgCjl+nYY+7PokIkPhT/GBrxjYsTTL4vPC+7iby6kp083k9fVq7/ILi5IuuL
ghtv8txmVpXAuvZYRR/4JeWlCp8qVLo09QuPDivUEUKv9eUvyoxdp9gNsZS7liU2pCbioG9i/nab
Qwki1ArfHNYPYH1hnqdcvNoLtfWL8OQ1hvfsncKIx9caSGVISCjgBH8uNMCqFTyIIvw8bvKGrFp+
t5tWVO53Nneqs2Jh+hUXg7Kvpi+H9D1aQ55csS46dAuGIoSF1HnNDw/nTKaNeBp8gkFqXPXlPEky
WJHi6nPcJlmwW/u44es7MpN+r+vlVC90eXA1Tyo2i6/qTMFP5bMhio95iTbixiY1XmtWJEZcwBFM
OamT2lAK5esQ+CZf+xBTo5LhlOdDukBHFOX1TLi0WPVQiKlX/othX8CkLgSEAxkPwx/5ONk0kx3F
j0MI+6z7hrn8QfhJaNOQV4qG89pPNZANowLBf5Z/8cfL06RIp20DmqfUJUOxdwnIgqPeQcai6QG8
FLHp4KQGYeJwl9w1vCEumSzPnLPFMlRGg3aYZrlQ8VjwwX60t2AuDKPp5ddm/qXqvumuYB6/Dh+J
szVhxgSyAGCIoCbfkL+Ab1VwkOhCeIJAZq3OLfMSDEdT9zpksXSlUIICT1q9jUq8e0s4ig5JG105
Bf/xXBsWBs1nSx8bfr0D33IcVbNeb4PxN9uIH2By8VzmdQIkzraZA2i0YPb/tLjorSA++mvgSbzO
GJaWKEjvpUVOFlDGEqgeXxS3v13nYwPK9vN+It7TdSqEkeKJ7iy7X7sRv96Vd0QIgci83ogmLqOw
vwd/bHlV/jbmZhmsg6G8U+QhtbN0fJxTXBdovD4l2Xm2CTRXRivh6irVQZDJjjH0wzRXCScm+Ixp
pvxSB5tbVggOs63iJvZxqBB3JKAwMA0CHYks0NXYSW/OSqyPKKkOgp7Rp7rVTR5z24hzW4oO6HDj
AUPSpwgNFxlKrUP5nUANNFwllEC2ztt3T/jLnYcJzzK+x3GLfuYz5th8V+JxM3gWTholKzHJWzQM
hj4x3WMqBT9YCRw8wChELW1mH7JeqanM/FnPMYjFXmEWu8viHJ3azbvBgcXiwMynQ2TDectuiZd3
5PTpwpX+TrU66xkeuLIf8TmkUDtF04JERCAj6/0FhELZSV0/tE7U0Zq7RZ9pCQ8bCWwet6MM77lH
68lrztPgD+mRK7wyu7NT0wm4lNzh7Ui2tGlMXoDuLhgJmlFCXTZ0ANGuCtr5A/0jKIVOlvxkuVrD
J9nHHDAF+9KF6qnWtJVfsBjVjCOtAQwmtLSvQs0319sITKB07ksKlYNPTdddQ3kksNx1Cnn25aQx
+/36QrwLK4+Lj37bNWNCP+yRXgA6z/RBKjZEEL8yoZhQKv2mK2OrKkbyUutqOS/MFQIG/IkSejK9
n4yJSFzobYf7WFjRMrilgJfXUFuTCaxWDElkrJU2MR5HJOLq27jedIdyPS319jCvjqO0Qt0st8vv
1zEIf4xtLpnBlBhaTUKPRaE9ZJHi7THJlM+OkvsofWJYs5Qj5+NQBlmWb/5u9WAv5+Rmy5upt4Vd
ugJsByEow/11Eqrur1fL+BYyQF2Aa9DSCIuGczj3qvMuUkv70mee859eBRj5Jg3NblbwIqTRdDvU
xXx/PieHcGB+7q6eQE6gAZJwlBOTPZxiFdRfC5Ki+NYrsowc6NAnGOEEMvF2dJEDEtGtg+eT/2mr
tiL2ss9EmrhH0HRq7dPNltFRPSUrg1GxKQhMMn9S7536B0DWwlbMnWPku3+aRLMiU+imZBA29rGU
HPH/d5nGPpchE6ThgFzvogmqZrdtgx4kDDS8SAPNuvTjiQ1hUGHmTXGBwC6DJ5Zp4ffh38cNNPRR
85F3vIqw9E2CNoLtBLDRErL0C3xYyCsYjzCW2Pdmh7CCT006niii3GDAYiuG62W6FgxU4ZNfqriT
Vl5PAjJ0Ci9Cm2YH88rp9rAeq+5ga+qInv+Vbtb0ZHiXSzS4qaQpGg1HXyFw6X68kmmwHogzJoxv
vQXF8zvwXMMJCZvfMdir7lWIQWSPZTmwh9yJ5doHLpsuIS94HI8BK94aZf2HYTBndj/FwJh5DZF3
fYDWICMuVRX2XMxI7XRiFvk6Rs52CiUA0VtgKu+0LdKz5kbo2qFlL9/S2LiRJi47pQTi39ptkhrP
q9qp9Eu6o3clRI/651k8Dfi7e6ZGYYt9stHofBRtAThGL20RIcSudYzdG1XEXuuL42n+Mk5tvep/
V+sxFkH/nSjLZX/XF38m5vVn5Km1gs2VsydGtxawamLE5xTTXSixqSXDEkDHw8Qa8fDdOHR107E/
SU51l5UxNH+O92IWtV/rV9Yl24UXbxwbi4JV/xgw+ezIkjd75F2tl4RGKHZcpXXOr6995V/WhzOZ
gE41tILEe9LLpZOMACoPk7WG+oDoHutTeqnqr7ku0+fIiA/HX0HAin5k027UFDv6C+16xodUVUqv
67OpdLjVBHicdaNniWSkJNCjS9D/Uz/SvSVWsvFyHdve/HI4b5yJhuVMl7LsuoA2KHEP3peUG193
5npp6N5pfNYv1XRF3H1D/m9HDOqgDOK5IcLw8vhjJ3k9TC/pnhSiSJLoIOGE6a4hl4p68lVKHNCQ
KZsuWkwOQzYNRViSbEZByXr7rb2svT1hsZQ1dp6gsQTkj9Cu078rTerFhOgmnBYJn8rOH+7xC8uF
x8+N38PW4+l2v5aMkI52ike2ovUymvOOfoI95quh6UcFqaGLOnsFp0+S1Gdei6TRrlnbEjs5VneX
msoPKIZDtDAHsy/akJIqXZPitRq9a3EtxvIyw/+umogW/aqv2BaisryxXeOtGFnAJuEpovdZbr3R
iVUIx9IgdsF9nRZ+vFs0mcs/CPsAeh3xrJS+clDSy1exqNvIBknP2EqqgPf2pNFLE2QivO9J/NJb
zheH91EqJohR0YE5Kxr3nCY8qe1ekLeLYsmTjcn37wjp1oi/jlgCYfHPs4E0HHhv/Z3R4h3Ct3FI
tepnv93FPbZ3N/7JOiN8OU/5SBF9PTBp+R467EawQm4nRdeOzcoABZzkX930LaWX7Y2RTEXeeXsY
cgQlsqKQue2iRxJ7jUlnqKGGdGf3xGfjWsWqEU+ua0RWMb1RJfnGR3IBr/XW2+k8eV1I7DijlDsK
PCxe0V93xQpmJ4SQyp8bookhL7cx/vzcMu5M5MZqcIEnGNQRM4sj+N54F1tCmdMwz5SqiDAyaGhr
6T+6B71VNBUXJ9qC5iE4MjRPnqKoyPb16Z4zIfJA6HVjsGN4U67wwdFS17KqaLUywBsB5YzdNmXs
UPvlzezqS4ZhgS7EOrMm6iKh958nsD5s/1KO238zbYAPVAvm64uJApjwkQsgktbK6UaRZF8Nc0o5
BRRbG+MEVYF6J9l7iBG9LTsWu+440OL3nO13UYE5c2CzT9BN5w1KkdN9TjjR8elYquaMdbQSYiRM
YLGlktAH5rUCYR9p1RQny1IzbJzxsSFFc2yF9JzknzMSYIUQs8462fZGrCfhYjOgvyb+0j6jMik6
hZsvDelvJZ24ITjfcta4Gmnve9bERRLLPrhSwPgE981ZmHgUyD4bRWcgSXl8dwCZKuZgJozkkZZu
cqVRqBectynnPpEevWhR4uy08atvB5NF0q+ccewlL6Djx+UOTCzC+0k22uvdP0C7IsnBkt3w48Lg
BtRfbgIyd9eIrJ3zSKLm0+qsT8KnVAJ9FT4BsaSujO74mxBn/vn4e/k2uiQPsS0vFbeOdZMESlH6
HHNt6oKMh8AcmV9PUF/XGRX8za7q3XJ6jj4w7A9EpPnQDBFn6PHev4bZPlsa7qXeBeS2iJX69nHH
IpEADHwj+5lF+OYvfziW2AxN8waC3wvbjvbyA5nSGLC/h0X4rkILNTVUgvku/Z7AqUmWWb/eSq8d
IsnUFVAWMZJt1UT2l35Z+ve+/9wU97Cq63OAE1KFk3+OnUDZEd6SbQ396MZO8dY+xkwOJqNxk0EG
aAtKCBx35+9MF+zUHwc+lRBfAnT76+cPUDuRmmnR3SG0vlA+dOZ+Vpe7kbp5MAtvtYUFUIRb8DcU
cVNL/anOfqHBRwzNKR77uagikBAEq5BlE1Pai9KRRv+uqjnyi4/pPhjovCLVMaP5C6fsQD2GszZd
jbeXls697TpNkfwKMnLoQXocKCuLcDfxWM+X4zmdopqAcmQmjoc+seeTzsatk/dvDcVxfAdwBky3
18/Adwmg9ii/kcT03PiKndASLPC57DjIjwSDdHRyRh0o78hIkzsFOLgpOudUG9RzJ5dKxXjEkxqe
ylarR+sU2Ovt3dTt0dEM7NGowBF/MjTlxwaSsi3G3EZYBkBfA2IMwP4P+baZh7Kvp0y3q4E/Mx+X
blfTlZq8BIYsexUfAovRPOx48+wT9vMR/oJ/Ogy0yFoIEDeb8J2DDNGT373Af7+vHrS4bjVtc8bi
F8RJ99Pq+0rmLhQpJ2XgWsZPlgmoaXx0ITRkw4NxTaYCq6RnlKW3H113Fc1yuq3XfFKyc0sReUqQ
uTSHXvVTxdl6l5hPdeB71mx9RYlHbtsBsT4l/Hvr2tof7LvYvSl/AKcRpbgCXZ6m6K/JvX/GIHnF
q21CuqTAqqv9VeCCrcNp/5IcmbJxBpMrxHzum6BnoIlG7eW2IzcXEU+00F+gkXoaoTrTxmwoyD07
1cVAh8duc19LIrsIughXh30aJrzo0Bvz1mbIM5xBwFgIf3t16jTH1DmGml9/cGyiCmxzfjiEmi31
7Vf8HumAk+maxV/2LdTj8elyUTq3LgtjYdgCp+bFkDfwE/NrzJU0/UozRw6u9fK3NKazuV68aHA0
SZfmBoV4sgzGbhrIConySDLyvsvtTvsoQphU7YvIvanEIp0JsPvyYWX0foulGRqSgceh42Ctzlkt
3P7oD4ZbtssOSsw2mIMya9C0QJmRvp7J8ehsFx6J8IwbyRwbFeVwPRl5xdNZYNtuNLaIzWU9fuxR
/U+20dILixL6AWJW6Ofh0QD4DSckIEQxF9LVeptnseZJPwstDTY9iyFVWnAdHNyZSG1gAyJbzNeI
WJSDdk+UqXdRDheMa4g8rjVP0izNC1AfxkpPeKqdvJ4fg1c3zjxjqbJ/EIaBmU1us0hb6pWiX+rx
j2S9UvbkbQouhbgjybKdb8uK1w3E2+TYGoysNPERjgkg3mysn0W73ZRIzGoPQ1ZfwpcyAno2BRmY
aYLFgKn7h7pFGSfwr1JZLix5wFUgf5wpnvhMoDvp/D+IUvrAVMzD2Yq2MxBWs2R0vSdDhcCPRTr4
3MvYphETMcVJU53LfToaKvvvIMWQ7jLlD9USYiXsb+15pAKnjHZN4vWEZQ/AT7+DRMY8fdx6sBj5
sVOkYctMMiovSLHYNxl10XzRARPw9z70CpIATCTlBzSGtTpd2LaVha86QIYFmNRGJCCu4y6R4bVZ
jZ+k51H/5l5FKgWk4msj+hg/0NNJbX6tmIyV4vsUpnaDlhi0MhlcVDOhsEd1cZLe+Xx5Yv6+yEtV
PEIQgj5t0jRCVjl8E05PTAx505nnOg9arSSG/JX23NwGiKbyrGsAuakQj1DBKWf4bF1w+qxDQa3L
SSyNqvgXXT1s1I2F6yI5xBsKrZFqSC25WcF6kzqpx+hr6mdKP+iYSFXq4LPmnJBqDZVt44r+xDaa
BJxlTRQq1yCvSZOYYTYKKPblGHRfjcyxpKe86Afkkh1kYv3i+9qiO6Xl6fu3JNbk6qpDLIHMshGK
oyXv94CC7ocNEmyGTfa7hD0BFeti5Bqi72/3gwu9r79Z0JPiXeLkC1NFE4dWsH8/TM9+6CEGyC3K
/IgcrO5xnDByBakmmCtgjB3jbbBIz2g4yoFxKGa7XYj6pGZ6MOuQDEV1x1gvEKLSZIbzvyD6cYae
d7NuEV9aCUpBawKq2Lq20L/hSgsGp5XV8IBgjpVbxiGzehEpLs1jThMTjvzThFmRZW0w9SrYg95h
eRfdG+qydZDHDe6CpgVpUDir8yqGTTmxNiB2wbFJ22BPMcH7Lmo9IeyRnHdddqYyrD06kQhuqTu+
2IRxz+soLOE8tpd5TPvMRbcg0uMVekJ3pyBfJHd38FVEfAca5xpS+mb9YNTVu5o1KhXMOutPBXDX
XcZh+kxULADs3aqFCPDl2VM+FOo+p5CIgOXy4+Q4vLn5bwR/wXYey94za1EWMoz8NBx66XB5iLAP
PbQ/+vlFnmpwNDWNkwwrI1zm4Vnf2z5FWf2eALc2vbbCtH4p2faOWpF72qxC9ncjE7LQvR+ZitHI
8C0n8+tuSTMSPyUclNAlc99o8nOj8TQA3pcExdn5fEjaej4xzsBEygILPmT3Ti9pLZlspScURomB
yDGEvNNxLakorqXvorLTLNgPqzuWgH0PMQhzN+R7Fh44XaB40B4UkrCkooNFzruf3YdjRvx4zPpZ
lXtHpogn9gWBif4mr4ZImhpIo1/X1ZvYIaeRcVAaZqkPTQDAA/lmicej+BrCN4ktwMjQcFlS5keY
uT6NFJbhQET4sCkRaUYUmPEb8NnMqhf5GGX161V1rBpz+BxTyqUB2Ly69MTqWAaRFoSk1RDNoNJZ
rOGqlWHTxhAhu9P3dNzf1MNOLizP+Bo3ANoVb2xtnux9tub1brYW9dqvM5AP4ZX0g8NNnZOqpowQ
d2WgCSMMv7P6uPcptBxim+6+S2c/vrCQjPb9B2VLP8aDM1hqYi8jjS3mL13c+9rMMXb7sAzx8Uyy
sz9eQU4EsJPBGytBPBdseu8SJT87ou63sCTUFbUhBoCUKaf/FExG6XuHZdMOmvOZMmPo+Sf1KNA0
YCYAk+UsVqzDRaZ6eJP6RHcxAoDNyzckQaPzTMggmYcVzmHsEPl1n31Hsj/bRlsFQ2z6LdSFNfMy
A8z0d08Gd8yHCPX8Pgz1wqjVupZy6gdUUQE+Abkc/6gbovVZdT4QF4BhajJ848nKJHTMxGRRAkrq
u4Gr0aIZ7QhhxH3y1RgNxDwHw3hygRRfLI2A0bAzKQQRHRK3txDLwlFQwu901s32GPC2BR/YSzb7
k5lgjT8H7UCU8HdvL5ACScR2rdLG7ED3ZHdKLKabK+2dnYUeYL4yyJugFPclHltIw8dZ8V9bRUbn
MY848iD1lY1RitMYylL4L6UIDoQgX8pUS8UcVNyGUUys+h5PSDTQo+wzzT6qf4dVyvSkQe73y9hr
tjJQB1NNcM2fVA2n/ro78iRKijHh9M46+8ZUe0dbt1MCenr9jsxbZJ5fcJWDqWMDhvDyr0fyhJL2
U7vftjbC52fFDJnp+6NOtZMag5LcLy+FHoxEDwBx/nDX5IIAJxnXlrb8ubu533UTEWkwDyVzG4QL
B/GIGAl1v435q6VwgfHIAU0qilJtP2hQkcCdwgA//gLQ6QA/mvUMaLY1sUhhhzUg75YoO3Fg8QOp
a7e9HJ9EFakf/8c8gkh6V/wX9e3u7hofJQyElq1071VLdfmg1yas5nzG59fLgJTNioiLiojqjiys
IruIRGiGymYKckVRTtv32w+6WMOe+5hk49xrIDSpj00c2OmW04l4PhiFz8Nir/z/DBCtAieTYIc7
0s0j9Ubr/M+rbo9atjw7ETcdWmPnm6XMuuN12UfXbYJ6E+dn/BUDJ3a5OA50q7IOd4A0JrG1I2wo
ZzHoXMdWI14ErfejkVRljxjWceqnsCBPON8aH8geH0yCjobGky+GfN4KURafEdZvWRy3DDHBb91p
YGSWP7aQlMvV8XDzPgBz6h606FG+ib9d8coRQcctr91zaIOkYn1X1NHkgxBb1J9GvJziLQCx0utl
1gbmnWYkF+8SPsNFvMGlX0bXhuthjmfTkKgR7Ig1fZi0cHON9hJKueUgJNPJhC4mcpq/gE8s1dCM
q97yfCr8kKQiMiYMfeY/boPhOYvEQzcLR8hPfix6bRTk5jtfXijNZ3VoRHSR5++H6jjfWjQopNZ7
PRuLEEu4eXiAam2yTfeHB5s7SlOvNLfoTTfxYak4IsxnwarGvY3zFW0F7KRdyNNObo7XEIL+ibSJ
AbjuTg9bSfz8T5yTYOvAl8QOBIXD72uMtJ1MdmJaaYuWar6AXUxal/hCSp8Ho/KUmx+nJyhFQ4VO
asidPPgIJWKWbvltPQohJnvu/58W/jJ5srpKg8OOb3NcB0xgmlwv4aVKYfA1EGtxnMw49XR9mt9M
1WQSy6ejCiCDsR92xlJsPA6MGAdam/VDfbkE4+4Na1OyJ8EGlkK8r4tNvTYWqmF4x4Pn3ERvc6XQ
8fnWDRHRF89HysmscjMwroXmvo4jXq/evH+rqNl30s4RbiAe7Icsd0R6d9saVEJogvSh+S0fg8+k
vF7y3Ro9dcO7XnlSksuxC2MiDtWpXG6yFycJPBN1l3KmtcetbX38rBW/GpAZYGbNuEJUNXncoxei
WnUZFUMI+CwXv1UbNZRfx668qQbK0PJWCQvzGueeFEUNCbWhC/s6cFGDaqAP1CCZMiau8XDq6hBs
7Two0hXuZuJSF/i0IbDMPlQRTJmWgSlCAUb7j3ZHS7zxfjzrZZ3Enmv4ul8imF/ZDcXwKHxONkb6
vXkFiFdx8e0Q2vR1mvKaXmRPBBbV6BPz0S+Hv5eUIDcwSfn1QBuINxU6Cb34yAYtU0s+Ly548KHO
VLFE8HuE2HNiNxw+7p8varNcI0B+fP5VPr305H/KaEg7uHZC/Pmp6jhaty6lFHYIMW0wLIIA+CLY
dEo7yw6gy2QBuvhb1AEHcnRvG5b2XG3WSjYXn4bVK71pDz+TzMKf2mToniuLBXfiFDWReW23LK20
67dfrVOp1SNNtOsq5kjQ5JxXs3p/uMCyQDFCPPZfV5oLM1s+iwBip/BJiv4jCJ4q2VRjKVauRfOu
tkyN6BfCKVORmTjQFmUYqcwMQSF/5dhGNap5KK+HIyKdAg0TcGySZ6OMOKwCprI2qtxb+BCSefqR
PdRPMAGYDTqNT6NJhaUfS7klHB3dvcSuFBWhDUyHrTC9tarI+yVJ0BIV9LYOXHNWrfquSU8IAkGL
1FrcLzX3/rxuxA9oawCH9JDI+oSrDaURoyTUWD+hrx48JY2gpxNNHfwhRrCrajQz122ypl0TTjTo
lpg7HAPPYtNASsDb37pM+Z16VoBSwykv+mXf3xafLg71Q9y7/E0HHJFRd3clgKg5qtVULj2xO2S2
4F+hSdCEboM2UaQKJDMIGnlOM7GquDhTPX6z32V5lDolLflTBY2pIchI/EWqfAb/Md2Ij/lF62pB
NAdni6zuSABN82m37UKaagvdMIRbmlD46GnWIcSSIGQ9OGQMgPq2uy6sMe3ajBx6flXgLooJFzjK
pA1ePfYW1z2ilg1+0rmH0o59fCRnif34Qif6fZDyvdVMLhIX470n3fFgYE7gmvLgu9asNoZ57AGK
guzAh4AcNtCmEp+bmhl6zDR8nBvTCLJDGlNOpxKJ2omFFkIZ4hmLc4QQn+NNyWDW7+4B3BUheY9q
YNqW2LAOLqIQELyfepz+xcT20z/3BgB+ado6iO9wz1bBSshVi3wMg6oG308TuZ05KCisJYyO/Dya
atPzFI69Dn9S6QLEIn4O3zVFgTsdrb2srFGPwR0JA6htrSQmtCycgTjpe5qgMGALRohUuzX6A09e
+0qPyVvzWK/+DyXf6QY5Yce+S9jzG+vV9ZGTynWuCQ756rU3R5AEx3J+rx/TZiouln7hTP2/Zabl
uK+NXtFlhgWQJCfmvl2AiyMZrP5VmSvx3x6R8DImHp8rpFPNzVCuznG5FDmFXmy792NgbtjqWyHc
1cq2p8ah9pIE0tjkCvydeHj3IvWmes5jH05Nleq+gZNJ0RNwV+TRsl+eR7ifqf+ZYBTNGKl1aFy/
FtcTIasI8U7CSzL21Aa81vJ8lbGvH1USfc2mDK1zspK4oP7h8SpuPUb1Wi7sv2bN8DQvevWpwLvy
kIoWMO6L4xKFOJhdSyCxfbYiBcRs7k7evH4FfGNlBHn4zhVpCJI1kcbl3epx5w4Ih3uMDi9LtKCg
FXYKa3N5/pgqHWmgFRchnr8wg1WSSgGsBuEOILIIUbYC2UyidoOHVcF8ByL5zDt0uYslp4bkJ1SE
NupB3EBKDFgJGeZTkBXY3LDyDBRH59J984oGNzq8c42wU2FVMBpaymzHzNCzx5o500/1ZUV00zw0
995Z9joBhdVaIdB4cJ1DTnSd8/Vk/KmgPcUgeKNhrT9BX+K77jByGtA8lyX8Qp2vXZcqbURiYPwb
wsUD2KYE98Yh6fW+ZirvTYqy1rBvooNITtkCt2220eHj3L/bNc1VPLNtRpVrpOHV+qg+jw/dCEH0
F55Gucm4OuQqMjfWFNNOer5XMazRrt8KDuEF4p5Yfa1iusLmckzuzcIpKPhE198OGK+zTle5fAUP
21jyjtd23IHSR1sC4B3Im5TtGcyxF8XSJRUBjfcJ9I21GhJknynLyHRzbLp+I5AwuZ6AOrzK48GI
nlMfOz5ioBjMpLtYjwHO1wWR2TJSZV4Kj0LJ8GXMUoXBxFlIlULd48EffRhVZuSfsXMSW7q8JYXa
0m2av9dA+KPqaBAUM5JYvfsOszHwOy6jevEnMtgGu8f2jR50GiiWzp6sqGolha1JGSkwiWFr7v+Z
rhXD7n8SSN2gbOh9zuCMiwcayPLLxdpQinZXJx/e0JjeMJY8+1DARkE0EbKulo2R56k9oWi2Mkqo
u36b+msvdBd5D/9qDREyKvohxPZwyDrIuNWy9NlgNSAW0KgJs4YIgXxWoMAbNWAkPmJjBjDPGjSO
9tmR2YNubQhT7cIWRnSW37mJawhamiOH9Ydyh+8VXZP2tKVOS0gVHir3xYceoU0lmem4HZKBw4k2
KH4ouYDB5cWZIvqLhozfyAfV+RyhgIT1QUIhYuR9dJCVGFIVGn7mveMl7vasCIDjxWmr8fXFDhly
g10B43LA57epbkYVu6AE8gPl0TTRXhEB2eKO4IGIEXEKX0lpBhWsIQy1pCQZZxNUmncprV1gAUiF
0ncFUJwbhRwsy63PwnknYXaAZBQEZY01YJgm2thZNCKqw16DcLZ8E5n33KSWBJ8+OZIgh8Tv6W0b
/Z65EvTnldciqhfcm+aFpbyDl0q/+WM6toJVcUoQ9baCUufjJ8cD8I7vMkjoIfMGSLuzZkcxMMkZ
KJcvMvs0fRPB6Tb/xt9LhNV+fiWbzmjnRtbHGtfnFyrcA+xbEe9c04rXB55+/BbzKHRMd8OHmfBI
Z7Dphlc8131Sl1WRuuvp0whx+JQMQufnwp4AgmXbngIjaa9ikELbPZLXBNVKf5X7Ug/EUiqU7mTw
HxV4z3KGj7+RNtYzYUwYL/Ue0wpVgAXJQAkqSFVXbe+NWgrfHRbu1ckq/lohdvOiXz5Lgdvlzz6K
TY+2SGYzTry8SavZU7dX70fDRdMSCmQL9eQpWKHkqZdjRjCXFqRbTiqZDkmt26FEUHdSS5YcZGMD
Lu9MN3IPW6j45wv16aC/Oj/tGeF0s8VvkiQ+hRyBF0g39ipMOy/vrT+2acvUiou/tPdHkHiCZgAZ
khctY5TH94Q7G1UKvmz49XrHQDeOdmuSdZ7XKEwHP2AY4GHbp21AB9SNvWi8ujFDY1YZoay5UQP9
F88XBbpLy2IhL34ySF3xcU8BvbZLGCZOtJNzF8JeHHdCs7G9dtxtwzA6bo6M+FO8f2IwisZWEGd6
0iWRn3/pNvIf14TV/YIoaAPP0voARjj5WVzjUsN8ZjOmo8EMp5c7nGIODoPArdwwxYk9X81PhCwA
0Q5DElrxz4gObYQcyLebN4jO8KzZ3YixhvsiS3JUrYeXT1FIxYOTDksAL9CrxHKrItTFrAdiyfI0
ehIQrG978Kj/lZLFdNs/D0+eWbHgElKWMC8lnbE4EM3GaglMP4+m1oiC9dVvp/EiOaPPm7B8YFaO
CTvUmO/meiMVqrHCMqUxY5v1u7NOp9mC5CSpncAgarNH9m5OU9do+PBwKy0qBlPjQbPtrPo/k7PR
x8ipOxg7Ly+5UDZLU0U52uzGndcYPVHfvp9K26QZBSMmz6RyCMzjLcGXqk40OpqX3YGomMRBOn2d
v0HE3gjZQOwZ6UvGcW7tPfCO/ZEMvtFaWYtThS4PKV5DNNvl3NJvZKPYJ6EzxUmGm7PFOuMoS2iR
rfF24cKuRVloiY2qxdDygIvGQU1werU9t3wW6S9LAR/Ae2RnkxJ/iKA0sMN3zUKGU7i2M+12/SW6
V1mDMh7wYbClwmea0vzL6rLDMvTY9kFKOC/wXTJ9FB0Eo4grRBfTCUoKfwibobD0OOifDoi1pmgM
XkG4hjPEXRbbPQ/wv1SKK8ItDPIP2O1fTEDhDL9/aHnon6U219ekn4cXk41KIQb8TCrryzUqnaVB
XwF2sSlaCIOw5WYctWjB+wiBTAE84KYeVJtFSDPJGRDZSsU+ON47bQ/yRnksAZE154a/NiTTH4rH
hu482Hq48Crv2mWSkjVGF3m5TMFoZsEWwttnH/avto34UjqMgBvyy2Lsn9zmSfvOwMdQqBkg081k
BaGZNJNRv1VVRgVyrCUNY8Km8URIx3KU7SCfqTy+///iE8djEW5gjT8Pf/Iqc3ppdtKbFQfudsdz
meRyCaTBzQqNHWRCwm9V1pbhzr8sHCyDbo6nGEmSRMQPD+xGGOkq/Yg/LC9RPRF5ImK1LiM1EDon
58JXMZPw0kErr5ABP8LObAf7HnZKrDNS2Me+R92FYjYxSMBE2D0D1ghfT93EwUuFqmkcW5hKIVqV
OLewgNYKn70lsf8Oy8NWoz3ORhEpk6JWoQd3+COX4/bz1ZxPlfbmhv+SikyYy8ZFrJC5zIw4hy/7
aoxsP78B3RabT2+gaZepiv+apW/c4lo0waX1AkVEjiviogaHz4we5HK9/ER5qUgaLHwqzJGvSxAI
CHnQoeFEJivUsPtZttLE4r/BQk4NO4YKbsTTZEAcinLLaJkhxBqUxE5T7bY8GVDzCMNLFbpkSAOV
WhzQ++G52LwXtBEoQhlE0PQKvrX1Lp7HjC0cOVBzsmlI5pWxrKSycSUbnmKbmwHQh6+MquY0bbpb
hZVWutJlhWzyVSPFHAMGiyUTXjg4HgLwheQTPT6O0V8jphLTx79zCzAn0Sem+a2S5w45br+bKPCb
zgRE+fqoepIJgQ/qvU8qWCOm8H+93Ag7GRHIcHvIB+wQyzmtpiRI0jYXcuX+mYOQnL7MgxuGjpoa
lEF0Ohl0oU4ugI4vdM3AdIE4aK4jRufvIO+mH5+FkiVJZkjF+eURDrIrYzt5OJi/gPBoUUwUgzfD
a9tp0EJj7J3/sim9VLnmk4cOz3eeSfbBKF+XztsxbFytdDpA9QqV87v04+HUlC7cGhjRwFQK0/X6
G/v38er6dnDUT8eXfMU9OF85j5euhMUmVJarLcGDQnhviJXy/15hR8ShDfGLLKrYSm04jAGJQD3r
EcZPe7LKDwFs8VnHvH3Ho5yOrwY7HoLTdbZ/erlJ6W1HM3FxRKiLO1SH1qMIEqr+NSvqs1G8aFIb
hhNlpZWHP7n9IpBhyDTM9FL7fVXh0+JsxSOIK0SeoEN4GlwZKIK59TyI+XElDLTTmOVeUt5LfU7R
6Ux74Al25aqPhkU7oglRKdILBCHdu5tSPPqhTxRULNKr6sYfvPt6U//aZI1lXYPfa5ToBlaQgln+
Mi+DinrwhnZO5jMsBHxKw1iNGAimm/oFMC+w/xPxNqxovibRupqXqW/4lapoccR1m7ZNpsO0JLSY
S2zXLgfInqhfX98+Q/eB2oeqsaYw2daOQu7wChMtWja4XU9in479OB9cGo4+HD9qG61rNhjtLVD3
SRT0mO8BwVqWKdFFCSqesyUG43U/GxSGAxGYg7NzSZvqtVWWQRCIMbsu2kGZmff/9fDsJ9NbWMIL
BIn47cbdJ5VFOEvVK0oeqhem7SHQcsYhDNKyqIv11pcaOaInPjgeqw9owpV4OlIYv5A/lwnA8Jq8
yP1Hco+tFNZnKAJ86+6vKZtTOHp65t14Jl4tBSAOJ5eP9AWKoG+TTaFLH9+pHRPtPhML5cqoufnv
i/zBJiXrKDKQkqL5Sn36q1vZk+76GLGPMgfy78CUYrK9Dhro8ev2NeJroJwyBfV4UbaLH5aon6CU
0L0erTpQzkJ6P7tll8+hrIKMf+pAZv2ZPuHDtX7bDBTRHmE2hRCqv5fcfbwbf/CcXtyNSYNlmTCD
hOZy9Zmg961I1ItzK0wv2cODQ9KZi0o1W23f3v8L9/dUwxvUAbSqNDA6DgI2pRyeh+IEfbmcmPxo
6deHPqAfHgoqM66GgQF+ofI/MgW2YmkzgrY3eQIluwr9CRCWVS+dV7VTIXEUhVz5Okml8heK0WQP
lwJeplnJMc6ePf9WN4e9xO9ZUfyiGKWU/hUN4pjxrg8M2vneMuwF7BlL7GsTmWHn+pzQL6YuXRQV
e04v20nFVh0457OIS1JTeMUtvqmzatY9vEdwENDMq7JtxRekouA0lmBPP0iTDM49WTF3HLXsL2JJ
eGJl1H0w6Q+s9RAW6XBOquqxr/J+RwTVnj/KpdOLZPgm3g5V8aZyIP8sFVcLd5fgZK4byvZ6ZCL/
+1lJzx9ecYGUU2y+UpipiFBF7dAexKcI7LQLdDFN9UxAZj4H5sIEzZlOwiw3YsT0hrNKcD3XX1Kp
4MHosPM3BbFplZ3cH/7KpKUNqHVWTEweLaHW2PuNTTdzk03T5EZ/OfPKoVCBm+PleUWdLSFOIl9Q
dbyiDGYMWnlvu7Qbwn06qbhwYK3Qq3WUydWwwaeBY5H40A8wpXON1W63X8ZNy/KFV/cYwsSwugey
eYWXEQZ/CWYlQyXaG/bZK1S3zFRippk/Itsrh0fe2tQNGeFkn5mViam+nU9IMsWMjy7eTHKNZOyU
MOcVDmCUvjpuqia0BaXqLJn4kzYYfN7MIKbxcVj+zFS7+WwqFCAE8V7crzW0ieou2VF60EZTxIDZ
CJncxByLSgW0oH465TNXuWjZRqUnwhu8LFb2ehambtcFRnDqX8uWf+ez4V86D8FOrfaDbWNyq2Hk
bW1Q99HnpKgFe3vBdep7GX4ddA9bTnox70cKqiqM44eikMd2T1UDsEJ9H+CitkpvfB/wia+D69BS
MQ1CciPcwbrrglrf/XpVdjISvtZH4QKfVyfWlhOQxqvvvj2NR5+KHzvoZDNoLvIoUQGkSlF5uN5+
VReRKw8r3QKiGzeRu2HK1W9FzN1BDxPIB4tSF1haaWJf34OjZd3m2rpgT0PaZPSDW6RNMnxSXHiz
6Ai9p0P22aSxydeUxviCEDAgaJgyOTiz5BD5AK5ygXVnYLghPuiIvZqFae4pLhWvrHzUI+Tg5bUT
+eQnUS7llS9cbY8JgpSstNUvWXXbf4ZgJbrYc74Vg8MSb1EQejwBWMYpkamqG58TfT8V/U4/k42D
cWeLNBBCyZvyoOWHbTK04hmM+ZqMQth0y9HY6lSm+J/IuMX4MA1Gs3ZbAIN3qFLOA+f+XZvZsIW2
7T0gmtxidIVSEpHFgyO4LyfPlHye9j2Mj8xuxfLsnLJA2CHMB44ui3VhdvIu/bIp/RerAoJWHzgq
ueIf5sp6rSl5Sc/yBHxEJRYlDdhUMQuQ2aSM6UaAPuCBcnxvNcxbF0rv0NZwyziEnls2AQzEpBmE
0rSCfHYnDu7nyRLY/5k/77jPWnMLR13CrPFbZHW4xmfB/xy9TDgHMYZ2L4tSUVKN9a/dhOMOiU9y
7nN9KTD/JHQIFtqItPW0k8gJQ+ACOGfaw37b3WWb4bhRU5ymJv9FHmAoAnC6vymYyGyvAwYJhhcF
mrLnWNpa8M6T+JKggK+vhvzCpA5iRdmBkzWCYlZwhUJEst4BMQ0+j8cY0kKQDCtbMYkYC43CKX15
5S/Lajvt8u4Ebe70gvgN3IxlBjnKHWFz+eTCuRKfZkDJ+mc3KmW6cdRt36SCNi3YUV2KWk7sOHRb
flbYH2UDk00bXzAM4BkTmiZeAZu3LZw4ePA2KMDC2H7jiFZKh5WOoT2Sfxkuw2I5eiH6SZIvBQWF
rYGRI0zh9lR4AjTn4fkfG0MJum1ZW05xlWn4EaxycfCXCYqAy8wh8diJDkXiYjhq/wgJ216P4Vg0
fw30OKqvdL9dkA0Q3d4siUXlNUJlqPZ/cS8bEiNsPkaF4kF3fany80axB0MczsE5X4jL5l8zWB3q
D/HfQendFIdjN1Pdn3mAvAU424PFUaDi0lbL837t/9QdWl/uv7d55aKL4SXgYQ2Sl1g6XRZvDpcs
BX/FTUYwxEgtGPo+uQbJNhF53Fey0Kpr7UY0zsA1PEHkjy/Y1DUxBD5/Jle+Nwcblti9n+Savuz6
TdNpjf3AKUvKlQOefhVPllz+xQXrOPh9lwng0NpcRG5W9kKwS0dYHjfnsKdTy5PedmO+0d35mRNV
dWGb/MXOcSPS4g4ttOLLE7oxYTkrD+SwRFIDJxcvwBCcw2PevO9c5s3VAEvvfLf/wjRSQLRrE2XD
/sWDSwDNBafzUudU6BuffAQ3fuqYOJF986alu2BwM8sqVMFVK49iMC8GiM9XdOKC6+O4o5m66mf0
vaPOF59QEtPe4x59mYRZW1+1cZu1wT+XmTNzLu+EA7p+OC/gz74zQIyHdaX5V7c1KNP3BbFe3qhy
YHpkCMfD4c4ajhB7nRNMWGoQQKTF/LAo8ii/kWnoc/aL4DVyzHMvmz1psnjiaQBarLf7UeY4m5Ak
vPUVqf9d4998ODbV0t1nJQwEeJy5CeI6WfVEKN1sT1p/hamzjg2VvO37ukhKwN4VR6SV7KLaLcXE
w4kI83KL24+HJWzzo/vNDygsr+MzayGdU0gPnxYZtTNR7ZDU+QgpC/myNo+JECYzpvioo7CBDbtx
68SWw7W5skHZWvI+A/vHhiRkZfidhb+i/bH/ppA533dMV3C4cBefd3/RHC/ozTkUXz5Ak4zoJJ36
KWatAveestpoblBfRYJqjSoD/7nRRFg5WzFjclbdyLBjPh1qnFNelJFANw9YMKJ1JFvjOLp9V4zk
uviEV3G5HMA5vT0le9D1t4L355tUn2q1+pVWqc7cRakCKoyw3AUiSWzh5Gtf7RDX+OROhENtsnUj
KoRGw2OtsGXspelklYKXQkEOi9nDxuHNuAR8tX39ZMyqlKsp1TB8gWMRPmyam3e8h2YsaUAic5K+
MZ8gttPNDk+/9gmFjrUzXiI8P0T+3Jx1jGFhuKxNVc8PoEtNlcxH7VxKYELs4DD1KYXNkPWDA+VS
8XLMVmg524Yw1mMgpNx4y+z7NQJHLaZxvY/u2IiDEwqN4QYmD4zwqn+c3wh7SQwv3C3o8EA3s8uc
ONemjc1aInrzw2uhO0I/sKDiKhSwMS4XsnWyR3FiOc9HkEJsXNxOON0U8agZiYSPeIWDN+BvtYz5
pdp3tFFL/XAli8RsTuJ8r2GxI08ruuErb1CLz4CaPfVQVgxLB5P+Ywx5iKSiwyKNSIc+AGfGJ1Ob
BpI2kcSGXsR5n0m7AxuglrEwppyPtQLjlDLLVKu2XA6v1gEcSoDFvVD1vWGpzXgTnVypJcodKWQ6
hX+17VZADp5GDlG0NbGu2thKigJOQIcSCyB8lMNYPmZO/cnkYTeti4QZ9E/vsv7sFXpylZgPa4yQ
Nlpb0Ds1OBQ4nuTsEm8Ft1sGULFPGpAma9M8nVy1wgeN+SZ3zvsAassm/7EZce1QQJ3WKGRzZH16
ubT25Him0xg+aseCdioko7/p57ToskYkcy83O9Ab2xSD74WvszRmrf6O734nCk+zZa9TlmwkoZqO
95yPeyZDNCmFrPuamjQFpxrSAg0NIVfPJq0uxAaKD3nvLesoxmyzOm+XFVaAVHV9eU6l2B2nLPVp
qlz/89YHR+gSWi56PPwU5OZ69w1YDpfgoqv1GMpPcBM1jF+lmcUtP5wohCrcPPMBWTo0XOglE0W8
qeFoEq4FeB8Fxx/QbbV2i6EEWJTcO8sciCnSbkUKqNguhOZrvT3xvXx3F9fcpHAG85IDfXdxDAYq
U3MsldhtRzQ2JXRGn2gWvCr6Ce0iVzmtyfl+xh1IKqBh0WcRMA3yO4UMTotN20yEoNES4yTZG5Vb
Fqb/B0jF8auh91phzyieZuBe84TzvjaXGMtQDwoknqfh5axQNYEw+Tpt6p51FT08f9lAb69UMlBK
4CHES7EHaLylUkCY2I4WA6TExjpugpWFSzsSywZTO+2z3c+MGu/moiSkLbduYE6UYcREMrR4d35/
O6y4bY7NMZiuUIKOQI41eNapWsuPgZ6k3HPMOA9V2sfSQ5Of/MubfoVB4DgM+RtpIXGqiNHbxD2F
o7c7uFe9OgOI7qC+dEdzl3fLBOui2vh55Ozso9Z92RaRLhzrwYsCV7yCXfStG4PVppE1lSOpCtJ+
ZmUTDFOnNM/9tdShu12pKjgo96HiRtnxTvTlKQZ7lD93y5MeHbw04os5V5awjcD939bPv0AnXAJ3
THJqAIOYgkBL/ma6vIfhH9a6V1wRWVhwnpzlG97wTB/ryjN7RdtQYM5oGOEt3VXsi9zv5gYMhMEa
wDBFVX5Zgr+IWXm+V6Cr7cAJ3lwvJ97ydPqnZ5BBjn4pD0/6oQ6AYHvHC85KjHg3shgzKe/eN/mS
oAmt+1a/pCrwoR6XcAd11hhKVomhlRpex+oL3qKxUuCGd6PmpmhH9WbdvwBCItNeMV23uFe78jiG
IaGIHAFeTbgwIRIHugkmLZ/UanoKui32jKKnDOLEAwq6TPlCEh1O0N4lJqygfGjwOSZa8nZfgqac
X/11zmKOrGuVBRG1/FEUE9lm7C/k5uyjp+RYCrwsOhsP4c3QklwBCrboH8l5r+FITjsEcQPlXn/w
OfjorVrh6yEb4BzHmoQ6DG6RDtPgknp7BEl66DpzsESkFNYdpG855oRwWbvCz1R40fd0pAOEuCrd
BG9uHDhGlfFuPxFOQbyxZ+qDJkQCoq77NsMk9zzDdOKCJ437MjHhmv+NK1AecokMXOIB7fHj20NL
sA3EHM/myFqTKP9GvikAdK9j9O5KI36O8ISA4mmFyJ9qGWV9vmL5A9/8mttfDUlYsyR3trretcZ5
sLxH0HlWSiDUbriW6lymlLklO8npVnqwYiPae2IGyIOY2Cfn/2cHCdhSbmsz/T3RWub7hS0arSQd
ohy9d/0Sl5fl7ruCa59O2iSMi7Ee2Pz1VHuxtAVy8b623Vo2/0Kq4YCTJ9w1PbZpGjg+9dzTCHf5
X9WuL4UT1gJW1jHeGFeuv2Ozu3FbHKFDbljtZL5tQdMNTnh7CbOt+uDsvK92BOg+ZvmD3CFcyRzo
gNJy8nWiaXeGQH4Zjk8cFgR8E0c2IzBKIk0pkwGHNpjLcu9CMJOQK+hA2/L5E9Rk3tok110vZj0Q
aeahPSSbhBCEd9JL2ut13Dxu4u+lxqoU/CZergdHWMmfnvulY9C2c0c74B1BPd7T/fdfurlmbRDa
oUG8bokoNSHFs5cR6iqYn1PYqqQLfUjwvPqFu6pVZhEDiAk2AacqsUunwvenl3UOOYZFl8CNjCxz
8XDpZnCZjpxGa371gtXNC98DGqlhFLK7SVB1bp6rGdowtmRDjtMM0Zh4SwsHxmdiDn3pYdhix95F
0zY6cUHEbtg4MjxZ17E5FhiutRxA+Su2b2M50Hu/kvHxSGxU5XoE2Rh3TIyNFcD5txGNqmvMTLw6
Ngzgc2xoETa3bZB/IXprJ7zwuJlWOvzyyTtTmJAuZ7spCAb/bBArEDmiLPgC2HLebd74k+rR6Yq9
IUxxYCYJgfDFOrYNLVy4J/FZFL1QUP2M7nqf/rSxE3M8xTZkM+tC1513/Fd4lwVOEObmcixkvsxc
meZIsfH8N7x8WBjWdRru5fQCp5YcOgN494jM9uMtuoEB5Qnz/R6Ht7XxjPfxPsD01gZCZKz7UFgc
LAnwDFWK9hdqcTQ7yCxI1HNTC3Mgae045J5izj5JOrO6d6aPl9eDeG/+UW26nZYyKjaC9+GtksbY
Yqyl+/9M4KbxD4t1yuHg7U5uMj1IOnqGOOZeJ3kE7SwQGUGV7n5wffeZNmid4i9iy+387pxqFlA/
rtOtgcT9HaCTo48lE5+ga6JgIKtznx4URwePa9u4XCnhIIF9N67RQL1Hj5oK8bU1864YcVwHimJv
5nEUxglu7ySE3PNs8+eczt5iL5DVzgPjx4Rv/KMZVoUSKDl1mYG0Q67HZXr8o6GFR3lCY66tKLae
bhqJxGNemxM7zbbw29WQxVGNCSOFG3tY/zEM+9XTg+ykuWMLfuBslYy+07FuH4ALF7oKF2wCjZmQ
DF9WSp4O+bksyxLo/twyUYz9xIA3knA3R7Y2hAv2I5wMYuFVJKA3tZtRXv97p1Dv4aUfK1XbND5b
2TU++wG+/h9VamDLYKKknngbUBkh8tVSQ0zc3XYc80Wj5AN+7k1zdGxC2HYLjsQGXoTRCFxR+sh5
7gJJI3+A+aHxSfKG9i/DYyA01U5PV4A6MJ5Rsg+mBWd7ivyih/bxwBhZrYvxlN+l3uJv5xxF8gWU
t9dMOpgWyGv3FGdumqgukVAo/v6s5hFCMdND5DnzY+OLws4IAQ3mZYeG3w1U6pmBeNwqI+ky5sav
I5S3/wfeEPFq2vSnF8XyNiZK6nYH7pkCxEu62elz0/7BnUF64qbEN5DwUySuLIiXm/Jnqpyk1/o0
t1aoIVDlqp9WKWUu7fzi0qb+CSaThi71q24XBTH/KWGkBRSCX8xFBpVBjJBvPhNUqQhnq2v0wtiO
iW5ObgG84fgeZvRXCuwzfx/yy8elkzyDRqd1wZLvjQmQ5LIsiGnP8sX1vkX32q74nMfR8DGjmINS
nveYtYql+jDJqR79LyiC6ZlIwv7Q49U3byho+sMymckxU1116oAHnDfjrjj8Z6RFtrwpODt5n/L0
ADFX2SatXEklIEYsPo2p8SF+X4k65pTnO9Y5a34d7EyV0GeIv2RUqwaToZuxkKnNzGsY0MKc2vrt
v4WXaFJlxx9zEPZPYhq7IzuOlEfRWsJTT2AdombPOb0OcAlEfdWFFrciyhsgwg8JetlzvX71ZKmf
+y9BfmbVChoAE3+MVSCAkJdHY79LDRHF/XftNi631tFWqfVH80Qb0SIy/I5Q0tEtvwXi97c8tKeN
axgn2LP7OGEoLK55iT/RFhnp046B6eMtcdf3sfS7e7w26DM9MHffQ2X0a/JcSx94hOXaX2EDAHQL
33HP+NYm/oSRMFKW41e/wZAm6J3NpveWZLkye9dL/imf9ngMR1wL93CSbqMGn2bUZUhSoLxw3Its
Y3wNc7oZT1H8g6phF/4OgyoQI3NauJEGkifb9rRHIE52wzW2knGe4Dlixm2pekDP/ZFRMmKmDyAX
XFRF2MLIeqk1Z903s8+k42bdyNQqDJKi9133JL5FDbEuw4zdvVqOtjLP5D1WvjbJ7zU/7f6WCpq3
jnzg6MzFRIQSIdsT22q6+1Bb3IrFGK42g8Nr9Wt9+Ec2x+cvZHhtpv8nlXuCrNDL2ERCoIshYqhj
fnoHawTzvTxKn/Y77K8XPgNsqKb4Y0IGdzXFuePLiA+Lxziwirr5D/w2G5h14GLA/Ve+2tGcxsn8
6hjpIL56xFj2H/Csy7g1kAESsJKo/2IO7xzCXNXfouFe3vQYyhyysOMU4jEqeq29fqEM5BL6iEhQ
K2rVTJjOjA342DM8VAglJaw5A533xKtIs21VC2MU2KBwKszVKVBFT0sttXiAiazDDOlDOVjJm2SZ
6xOES4za76HmcxYop4qPTnar6YG1XOHhPOBS7swXpkmZrd2nQ/e6kfHj0BXCmZvxQxlChZMDr0r5
qRz/h3fnC6Rs4qf9fuaHsqd4RD2+lTEJLpNbeiS9FAt6lkCJXAor21nLDbEyjWoMW9+MY4cg1d8M
oKq9Gq2vsScwtzGoSK8htUSulrQLgv8IJN+eFnT/6SZFIRyt51ouzxum2o7z2TOG8lWuz84TvAEb
RyhPt9BponTmVm87NNzz/F+RYBVvPqniie+Ug3nSO7uboeF90BS5V0SVveVyObnY0e7wDrJ87iCp
12ZdePf37LXJAONNGQIP1jye4AxUslxA9hhZd2RUlFIpAM7cMseGcMHi+U/291+PUmJvgGGIfIOr
LHbQ7umpFDR79EhLs/y4YmqTPEA9JTpUblTU7HAgE8H9PC6nb+Jox2+1VUi6y30kgDTBfC0ZKoZ1
17HhL0S6B3ZJhoCL6z8Net1HbYAEm/FUp6GB5SedJW9uqlSOF7KSZnbgJJUdPSrTpRCsRRjvz/ft
uQjbTenH180zoON1jqIK7X3ieu9z78gYWr+h0QEEGw01X1sUQDu0u+tLaBHSeZ3s5EpZGDZu4qEW
zDSm9dtDqnfulGMuuLtIdC+bOubowSsHGoxINnVnV0oktsB6Q086IiBn2TMhxXenzAQwD/FgsCsm
nGZfeI8nc96LW+yXuIMbiTQG
`protect end_protected
