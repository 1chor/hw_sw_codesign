-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
JJbjxg8xyYS3Z+FG7uMsZs9DmNZAmmb5iwOMKS4rYETv/3W3ZEFnRC14dZ6oFfxR
Z2HCVh+jNRkFXX97oLn5RqHOjJh6DyVSxhbjL7OBWRoWTvT/g/bHTxPu2JZnReFE
2WJy/4LSrdwbVTyyTVaejw7x57VqoKk3tJCIQMhORyM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8352)
`protect data_block
JgCQccAWZmai/CFTjtavq2iSN2HmBe7DdZOqEjJMwQP7BN37ZKd62cNZk1LX2Ck/
mNRBzmm5cVLxjsaGoFF0c80iPA1RA9mAMhHI4C7PISXYNxj1qjUofFkzyriYOS8l
aGyMVPbLobuYl8HuAo6a9+1VpnFrnJStd662sHYsNMqNnaAev7ClFZOc+7szFFDp
H0AR499GDoo/yaGa8uZR8w7rEzRv2ZXk8Pktmd80kb28/BQ+oKAsSmnB/8Xfydpf
ANNvn0NTqfzPY2WEI0Wvji1p1qj6YU8NlWFjH94rWRhoFoZoZpW1KJFGnrQTBCkF
qgsiqKQ5OQfHLNXePfyaKjz11EpkU5RHQRxeuvNIrWx2qUuKuJqsFCwsphgfeBtr
e/n/7yZBYp9rLaN7CU+DVAqihd1Jhfd76id63ofENkY/xi0h6qWsz57R5wHi4s1i
bnMSv7N0sakRpBIHEpWggCZmOLFupZ/3JuTg7i7tLiaqbFn7bmDOqwsxb1wvOe8v
WXIRmGoHlOFU9qAXVak+F7ax6MMCDPJWHPRo/2UXPL7dO0d2VWsWGW3HSFHfqKb+
OPtTBeJzvhadit1Tr0H0M6X+4usXi/PxMl/fDDlT6FJ3SyPmFVTaGLomQFeSqjBL
fNN8TUI9eaIPHFlU6j3MrMcPIm7fzxaO2xDtkTKubZPhqrURd8Og4Fkm804/Wsns
JjIR7JHddrSvDQgSGFzxkAqCt6ZEIiQmKD6a/f9xtaRDBFpHQD80w2uNbqJeqZyd
By27PEtmpTfWC+myq54Mh+lh6isjFsipIGy7kZ+oI8fOXLmlZohqZ8dUU5gvRJzY
P0uynymT9xi10fMX2hLRvSohPIAipKA3KyrnVF5gltPOCipN0OXRDJQ8GXVyTv2E
lIUkB0BrJg8Nvy3L4mRDSJILq9xbayf401Qe12GeKEZV5mWvSZMuUHISKnfsQMiv
9TLU9H9/qFgjiJMHycS4dfvyr6JpnqoV7SrpgvWD5dVy6V+JWePt20PYuZVE/ux2
hEDq9m4DwcYkx0PkHK/l7GFPG9lSTRFOmmGd7YiZZObR9XTKvcw2/+P+kXnmZlta
qI/fqvCEPSo5Io3r1NuScAwQkLqdjriQrQNAaj6TknhSlBPTMY25tIYFDiaCt9q0
/3hxRBDp0/hpf80+H+/XKX2GW9dqfnygoov4LxDhtns750WzYJCcMlHIqgfkefBu
viyvAROuNofwcE2++pxH2HfdS3GoWjZxDbuaARhQLFL1MQ9ngd6s0CXDCgyEEyKf
6UL3wFzfIM9RF+7SvIE6MFEoRU0iRmXXrWlDqjONQl91e3lIYVP/vJz34C+XC7im
O8wQsykLCKjIKQf82QmAiCaEVdWLMPMfafCMAX5l+23m14+Iqeu92GiuZUbkPQuD
PUS4qbHzPrHkqmiy+43JLZMP2oAF1RMUNLC8n7oiG8/XTMDE010qEkF9TU0pdfq3
TRLLbZRWilNtl8SQRAOciqaSeMNSjAKt6/cTDVnrbaqNim8gmaWXNxBQ2ZFiSVaD
DCMXvee8hvfZbiStmq7FlxL8An7+LRc8fNlt85lRUVPQW+TKcyTQhpICC8VFbQAa
qQ4pcDOEiVA7x9Sz+d0drh1PWw2s3TuJYG61wr7t/kGPGUHoGpXGLT3g/5farTGy
PK1Mq6kJYw+0K2puG+3G4aedAncuODgwN+Gt5WnWb9J2pI9rBVH2n7cGJOinXfz4
+T5IpuxhaqCzm27XGZRwIaedV5m3wPI2m1iORo7QI1NGVxt9ZnZ/etk/GnGOpJyS
7WRu+Namm4B2bDM+8ZzAT6QpR5MNejbMm3pCmUAcex3iqNzuyRi0p/7rZnCAC0Fm
dhM3JmuBvIknlnCiM6wN5GYB3aXtphs1F0O0ttOAA6uf1qDSxyxKFsyqmSQ3Ggv9
pCw+A+BiflqG4sIaK8GxnlH8cy4on5vlRaFZO8qAfFORdh9roEqfSpB/exS//4sc
VEptQKCy8tElj5xykzkk3q5XzrxnCAPzv5M+7REnaOm/HB3KgrbMwhQumOmPEqhy
79jpMAXCuHO4GCN8ynxXRrRlevjA98lhuzJCoGO+hiLuJvB+uJMEiHORsRpe1alB
IokzDGwqHg/fXEnzxENgmET4rvHEyjtqQd6BDgTfYB96mKOMEHGA3sLAC78C/Mxm
60o7Or1rEaWc6+ZcRNAZkA568p/P1sgTSM77SATCmk8ICEKIllHn2hd/H9ngBdSQ
BhyrJgu7nhJZX4AiLAv6wxPWqFJ56IQaLAXpvw4j1KG3e0W+VRuoXoPbrUhuh3CU
HCQrprruOw2AGWc5LBsoSltt4wpXhI2fGqzIzG8yk3pVrM+3TlaklChGwbKijgae
/UU7LGxxKtC1HGdQvOij6sRzBUzFVdDCPsBZuA/IU81t++djSMejso23oMfa/pL7
imq3XtP1w5Wf2MkRCMwTiY88/0vu3xxMQBscsqSETbANgXqh9dcWd8PkNrzBv+ln
TjX8vusrUTUOB9M9ZImhLuDedcAQ3pdj1cab9SED4KJvMgK9goQPlVuBAr13zkoI
t4q1OL4pONqcrOv7GqR2zhhO5Q1FCXOX+XF5S3e3ASVVwrND0XVcg0cntJoTfuU+
o2rMUpUmnvsBBmTV23FLPvoOHMBMuXwg3HZz2R1ekgrje8NJz3oPNCj6vrkjZZl3
pL17sRQ9XUj+UiTq7ws7uprQ/bziRFXxxsMNfhlQRHXaLvrZvMNn2xEfQhOdC0J+
0KTELaTsY4L4ylHCKPf4PAPJg04A6LBuVz3+tc/4UEqmwX9juQ/IWi1HOermcQnD
d6Ol9e0muiWNqmbdGszvjB862g0sBkPGUEH1KvN768jOCRFc2x2D17KBhnmbOycz
r5fVy+kPRUlHuC1T/cFTRKiKPSU96BL/lflqNKczU1pvXRU7pD1Uynm9ZCXGrDLq
4K9+HlNNAZklicq4BScA0fdn1yQT1lD+EuTMSiHkY2TyuPAfcqM9uAVhd+vstfXi
sbGUviChaZRsKzVTPzmS2cr3IkFwdf6Gw8p/Rpe/orQPbKsjIrNYkc7DxEzmxdwQ
iqQTngOekKfv1BLlvKTiy1Evpm25/CKxKtJfryNZ2yfdJKYiymWEcdoWrNe9Lgrb
UGp+tgxkejsmiavqcaJqKTaasj+L5L5QsYGQ7NGQjtd0HBr9NBqBDgisGgzvSsPI
wj2AIej4nu7GfknTBM1SH+PtBpUnKAdU070K62vAVORGS7wVA2MiCjpiGWrunNfE
qnsgcLDEsilhiAme8/0K0GNN+NRm+eCnTqgiSYwtyntY/Pm3HxKHly60wNjFRbRg
g+DMC2l7GgCVOa33a12awcoGj2ve9qgCv5PjGN+pGToLIBaHhAXf+XEmCatmw+Bg
jNprYO4aVH7WdRLv5m3L+NMZBJvfyFu6Mc1IZfsjjuo6c1DPdiWd9nXhfwI6bTd9
R8CxcOrWDm7IQD8yLSRPWxluyrw2hgx8+XYXHdy+2JOeU6K3q0vs8dulDrpfmnc0
YndorJJDx4a7SZNktPG8lU6PeaIlthPArU7cGT+iV8emEyAdSraCXzJfW8X4FQWa
Rlzsg+c4Dc/ICvBPCqXJeP9oCTq/Jx+pRa7PSB8cPwmN3BzkiMVuZmnKn4TtZY8d
uif5U/BHaWTY5KOKjObvyCmvRFvE5kjOWtERYxQ+fphxhFxm7MOP47QXof39s9ii
S1tjC/CtLlC6Z9uPoxm0Qh6EA98yR2c0Fmv2Q1bQrYmUJsKQ2MNFAD269TfU4Aie
sPcFcoMsvUok1A0ulTW4HXaiVRE6/0lP4fhDKE1kZaKpTa0RG5DsPfzoqfNwz0JL
MbNZ9rSCp/ta89w1cB5NXn3WFvb4t+t5VnCFtMhTpuJKxLZtuHuOvD9YniJ4BK0F
qBfQ0TSbiWFlVGfCnuzCMZ/yRNDNBu8YXwvRpdMhRyKWnLnFje4Etjllelc6X9Gy
IndAbLt5jntxPZtSuoDXyb1spajidacXf2te9Ao/nOa8tKiVXZFgVBxYLuRo3QQ5
kjP45r8NAwvCm03n1S1ymPEg6Dj2KJSYcYkjzocSJqJlVYbYVBfM1RgCv7Ifhyy3
c2YZvT41LfDR1zmaGzuYJPAm1YUAihMd2RRcfeJ/RPyDZUFShd7xhu/CKNME8K0L
lndqrx/auS7RRLxqJhdjVpJOgz9EoEPYdsTeHRVmqroudIAeHNFAS6wbO8hKeqgB
7fxBo1FCQgy8nxNpRq3Gj7qnjfDdaw1yDM1SjLo7fh6GyjK+stNSd5erhZNGJOuo
Ctz6oBydEcbyIwIN+VcFB4cu6N2CvMFVX91/NWdtnMT6LNLKAixmThMYS+idB/Nf
NGG7S39/Ut5pn/LO6ACyOnfZXPU+3hhmc0aiaQxDYxBjY+s5JNh9LJpnAnBELbwc
wpAEUoqVqyfYn7nx7x2Gv09eWmljOAn6qZF9nNXuKcHRxRtNqM8rMDk+TKfuVGC6
BnGyV2AVb8JK5nXOrmXvOa7kyCQN/Usd1TojtQGVh/yLTBiGL6U7X0CJK23QPX9d
9TUXjGqq/v1Z55CUqq8nCxj7z1rlyzLulraNfa8YPUcFpx6PppkCtLwYtMsQUmxp
Eafw7brwDtPGpDHhhaUvfanFOnjnFHHGksJT5UQWfD5SE+BehP9StyyjP+sqtqe6
sNAV4mdAEsHj99pepKGJV9Ul+wBzYaUneeGbiQ+Sn7tm9h/b8z16Og+02wPLI+ZJ
MRMK8IrWWSejVP4NGc7lqeHQLhzgkSqXHaaIxUwm5phGc2WuZ5HW8BuleVcybeG2
ofBlAWJaKZ+B1ucUvkAb5agjLbllE7NG9AGqksTkp1u8sZNbtJKKMX9KZrfiMNmd
lqmVlsKvRTlvY7QgZ5X/tUwRv4KMssDW1vAwOMB8kOi1lousr+IsaudxjivC6ri7
aTAsWSqrXJn7KCmN7r0gsw8+XLumI51HDk1pfogL0NahPNu1P7fCTPAM4hzftMNB
BxEhZid04lTw+J9ib3jIjlg3TpJjW6V1ZmECz8sPQI/gyLQ+PqVeOLNxEGB88wmh
bJxQZkQMA2cVAZnLhqjWc2FOnHIsHk+l8Z4wBk1h7vcy4b2UHj4wzsg92CeBD5PI
4n4ADQhYjq34QCypidlw0N/C6Tyxv7qKWM1nrl1xyfuBqYFDJ/oP2FdP4xKvwsjD
FD3DcjbTSqvBtUznvrPZpY82MGVA5WF+dO5T4SovJj4oQt3WOLFxWoXHd0yiIGiC
UWT21c0Ezrwc6VVXJ06cpWcTrRftYa4P6MeZi34pvnABSgGn+qN0QRM3FTVG88lq
cdfFpIxcqA3eOnnZuicTrl72Hp6+kovmWtwDTgrDQD/s6Udi2CK6evxtkD1rFczO
NtAgMYykogAzsmKpdPmfH++n376t6wqicGPhPEwgUxew83nCnrzLLrrFZHphYupN
N19Drt531Pk1SVU6g8o2jXB1IaTK44Hyi6iNysBm+aZEPyIJvFO/ngSfufeIaCk8
Ev0GFucSzdXDmjCGtb1BZ4Z5pCX55jBUyxsjjksaNXWynZQ3vB+ZtHdDECeM7abN
B764Z1EKOhup0TBcyxw1RDf4zbx7+ogFbYvaOEACeeGMavOSwFMEabNvQTqxRiaI
fMfFMJhdvT4SxjAXhKuaf3d6RYNAP4cLBf5zEzLHm0+xfYdPi6ATDEIabY2kXAj8
h6N/qOarjVCbtQrY4zrUZxJ5xW6UZ4nkTzmWFgfoPUJh0K/Ks2VyLXG9Yquq0sXf
c5TbBb/gM71E6vKBI8s9BfpAsAPzgpgH5bomZXaaA5gUZ6q6m1/4QpZCVSUDKaxm
xEOFpHovm4BkDWIVYUzu5bAHUJ5gEWQjDu6NqWRofMiWMMOvnrIOL91us5aK00sF
XrxR8T94mdfGZFAaEu0Li0ks2YnUC2ZT/GxzX99qfJEeOa87CzN1kGqak8cKSOuz
VonVqzrEbDShQmeZsFuH8YR5RaHSix9TR1yTsUfxfIeHOEtjXnDdaycBsld6wmbT
qYVZ5oLqRv86WmUpaKzQ11/46I4nDTuUWZXcCgqpaFElK4Xiztmx0ez22ypCw33i
xKcrwTUYSu1xOqnu4GVjtwva52FBLbDG6krRUIkbZhY+BA0AbWK2mzcDHkz054O/
ohxxTCJjc+b57ktqFaY1vybpMboAK9UXEf0VLCwwkN0IG85z0CsIWlJ4xE7RiK9z
Hx+i1WaSHabWheQAwaR2y+3GkZawuWnDxvkmtL/c4iAjvh8jzIo2HyzCzZm1F+oq
LtpnWb6UPx0L4tfgTfA27S+86dD6FjKiEVwgot0QMDH9vY7yItaXclmVdhxpYNFC
7OdD9Te2cR5b0kS8znSL54R0rRAeKHRbNNW6YrGvrGv8v+hDjKmnIcwgpU5e80Ic
3BBiZV+JcqIXcUIa5FFzlWjkZ/LFuLDFEKvhk+9VyAsEF4Cjp/a1Bw4UNhsfqcOb
kG7uzJVX+jQXHmer9n57oA34ee/oXiZCmpMQOuxF2/PQ1hE5OCobg1KLlHIQ3I0v
pA3LKlC1YyuU7PiTKZs7K9zOxrSlQTYslXqV7vjeRDEslTz66Gjzt2HZP3WzVJU1
pIpoUvmCv1YGd42/DnzOfECpx88uoC7W2flD9H9Y364eYtmEWrGuykOYpX/tUhBM
owYX25mG073NPn+XrlM+kzmvzVt/yshTISFdSaqeZDDJgjTfUGkfDL6Wczk/6qAX
7x9yBFANASlBKt76l7ZrgA1oaUIqgasvtfCwKctVqHfAQqZrxJZAPKEnk5zPTD4C
8/vfthtQJF0cUxP5LIQje3dQbkh/EeRyp1sYbE6Xxr9hWYREwYYQbBSehT8ta228
NjaPvVF3cx4MQV5H4j7iHn4geB8HJ3xB1BLJoWwZngvNYRCKC1hg//Z5RLc3KZlh
XrVBekYWMo1esklsJtup19njeH917qooT9fUxmqjbAuZHI06E3Z4/bLHMk4Tm3rp
fo7foFJnf7snjqxzF9HzsqEPwZeEgfRplEDRj5h5AgvAh0043+3WeLupLHjt1rB6
1H2lMoxfMS2ExeQtEMLIvR4+At3yhBH9rmrVwkJrBwLKwdvp1Tll0UXaOIl4Dw78
UL364qfDjlCRFxBIaJmNEkI0Az5RG4CDFW4oP99LyTomQWLgE1Tdf+i89qYp9cyv
hHQrN7EkHcBau8DQcrEICwjHV097ip+IYLRvUdsLxWuGQZvYCQ7ZpVxy80Z6PnXB
w23ndZNRGmD45wtJvKnT6S2enrUR2veLBWJuqwcmfvbtmxciPsPH75i8mUrVeGhd
StT1SLWDExYNiyWtZmal2YJNDSlSE3U6k2VxSs9YV1lh3OWU0VI2ooSZVMqJAI7Z
ZRsEd7wtMNf4sSTbl9pogYQoeA65Wl/0Eg+dayrADTBKfqzyY8GjWR1EdDRRvKGs
KljXjp1ZRPonE3LkkHmtMtdZog3bdrxhPmThn2JHY/Fdxqf/aiVeJ7mlSsUiKeHy
OlY8dvvNn5wRzvZlF7Wds30FeMLrsQ9CcFxOFDbIh1FiXNi6K1INyB9mcO2eddpn
IqYdXZNX62hbmzWXcg6KHyeVSZnH5CbUN/CGp99EAqPqBns4GdwMs+b0N2p2OEzT
qLfv0qze3Hr8/0jdRQI0mljbOmighZzmNubiG5YEMhPvpeGLbAuEhv3PdPc+hWhF
/L03Fo3yr3M+NXF+6LRw1DKjtpdxOpQ4Bj2NvPqUVvQjnGB9tVeD9YbxCydm6P1O
8eYV4dFIlsDRJCbalcZgva9mq+JjQgQccpbpO0aX/0tQyrAwsEP4IED2klwWzf7p
bNJ9RUzt9pbw4ajcTdKMv8qqaXKgea2hDqOb3JC4yxkpN/0DS+6Ikaco4CT5exmD
McmRUndz1C8TTDkHPb7sgK6wCOmixKKwWIyixiad100EE3YssppJqP2zs4AdA8vV
wj/RdLQuitYG9P5mpNorEaJHaeOwDkJTl5SfevjO4bNl5QLhshrV+3+CU00MlXeW
2wsmc+4PGYapvZRg+S72uV6OScXrISNIlcKGjS2tbu0xiclXkohvlo/ioox7VR5V
4jP57USTOW7YCj0lxnMux703Opb0xUUYNn/odewEKtLIyxe+420SG+eDDXTeuX+O
0tpUhRLFKcnE0C9KpFB/Evdovu8gBz9P6t0K/BMoOkKyRsj1dmAkuQibhA8kQc/i
cU0O5nuOJrUokyMSbGp0DhOnwltftezjiJkVKm4SZoIZlUTKbXCA16uSFNlNh/Au
Pf9aPovWkBYQeByCa68lLeri3W8XBEgFvgcy4cdOxHra/VkpES12TA/915mbcB+6
ReKuTpq11iLpDZZbuNaFIk0XKOD8LijLmfWdHvxRldrIwSwaWFwkNi80doc0Q0Ky
RD2vLqDN8C72ZN0yAPdhvt9AYeY1nQKGYFCDJfWfx0VgljNB4NXgDkIltl+hhG8X
mgpwuW0tM98wIobvyidGfNnkfR5yT+3B6RBn4Pq3QljNSRuOQvkZq9YQnoRwhe7L
+otrRX70g/AIfiaasXeEoIyS+8FBDheBbNF40Qewo0MyZj3ChH/QKFKcTqmulJml
9GRXqIJqGbUmUXH5o7XBkw1jGJgokl3ahGHEJAxB0D+wgPvfuzTSZSR6dja2ZI1A
eHSZchSnHO7xD5EV6DCT182gwI1yEijad8WV0RvAkgQrW8vAT2Tev6IcQOi3mRPr
uxi0X8wHLh9I7TaF88iId9w6RHG7+myAAAhwWJrwCkGy3X46fy7FV43aQQT/cLp2
qaNyUmSFFsJYLS391zFjuMsnEH86ClAD33akLoKhT6LwhYNtLEjUGJDaHuJ+oGpJ
zhvF2KI7z4PogXukDA8gFdHfVe37WDobC0nF45RzjKVc0dea1i1FHPOZuoOSUd6l
sPPpB5NHpTJ+WXWGEmwdBHagyAuIq0pXCwg/n5dwnpQNxeLIrR/LuBldCKx5fAZK
pLCAm625drqzhFcAsIfemA+rW3Woy1InURZU9jXdaIQp9bhRELLX8Ajzmucrq+fF
ZZ7+wK74vgMMaS9v+fWkiOtS3Hui2JCo1GWgso6zLBaH22ehxTzMFF2kR/lOjQPt
urCxzwnsB/WuuWBBG7SoE+cfTstkFBEQkpYyufdITdFOyYJ2SnSP0k8S+IBvGamX
ZJkDhwUPRR/n3i8gF+DrANL8ZbHaXhWLvoSod70L4ESGIb5L528757y0jhIAZLNw
Gw8p+qDh7iWUfLPb9MWSeVy3G+k6pOt/fHOl+oq8DHF0DESIyUNdm5nnOXvyM2ia
f/wVL9ZgfSWfvbG3y/uesEAASK0dnhIU8DkNcO/Pkt2xtKyuzrCO1SIRh+KGw7IC
jHX3kEoi9kNBayeKYqi9NoPEAYl8smEu+Torqm8SQGmOzkGhQ0TuhswH3Xxt1D/C
qTPCg3rQLI4ackcsRDEIEWYOhbpaiqlxV166uzpaL/vw8F5TZ7bKKfYv2hAV6Bls
SSwInt4B3TX7OyjtosI2ioItI4A1ENb5a3PSGKJsgBFx0kbI/xiDyEzS71OLsgjy
CO6TjOea8nPWxhwnJO7DAiTkP0kOZgo1BrecMBrvLFF1EFFSj2WicygMcPHSj7WY
CKiT00llodbk3pbhIkoBYgcHKsRMenR5JCVt8c8iOXQ8OE7iQHC6nBDhAlYWueIe
ey79sJe+NBvzosVIDtWdj4ADC9oJM3bmgT5zSoP0bYeKCOw2HxFCrApX9b99yCoM
+kQlP/zqoE8ahjzyM2GeHjtgol6RMm3SyVOd8cp7TdiE9SHCNRJrMTpQb1/guuZA
6zOCdwZ0WfbTUm5Mad3FuJad3graZECILahj9Q5awhmIf8mly25tqBbIFE55ZSDB
qQfsnTBMuzpnboGEZJalbUt9KqeeJutiK3SIyAnuTIDl2d8tbONaEGpJt084gxJF
h0kus0HamZ2/eTZl7gdIqPC/YAIswuchCBv2WAOGTb7XnzVB8AktueU660GvCufT
faPtHldQ+IKD6Cq0MkNrP2wgqcS9aTeHuCa9yFxvK0H4YbbH7lst5gP4skiUKGZZ
q1llUDb756yFSap7BFBTOZOrq9oovytPLt0mQkxAZwQ3kVpMod21hzPkfovDyuoU
5dFLUef6wIWwd4e96RoHDsONsKu1IUE8dzWTe0GpYJl0PK4uclpBdtUcS2RF99Z3
BxbtVKbR4xikLUpFHPqG1PRl9hkqd1O/x+dqWbLTZguItikUjX1NwOfP1JHMdZ1w
21gwfiXDThv21fSR+4kWJai1q1sYSlutif9cqZUr1yQYKGQb2SZtjgHsVulymOX9
IFoYGOR2td3IKoxqiovValSx6I8dHN4MO0P8hxCJOhXqBBLLKCJI+QJIfSxuJx1h
MKzPWzqvBh8YG72e9dd/estbfw+ELraSepobBxHoWtesCNQ8JT363xQ7bIq1UdbM
hTiPcUP4XBpTvNsSECPZzlmQEh7YTozSeOa4vm6u0ODn39IjYhGAEcRoyOWMCHHp
nRXnlUbYC7JIqbz4XFdmnNEda1MAfZdL9JSDKsIwtKN0C9Lq1f5E1ZT6zRsP9WUV
9Fd5w0St5sh1truTvR4LWsKFd3fpb36Z2+hubMl3lZ9o6thv4cGP7fJeHHRnx+qo
TgY/n5evCmHMVMD/U1J1Eaz/Aqkxo8GbPLI/J4Z94gfaoiF13EBOVEvfELWQT9QL
cSlb2SSImkgbt+9h16fixVyAsjGaD8v+X+4u+bJlDo4+rsHw6jlVLYBoXZd25SoB
nGG0a+mOeSGwYOAWC+sf1mqPRg+zDgElMh96/ZsmDiQEpkIogQkr3npTsqptviEo
A/4SQ8kgDmgVzLHSWOfHe12WalCibZKIuDEZH6LVL6GyA6r2eBE31fDyZfG4eSIo
Oyvi5QI5IdzK7BNWVVbvSgphtkWMjAG/f98EmvMJGAm97RnTT6t02EKD0Wc++Rt0
e2ehTVZm7KQcDC4lbpH/y7KzE7Hk5mPlwTUfagPhMQCg8P4rFlCF9Hy+4zjg8YaS
kx3CRcygy9kaTvnROLMUviUFkQOwCIIp+ptDtshRHRw3Gfuy3IpdkPwgMeqqvpIW
F0CY0kP/c0FzezASWV7Qka/k9MK8QzZfxqBpwYv+auVMxaRYxDEb41CAIdhCfrw1
`protect end_protected
